

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238;

  NAND2_X1 U3466 ( .A1(n6041), .A2(n6043), .ZN(n6031) );
  AND2_X1 U3467 ( .A1(n6085), .A2(n3489), .ZN(n6041) );
  AND2_X1 U34680 ( .A1(n6007), .A2(n5211), .ZN(n6994) );
  OR2_X1 U34690 ( .A1(n6769), .A2(n5206), .ZN(n6107) );
  AND2_X1 U34700 ( .A1(n4068), .A2(n4067), .ZN(n7026) );
  CLKBUF_X2 U34710 ( .A(n4332), .Z(n3447) );
  CLKBUF_X2 U34720 ( .A(n3698), .Z(n3434) );
  CLKBUF_X2 U34730 ( .A(n3680), .Z(n4679) );
  CLKBUF_X2 U34740 ( .A(n3856), .Z(n3798) );
  INV_X1 U3475 ( .A(n4097), .ZN(n3511) );
  AND2_X1 U3476 ( .A1(n3830), .A2(n3720), .ZN(n3748) );
  NAND4_X1 U3477 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n4246)
         );
  NAND2_X2 U3478 ( .A1(n3578), .A2(n3665), .ZN(n3666) );
  CLKBUF_X3 U3479 ( .A(n4658), .Z(n3457) );
  AND2_X1 U3480 ( .A1(n5005), .A2(n4821), .ZN(n3693) );
  AND2_X1 U3481 ( .A1(n4810), .A2(n5019), .ZN(n3680) );
  AND2_X1 U3482 ( .A1(n5005), .A2(n5032), .ZN(n3698) );
  AND2_X1 U3483 ( .A1(n4821), .A2(n3587), .ZN(n4332) );
  NAND2_X1 U3484 ( .A1(n4125), .A2(n4202), .ZN(n4898) );
  INV_X1 U3485 ( .A(n7008), .ZN(n6998) );
  AND2_X1 U3486 ( .A1(n6007), .A2(n5218), .ZN(n7008) );
  AND2_X1 U3487 ( .A1(n4789), .A2(n4788), .ZN(n4874) );
  AND2_X1 U3488 ( .A1(n4404), .A2(n4398), .ZN(n5836) );
  INV_X1 U3489 ( .A(n7015), .ZN(n7006) );
  INV_X1 U3490 ( .A(n7017), .ZN(n6999) );
  XNOR2_X1 U3491 ( .A(n4204), .B(n3513), .ZN(n6128) );
  AND2_X1 U3492 ( .A1(n6198), .A2(n4005), .ZN(n3433) );
  NAND2_X2 U3493 ( .A1(n4001), .A2(n4000), .ZN(n6211) );
  NAND2_X2 U3494 ( .A1(n6256), .A2(n3999), .ZN(n4001) );
  AND2_X2 U3495 ( .A1(n3719), .A2(n4246), .ZN(n3726) );
  XNOR2_X2 U3497 ( .A(n3795), .B(n3797), .ZN(n5972) );
  NAND4_X4 U3498 ( .A1(n3655), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3718)
         );
  AND4_X2 U3499 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(n3654)
         );
  NAND2_X2 U3500 ( .A1(n3923), .A2(n3922), .ZN(n3924) );
  INV_X4 U3501 ( .A(n6368), .ZN(n6369) );
  CLKBUF_X2 U3502 ( .A(n7193), .Z(n7197) );
  NAND2_X1 U3503 ( .A1(n3897), .A2(n3896), .ZN(n5042) );
  NAND2_X2 U3505 ( .A1(n3830), .A2(n4098), .ZN(n4103) );
  AND4_X1 U3506 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n3690)
         );
  BUF_X1 U3508 ( .A(n3705), .Z(n3459) );
  AOI21_X1 U3509 ( .B1(n6017), .B2(n6254), .A(n4734), .ZN(n4735) );
  XNOR2_X1 U3510 ( .A(n3571), .B(n4723), .ZN(n6017) );
  NAND2_X1 U3511 ( .A1(n3539), .A2(n3538), .ZN(n6205) );
  AOI21_X1 U3512 ( .B1(n6134), .B2(n6102), .A(n6086), .ZN(n7214) );
  INV_X1 U3513 ( .A(n6750), .ZN(n7211) );
  NAND2_X1 U3514 ( .A1(n3992), .A2(n5844), .ZN(n3444) );
  CLKBUF_X1 U3515 ( .A(n3504), .Z(n3454) );
  AOI21_X1 U3516 ( .B1(n3549), .B2(n3551), .A(n3547), .ZN(n3546) );
  AOI21_X1 U3517 ( .B1(n4751), .B2(n6873), .A(n4750), .ZN(n4752) );
  NOR2_X1 U3518 ( .A1(n5445), .A2(n4362), .ZN(n5672) );
  OAI21_X1 U3519 ( .B1(n5743), .B2(n3551), .A(n5733), .ZN(n3550) );
  NOR2_X1 U3520 ( .A1(n3556), .A2(n3553), .ZN(n3552) );
  OAI21_X1 U3521 ( .B1(n6128), .B2(n6794), .A(n3480), .ZN(n3506) );
  AND2_X1 U3522 ( .A1(n4771), .A2(n4770), .ZN(n4772) );
  INV_X1 U3523 ( .A(n3990), .ZN(n3551) );
  OAI21_X1 U3524 ( .B1(n3471), .B2(n4743), .A(n4742), .ZN(n4204) );
  NAND2_X1 U3525 ( .A1(n3471), .A2(n4208), .ZN(n4742) );
  NOR2_X1 U3526 ( .A1(n6056), .A2(n6045), .ZN(n6044) );
  NOR2_X1 U3527 ( .A1(n6056), .A2(n3520), .ZN(n4768) );
  OAI21_X1 U3528 ( .B1(n4283), .B2(n4221), .A(n3947), .ZN(n3948) );
  OAI21_X1 U3529 ( .B1(n4283), .B2(n4419), .A(n4282), .ZN(n4848) );
  NAND2_X1 U3530 ( .A1(n3961), .A2(n3960), .ZN(n3982) );
  NAND2_X1 U3531 ( .A1(n4260), .A2(n4875), .ZN(n4878) );
  NOR2_X1 U3532 ( .A1(n5857), .A2(n4884), .ZN(n6378) );
  CLKBUF_X1 U3533 ( .A(n4244), .Z(n3463) );
  AND2_X1 U3534 ( .A1(n4235), .A2(n4234), .ZN(n6818) );
  NAND2_X1 U3535 ( .A1(n4913), .A2(n7096), .ZN(n3897) );
  CLKBUF_X1 U3536 ( .A(n4913), .Z(n5387) );
  NAND2_X2 U3538 ( .A1(n6706), .A2(n4868), .ZN(n6156) );
  NAND2_X1 U3539 ( .A1(n3864), .A2(n3863), .ZN(n3876) );
  XNOR2_X1 U3540 ( .A(n5022), .B(n5020), .ZN(n4913) );
  MUX2_X1 U3541 ( .A(n5203), .B(n4869), .S(n4870), .Z(n4788) );
  OR2_X1 U3542 ( .A1(n3880), .A2(n3879), .ZN(n5022) );
  XNOR2_X1 U3543 ( .A(n3880), .B(n3878), .ZN(n4975) );
  AOI21_X1 U3544 ( .B1(n5972), .B2(n7096), .A(n3813), .ZN(n3829) );
  NAND2_X1 U3545 ( .A1(n3884), .A2(n3883), .ZN(n5020) );
  NAND2_X1 U3546 ( .A1(n3848), .A2(n3847), .ZN(n3878) );
  OAI22_X1 U3547 ( .A1(n4773), .A2(n3755), .B1(n3754), .B2(n4862), .ZN(n3756)
         );
  AND2_X1 U3548 ( .A1(n4117), .A2(n4116), .ZN(n4896) );
  AND4_X1 U3549 ( .A1(n3484), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3745)
         );
  NOR2_X1 U3550 ( .A1(n4073), .A2(n3501), .ZN(n3500) );
  AND3_X1 U3551 ( .A1(n3790), .A2(n3789), .A3(n3788), .ZN(n3793) );
  NAND2_X1 U3552 ( .A1(n3850), .A2(n3849), .ZN(n4063) );
  CLKBUF_X1 U3553 ( .A(n3739), .Z(n3448) );
  OR2_X1 U3554 ( .A1(n4203), .A2(EBX_REG_1__SCAN_IN), .ZN(n4108) );
  OR2_X1 U3555 ( .A1(n4030), .A2(n4103), .ZN(n4812) );
  NAND2_X1 U3556 ( .A1(n4791), .A2(n4202), .ZN(n4195) );
  AND2_X1 U3557 ( .A1(n4075), .A2(n4099), .ZN(n3754) );
  INV_X1 U3558 ( .A(n4044), .ZN(n4052) );
  AND2_X1 U3559 ( .A1(n3747), .A2(n3746), .ZN(n3749) );
  NAND2_X1 U3560 ( .A1(n4035), .A2(n4944), .ZN(n4862) );
  NAND3_X1 U3561 ( .A1(n4755), .A2(n4097), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4044) );
  OR2_X1 U3562 ( .A1(n3786), .A2(n3785), .ZN(n3983) );
  CLKBUF_X1 U3563 ( .A(n4246), .Z(n4868) );
  OR2_X1 U3564 ( .A1(n3774), .A2(n3773), .ZN(n3866) );
  OR2_X1 U3565 ( .A1(n3808), .A2(n3807), .ZN(n3865) );
  AND2_X1 U3566 ( .A1(n4246), .A2(n3718), .ZN(n4091) );
  OR2_X2 U3567 ( .A1(n3679), .A2(n3678), .ZN(n3830) );
  NAND2_X2 U3568 ( .A1(n4098), .A2(n4097), .ZN(n5221) );
  NAND4_X2 U3569 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n4097)
         );
  AND4_X1 U3570 ( .A1(n3589), .A2(n3590), .A3(n3591), .A4(n3588), .ZN(n3592)
         );
  AND4_X1 U3571 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3716)
         );
  AND4_X1 U3572 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3653)
         );
  AND2_X1 U3573 ( .A1(n3621), .A2(n3449), .ZN(n3633) );
  AND4_X1 U3574 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3632)
         );
  AND4_X1 U3575 ( .A1(n3664), .A2(n3663), .A3(n3662), .A4(n3661), .ZN(n3665)
         );
  AND4_X1 U3576 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3691)
         );
  AND4_X1 U3577 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3631)
         );
  AND4_X1 U3578 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3612)
         );
  AND4_X1 U3579 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3578)
         );
  AND4_X1 U3580 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(n3611)
         );
  AND4_X1 U3581 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(n3613)
         );
  AND4_X1 U3582 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3717)
         );
  AND4_X1 U3583 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), .ZN(n3714)
         );
  AND4_X1 U3584 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3634)
         );
  AND3_X1 U3585 ( .A1(n3622), .A2(n3620), .A3(n3619), .ZN(n3449) );
  AND4_X1 U3586 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3652)
         );
  BUF_X4 U3587 ( .A(n4674), .Z(n3469) );
  BUF_X4 U3588 ( .A(n4658), .Z(n3456) );
  BUF_X2 U3589 ( .A(n3673), .Z(n4698) );
  BUF_X2 U3590 ( .A(n3855), .Z(n3776) );
  BUF_X2 U3591 ( .A(n3672), .Z(n4697) );
  AND2_X2 U3592 ( .A1(n4809), .A2(n5005), .ZN(n3465) );
  OR2_X2 U3593 ( .A1(n7116), .A2(n6401), .ZN(n6398) );
  AND2_X2 U3594 ( .A1(n4809), .A2(n5005), .ZN(n4485) );
  AND2_X2 U3595 ( .A1(n4810), .A2(n3587), .ZN(n4658) );
  AND2_X2 U3596 ( .A1(n5032), .A2(n5019), .ZN(n3470) );
  AND2_X2 U3597 ( .A1(n5032), .A2(n5019), .ZN(n3660) );
  AND2_X2 U3598 ( .A1(n3510), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4809)
         );
  AND2_X4 U3599 ( .A1(n4821), .A2(n5019), .ZN(n3681) );
  NOR2_X1 U3600 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5203) );
  AND2_X2 U3601 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4821) );
  NOR2_X2 U3602 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3587) );
  NAND2_X1 U3603 ( .A1(n5847), .A2(n3438), .ZN(n3435) );
  NAND2_X1 U3604 ( .A1(n3435), .A2(n3436), .ZN(n5945) );
  OR2_X1 U3605 ( .A1(n3437), .A2(n3443), .ZN(n3436) );
  INV_X1 U3606 ( .A(n3441), .ZN(n3437) );
  AND2_X1 U3607 ( .A1(n5845), .A2(n3441), .ZN(n3438) );
  NAND2_X1 U3608 ( .A1(n6198), .A2(n4005), .ZN(n3439) );
  NAND2_X1 U3609 ( .A1(n6198), .A2(n4005), .ZN(n3440) );
  NAND2_X1 U3610 ( .A1(n5837), .A2(n4404), .ZN(n5868) );
  OR2_X1 U3611 ( .A1(n3442), .A2(n3552), .ZN(n3441) );
  INV_X1 U3612 ( .A(n3554), .ZN(n3442) );
  AND2_X1 U3613 ( .A1(n5844), .A2(n3554), .ZN(n3443) );
  AND2_X2 U3614 ( .A1(n6000), .A2(n4810), .ZN(n3672) );
  INV_X2 U3616 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3581) );
  OR2_X2 U3617 ( .A1(n3967), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5606)
         );
  AND2_X1 U3618 ( .A1(n3874), .A2(n3873), .ZN(n3450) );
  OR2_X1 U3619 ( .A1(n4739), .A2(n4738), .ZN(n3451) );
  NAND2_X1 U3620 ( .A1(n3451), .A2(n4737), .ZN(n4740) );
  OAI21_X1 U3621 ( .B1(n3440), .B2(n4009), .A(n6174), .ZN(n3452) );
  OAI21_X1 U3622 ( .B1(n3439), .B2(n4009), .A(n6174), .ZN(n3453) );
  OAI21_X1 U3623 ( .B1(n3439), .B2(n4009), .A(n6174), .ZN(n4739) );
  NOR2_X2 U3624 ( .A1(n5891), .A2(n5925), .ZN(n5917) );
  AND2_X1 U3625 ( .A1(n3923), .A2(n3922), .ZN(n3455) );
  NAND2_X1 U3626 ( .A1(n5483), .A2(n3988), .ZN(n3504) );
  NAND2_X2 U3627 ( .A1(n6263), .A2(n3997), .ZN(n6256) );
  INV_X2 U3628 ( .A(n3666), .ZN(n3720) );
  AND2_X2 U3629 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5019) );
  AND2_X2 U3630 ( .A1(n3509), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n6000)
         );
  NOR2_X2 U3631 ( .A1(n5918), .A2(n3564), .ZN(n6100) );
  XNOR2_X1 U3632 ( .A(n3982), .B(n3970), .ZN(n4300) );
  NAND2_X1 U3633 ( .A1(n4811), .A2(n7096), .ZN(n3502) );
  AND2_X2 U3634 ( .A1(n6000), .A2(n5032), .ZN(n3458) );
  BUF_X8 U3636 ( .A(n3705), .Z(n3460) );
  AND2_X2 U3637 ( .A1(n3587), .A2(n5032), .ZN(n3705) );
  AND2_X2 U3638 ( .A1(n4034), .A2(n4097), .ZN(n3821) );
  XNOR2_X2 U3639 ( .A(n3924), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5137)
         );
  NAND2_X2 U3640 ( .A1(n3503), .A2(n4004), .ZN(n6198) );
  AND2_X2 U3641 ( .A1(n3511), .A2(n4034), .ZN(n4035) );
  AND2_X1 U3642 ( .A1(n3512), .A2(n4034), .ZN(n3737) );
  INV_X2 U3643 ( .A(n4098), .ZN(n4034) );
  INV_X2 U3644 ( .A(n3718), .ZN(n3746) );
  NOR2_X2 U3645 ( .A1(n4853), .A2(n4855), .ZN(n4845) );
  INV_X4 U3646 ( .A(n6368), .ZN(n3461) );
  INV_X2 U3647 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3510) );
  NOR2_X2 U3648 ( .A1(n6031), .A2(n3569), .ZN(n4764) );
  OAI21_X2 U3649 ( .B1(n6737), .B2(n6740), .A(n6738), .ZN(n5847) );
  OAI21_X2 U3650 ( .B1(n5945), .B2(n3996), .A(n3995), .ZN(n6263) );
  BUF_X1 U3651 ( .A(n4914), .Z(n3462) );
  XNOR2_X1 U3652 ( .A(n3875), .B(n3876), .ZN(n4244) );
  AND2_X1 U3653 ( .A1(n4809), .A2(n5005), .ZN(n3464) );
  BUF_X8 U3654 ( .A(n3699), .Z(n3467) );
  AND2_X2 U3655 ( .A1(n5005), .A2(n4810), .ZN(n3699) );
  BUF_X8 U3656 ( .A(n4674), .Z(n3468) );
  AND2_X1 U3657 ( .A1(n4809), .A2(n3587), .ZN(n3856) );
  AND2_X2 U3658 ( .A1(n3582), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4810)
         );
  AND2_X4 U3659 ( .A1(n6000), .A2(n5032), .ZN(n3700) );
  NOR2_X4 U3660 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5032) );
  AND2_X4 U3661 ( .A1(n3581), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5005)
         );
  OR2_X1 U3662 ( .A1(n7026), .A2(n7073), .ZN(n4780) );
  OR2_X1 U3663 ( .A1(n4755), .A2(n7096), .ZN(n3849) );
  AOI21_X1 U3664 ( .B1(n3469), .B2(INSTQUEUE_REG_14__0__SCAN_IN), .A(n3709), 
        .ZN(n3715) );
  NAND2_X1 U3665 ( .A1(n3747), .A2(n3830), .ZN(n3512) );
  INV_X1 U3666 ( .A(n5203), .ZN(n4689) );
  AOI21_X1 U3667 ( .B1(n6174), .B2(n3536), .A(n3487), .ZN(n3535) );
  INV_X1 U3668 ( .A(n3491), .ZN(n3536) );
  NAND2_X1 U3669 ( .A1(n3544), .A2(n3541), .ZN(n3540) );
  NAND2_X1 U3670 ( .A1(n3545), .A2(n3542), .ZN(n3541) );
  NAND2_X1 U3671 ( .A1(n4975), .A2(n7096), .ZN(n3864) );
  OR2_X1 U3672 ( .A1(n6369), .A2(n3998), .ZN(n3999) );
  INV_X1 U3673 ( .A(n4767), .ZN(n3519) );
  NAND2_X1 U3674 ( .A1(n6205), .A2(n6206), .ZN(n3503) );
  NAND2_X1 U3675 ( .A1(n4094), .A2(n4093), .ZN(n4233) );
  INV_X1 U3676 ( .A(n3830), .ZN(n4944) );
  AND2_X1 U3677 ( .A1(n3926), .A2(n3938), .ZN(n3576) );
  INV_X1 U3678 ( .A(n3939), .ZN(n3938) );
  INV_X1 U3679 ( .A(n6058), .ZN(n3557) );
  INV_X1 U3680 ( .A(n4671), .ZN(n4711) );
  AND2_X1 U3681 ( .A1(n4394), .A2(n3573), .ZN(n3572) );
  AND2_X1 U3682 ( .A1(n4393), .A2(n5749), .ZN(n4394) );
  NAND2_X1 U3683 ( .A1(n5672), .A2(n4392), .ZN(n4404) );
  XNOR2_X1 U3684 ( .A(n3925), .B(n3926), .ZN(n4277) );
  INV_X1 U3685 ( .A(n4689), .ZN(n4716) );
  INV_X1 U3686 ( .A(n3994), .ZN(n3556) );
  INV_X1 U3687 ( .A(n5877), .ZN(n3553) );
  OR2_X1 U3688 ( .A1(n3492), .A2(n5871), .ZN(n3516) );
  NAND2_X1 U3689 ( .A1(n3577), .A2(n3735), .ZN(n4214) );
  NAND2_X1 U3690 ( .A1(n4097), .A2(n3720), .ZN(n3735) );
  INV_X1 U3691 ( .A(n3550), .ZN(n3549) );
  NAND2_X1 U3692 ( .A1(n3874), .A2(n3873), .ZN(n3903) );
  NAND2_X1 U3693 ( .A1(n3871), .A2(n3476), .ZN(n3495) );
  NAND2_X1 U3694 ( .A1(n3502), .A2(n3479), .ZN(n3836) );
  OR2_X1 U3695 ( .A1(n3895), .A2(n3894), .ZN(n3919) );
  NAND2_X1 U3696 ( .A1(n3837), .A2(n3836), .ZN(n3875) );
  NAND2_X1 U3697 ( .A1(n3446), .A2(n3843), .ZN(n3880) );
  NOR2_X1 U3698 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4927), .ZN(n4966) );
  AOI22_X1 U3699 ( .A1(n4332), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3674) );
  NOR2_X1 U3700 ( .A1(n3639), .A2(n3638), .ZN(n3655) );
  AND2_X1 U3701 ( .A1(n6107), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6007) );
  OR2_X1 U3702 ( .A1(n6149), .A2(n6250), .ZN(n3566) );
  OR2_X1 U3703 ( .A1(n6979), .A2(n4689), .ZN(n4519) );
  NAND2_X1 U3704 ( .A1(n7121), .A2(n4866), .ZN(n7125) );
  INV_X1 U3705 ( .A(n3569), .ZN(n3567) );
  AND2_X1 U3706 ( .A1(n6068), .A2(n3559), .ZN(n3558) );
  AND2_X1 U3707 ( .A1(n4000), .A2(n4002), .ZN(n3545) );
  AND2_X1 U3708 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n4272), .ZN(n4278)
         );
  OR2_X1 U3709 ( .A1(n6152), .A2(n6151), .ZN(n6358) );
  AND3_X1 U3710 ( .A1(n3980), .A2(n3971), .A3(n3983), .ZN(n3981) );
  OR2_X2 U3711 ( .A1(n5930), .A2(n5921), .ZN(n6152) );
  OR2_X1 U3712 ( .A1(n6369), .A2(n6845), .ZN(n3995) );
  NAND2_X1 U3713 ( .A1(n4896), .A2(n4894), .ZN(n4895) );
  INV_X1 U3714 ( .A(n3834), .ZN(n3497) );
  AND3_X1 U3715 ( .A1(n4807), .A2(n4806), .A3(n4805), .ZN(n7047) );
  INV_X1 U3716 ( .A(n4966), .ZN(n5256) );
  AND2_X1 U3717 ( .A1(n6107), .A2(n5207), .ZN(n7016) );
  NAND2_X1 U3718 ( .A1(n6706), .A2(n6016), .ZN(n6154) );
  OR2_X1 U3719 ( .A1(n6749), .A2(n6709), .ZN(n6755) );
  NAND2_X1 U3720 ( .A1(n7121), .A2(n7062), .ZN(n7033) );
  INV_X1 U3721 ( .A(n4242), .ZN(n4243) );
  INV_X1 U3722 ( .A(n4205), .ZN(n3513) );
  XNOR2_X1 U3723 ( .A(n4016), .B(n4015), .ZN(n4736) );
  OAI211_X1 U3724 ( .C1(n3433), .C2(n3533), .A(n3531), .B(n3527), .ZN(n6279)
         );
  OR2_X1 U3725 ( .A1(n3537), .A2(n3534), .ZN(n3533) );
  NAND2_X1 U3726 ( .A1(n3529), .A2(n3528), .ZN(n3527) );
  NAND2_X1 U3727 ( .A1(n4233), .A2(n4207), .ZN(n6794) );
  INV_X1 U3728 ( .A(n6794), .ZN(n6873) );
  INV_X1 U3729 ( .A(n4812), .ZN(n3501) );
  AND2_X1 U3730 ( .A1(n7043), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4024)
         );
  OR2_X1 U3731 ( .A1(n3937), .A2(n3936), .ZN(n3945) );
  NAND2_X1 U3732 ( .A1(n4034), .A2(n3723), .ZN(n3753) );
  OR2_X1 U3733 ( .A1(n3862), .A2(n3861), .ZN(n3867) );
  INV_X1 U3734 ( .A(n3733), .ZN(n4030) );
  AOI22_X1 U3735 ( .A1(n3673), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U3736 ( .A1(n3673), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U3737 ( .A1(n3660), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U3738 ( .A1(n3673), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3675) );
  AND2_X1 U3739 ( .A1(n3470), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U3740 ( .A1(n3445), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3850) );
  OR2_X1 U3741 ( .A1(n4044), .A2(n4221), .ZN(n4053) );
  OR2_X1 U3742 ( .A1(n4057), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4083)
         );
  AOI22_X1 U3743 ( .A1(n4674), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3588) );
  NAND2_X1 U3744 ( .A1(n3570), .A2(n4762), .ZN(n3569) );
  INV_X1 U3745 ( .A(n6033), .ZN(n3570) );
  NOR2_X1 U3746 ( .A1(n6218), .A2(n3560), .ZN(n3559) );
  INV_X1 U3747 ( .A(n6088), .ZN(n3560) );
  NOR2_X1 U3748 ( .A1(n3563), .A2(n3562), .ZN(n3561) );
  INV_X1 U3749 ( .A(n5870), .ZN(n3562) );
  INV_X1 U3750 ( .A(n3493), .ZN(n3563) );
  NAND2_X1 U3751 ( .A1(n4363), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4399)
         );
  NOR2_X1 U3752 ( .A1(n3574), .A2(n3575), .ZN(n3573) );
  INV_X1 U3753 ( .A(n5196), .ZN(n3574) );
  OR2_X1 U3754 ( .A1(n4873), .A2(n4874), .ZN(n4877) );
  OR2_X1 U3755 ( .A1(n6045), .A2(n3521), .ZN(n3520) );
  INV_X1 U3756 ( .A(n6030), .ZN(n3521) );
  AND2_X1 U3757 ( .A1(n6181), .A2(n4008), .ZN(n6174) );
  OR2_X1 U3758 ( .A1(n5448), .A2(n5198), .ZN(n3518) );
  NAND2_X1 U3759 ( .A1(n3461), .A2(n3986), .ZN(n3987) );
  NAND2_X1 U3760 ( .A1(n3977), .A2(n3976), .ZN(n3978) );
  AND2_X1 U3761 ( .A1(n4850), .A2(n4906), .ZN(n4905) );
  NAND2_X1 U3762 ( .A1(n3844), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3848) );
  INV_X1 U3763 ( .A(n3462), .ZN(n5173) );
  INV_X1 U3764 ( .A(n4811), .ZN(n4974) );
  NAND4_X1 U3765 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n3610), .ZN(n3667)
         );
  NOR2_X1 U3766 ( .A1(n7075), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4725) );
  CLKBUF_X1 U3767 ( .A(n4773), .Z(n4774) );
  NAND2_X1 U3768 ( .A1(n4214), .A2(n3745), .ZN(n3796) );
  NAND2_X1 U3769 ( .A1(n6316), .A2(n4190), .ZN(n6072) );
  OR2_X1 U3770 ( .A1(n5100), .A2(n3518), .ZN(n5676) );
  NOR2_X1 U3771 ( .A1(n4780), .A2(n4779), .ZN(n6613) );
  INV_X1 U3772 ( .A(n4280), .ZN(n4720) );
  AOI21_X1 U3773 ( .B1(n4719), .B2(n4718), .A(n4717), .ZN(n4753) );
  NOR2_X1 U3774 ( .A1(n4651), .A2(n4650), .ZN(n4652) );
  AOI22_X1 U3775 ( .A1(n4649), .A2(n4648), .B1(n5203), .B2(n6050), .ZN(n6043)
         );
  AND2_X1 U3776 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4614), .ZN(n4615)
         );
  INV_X1 U3777 ( .A(n4613), .ZN(n4614) );
  AND2_X1 U3778 ( .A1(n5203), .A2(n6078), .ZN(n4610) );
  NAND2_X1 U3779 ( .A1(n4534), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4535)
         );
  NOR2_X1 U3780 ( .A1(n4535), .A2(n4547), .ZN(n4578) );
  NAND2_X1 U3781 ( .A1(n6144), .A2(n3565), .ZN(n3564) );
  INV_X1 U3782 ( .A(n3566), .ZN(n3565) );
  NOR2_X1 U3783 ( .A1(n4501), .A2(n6252), .ZN(n4502) );
  AND2_X1 U3784 ( .A1(n4502), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4534)
         );
  NOR2_X1 U3785 ( .A1(n4468), .A2(n5940), .ZN(n4469) );
  NAND2_X1 U3786 ( .A1(n4469), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4501)
         );
  AND2_X1 U3787 ( .A1(n4437), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4452)
         );
  NOR2_X1 U3788 ( .A1(n4399), .A2(n5759), .ZN(n4400) );
  NAND2_X1 U3789 ( .A1(n4400), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4421)
         );
  NOR2_X1 U3790 ( .A1(n4347), .A2(n4331), .ZN(n4363) );
  NAND2_X1 U3791 ( .A1(n4330), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4347)
         );
  NOR2_X1 U3792 ( .A1(n4315), .A2(n5242), .ZN(n4330) );
  NAND2_X1 U3793 ( .A1(n4296), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4315)
         );
  CLKBUF_X1 U3794 ( .A(n5096), .Z(n5097) );
  CLKBUF_X1 U3795 ( .A(n4846), .Z(n4847) );
  AND3_X1 U3796 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n4272) );
  AOI21_X1 U3797 ( .B1(n4277), .B2(n4431), .A(n4276), .ZN(n4855) );
  CLKBUF_X1 U3798 ( .A(n4853), .Z(n4854) );
  NAND2_X1 U3799 ( .A1(n3482), .A2(n3496), .ZN(n6719) );
  NAND2_X1 U3800 ( .A1(n6707), .A2(n3835), .ZN(n3498) );
  NAND2_X1 U3801 ( .A1(n3535), .A2(n3534), .ZN(n3532) );
  NAND2_X1 U3802 ( .A1(n3535), .A2(n3530), .ZN(n3529) );
  NAND2_X1 U3803 ( .A1(n3537), .A2(n3534), .ZN(n3530) );
  OR2_X1 U3804 ( .A1(n3535), .A2(n6175), .ZN(n3528) );
  INV_X1 U3805 ( .A(n6175), .ZN(n3534) );
  INV_X1 U3806 ( .A(n6174), .ZN(n3537) );
  NAND2_X1 U3807 ( .A1(n3433), .A2(n3491), .ZN(n6182) );
  NAND2_X1 U3808 ( .A1(n3543), .A2(n3494), .ZN(n3538) );
  AND2_X1 U3809 ( .A1(n6137), .A2(n6090), .ZN(n6316) );
  NOR2_X1 U3810 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  NAND2_X1 U3811 ( .A1(n3508), .A2(n3507), .ZN(n6136) );
  INV_X1 U3812 ( .A(n6105), .ZN(n3507) );
  INV_X1 U3813 ( .A(n6104), .ZN(n3508) );
  NOR2_X2 U3814 ( .A1(n6358), .A2(n6359), .ZN(n6357) );
  OR2_X1 U3815 ( .A1(n3516), .A2(n3515), .ZN(n3514) );
  INV_X1 U3816 ( .A(n5927), .ZN(n3515) );
  AOI21_X1 U3817 ( .B1(n3555), .B2(n3994), .A(n3481), .ZN(n3554) );
  INV_X1 U3818 ( .A(n3993), .ZN(n3555) );
  NOR2_X1 U3819 ( .A1(n5872), .A2(n3516), .ZN(n5928) );
  NAND2_X1 U3820 ( .A1(n3444), .A2(n5877), .ZN(n5876) );
  INV_X1 U3821 ( .A(n6835), .ZN(n6350) );
  INV_X1 U3822 ( .A(n5734), .ZN(n3547) );
  OR2_X1 U3823 ( .A1(n5100), .A2(n5198), .ZN(n5447) );
  NAND2_X1 U3824 ( .A1(n5606), .A2(n3526), .ZN(n3523) );
  INV_X1 U3825 ( .A(n3949), .ZN(n3526) );
  NAND2_X1 U3826 ( .A1(n4123), .A2(n4122), .ZN(n4858) );
  INV_X1 U3827 ( .A(n4856), .ZN(n4122) );
  INV_X1 U3828 ( .A(n4895), .ZN(n4123) );
  AOI21_X1 U3829 ( .B1(n4267), .B2(n3971), .A(n3902), .ZN(n5344) );
  NAND2_X1 U3830 ( .A1(n4899), .A2(n4791), .ZN(n3522) );
  INV_X1 U3831 ( .A(n5221), .ZN(n4791) );
  NAND2_X1 U3832 ( .A1(n4233), .A2(n4822), .ZN(n5878) );
  INV_X1 U3833 ( .A(n3793), .ZN(n3791) );
  NAND2_X1 U3834 ( .A1(n3838), .A2(n3764), .ZN(n3839) );
  NAND2_X1 U3835 ( .A1(n3763), .A2(n3472), .ZN(n3764) );
  INV_X1 U3836 ( .A(n3736), .ZN(n5969) );
  AND2_X1 U3837 ( .A1(n3463), .A2(n4979), .ZN(n5507) );
  NOR2_X1 U3838 ( .A1(n5174), .A2(n5173), .ZN(n5261) );
  INV_X1 U3839 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7043) );
  NOR2_X1 U3840 ( .A1(n5993), .A2(n4974), .ZN(n5389) );
  AOI21_X1 U3841 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7043), .A(n5256), .ZN(
        n5689) );
  AND2_X1 U3842 ( .A1(n5018), .A2(n5017), .ZN(n7059) );
  INV_X1 U3843 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5759) );
  INV_X1 U3844 ( .A(n7009), .ZN(n6980) );
  AND2_X1 U3845 ( .A1(n7001), .A2(n5208), .ZN(n6120) );
  XNOR2_X1 U3846 ( .A(n4111), .B(n4899), .ZN(n6122) );
  AND2_X1 U3847 ( .A1(n6007), .A2(n5222), .ZN(n7015) );
  INV_X1 U3848 ( .A(n6154), .ZN(n6702) );
  INV_X1 U3849 ( .A(n6266), .ZN(n7202) );
  AND2_X1 U3850 ( .A1(n6015), .A2(n5934), .ZN(n7236) );
  NAND2_X1 U3851 ( .A1(n4867), .A2(n7125), .ZN(n6015) );
  OAI21_X1 U3852 ( .B1(n4864), .B2(n4863), .A(n7092), .ZN(n4867) );
  NOR2_X1 U3853 ( .A1(n6631), .A2(n6613), .ZN(n6620) );
  NAND2_X1 U3854 ( .A1(n4001), .A2(n3545), .ZN(n6224) );
  CLKBUF_X1 U3855 ( .A(n5837), .Z(n5838) );
  INV_X1 U3856 ( .A(n6755), .ZN(n6269) );
  INV_X1 U3857 ( .A(n7033), .ZN(n6751) );
  NAND2_X1 U3858 ( .A1(n5466), .A2(n5465), .ZN(n3525) );
  NAND2_X1 U3859 ( .A1(n3834), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4880)
         );
  NAND2_X1 U3860 ( .A1(n3497), .A2(n3835), .ZN(n4881) );
  INV_X1 U3861 ( .A(n3463), .ZN(n5106) );
  AND2_X1 U3862 ( .A1(n5038), .A2(n5256), .ZN(n6399) );
  OR2_X1 U3863 ( .A1(n5215), .A2(n5025), .ZN(n7036) );
  NOR2_X1 U3864 ( .A1(n5536), .A2(n5303), .ZN(n5584) );
  NOR2_X1 U3865 ( .A1(n5397), .A2(n5303), .ZN(n5441) );
  INV_X1 U3866 ( .A(n5335), .ZN(n5569) );
  INV_X1 U3867 ( .A(n5334), .ZN(n5434) );
  AND2_X1 U3868 ( .A1(n5304), .A2(n5303), .ZN(n5433) );
  NOR2_X1 U3869 ( .A1(n6506), .A2(n5256), .ZN(n5694) );
  INV_X1 U3870 ( .A(n7222), .ZN(n5642) );
  NOR2_X1 U3871 ( .A1(n6558), .A2(n5256), .ZN(n5720) );
  NOR2_X1 U3872 ( .A1(n6450), .A2(n5256), .ZN(n5715) );
  NOR2_X1 U3873 ( .A1(n6448), .A2(n5256), .ZN(n5700) );
  INV_X1 U3874 ( .A(n5806), .ZN(n5704) );
  NOR2_X1 U3875 ( .A1(n6504), .A2(n5256), .ZN(n5705) );
  INV_X1 U3876 ( .A(n5813), .ZN(n5709) );
  NOR2_X1 U3877 ( .A1(n6507), .A2(n5256), .ZN(n5726) );
  NAND2_X1 U3878 ( .A1(n5176), .A2(n5303), .ZN(n7217) );
  INV_X1 U3879 ( .A(n5720), .ZN(n5826) );
  INV_X1 U3880 ( .A(n5715), .ZN(n5798) );
  NOR2_X1 U3881 ( .A1(n5119), .A2(n4944), .ZN(n5799) );
  INV_X1 U3882 ( .A(n5710), .ZN(n5805) );
  NOR2_X1 U3883 ( .A1(n5119), .A2(n3614), .ZN(n5806) );
  INV_X1 U3884 ( .A(n5705), .ZN(n5819) );
  INV_X1 U3885 ( .A(n5726), .ZN(n5791) );
  OR2_X1 U3886 ( .A1(n4990), .A2(n4915), .ZN(n5357) );
  INV_X1 U3887 ( .A(n5694), .ZN(n5784) );
  INV_X1 U3888 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7096) );
  NOR2_X1 U3889 ( .A1(n7026), .A2(n7084), .ZN(n7087) );
  INV_X1 U3890 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7077) );
  INV_X1 U3891 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7084) );
  INV_X1 U3892 ( .A(n4760), .ZN(n4761) );
  OAI21_X1 U3893 ( .B1(n5968), .B2(n6154), .A(n3580), .ZN(n4760) );
  OR2_X1 U3894 ( .A1(n6275), .A2(n6154), .ZN(n4771) );
  OAI21_X1 U3895 ( .B1(n6755), .B2(n5227), .A(n4733), .ZN(n4734) );
  OAI21_X1 U3896 ( .B1(n6279), .B2(n7033), .A(n6180), .ZN(U2957) );
  OAI21_X1 U3897 ( .B1(n4736), .B2(n6878), .A(n3505), .ZN(U2987) );
  INV_X1 U3898 ( .A(n3506), .ZN(n3505) );
  INV_X1 U3899 ( .A(n4749), .ZN(n4750) );
  NAND2_X2 U3900 ( .A1(n3746), .A2(n3820), .ZN(n3747) );
  NAND2_X1 U3901 ( .A1(n3720), .A2(n3473), .ZN(n3736) );
  AND2_X1 U3903 ( .A1(n6085), .A2(n3559), .ZN(n6067) );
  OR2_X1 U3904 ( .A1(n5918), .A2(n6149), .ZN(n6148) );
  NAND2_X1 U3905 ( .A1(n5868), .A2(n5870), .ZN(n5869) );
  NAND2_X1 U3906 ( .A1(n3927), .A2(n3576), .ZN(n3962) );
  AND2_X2 U3907 ( .A1(n4809), .A2(n6000), .ZN(n3673) );
  OR3_X1 U3908 ( .A1(n6056), .A2(n3520), .A3(n3519), .ZN(n3471) );
  NAND2_X1 U3909 ( .A1(n6085), .A2(n6088), .ZN(n6087) );
  OR2_X1 U3910 ( .A1(n3762), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3472)
         );
  AND3_X1 U3911 ( .A1(n4755), .A2(n3746), .A3(n4246), .ZN(n3473) );
  OR2_X1 U3912 ( .A1(n3775), .A2(n3849), .ZN(n3474) );
  NOR3_X1 U3913 ( .A1(n5100), .A2(n4145), .A3(n3518), .ZN(n3475) );
  AND2_X1 U3914 ( .A1(n3870), .A2(n3872), .ZN(n3476) );
  NOR2_X1 U3915 ( .A1(n5918), .A2(n3566), .ZN(n3477) );
  NAND2_X1 U3916 ( .A1(n6085), .A2(n3558), .ZN(n6057) );
  OR2_X1 U3917 ( .A1(n6029), .A2(n4741), .ZN(n3478) );
  BUF_X1 U3918 ( .A(n3667), .Z(n4755) );
  INV_X1 U3919 ( .A(n3667), .ZN(n3614) );
  AND2_X1 U3920 ( .A1(n3793), .A2(n3474), .ZN(n3479) );
  AND2_X1 U3921 ( .A1(n3579), .A2(n4243), .ZN(n3480) );
  AND2_X1 U3922 ( .A1(n3461), .A2(n5899), .ZN(n3481) );
  OR2_X1 U3923 ( .A1(n6707), .A2(n3835), .ZN(n3482) );
  OAI22_X1 U3924 ( .A1(n6214), .A2(n6213), .B1(n6368), .B2(n6212), .ZN(n6239)
         );
  AND2_X1 U3925 ( .A1(n3725), .A2(n3740), .ZN(n3483) );
  AND2_X1 U3926 ( .A1(n3727), .A2(n4812), .ZN(n3484) );
  AND2_X1 U3927 ( .A1(n4135), .A2(n4134), .ZN(n5198) );
  NAND2_X1 U3928 ( .A1(n6357), .A2(n6146), .ZN(n6104) );
  AND2_X1 U3929 ( .A1(n5096), .A2(n5196), .ZN(n3485) );
  INV_X1 U3930 ( .A(n6878), .ZN(n6857) );
  NAND2_X1 U3931 ( .A1(n5742), .A2(n3990), .ZN(n5732) );
  NAND2_X1 U3932 ( .A1(n3548), .A2(n3546), .ZN(n6737) );
  NAND2_X1 U3933 ( .A1(n3525), .A2(n3949), .ZN(n5604) );
  NAND2_X1 U3934 ( .A1(n5876), .A2(n3993), .ZN(n5896) );
  INV_X1 U3935 ( .A(n5445), .ZN(n5492) );
  NOR2_X1 U3936 ( .A1(n6175), .A2(n4012), .ZN(n3486) );
  AND2_X1 U3937 ( .A1(n4519), .A2(n4518), .ZN(n6144) );
  AND2_X1 U3938 ( .A1(n3461), .A2(n6280), .ZN(n3487) );
  INV_X1 U3939 ( .A(n3544), .ZN(n3543) );
  OAI21_X1 U3940 ( .B1(n4000), .B2(n3494), .A(n6368), .ZN(n3544) );
  AND2_X1 U3941 ( .A1(n4753), .A2(n3567), .ZN(n3488) );
  AND2_X1 U3942 ( .A1(n3558), .A2(n3557), .ZN(n3489) );
  INV_X1 U3943 ( .A(n4284), .ZN(n4327) );
  INV_X1 U3944 ( .A(n4327), .ZN(n4721) );
  NOR2_X1 U3945 ( .A1(n4974), .A2(n4975), .ZN(n3490) );
  NAND3_X1 U3946 ( .A1(n3733), .A2(n4091), .A3(n3666), .ZN(n4075) );
  NOR2_X1 U3947 ( .A1(n4858), .A2(n4849), .ZN(n4850) );
  NAND2_X1 U3948 ( .A1(n4905), .A2(n5099), .ZN(n5100) );
  NAND2_X1 U3949 ( .A1(n4245), .A2(n4280), .ZN(n4873) );
  NAND2_X1 U3950 ( .A1(n6369), .A2(n4006), .ZN(n3491) );
  OR2_X1 U3951 ( .A1(n5872), .A2(n5871), .ZN(n3517) );
  AND2_X1 U3952 ( .A1(n5985), .A2(n5986), .ZN(n4894) );
  NAND2_X1 U3953 ( .A1(n4156), .A2(n4155), .ZN(n3492) );
  NAND3_X1 U3954 ( .A1(n4436), .A2(n4435), .A3(n4434), .ZN(n3493) );
  INV_X2 U3955 ( .A(n6742), .ZN(n6254) );
  OR2_X1 U3956 ( .A1(n4003), .A2(n6353), .ZN(n3494) );
  INV_X1 U3957 ( .A(n4240), .ZN(n3542) );
  INV_X1 U3958 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3509) );
  NOR3_X2 U3959 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n4987), .ZN(n5152) );
  NAND2_X1 U3960 ( .A1(n6719), .A2(n3495), .ZN(n3874) );
  NAND2_X1 U3961 ( .A1(n3498), .A2(n3834), .ZN(n3496) );
  NAND2_X1 U3962 ( .A1(n3871), .A2(n3870), .ZN(n6720) );
  NAND2_X1 U3963 ( .A1(n3499), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U3964 ( .A1(n3728), .A2(n3500), .A3(n3727), .A4(n3483), .ZN(n3499)
         );
  INV_X1 U3965 ( .A(n3760), .ZN(n3844) );
  NAND2_X1 U3966 ( .A1(n3502), .A2(n3474), .ZN(n3792) );
  NAND2_X1 U3967 ( .A1(n3549), .A2(n3504), .ZN(n3548) );
  OAI21_X1 U3968 ( .B1(n5743), .B2(n3454), .A(n5742), .ZN(n6827) );
  NAND2_X1 U3969 ( .A1(n3454), .A2(n5743), .ZN(n5742) );
  NAND2_X4 U3970 ( .A1(n3691), .A2(n3690), .ZN(n4098) );
  OR2_X2 U3971 ( .A1(n5872), .A2(n3514), .ZN(n5930) );
  INV_X1 U3972 ( .A(n3517), .ZN(n5894) );
  AND2_X2 U3973 ( .A1(n4111), .A2(n3522), .ZN(n5986) );
  NAND3_X1 U3974 ( .A1(n3524), .A2(n5605), .A3(n3523), .ZN(n6733) );
  NAND3_X1 U3975 ( .A1(n5466), .A2(n5606), .A3(n5465), .ZN(n3524) );
  OR2_X1 U3976 ( .A1(n3439), .A2(n3532), .ZN(n3531) );
  NAND2_X1 U3977 ( .A1(n4001), .A2(n3540), .ZN(n3539) );
  NAND2_X1 U3978 ( .A1(n5868), .A2(n3561), .ZN(n5891) );
  NOR2_X1 U3979 ( .A1(n6031), .A2(n6033), .ZN(n4763) );
  NAND2_X1 U3980 ( .A1(n3568), .A2(n3488), .ZN(n3571) );
  INV_X1 U3981 ( .A(n6031), .ZN(n3568) );
  NAND2_X1 U3982 ( .A1(n5096), .A2(n3572), .ZN(n4397) );
  NAND2_X1 U3983 ( .A1(n5096), .A2(n3573), .ZN(n5445) );
  INV_X1 U3984 ( .A(n5446), .ZN(n3575) );
  NAND2_X1 U3985 ( .A1(n3927), .A2(n3926), .ZN(n3940) );
  INV_X1 U3986 ( .A(n3962), .ZN(n3961) );
  AND2_X1 U3987 ( .A1(n3732), .A2(n3734), .ZN(n3577) );
  NOR2_X1 U3988 ( .A1(n4230), .A2(n4732), .ZN(n3579) );
  AND2_X1 U3989 ( .A1(n4759), .A2(n7092), .ZN(n6706) );
  INV_X1 U3990 ( .A(n6706), .ZN(n4769) );
  AOI21_X1 U3991 ( .B1(n4293), .B2(n4431), .A(n4292), .ZN(n4904) );
  INV_X1 U3992 ( .A(n4904), .ZN(n4294) );
  OR2_X1 U3993 ( .A1(n6706), .A2(n5961), .ZN(n3580) );
  INV_X1 U3994 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4015) );
  NAND2_X1 U3995 ( .A1(n3820), .A2(n4098), .ZN(n4221) );
  INV_X1 U3996 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4010) );
  INV_X1 U3997 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3835) );
  INV_X1 U3998 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7054) );
  INV_X1 U3999 ( .A(n3866), .ZN(n3775) );
  OR3_X1 U4000 ( .A1(n4041), .A2(n4040), .A3(n4039), .ZN(n4047) );
  NAND2_X1 U4001 ( .A1(n3698), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3649) );
  NAND2_X1 U4002 ( .A1(n3468), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3643)
         );
  OR2_X1 U4003 ( .A1(n3959), .A2(n3958), .ZN(n3972) );
  AOI22_X1 U4004 ( .A1(n3693), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4658), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3586) );
  INV_X1 U4005 ( .A(n4221), .ZN(n3971) );
  OR2_X1 U4006 ( .A1(n6369), .A2(n5899), .ZN(n3994) );
  OR2_X1 U4007 ( .A1(n3916), .A2(n3915), .ZN(n3942) );
  INV_X1 U4008 ( .A(n4393), .ZN(n4362) );
  OR2_X1 U4009 ( .A1(n4715), .A2(n6022), .ZN(n4729) );
  OR2_X1 U4010 ( .A1(n4609), .A2(n4608), .ZN(n4613) );
  INV_X2 U4011 ( .A(n4203), .ZN(n4191) );
  AND2_X1 U4012 ( .A1(n4154), .A2(n4153), .ZN(n5871) );
  AND2_X1 U4013 ( .A1(n4121), .A2(n4120), .ZN(n4856) );
  INV_X1 U4014 ( .A(n4053), .ZN(n4066) );
  NAND2_X1 U4015 ( .A1(n4615), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4651)
         );
  OR2_X1 U4016 ( .A1(n6369), .A2(n6300), .ZN(n4004) );
  AND2_X1 U4017 ( .A1(n5398), .A2(n5764), .ZN(n5401) );
  INV_X1 U4018 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5534) );
  OAI21_X1 U4019 ( .B1(n5828), .B2(n7084), .A(n5775), .ZN(n5827) );
  AOI21_X1 U4020 ( .B1(n6766), .B2(n4911), .A(n7087), .ZN(n4927) );
  NOR2_X1 U4021 ( .A1(n4421), .A2(n4420), .ZN(n4437) );
  INV_X1 U4022 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5242) );
  INV_X1 U4023 ( .A(n6994), .ZN(n7010) );
  INV_X1 U4024 ( .A(n4753), .ZN(n4754) );
  NAND2_X1 U4025 ( .A1(n4452), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4468)
         );
  AND2_X1 U4026 ( .A1(n4278), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4285)
         );
  NAND2_X1 U4027 ( .A1(n6368), .A2(n4010), .ZN(n4738) );
  AND2_X1 U4028 ( .A1(n6868), .A2(n5904), .ZN(n5857) );
  INV_X1 U4029 ( .A(n5567), .ZN(n5120) );
  INV_X1 U4030 ( .A(n4915), .ZN(n5303) );
  OR2_X1 U4031 ( .A1(n5174), .A2(n3462), .ZN(n5502) );
  NAND2_X1 U4032 ( .A1(n5261), .A2(n4915), .ZN(n5830) );
  AND2_X1 U4033 ( .A1(n3463), .A2(n4963), .ZN(n5176) );
  OR2_X1 U4034 ( .A1(n4927), .A2(n7082), .ZN(n5119) );
  NAND2_X1 U4035 ( .A1(n7121), .A2(n6757), .ZN(n7122) );
  INV_X1 U4036 ( .A(n4743), .ZN(n4744) );
  NAND2_X1 U4037 ( .A1(n4742), .A2(n3478), .ZN(n4745) );
  AND2_X1 U4038 ( .A1(n6107), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7009) );
  AND2_X1 U4039 ( .A1(n6107), .A2(n5212), .ZN(n6974) );
  AND2_X1 U4040 ( .A1(n6107), .A2(n5228), .ZN(n7017) );
  INV_X1 U4041 ( .A(n6015), .ZN(n7235) );
  INV_X1 U4042 ( .A(n7125), .ZN(n7196) );
  AND2_X1 U4043 ( .A1(n4285), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4296)
         );
  INV_X1 U4044 ( .A(n4780), .ZN(n7121) );
  INV_X1 U4045 ( .A(n4925), .ZN(n5538) );
  NOR2_X1 U4046 ( .A1(n5536), .A2(n4915), .ZN(n5583) );
  NOR2_X1 U4047 ( .A1(n5397), .A2(n4915), .ZN(n5440) );
  AND2_X1 U4048 ( .A1(n5507), .A2(n4915), .ZN(n5567) );
  NOR2_X1 U4049 ( .A1(n5387), .A2(n5687), .ZN(n5302) );
  NOR2_X2 U4050 ( .A1(n5502), .A2(n4915), .ZN(n5833) );
  AND2_X1 U4051 ( .A1(n5176), .A2(n4915), .ZN(n7222) );
  AND2_X1 U4052 ( .A1(n5387), .A2(n5764), .ZN(n5306) );
  NOR2_X1 U4053 ( .A1(n6560), .A2(n5256), .ZN(n5581) );
  NOR2_X1 U4054 ( .A1(n6503), .A2(n5256), .ZN(n5710) );
  NOR2_X1 U4055 ( .A1(n5119), .A2(n6016), .ZN(n5776) );
  NAND2_X1 U4056 ( .A1(n7122), .A2(n7118), .ZN(n6769) );
  INV_X1 U4057 ( .A(n7016), .ZN(n7001) );
  NAND2_X1 U4058 ( .A1(n6015), .A2(n4872), .ZN(n5916) );
  INV_X1 U4059 ( .A(n6613), .ZN(n6633) );
  NAND2_X1 U4060 ( .A1(n4233), .A2(n4102), .ZN(n6878) );
  INV_X1 U4061 ( .A(n5776), .ZN(n5560) );
  AND2_X1 U4062 ( .A1(n4921), .A2(n4920), .ZN(n5384) );
  NAND2_X1 U4063 ( .A1(n4916), .A2(n4915), .ZN(n5594) );
  AOI22_X1 U4064 ( .A1(n5773), .A2(n5769), .B1(n5768), .B2(n5767), .ZN(n5835)
         );
  INV_X1 U4065 ( .A(n5799), .ZN(n5714) );
  INV_X1 U4066 ( .A(n5581), .ZN(n7227) );
  INV_X1 U4067 ( .A(n5700), .ZN(n5812) );
  AND2_X1 U4068 ( .A1(STATE_REG_1__SCAN_IN), .A2(n7105), .ZN(n7116) );
  OAI21_X1 U4069 ( .B1(n6160), .B2(n6156), .A(n4772), .ZN(U2830) );
  INV_X1 U4070 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4071 ( .A1(n3700), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3680), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4072 ( .A1(n3660), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4073 ( .A1(n4485), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4074 ( .A1(n3466), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4075 ( .A1(n3856), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3459), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4076 ( .A1(n3673), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4332), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3589) );
  AND2_X4 U4077 ( .A1(n4809), .A2(n5019), .ZN(n4674) );
  NAND2_X4 U4078 ( .A1(n3593), .A2(n3592), .ZN(n3820) );
  NAND2_X1 U4079 ( .A1(n3465), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3597) );
  NAND2_X1 U4080 ( .A1(n3856), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4081 ( .A1(n3693), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3595) );
  NAND2_X1 U4082 ( .A1(n4658), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4083 ( .A1(n3698), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3601) );
  NAND2_X1 U4084 ( .A1(n3466), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3600) );
  NAND2_X1 U4085 ( .A1(n3700), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3599) );
  NAND2_X1 U4086 ( .A1(n3680), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3598)
         );
  NAND2_X1 U4087 ( .A1(n3672), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U4088 ( .A1(n4674), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3604)
         );
  NAND2_X1 U4089 ( .A1(n3855), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3603)
         );
  NAND2_X1 U4090 ( .A1(n3459), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3602) );
  NAND2_X1 U4091 ( .A1(n3673), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3609)
         );
  NAND2_X1 U4092 ( .A1(n3660), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3608)
         );
  NAND2_X1 U4093 ( .A1(n4332), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U4094 ( .A1(n3681), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3606)
         );
  AND4_X1 U4095 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(n3610)
         );
  AND2_X2 U4096 ( .A1(n3820), .A2(n3614), .ZN(n3733) );
  NAND2_X1 U4097 ( .A1(n3660), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3618)
         );
  NAND2_X1 U4098 ( .A1(n3673), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3617)
         );
  NAND2_X1 U4099 ( .A1(n4332), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3616) );
  NAND2_X1 U4100 ( .A1(n3681), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3615)
         );
  NAND2_X1 U4101 ( .A1(n3698), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3622) );
  NAND2_X1 U4102 ( .A1(n3467), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3621) );
  NAND2_X1 U4103 ( .A1(n3700), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3620) );
  NAND2_X1 U4104 ( .A1(n3680), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3619)
         );
  NAND2_X1 U4105 ( .A1(n3672), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3626) );
  NAND2_X1 U4106 ( .A1(n3468), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3625)
         );
  NAND2_X1 U4107 ( .A1(n3855), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3624)
         );
  NAND2_X1 U4108 ( .A1(n3460), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3623) );
  NAND2_X1 U4109 ( .A1(n4485), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U4110 ( .A1(n3856), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4111 ( .A1(n3693), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3628) );
  NAND2_X1 U4112 ( .A1(n3456), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3627) );
  NAND2_X1 U4113 ( .A1(n3672), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4114 ( .A1(n4332), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4115 ( .A1(n3673), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3635)
         );
  NAND3_X1 U4116 ( .A1(n3637), .A2(n3636), .A3(n3635), .ZN(n3639) );
  NAND2_X1 U4117 ( .A1(n3464), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U4118 ( .A1(n3856), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3641) );
  NAND2_X1 U4119 ( .A1(n3681), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3640)
         );
  NAND2_X1 U4120 ( .A1(n3693), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3647) );
  NAND2_X1 U4121 ( .A1(n4658), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3646) );
  NAND2_X1 U4122 ( .A1(n3466), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4123 ( .A1(n3700), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3644) );
  NAND2_X1 U4124 ( .A1(n3855), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3651)
         );
  NAND2_X1 U4125 ( .A1(n3680), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3650)
         );
  NAND2_X1 U4126 ( .A1(n3459), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4127 ( .A1(n3856), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3693), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4128 ( .A1(n3467), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3680), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4129 ( .A1(n3672), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4130 ( .A1(n4485), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4131 ( .A1(n3698), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3458), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4132 ( .A1(n3855), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4332), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3661) );
  INV_X1 U4133 ( .A(n3820), .ZN(n3724) );
  NAND3_X1 U4134 ( .A1(n4091), .A2(n3720), .A3(n3724), .ZN(n4099) );
  NAND2_X1 U4135 ( .A1(n3754), .A2(n3736), .ZN(n3692) );
  AOI22_X1 U4136 ( .A1(n3467), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4137 ( .A1(n3693), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4138 ( .A1(n3465), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4139 ( .A1(n3700), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3680), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3668) );
  NAND4_X1 U4140 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3679)
         );
  AOI22_X1 U4141 ( .A1(n3672), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4142 ( .A1(n3855), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3676) );
  NAND4_X1 U4143 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3678)
         );
  AOI22_X1 U4144 ( .A1(n3467), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4145 ( .A1(n3700), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3680), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4146 ( .A1(n3457), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4147 ( .A1(n3672), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4148 ( .A1(n3856), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4149 ( .A1(n3465), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3693), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4150 ( .A1(n3660), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4332), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3686) );
  NAND2_X1 U4151 ( .A1(n3692), .A2(n3737), .ZN(n3732) );
  NAND2_X1 U4152 ( .A1(n4485), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3697) );
  NAND2_X1 U4153 ( .A1(n3856), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3696) );
  INV_X1 U4154 ( .A(n3693), .ZN(n3885) );
  NAND2_X1 U4155 ( .A1(n3693), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3695) );
  NAND2_X1 U4156 ( .A1(n3457), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3694) );
  NAND2_X1 U4157 ( .A1(n3698), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U4158 ( .A1(n3467), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4159 ( .A1(n3700), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3702) );
  NAND2_X1 U4160 ( .A1(n3680), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3701)
         );
  NAND2_X1 U4161 ( .A1(n3672), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3708) );
  NAND2_X1 U4162 ( .A1(n3459), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3707) );
  NAND2_X1 U4163 ( .A1(n3855), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3706)
         );
  NAND3_X1 U4164 ( .A1(n3708), .A2(n3707), .A3(n3706), .ZN(n3709) );
  NAND2_X1 U4165 ( .A1(n3673), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3713)
         );
  NAND2_X1 U4166 ( .A1(n3660), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3712)
         );
  NAND2_X1 U4167 ( .A1(n4332), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3711) );
  NAND2_X1 U4168 ( .A1(n3681), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3710)
         );
  NAND2_X1 U4169 ( .A1(n3732), .A2(n3511), .ZN(n3728) );
  NAND2_X1 U4170 ( .A1(n3724), .A2(n3718), .ZN(n3719) );
  OAI21_X1 U4171 ( .B1(n4755), .B2(n3747), .A(n3726), .ZN(n3739) );
  INV_X1 U4172 ( .A(n3739), .ZN(n3721) );
  NAND2_X1 U4173 ( .A1(n3721), .A2(n3748), .ZN(n4073) );
  INV_X1 U4174 ( .A(STATE_REG_1__SCAN_IN), .ZN(n3722) );
  XNOR2_X1 U4175 ( .A(n3722), .B(STATE_REG_2__SCAN_IN), .ZN(n7101) );
  INV_X1 U4176 ( .A(n7101), .ZN(n3723) );
  NAND2_X1 U4177 ( .A1(n3753), .A2(n3724), .ZN(n3725) );
  NAND2_X1 U4178 ( .A1(n3747), .A2(n4755), .ZN(n3740) );
  NAND2_X1 U4179 ( .A1(n3726), .A2(n3614), .ZN(n4071) );
  NAND2_X1 U4180 ( .A1(n3821), .A2(n4071), .ZN(n3727) );
  NAND2_X1 U4181 ( .A1(n3844), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3731) );
  NAND2_X1 U4182 ( .A1(n7077), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4089) );
  NAND2_X1 U4183 ( .A1(n7077), .A2(n7084), .ZN(n7075) );
  MUX2_X1 U4184 ( .A(n4089), .B(n4725), .S(n7043), .Z(n3729) );
  INV_X1 U4185 ( .A(n3729), .ZN(n3730) );
  NAND2_X1 U4186 ( .A1(n3731), .A2(n3730), .ZN(n3795) );
  NAND2_X1 U4187 ( .A1(n3733), .A2(n4098), .ZN(n3734) );
  NOR2_X1 U4188 ( .A1(n7075), .A2(n7096), .ZN(n3744) );
  OAI21_X1 U4189 ( .B1(n3736), .B2(n3830), .A(n3511), .ZN(n3738) );
  NAND2_X1 U4190 ( .A1(n3738), .A2(n3737), .ZN(n3743) );
  NAND2_X1 U4191 ( .A1(n3740), .A2(n3830), .ZN(n3741) );
  OAI21_X1 U4192 ( .B1(n3448), .B2(n3741), .A(n4098), .ZN(n3742) );
  AND2_X2 U4193 ( .A1(n3795), .A2(n3796), .ZN(n3840) );
  INV_X1 U4195 ( .A(n4071), .ZN(n3750) );
  INV_X1 U4196 ( .A(n4070), .ZN(n3752) );
  NAND2_X1 U4197 ( .A1(n3752), .A2(n4097), .ZN(n4773) );
  INV_X1 U4198 ( .A(n3753), .ZN(n3755) );
  NAND2_X1 U4199 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3756), .ZN(n3761) );
  INV_X1 U4200 ( .A(n4725), .ZN(n3758) );
  NAND2_X1 U4201 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3845) );
  OAI21_X1 U4202 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n3845), .ZN(n4960) );
  INV_X1 U4203 ( .A(n4089), .ZN(n3757) );
  OAI22_X1 U4204 ( .A1(n3758), .A2(n4960), .B1(n3757), .B2(n5534), .ZN(n3762)
         );
  INV_X1 U4205 ( .A(n3762), .ZN(n3759) );
  OAI211_X1 U4206 ( .C1(n3760), .C2(n3582), .A(n3761), .B(n3759), .ZN(n3838)
         );
  INV_X1 U4207 ( .A(n3761), .ZN(n3763) );
  XNOR2_X2 U4208 ( .A(n3840), .B(n3839), .ZN(n4811) );
  AOI22_X1 U4209 ( .A1(n4485), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4210 ( .A1(n3700), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4211 ( .A1(n3776), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4212 ( .A1(n3468), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4332), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4213 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3774)
         );
  AOI22_X1 U4214 ( .A1(n3798), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4215 ( .A1(n4696), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4216 ( .A1(n3673), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4217 ( .A1(n4697), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4218 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3773)
         );
  NAND2_X1 U4219 ( .A1(n4052), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3790) );
  OR2_X1 U4220 ( .A1(n3850), .A2(n3775), .ZN(n3789) );
  INV_X1 U4221 ( .A(n3849), .ZN(n3980) );
  AOI22_X1 U4222 ( .A1(n4697), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4223 ( .A1(n4485), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4224 ( .A1(n4696), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4225 ( .A1(n3468), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4226 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3786)
         );
  AOI22_X1 U4227 ( .A1(n3467), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4228 ( .A1(n3434), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4229 ( .A1(n4698), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4230 ( .A1(n3460), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4332), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4231 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3785)
         );
  INV_X1 U4232 ( .A(n3983), .ZN(n3787) );
  NAND2_X1 U4233 ( .A1(n3980), .A2(n3787), .ZN(n3788) );
  NAND2_X1 U4234 ( .A1(n3792), .A2(n3791), .ZN(n3794) );
  NAND2_X1 U4235 ( .A1(n3794), .A2(n3836), .ZN(n3815) );
  INV_X1 U4236 ( .A(n3796), .ZN(n3797) );
  AOI22_X1 U4237 ( .A1(n3798), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4238 ( .A1(n3434), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4239 ( .A1(n3673), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4240 ( .A1(n3776), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4332), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3799) );
  NAND4_X1 U4241 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3808)
         );
  AOI22_X1 U4242 ( .A1(n3465), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4243 ( .A1(n3467), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4244 ( .A1(n4697), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4245 ( .A1(n3469), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4246 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3807)
         );
  XNOR2_X1 U4247 ( .A(n3983), .B(n3865), .ZN(n3809) );
  NOR2_X1 U4248 ( .A1(n3809), .A2(n3849), .ZN(n3827) );
  INV_X1 U4249 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3812) );
  AOI21_X1 U4250 ( .B1(n3614), .B2(n3983), .A(n7096), .ZN(n3811) );
  NAND2_X1 U4251 ( .A1(n3445), .A2(n3865), .ZN(n3810) );
  OAI211_X1 U4252 ( .C1(n4044), .C2(n3812), .A(n3811), .B(n3810), .ZN(n3826)
         );
  AND2_X1 U4253 ( .A1(n3827), .A2(n3826), .ZN(n3813) );
  NAND2_X1 U4254 ( .A1(n3980), .A2(n3983), .ZN(n3814) );
  NAND2_X1 U4255 ( .A1(n3829), .A2(n3814), .ZN(n3816) );
  NAND2_X1 U4256 ( .A1(n3815), .A2(n3816), .ZN(n3819) );
  INV_X1 U4257 ( .A(n3815), .ZN(n3818) );
  INV_X1 U4258 ( .A(n3816), .ZN(n3817) );
  NAND2_X1 U4259 ( .A1(n3818), .A2(n3817), .ZN(n3837) );
  NAND2_X1 U4260 ( .A1(n3819), .A2(n3837), .ZN(n4914) );
  NAND2_X1 U4261 ( .A1(n4914), .A2(n3971), .ZN(n3825) );
  XNOR2_X1 U4262 ( .A(n3866), .B(n3865), .ZN(n3822) );
  INV_X1 U4263 ( .A(n3821), .ZN(n6773) );
  OAI211_X1 U4264 ( .C1(n3822), .C2(n6773), .A(n3748), .B(n3820), .ZN(n3823)
         );
  INV_X1 U4265 ( .A(n3823), .ZN(n3824) );
  NAND2_X1 U4266 ( .A1(n3825), .A2(n3824), .ZN(n3834) );
  OR2_X1 U4267 ( .A1(n3827), .A2(n3826), .ZN(n3828) );
  NAND2_X2 U4268 ( .A1(n3829), .A2(n3828), .ZN(n4915) );
  OR2_X1 U4269 ( .A1(n4915), .A2(n4221), .ZN(n3833) );
  NAND2_X1 U4270 ( .A1(n3445), .A2(n3830), .ZN(n3868) );
  OAI21_X1 U4271 ( .B1(n6773), .B2(n3865), .A(n3868), .ZN(n3831) );
  INV_X1 U4272 ( .A(n3831), .ZN(n3832) );
  NAND2_X1 U4273 ( .A1(n3833), .A2(n3832), .ZN(n6708) );
  NAND2_X1 U4274 ( .A1(n6708), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6707)
         );
  INV_X1 U4275 ( .A(n3839), .ZN(n3842) );
  INV_X1 U4276 ( .A(n3840), .ZN(n3841) );
  NAND2_X1 U4277 ( .A1(n3842), .A2(n3841), .ZN(n3843) );
  INV_X1 U4278 ( .A(n3845), .ZN(n7050) );
  NAND2_X1 U4279 ( .A1(n7050), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U4280 ( .A1(n3845), .A2(n7054), .ZN(n3846) );
  AND2_X1 U4281 ( .A1(n5277), .A2(n3846), .ZN(n4922) );
  AOI22_X1 U4282 ( .A1(n4725), .A2(n4922), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4089), .ZN(n3847) );
  AOI22_X1 U4283 ( .A1(n3465), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4284 ( .A1(n3457), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4285 ( .A1(n3700), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4286 ( .A1(n4698), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3851) );
  NAND4_X1 U4287 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3862)
         );
  AOI22_X1 U4288 ( .A1(n4697), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4289 ( .A1(n3467), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4290 ( .A1(n3798), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4291 ( .A1(n3447), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4292 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  AOI22_X1 U4293 ( .A1(n4063), .A2(n3867), .B1(INSTQUEUE_REG_0__2__SCAN_IN), 
        .B2(n4052), .ZN(n3863) );
  NAND2_X1 U4294 ( .A1(n4244), .A2(n3971), .ZN(n3871) );
  NAND2_X1 U4295 ( .A1(n3866), .A2(n3865), .ZN(n3899) );
  INV_X1 U4296 ( .A(n3867), .ZN(n3898) );
  XNOR2_X1 U4297 ( .A(n3899), .B(n3898), .ZN(n3869) );
  INV_X1 U4298 ( .A(n3868), .ZN(n4215) );
  AOI21_X1 U4299 ( .B1(n3869), .B2(n3821), .A(n4215), .ZN(n3870) );
  INV_X1 U4300 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3872) );
  NAND2_X1 U4301 ( .A1(n6720), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3873)
         );
  NAND2_X1 U4302 ( .A1(n3903), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5341)
         );
  INV_X1 U4303 ( .A(n3875), .ZN(n3877) );
  NAND2_X1 U4304 ( .A1(n3877), .A2(n3876), .ZN(n3905) );
  INV_X1 U4305 ( .A(n3878), .ZN(n3879) );
  NAND2_X1 U4306 ( .A1(n3844), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3884) );
  INV_X1 U4307 ( .A(n5277), .ZN(n3881) );
  NAND2_X1 U4308 ( .A1(n3881), .A2(n7060), .ZN(n5437) );
  NAND2_X1 U4309 ( .A1(n5277), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3882) );
  NAND2_X1 U4310 ( .A1(n5437), .A2(n3882), .ZN(n4977) );
  AOI22_X1 U4311 ( .A1(n4977), .A2(n4725), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4089), .ZN(n3883) );
  AOI22_X1 U4312 ( .A1(n3465), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3889) );
  INV_X2 U4313 ( .A(n3885), .ZN(n4696) );
  AOI22_X1 U4314 ( .A1(n4696), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4315 ( .A1(n3467), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4316 ( .A1(n3700), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3886) );
  NAND4_X1 U4317 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3895)
         );
  AOI22_X1 U4318 ( .A1(n4697), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4319 ( .A1(n3776), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4320 ( .A1(n4698), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4321 ( .A1(n3447), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4322 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3894)
         );
  AOI22_X1 U4323 ( .A1(n4063), .A2(n3919), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n4052), .ZN(n3896) );
  XNOR2_X2 U4324 ( .A(n3905), .B(n5042), .ZN(n4267) );
  NAND2_X1 U4325 ( .A1(n3899), .A2(n3898), .ZN(n3920) );
  INV_X1 U4326 ( .A(n3919), .ZN(n3900) );
  XNOR2_X1 U4327 ( .A(n3920), .B(n3900), .ZN(n3901) );
  AND2_X1 U4328 ( .A1(n3901), .A2(n3821), .ZN(n3902) );
  NAND2_X1 U4329 ( .A1(n5341), .A2(n5344), .ZN(n3904) );
  NAND2_X1 U4330 ( .A1(n3450), .A2(n5345), .ZN(n5342) );
  NAND2_X1 U4331 ( .A1(n3904), .A2(n5342), .ZN(n5136) );
  INV_X1 U4332 ( .A(n3905), .ZN(n3906) );
  NAND2_X1 U4333 ( .A1(n3906), .A2(n5042), .ZN(n3925) );
  AOI22_X1 U4334 ( .A1(n3465), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4335 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3456), .B1(n4696), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4336 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3467), .B1(n3434), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4337 ( .A1(n3458), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3907) );
  NAND4_X1 U4338 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3916)
         );
  AOI22_X1 U4339 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4697), .B1(n3468), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4340 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3776), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4341 ( .A1(n4698), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4342 ( .A1(n3447), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3911) );
  NAND4_X1 U4343 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3915)
         );
  NAND2_X1 U4344 ( .A1(n4063), .A2(n3942), .ZN(n3918) );
  NAND2_X1 U4345 ( .A1(n4052), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3917) );
  NAND2_X1 U4346 ( .A1(n3918), .A2(n3917), .ZN(n3926) );
  NAND2_X1 U4347 ( .A1(n4277), .A2(n3971), .ZN(n3923) );
  NAND2_X1 U4348 ( .A1(n3920), .A2(n3919), .ZN(n3944) );
  XNOR2_X1 U4349 ( .A(n3944), .B(n3942), .ZN(n3921) );
  NAND2_X1 U4350 ( .A1(n3921), .A2(n3821), .ZN(n3922) );
  INV_X1 U4351 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4118) );
  OAI22_X2 U4352 ( .A1(n5136), .A2(n5137), .B1(n3455), .B2(n4118), .ZN(n5466)
         );
  INV_X1 U4353 ( .A(n3925), .ZN(n3927) );
  AOI22_X1 U4354 ( .A1(n4696), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4355 ( .A1(n4698), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4356 ( .A1(n3467), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4357 ( .A1(n3776), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4358 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3937)
         );
  AOI22_X1 U4359 ( .A1(n3434), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4360 ( .A1(n4485), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4361 ( .A1(n4697), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4362 ( .A1(n3660), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4363 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3936)
         );
  AOI22_X1 U4364 ( .A1(n4063), .A2(n3945), .B1(INSTQUEUE_REG_0__5__SCAN_IN), 
        .B2(n4052), .ZN(n3939) );
  NAND2_X1 U4365 ( .A1(n3940), .A2(n3939), .ZN(n3941) );
  NAND2_X1 U4366 ( .A1(n3962), .A2(n3941), .ZN(n4283) );
  INV_X1 U4367 ( .A(n3942), .ZN(n3943) );
  NOR2_X1 U4368 ( .A1(n3944), .A2(n3943), .ZN(n3946) );
  NAND2_X1 U4369 ( .A1(n3946), .A2(n3945), .ZN(n3974) );
  OAI211_X1 U4370 ( .C1(n3946), .C2(n3945), .A(n3974), .B(n3821), .ZN(n3947)
         );
  INV_X1 U4371 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5610) );
  XNOR2_X1 U4372 ( .A(n3948), .B(n5610), .ZN(n5465) );
  NAND2_X1 U4373 ( .A1(n3948), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3949)
         );
  AOI22_X1 U4374 ( .A1(n3465), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4375 ( .A1(n4696), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4376 ( .A1(n3467), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4377 ( .A1(n3700), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3950) );
  NAND4_X1 U4378 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3959)
         );
  AOI22_X1 U4379 ( .A1(n4697), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4380 ( .A1(n3776), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4381 ( .A1(n4698), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4382 ( .A1(n3447), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4383 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3958)
         );
  AOI22_X1 U4384 ( .A1(n4063), .A2(n3972), .B1(n4052), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3963) );
  INV_X1 U4385 ( .A(n3963), .ZN(n3960) );
  NAND2_X1 U4386 ( .A1(n3962), .A2(n3963), .ZN(n4293) );
  NAND3_X1 U4387 ( .A1(n3982), .A2(n3971), .A3(n4293), .ZN(n3966) );
  XNOR2_X1 U4388 ( .A(n3974), .B(n3972), .ZN(n3964) );
  NAND2_X1 U4389 ( .A1(n3964), .A2(n3821), .ZN(n3965) );
  NAND2_X1 U4390 ( .A1(n3966), .A2(n3965), .ZN(n3967) );
  NAND2_X1 U4391 ( .A1(n3967), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5605)
         );
  INV_X1 U4392 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3969) );
  NAND2_X1 U4393 ( .A1(n4063), .A2(n3983), .ZN(n3968) );
  OAI21_X1 U4394 ( .B1(n3969), .B2(n4044), .A(n3968), .ZN(n3970) );
  NAND2_X1 U4395 ( .A1(n4300), .A2(n3971), .ZN(n3977) );
  INV_X1 U4396 ( .A(n3972), .ZN(n3973) );
  OR2_X1 U4397 ( .A1(n3974), .A2(n3973), .ZN(n3985) );
  XNOR2_X1 U4398 ( .A(n3985), .B(n3983), .ZN(n3975) );
  NAND2_X1 U4399 ( .A1(n3975), .A2(n3821), .ZN(n3976) );
  INV_X1 U4400 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6807) );
  XNOR2_X1 U4401 ( .A(n3978), .B(n6807), .ZN(n6732) );
  NAND2_X1 U4402 ( .A1(n6733), .A2(n6732), .ZN(n6731) );
  NAND2_X1 U4403 ( .A1(n3978), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3979)
         );
  NAND2_X1 U4404 ( .A1(n6731), .A2(n3979), .ZN(n5485) );
  AND2_X4 U4405 ( .A1(n3982), .A2(n3981), .ZN(n6368) );
  NAND2_X1 U4406 ( .A1(n3821), .A2(n3983), .ZN(n3984) );
  OR2_X1 U4407 ( .A1(n3985), .A2(n3984), .ZN(n3986) );
  INV_X1 U4408 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6801) );
  XNOR2_X1 U4409 ( .A(n3987), .B(n6801), .ZN(n5484) );
  NAND2_X1 U4410 ( .A1(n5485), .A2(n5484), .ZN(n5483) );
  NAND2_X1 U4411 ( .A1(n3987), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3988)
         );
  XNOR2_X1 U4412 ( .A(n6369), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5743)
         );
  INV_X1 U4413 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3989) );
  OR2_X1 U4414 ( .A1(n3461), .A2(n3989), .ZN(n3990) );
  INV_X1 U4415 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4140) );
  NAND2_X1 U4416 ( .A1(n3461), .A2(n4140), .ZN(n5733) );
  OR2_X1 U4417 ( .A1(n6369), .A2(n4140), .ZN(n5734) );
  INV_X1 U4418 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6834) );
  NOR2_X1 U4419 ( .A1(n6369), .A2(n6834), .ZN(n6740) );
  NAND2_X1 U4420 ( .A1(n6369), .A2(n6834), .ZN(n6738) );
  INV_X1 U4421 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3991) );
  OR2_X1 U4422 ( .A1(n3461), .A2(n3991), .ZN(n5845) );
  NAND2_X1 U4423 ( .A1(n5847), .A2(n5845), .ZN(n3992) );
  NAND2_X1 U4424 ( .A1(n6369), .A2(n3991), .ZN(n5844) );
  XNOR2_X1 U4425 ( .A(n3461), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5877)
         );
  INV_X1 U4426 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4220) );
  NAND2_X1 U4427 ( .A1(n3461), .A2(n4220), .ZN(n3993) );
  INV_X1 U4428 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5899) );
  INV_X1 U4429 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6845) );
  AND2_X1 U4430 ( .A1(n3461), .A2(n6845), .ZN(n3996) );
  INV_X1 U4431 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4157) );
  NAND2_X1 U4432 ( .A1(n3461), .A2(n4157), .ZN(n3997) );
  INV_X1 U4433 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6377) );
  INV_X1 U4434 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6379) );
  AND3_X1 U4435 ( .A1(n4157), .A2(n6377), .A3(n6379), .ZN(n3998) );
  NAND2_X1 U4436 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U4437 ( .A1(n6369), .A2(n6351), .ZN(n4000) );
  NAND2_X1 U4438 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U4439 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6352) );
  NOR2_X1 U4440 ( .A1(n6323), .A2(n6352), .ZN(n4002) );
  NAND2_X1 U4441 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4240) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6332) );
  INV_X1 U4443 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4186) );
  INV_X1 U4444 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6233) );
  INV_X1 U4445 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6863) );
  NAND4_X1 U4446 ( .A1(n6332), .A2(n4186), .A3(n6233), .A4(n6863), .ZN(n4003)
         );
  INV_X1 U4447 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6346) );
  INV_X1 U4448 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U4449 ( .A1(n6346), .A2(n6364), .ZN(n6353) );
  XNOR2_X1 U4450 ( .A(n3461), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6206)
         );
  INV_X1 U4451 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6300) );
  INV_X1 U4452 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U4453 ( .A1(n3461), .A2(n6299), .ZN(n4005) );
  INV_X1 U4454 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4006) );
  NAND2_X1 U4455 ( .A1(n6182), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4014) );
  AND2_X1 U4456 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U4457 ( .A1(n6272), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4747) );
  AND2_X1 U4458 ( .A1(n6369), .A2(n4747), .ZN(n4009) );
  NOR2_X1 U4459 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4007) );
  OR2_X1 U4460 ( .A1(n6369), .A2(n4007), .ZN(n6181) );
  INV_X1 U4461 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6280) );
  OR2_X1 U4462 ( .A1(n3461), .A2(n6280), .ZN(n4008) );
  NAND2_X1 U4463 ( .A1(n3452), .A2(n4010), .ZN(n4013) );
  XNOR2_X1 U4464 ( .A(n6369), .B(n4010), .ZN(n6175) );
  NAND2_X1 U4465 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4011) );
  AND2_X1 U4466 ( .A1(n4011), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4012)
         );
  NAND3_X1 U4467 ( .A1(n4014), .A2(n4013), .A3(n3486), .ZN(n4016) );
  XNOR2_X1 U4468 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U4469 ( .A1(n4024), .A2(n4023), .ZN(n4018) );
  NAND2_X1 U4470 ( .A1(n5534), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4017) );
  NAND2_X1 U4471 ( .A1(n4018), .A2(n4017), .ZN(n4032) );
  MUX2_X1 U4472 ( .A(n7054), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4033) );
  NAND2_X1 U4473 ( .A1(n4032), .A2(n4033), .ZN(n4020) );
  NAND2_X1 U4474 ( .A1(n7054), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4019) );
  NAND2_X1 U4475 ( .A1(n4020), .A2(n4019), .ZN(n4051) );
  MUX2_X1 U4476 ( .A(n7060), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n4050) );
  INV_X1 U4477 ( .A(n4050), .ZN(n4021) );
  XNOR2_X1 U4478 ( .A(n4051), .B(n4021), .ZN(n4080) );
  INV_X1 U4479 ( .A(n4080), .ZN(n4048) );
  INV_X1 U4480 ( .A(n4024), .ZN(n4022) );
  OAI21_X1 U4481 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7043), .A(n4022), 
        .ZN(n4027) );
  INV_X1 U4482 ( .A(n4027), .ZN(n4031) );
  INV_X1 U4483 ( .A(n4023), .ZN(n4025) );
  XNOR2_X1 U4484 ( .A(n4025), .B(n4024), .ZN(n4079) );
  OAI21_X1 U4485 ( .B1(n4044), .B2(n4079), .A(n3820), .ZN(n4026) );
  AOI21_X1 U4486 ( .B1(n4063), .B2(n4098), .A(n4026), .ZN(n4037) );
  NAND2_X1 U4487 ( .A1(n4079), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4038) );
  INV_X1 U4488 ( .A(n4063), .ZN(n4028) );
  AOI211_X1 U4489 ( .C1(n4037), .C2(n4038), .A(n4028), .B(n4027), .ZN(n4029)
         );
  NOR2_X1 U4490 ( .A1(n4029), .A2(n4066), .ZN(n4036) );
  AOI211_X1 U4491 ( .C1(n4031), .C2(n4030), .A(n3445), .B(n4036), .ZN(n4041)
         );
  XOR2_X1 U4492 ( .A(n4033), .B(n4032), .Z(n4078) );
  NAND2_X1 U4493 ( .A1(n4063), .A2(n4078), .ZN(n4042) );
  AOI21_X1 U4494 ( .B1(n4034), .B2(n3820), .A(n4035), .ZN(n4043) );
  AOI21_X1 U4495 ( .B1(n4036), .B2(n4042), .A(n4043), .ZN(n4040) );
  AOI21_X1 U4496 ( .B1(n4053), .B2(n4038), .A(n4037), .ZN(n4039) );
  AND2_X1 U4497 ( .A1(n4043), .A2(n4042), .ZN(n4045) );
  OAI22_X1 U4498 ( .A1(n4045), .A2(n4048), .B1(n4078), .B2(n4044), .ZN(n4046)
         );
  AOI22_X1 U4499 ( .A1(n4066), .A2(n4048), .B1(n4047), .B2(n4046), .ZN(n4055)
         );
  NOR2_X1 U4500 ( .A1(n3581), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4049)
         );
  AOI21_X1 U4501 ( .B1(n4051), .B2(n4050), .A(n4049), .ZN(n4058) );
  NAND2_X1 U4502 ( .A1(n4058), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4057) );
  NOR2_X1 U4503 ( .A1(n4052), .A2(n4083), .ZN(n4054) );
  OAI22_X1 U4504 ( .A1(n4055), .A2(n4054), .B1(n4053), .B2(n4083), .ZN(n4056)
         );
  AOI21_X1 U4505 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7096), .A(n4056), 
        .ZN(n4065) );
  NAND2_X1 U4506 ( .A1(n4057), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4062) );
  INV_X1 U4507 ( .A(n4058), .ZN(n4060) );
  INV_X1 U4508 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4059) );
  NAND2_X1 U4509 ( .A1(n4060), .A2(n4059), .ZN(n4061) );
  NAND2_X1 U4510 ( .A1(n4062), .A2(n4061), .ZN(n4082) );
  NAND2_X1 U4511 ( .A1(n4063), .A2(n4082), .ZN(n4064) );
  NAND2_X1 U4512 ( .A1(n4065), .A2(n4064), .ZN(n4068) );
  NAND2_X1 U4513 ( .A1(n4066), .A2(n4082), .ZN(n4067) );
  INV_X1 U4514 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7105) );
  NAND2_X1 U4515 ( .A1(n7101), .A2(n7105), .ZN(n6771) );
  NAND2_X1 U4516 ( .A1(n4034), .A2(n6771), .ZN(n5210) );
  INV_X1 U4517 ( .A(READY_N), .ZN(n7124) );
  NAND2_X1 U4518 ( .A1(n5210), .A2(n7124), .ZN(n4069) );
  OR2_X1 U4519 ( .A1(n7026), .A2(n4069), .ZN(n4793) );
  MUX2_X1 U4520 ( .A(n4034), .B(n4071), .S(n3747), .Z(n4072) );
  NAND2_X1 U4521 ( .A1(n4072), .A2(n4097), .ZN(n4212) );
  AND2_X1 U4522 ( .A1(n3747), .A2(n3445), .ZN(n4074) );
  NOR2_X1 U4523 ( .A1(n4073), .A2(n4074), .ZN(n4095) );
  NAND2_X1 U4524 ( .A1(n4212), .A2(n4095), .ZN(n4077) );
  NAND2_X1 U4525 ( .A1(n4944), .A2(n3445), .ZN(n4076) );
  OR2_X1 U4526 ( .A1(n4075), .A2(n4076), .ZN(n7029) );
  NAND2_X1 U4527 ( .A1(n4077), .A2(n7029), .ZN(n4803) );
  NAND2_X1 U4528 ( .A1(n4098), .A2(n6771), .ZN(n4085) );
  AND3_X1 U4529 ( .A1(n4080), .A2(n4079), .A3(n4078), .ZN(n4081) );
  OR2_X1 U4530 ( .A1(n4082), .A2(n4081), .ZN(n4084) );
  NAND2_X1 U4531 ( .A1(n4084), .A2(n4083), .ZN(n7030) );
  AND2_X1 U4532 ( .A1(n7124), .A2(n7030), .ZN(n4798) );
  NAND3_X1 U4533 ( .A1(n4085), .A2(n3666), .A3(n4798), .ZN(n4086) );
  AND2_X1 U4534 ( .A1(n4803), .A2(n4086), .ZN(n4088) );
  NAND3_X1 U4535 ( .A1(n7026), .A2(n5969), .A3(n3971), .ZN(n4087) );
  OAI211_X1 U4536 ( .C1(n4793), .C2(n4070), .A(n4088), .B(n4087), .ZN(n4090)
         );
  OR2_X1 U4537 ( .A1(n4089), .A2(n7096), .ZN(n7073) );
  INV_X1 U4538 ( .A(n7073), .ZN(n7092) );
  NAND2_X1 U4539 ( .A1(n4090), .A2(n7092), .ZN(n4094) );
  INV_X1 U4540 ( .A(n4091), .ZN(n5933) );
  AOI21_X1 U4541 ( .B1(n5933), .B2(n4097), .A(n3666), .ZN(n4092) );
  NAND2_X1 U4542 ( .A1(n7121), .A2(n4092), .ZN(n4093) );
  AND2_X1 U4543 ( .A1(n4095), .A2(n3733), .ZN(n7062) );
  INV_X1 U4544 ( .A(n7062), .ZN(n4096) );
  NAND2_X1 U4545 ( .A1(n4095), .A2(n4035), .ZN(n4823) );
  AND2_X1 U4546 ( .A1(n4096), .A2(n4823), .ZN(n7024) );
  NOR2_X1 U4547 ( .A1(n4075), .A2(n4862), .ZN(n5024) );
  INV_X1 U4548 ( .A(n5024), .ZN(n4101) );
  OR2_X1 U4549 ( .A1(n4070), .A2(n5221), .ZN(n4865) );
  OR3_X1 U4550 ( .A1(n4099), .A2(n4862), .A3(n3614), .ZN(n4100) );
  NAND4_X1 U4551 ( .A1(n7024), .A2(n4101), .A3(n4865), .A4(n4100), .ZN(n4102)
         );
  NAND2_X1 U4552 ( .A1(n4944), .A2(n4097), .ZN(n4125) );
  BUF_X2 U4553 ( .A(n4103), .Z(n4202) );
  OAI22_X1 U4554 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5221), .ZN(n4205) );
  OR2_X2 U4555 ( .A1(n5221), .A2(n4202), .ZN(n4203) );
  NAND2_X1 U4556 ( .A1(n4125), .A2(n3835), .ZN(n4106) );
  INV_X1 U4557 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4104) );
  NAND2_X1 U4558 ( .A1(n4791), .A2(n4104), .ZN(n4105) );
  NAND3_X1 U4559 ( .A1(n4106), .A2(n4105), .A3(n4202), .ZN(n4107) );
  NAND2_X1 U4560 ( .A1(n4108), .A2(n4107), .ZN(n4111) );
  NAND2_X1 U4561 ( .A1(n4125), .A2(EBX_REG_0__SCAN_IN), .ZN(n4110) );
  INV_X1 U4562 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U4563 ( .A1(n4202), .A2(n5458), .ZN(n4109) );
  NAND2_X1 U4564 ( .A1(n4110), .A2(n4109), .ZN(n4899) );
  INV_X1 U4565 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U4566 ( .A1(n4191), .A2(n5994), .ZN(n4115) );
  NAND2_X1 U4567 ( .A1(n4125), .A2(n3872), .ZN(n4113) );
  NAND2_X1 U4568 ( .A1(n4791), .A2(n5994), .ZN(n4112) );
  NAND3_X1 U4569 ( .A1(n4113), .A2(n4112), .A3(n4202), .ZN(n4114) );
  NAND2_X1 U4570 ( .A1(n4115), .A2(n4114), .ZN(n5985) );
  MUX2_X1 U4571 ( .A(n4195), .B(n4202), .S(EBX_REG_3__SCAN_IN), .Z(n4117) );
  OR2_X1 U4572 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4116)
         );
  INV_X1 U4573 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U4574 ( .A1(n4191), .A2(n5224), .ZN(n4121) );
  NAND2_X1 U4575 ( .A1(n4125), .A2(n4118), .ZN(n4119) );
  OAI211_X1 U4576 ( .C1(n5221), .C2(EBX_REG_4__SCAN_IN), .A(n4119), .B(n4202), 
        .ZN(n4120) );
  MUX2_X1 U4577 ( .A(n4195), .B(n4202), .S(EBX_REG_5__SCAN_IN), .Z(n4124) );
  OAI21_X1 U4578 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4898), .A(n4124), 
        .ZN(n4849) );
  INV_X1 U4579 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U4580 ( .A1(n4191), .A2(n6880), .ZN(n4130) );
  INV_X1 U4581 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4126) );
  NAND2_X1 U4582 ( .A1(n4125), .A2(n4126), .ZN(n4128) );
  NAND2_X1 U4583 ( .A1(n4791), .A2(n6880), .ZN(n4127) );
  NAND3_X1 U4584 ( .A1(n4128), .A2(n4127), .A3(n4202), .ZN(n4129) );
  NAND2_X1 U4585 ( .A1(n4130), .A2(n4129), .ZN(n4906) );
  OR2_X1 U4586 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4132)
         );
  MUX2_X1 U4587 ( .A(n4195), .B(n4202), .S(EBX_REG_7__SCAN_IN), .Z(n4131) );
  AND2_X1 U4588 ( .A1(n4132), .A2(n4131), .ZN(n5099) );
  INV_X1 U4589 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U4590 ( .A1(n4191), .A2(n5241), .ZN(n4135) );
  NAND2_X1 U4591 ( .A1(n4125), .A2(n6801), .ZN(n4133) );
  OAI211_X1 U4592 ( .C1(n5221), .C2(EBX_REG_8__SCAN_IN), .A(n4133), .B(n4202), 
        .ZN(n4134) );
  MUX2_X1 U4593 ( .A(n4195), .B(n4202), .S(EBX_REG_9__SCAN_IN), .Z(n4137) );
  OR2_X1 U4594 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4136)
         );
  NAND2_X1 U4595 ( .A1(n4137), .A2(n4136), .ZN(n5448) );
  OR2_X1 U4596 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4139)
         );
  MUX2_X1 U4597 ( .A(n4195), .B(n4202), .S(EBX_REG_11__SCAN_IN), .Z(n4138) );
  AND2_X1 U4598 ( .A1(n4139), .A2(n4138), .ZN(n5677) );
  INV_X1 U4599 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U4600 ( .A1(n4191), .A2(n5595), .ZN(n4144) );
  NAND2_X1 U4601 ( .A1(n4125), .A2(n4140), .ZN(n4142) );
  NAND2_X1 U4602 ( .A1(n4791), .A2(n5595), .ZN(n4141) );
  NAND3_X1 U4603 ( .A1(n4142), .A2(n4141), .A3(n4202), .ZN(n4143) );
  NAND2_X1 U4604 ( .A1(n4144), .A2(n4143), .ZN(n5678) );
  NAND2_X1 U4605 ( .A1(n5677), .A2(n5678), .ZN(n4145) );
  NAND2_X1 U4606 ( .A1(n4103), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4146) );
  NAND2_X1 U4607 ( .A1(n4125), .A2(n4146), .ZN(n4149) );
  INV_X1 U4608 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4147) );
  NAND2_X1 U4609 ( .A1(n4791), .A2(n4147), .ZN(n4148) );
  NAND2_X1 U4610 ( .A1(n4149), .A2(n4148), .ZN(n4150) );
  OAI21_X1 U4611 ( .B1(EBX_REG_12__SCAN_IN), .B2(n4203), .A(n4150), .ZN(n5757)
         );
  NAND2_X1 U4612 ( .A1(n3475), .A2(n5757), .ZN(n5841) );
  MUX2_X1 U4613 ( .A(n4195), .B(n4202), .S(EBX_REG_13__SCAN_IN), .Z(n4151) );
  OAI21_X1 U4614 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n4898), .A(n4151), 
        .ZN(n5842) );
  OR2_X2 U4615 ( .A1(n5841), .A2(n5842), .ZN(n5872) );
  INV_X1 U4616 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U4617 ( .A1(n4191), .A2(n6931), .ZN(n4154) );
  NAND2_X1 U4618 ( .A1(n4125), .A2(n5899), .ZN(n4152) );
  OAI211_X1 U4619 ( .C1(n5221), .C2(EBX_REG_14__SCAN_IN), .A(n4152), .B(n4202), 
        .ZN(n4153) );
  MUX2_X1 U4620 ( .A(n4195), .B(n4202), .S(EBX_REG_15__SCAN_IN), .Z(n4156) );
  OR2_X1 U4621 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4155)
         );
  INV_X1 U4622 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6953) );
  NAND2_X1 U4623 ( .A1(n4191), .A2(n6953), .ZN(n4161) );
  NAND2_X1 U4624 ( .A1(n4125), .A2(n4157), .ZN(n4159) );
  NAND2_X1 U4625 ( .A1(n4791), .A2(n6953), .ZN(n4158) );
  NAND3_X1 U4626 ( .A1(n4159), .A2(n4158), .A3(n4103), .ZN(n4160) );
  NAND2_X1 U4627 ( .A1(n4161), .A2(n4160), .ZN(n5927) );
  OR2_X1 U4628 ( .A1(n4195), .A2(EBX_REG_17__SCAN_IN), .ZN(n4164) );
  NAND2_X1 U4629 ( .A1(n4103), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4162) );
  OAI211_X1 U4630 ( .C1(n5221), .C2(EBX_REG_17__SCAN_IN), .A(n4125), .B(n4162), 
        .ZN(n4163) );
  NAND2_X1 U4631 ( .A1(n4164), .A2(n4163), .ZN(n5921) );
  INV_X1 U4632 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U4633 ( .A1(n4191), .A2(n6155), .ZN(n4168) );
  NAND2_X1 U4634 ( .A1(n4202), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U4635 ( .A1(n4125), .A2(n4165), .ZN(n4166) );
  OAI21_X1 U4636 ( .B1(EBX_REG_18__SCAN_IN), .B2(n5221), .A(n4166), .ZN(n4167)
         );
  AND2_X1 U4637 ( .A1(n4168), .A2(n4167), .ZN(n6151) );
  OR2_X1 U4638 ( .A1(n4195), .A2(EBX_REG_19__SCAN_IN), .ZN(n4171) );
  NAND2_X1 U4639 ( .A1(n4103), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4169) );
  OAI211_X1 U4640 ( .C1(n5221), .C2(EBX_REG_19__SCAN_IN), .A(n4125), .B(n4169), 
        .ZN(n4170) );
  NAND2_X1 U4641 ( .A1(n4171), .A2(n4170), .ZN(n6359) );
  NAND2_X1 U4642 ( .A1(n4202), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4172) );
  NAND2_X1 U4643 ( .A1(n4125), .A2(n4172), .ZN(n4174) );
  INV_X1 U4644 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U4645 ( .A1(n4791), .A2(n6147), .ZN(n4173) );
  NAND2_X1 U4646 ( .A1(n4174), .A2(n4173), .ZN(n4175) );
  OAI21_X1 U4647 ( .B1(EBX_REG_20__SCAN_IN), .B2(n4203), .A(n4175), .ZN(n6146)
         );
  OR2_X1 U4648 ( .A1(n4195), .A2(EBX_REG_21__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U4649 ( .A1(n4202), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4176) );
  OAI211_X1 U4650 ( .C1(n5221), .C2(EBX_REG_21__SCAN_IN), .A(n4125), .B(n4176), 
        .ZN(n4177) );
  NAND2_X1 U4651 ( .A1(n4178), .A2(n4177), .ZN(n6105) );
  INV_X1 U4652 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6997) );
  NAND2_X1 U4653 ( .A1(n4191), .A2(n6997), .ZN(n4181) );
  NAND2_X1 U4654 ( .A1(n4125), .A2(n6233), .ZN(n4179) );
  OAI211_X1 U4655 ( .C1(n5221), .C2(EBX_REG_22__SCAN_IN), .A(n4179), .B(n4103), 
        .ZN(n4180) );
  AND2_X1 U4656 ( .A1(n4181), .A2(n4180), .ZN(n6135) );
  MUX2_X1 U4657 ( .A(n4195), .B(n4103), .S(EBX_REG_23__SCAN_IN), .Z(n4183) );
  OR2_X1 U4658 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4182)
         );
  AND2_X1 U4659 ( .A1(n4183), .A2(n4182), .ZN(n6090) );
  MUX2_X1 U4660 ( .A(n4195), .B(n4103), .S(EBX_REG_25__SCAN_IN), .Z(n4185) );
  OR2_X1 U4661 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4184)
         );
  NAND2_X1 U4662 ( .A1(n4185), .A2(n4184), .ZN(n6070) );
  INV_X1 U4663 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U4664 ( .A1(n4191), .A2(n6705), .ZN(n4189) );
  NAND2_X1 U4665 ( .A1(n4125), .A2(n4186), .ZN(n4187) );
  OAI211_X1 U4666 ( .C1(n5221), .C2(EBX_REG_24__SCAN_IN), .A(n4187), .B(n4202), 
        .ZN(n4188) );
  AND2_X1 U4667 ( .A1(n4189), .A2(n4188), .ZN(n6315) );
  NOR2_X1 U4668 ( .A1(n6070), .A2(n6315), .ZN(n4190) );
  INV_X1 U4669 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U4670 ( .A1(n4191), .A2(n6131), .ZN(n4194) );
  NAND2_X1 U4671 ( .A1(n4125), .A2(n6299), .ZN(n4192) );
  OAI211_X1 U4672 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5221), .A(n4192), .B(n4202), 
        .ZN(n4193) );
  AND2_X1 U4673 ( .A1(n4194), .A2(n4193), .ZN(n6054) );
  OR2_X2 U4674 ( .A1(n6072), .A2(n6054), .ZN(n6056) );
  MUX2_X1 U4675 ( .A(n4195), .B(n4103), .S(EBX_REG_27__SCAN_IN), .Z(n4197) );
  OR2_X1 U4676 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4196)
         );
  NAND2_X1 U4677 ( .A1(n4197), .A2(n4196), .ZN(n6045) );
  NAND2_X1 U4678 ( .A1(n4202), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4198) );
  NAND2_X1 U4679 ( .A1(n4125), .A2(n4198), .ZN(n4200) );
  INV_X1 U4680 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U4681 ( .A1(n4791), .A2(n6129), .ZN(n4199) );
  NAND2_X1 U4682 ( .A1(n4200), .A2(n4199), .ZN(n4201) );
  OAI21_X1 U4683 ( .B1(EBX_REG_28__SCAN_IN), .B2(n4203), .A(n4201), .ZN(n6030)
         );
  OAI22_X1 U4684 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n5221), .ZN(n4741) );
  INV_X1 U4685 ( .A(n4202), .ZN(n4208) );
  OAI22_X1 U4686 ( .A1(n4741), .A2(n4208), .B1(EBX_REG_29__SCAN_IN), .B2(n4203), .ZN(n4767) );
  OAI22_X1 U4687 ( .A1(n4898), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n5221), .ZN(n4743) );
  OR2_X1 U4688 ( .A1(n4070), .A2(n6773), .ZN(n7069) );
  OR3_X1 U4689 ( .A1(n4099), .A2(n4755), .A3(n4862), .ZN(n4206) );
  NAND2_X1 U4690 ( .A1(n7069), .A2(n4206), .ZN(n4207) );
  NOR2_X1 U4691 ( .A1(n7029), .A2(n4034), .ZN(n5010) );
  NAND2_X1 U4692 ( .A1(n4233), .A2(n5010), .ZN(n6868) );
  AOI22_X1 U4693 ( .A1(n3448), .A2(n4208), .B1(n3666), .B2(n5933), .ZN(n4211)
         );
  NAND2_X1 U4694 ( .A1(n3445), .A2(n4098), .ZN(n5213) );
  NOR2_X1 U4695 ( .A1(n5213), .A2(n3666), .ZN(n4801) );
  INV_X1 U4696 ( .A(n3748), .ZN(n4209) );
  OAI21_X1 U4697 ( .B1(n4801), .B2(n4898), .A(n4209), .ZN(n4210) );
  AND3_X1 U4698 ( .A1(n4212), .A2(n4211), .A3(n4210), .ZN(n4213) );
  AND2_X1 U4699 ( .A1(n4214), .A2(n4213), .ZN(n4814) );
  INV_X1 U4700 ( .A(n4862), .ZN(n4216) );
  AOI22_X1 U4701 ( .A1(n4216), .A2(n3746), .B1(n3733), .B2(n4215), .ZN(n4217)
         );
  NAND2_X1 U4702 ( .A1(n4814), .A2(n4217), .ZN(n4218) );
  NAND2_X1 U4703 ( .A1(n4233), .A2(n4218), .ZN(n5904) );
  INV_X1 U4704 ( .A(n6868), .ZN(n4219) );
  NOR2_X1 U4705 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4219), .ZN(n4884)
         );
  NAND2_X1 U4706 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U4707 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5880) );
  NOR2_X1 U4708 ( .A1(n4220), .A2(n5880), .ZN(n5900) );
  NAND2_X1 U4709 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5900), .ZN(n6386) );
  NOR2_X1 U4710 ( .A1(n6349), .A2(n6386), .ZN(n4223) );
  NAND2_X1 U4711 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6810) );
  NAND4_X1 U4712 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(INSTADDRPOINTER_REG_4__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6797) );
  NOR3_X1 U4713 ( .A1(n6801), .A2(n6807), .A3(n6797), .ZN(n6809) );
  NAND3_X1 U4714 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6809), .ZN(n6813) );
  NOR2_X1 U4715 ( .A1(n6810), .A2(n6813), .ZN(n5856) );
  NAND2_X1 U4716 ( .A1(n4223), .A2(n5856), .ZN(n6374) );
  NOR2_X1 U4717 ( .A1(n6374), .A2(n6351), .ZN(n4232) );
  NAND2_X1 U4718 ( .A1(n6378), .A2(n4232), .ZN(n4226) );
  NOR2_X1 U4719 ( .A1(n4221), .A2(n3445), .ZN(n4222) );
  AND3_X1 U4720 ( .A1(n3748), .A2(n5969), .A3(n4222), .ZN(n4822) );
  INV_X1 U4721 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6870) );
  OAI21_X1 U4722 ( .B1(n3835), .B2(n6870), .A(n3872), .ZN(n6778) );
  NAND2_X1 U4723 ( .A1(n6809), .A2(n6778), .ZN(n6815) );
  NOR2_X1 U4724 ( .A1(n6815), .A2(n6810), .ZN(n5859) );
  NAND3_X1 U4725 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5859), .A3(n4223), .ZN(n6375) );
  NOR2_X1 U4726 ( .A1(n6379), .A2(n6375), .ZN(n4231) );
  INV_X1 U4727 ( .A(n4231), .ZN(n4224) );
  OR2_X1 U4728 ( .A1(n5878), .A2(n4224), .ZN(n4225) );
  NAND2_X1 U4729 ( .A1(n4226), .A2(n4225), .ZN(n4227) );
  INV_X1 U4730 ( .A(n6352), .ZN(n6212) );
  NAND2_X1 U4731 ( .A1(n4227), .A2(n6212), .ZN(n6339) );
  NOR2_X1 U4732 ( .A1(n6339), .A2(n6323), .ZN(n6864) );
  NAND2_X1 U4733 ( .A1(n6864), .A2(n3542), .ZN(n6310) );
  INV_X1 U4734 ( .A(n6310), .ZN(n4228) );
  AND2_X1 U4735 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U4736 ( .A1(n4228), .A2(n6298), .ZN(n6292) );
  INV_X1 U4737 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4229) );
  NOR4_X1 U4738 ( .A1(n6292), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4747), 
        .A4(n4229), .ZN(n4230) );
  NOR2_X2 U4739 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5764) );
  AND2_X1 U4740 ( .A1(n5764), .A2(n7077), .ZN(n5212) );
  AND2_X2 U4741 ( .A1(n5212), .A2(n7096), .ZN(n6847) );
  AND2_X1 U4742 ( .A1(n6847), .A2(REIP_REG_31__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U4743 ( .A1(n5857), .A2(n5878), .ZN(n6790) );
  INV_X1 U4744 ( .A(n6790), .ZN(n4883) );
  INV_X1 U4745 ( .A(n5878), .ZN(n6816) );
  OR2_X1 U4746 ( .A1(n6378), .A2(n6816), .ZN(n4239) );
  INV_X1 U4747 ( .A(n6323), .ZN(n4238) );
  NOR2_X1 U4748 ( .A1(n5878), .A2(n4231), .ZN(n6345) );
  OR2_X1 U4749 ( .A1(n6345), .A2(n6352), .ZN(n4237) );
  OR2_X1 U4750 ( .A1(n5857), .A2(n4232), .ZN(n4236) );
  OR2_X1 U4751 ( .A1(n5904), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4235)
         );
  OR2_X1 U4752 ( .A1(n4233), .A2(n6847), .ZN(n4234) );
  NAND2_X1 U4753 ( .A1(n4236), .A2(n6818), .ZN(n6344) );
  AOI21_X1 U4754 ( .B1(n6790), .B2(n4237), .A(n6344), .ZN(n6333) );
  OAI21_X1 U4755 ( .B1(n6339), .B2(n4238), .A(n6333), .ZN(n6862) );
  AOI21_X1 U4756 ( .B1(n4240), .B2(n4239), .A(n6862), .ZN(n6318) );
  OAI21_X1 U4757 ( .B1(n4883), .B2(n6298), .A(n6318), .ZN(n6294) );
  AOI21_X1 U4758 ( .B1(n4747), .B2(n6790), .A(n6294), .ZN(n4746) );
  INV_X1 U4759 ( .A(n6318), .ZN(n6312) );
  OAI21_X1 U4760 ( .B1(n6312), .B2(n6790), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n4241) );
  AOI21_X1 U4761 ( .B1(n4746), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4241), 
        .ZN(n4242) );
  INV_X2 U4762 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7076) );
  NOR2_X2 U4763 ( .A1(n3718), .A2(n7076), .ZN(n4431) );
  NAND2_X1 U4764 ( .A1(n4244), .A2(n4431), .ZN(n4245) );
  NAND2_X1 U4765 ( .A1(n7076), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4280) );
  NAND2_X1 U4766 ( .A1(n4914), .A2(n4431), .ZN(n4250) );
  NOR2_X2 U4767 ( .A1(n4868), .A2(n7076), .ZN(n4284) );
  AOI22_X1 U4768 ( .A1(n4721), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n7076), .ZN(n4248) );
  AND2_X1 U4769 ( .A1(n4091), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4254) );
  NAND2_X1 U4770 ( .A1(n4254), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4247) );
  AND2_X1 U4771 ( .A1(n4248), .A2(n4247), .ZN(n4249) );
  NAND2_X1 U4772 ( .A1(n4250), .A2(n4249), .ZN(n4789) );
  AND2_X1 U4773 ( .A1(n3746), .A2(n4868), .ZN(n4251) );
  AOI21_X1 U4774 ( .B1(n4915), .B2(n4251), .A(n7076), .ZN(n4869) );
  INV_X1 U4775 ( .A(n4254), .ZN(n4271) );
  NAND2_X1 U4776 ( .A1(n5972), .A2(n4431), .ZN(n4253) );
  AOI22_X1 U4777 ( .A1(n4721), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n7076), .ZN(n4252) );
  OAI211_X1 U4778 ( .C1(n4271), .C2(n3510), .A(n4253), .B(n4252), .ZN(n4870)
         );
  NAND2_X1 U4779 ( .A1(n4873), .A2(n4874), .ZN(n4260) );
  NAND2_X1 U4780 ( .A1(n4254), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4259) );
  INV_X1 U4781 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4256) );
  NAND2_X1 U4782 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4261) );
  OAI21_X1 U4783 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4261), .ZN(n6727) );
  NAND2_X1 U4784 ( .A1(n5203), .A2(n6727), .ZN(n4255) );
  OAI21_X1 U4785 ( .B1(n4280), .B2(n4256), .A(n4255), .ZN(n4257) );
  AOI21_X1 U4786 ( .B1(n4721), .B2(EAX_REG_2__SCAN_IN), .A(n4257), .ZN(n4258)
         );
  AND2_X1 U4787 ( .A1(n4259), .A2(n4258), .ZN(n4875) );
  INV_X1 U4788 ( .A(n4261), .ZN(n4263) );
  INV_X1 U4789 ( .A(n4272), .ZN(n4262) );
  OAI21_X1 U4790 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4263), .A(n4262), 
        .ZN(n5247) );
  AOI22_X1 U4791 ( .A1(n5203), .A2(n5247), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U4792 ( .A1(n4721), .A2(EAX_REG_3__SCAN_IN), .ZN(n4264) );
  OAI211_X1 U4793 ( .C1(n4271), .C2(n3581), .A(n4265), .B(n4264), .ZN(n4266)
         );
  AOI21_X1 U4794 ( .B1(n4267), .B2(n4431), .A(n4266), .ZN(n4268) );
  INV_X1 U4795 ( .A(n4268), .ZN(n4892) );
  NAND3_X1 U4796 ( .A1(n4878), .A2(n4892), .A3(n4877), .ZN(n4853) );
  INV_X1 U4797 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7040) );
  INV_X1 U4798 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6581) );
  OAI21_X1 U4799 ( .B1(n6581), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7076), 
        .ZN(n4270) );
  NAND2_X1 U4800 ( .A1(n4721), .A2(EAX_REG_4__SCAN_IN), .ZN(n4269) );
  OAI211_X1 U4801 ( .C1(n4271), .C2(n7040), .A(n4270), .B(n4269), .ZN(n4275)
         );
  NOR2_X1 U4802 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n4272), .ZN(n4273)
         );
  NOR2_X1 U4803 ( .A1(n4278), .A2(n4273), .ZN(n5668) );
  NAND2_X1 U4804 ( .A1(n5668), .A2(n4716), .ZN(n4274) );
  AND2_X1 U4805 ( .A1(n4275), .A2(n4274), .ZN(n4276) );
  INV_X1 U4806 ( .A(n4431), .ZN(n4419) );
  NOR2_X1 U4807 ( .A1(n4278), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4279)
         );
  NOR2_X1 U4808 ( .A1(n4285), .A2(n4279), .ZN(n5652) );
  INV_X1 U4809 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5650) );
  OAI22_X1 U4810 ( .A1(n5652), .A2(n4689), .B1(n4280), .B2(n5650), .ZN(n4281)
         );
  AOI21_X1 U4811 ( .B1(n4284), .B2(EAX_REG_5__SCAN_IN), .A(n4281), .ZN(n4282)
         );
  NAND2_X1 U4812 ( .A1(n4845), .A2(n4848), .ZN(n4846) );
  INV_X1 U4813 ( .A(n4846), .ZN(n4295) );
  INV_X1 U4814 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4291) );
  INV_X1 U4815 ( .A(n4296), .ZN(n4289) );
  INV_X1 U4816 ( .A(n4285), .ZN(n4287) );
  INV_X1 U4817 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4286) );
  NAND2_X1 U4818 ( .A1(n4287), .A2(n4286), .ZN(n4288) );
  NAND2_X1 U4819 ( .A1(n4289), .A2(n4288), .ZN(n6888) );
  AOI22_X1 U4820 ( .A1(n6888), .A2(n4716), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4290) );
  OAI21_X1 U4821 ( .B1(n4327), .B2(n4291), .A(n4290), .ZN(n4292) );
  NAND2_X1 U4822 ( .A1(n4295), .A2(n4294), .ZN(n5098) );
  INV_X1 U4823 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4298) );
  OAI21_X1 U4824 ( .B1(n4296), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4315), 
        .ZN(n6901) );
  AOI22_X1 U4825 ( .A1(n6901), .A2(n4716), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4297) );
  OAI21_X1 U4826 ( .B1(n4327), .B2(n4298), .A(n4297), .ZN(n4299) );
  AOI21_X1 U4827 ( .B1(n4300), .B2(n4431), .A(n4299), .ZN(n5095) );
  NOR2_X2 U4828 ( .A1(n5098), .A2(n5095), .ZN(n5096) );
  AOI22_X1 U4829 ( .A1(n4697), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U4830 ( .A1(n3467), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U4831 ( .A1(n3434), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3458), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4302) );
  AOI22_X1 U4832 ( .A1(n3798), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4301) );
  NAND4_X1 U4833 ( .A1(n4304), .A2(n4303), .A3(n4302), .A4(n4301), .ZN(n4310)
         );
  AOI22_X1 U4834 ( .A1(n4485), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4308) );
  AOI22_X1 U4835 ( .A1(n4696), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4307) );
  AOI22_X1 U4836 ( .A1(n4698), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4306) );
  AOI22_X1 U4837 ( .A1(n3447), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4305) );
  NAND4_X1 U4838 ( .A1(n4308), .A2(n4307), .A3(n4306), .A4(n4305), .ZN(n4309)
         );
  OAI21_X1 U4839 ( .B1(n4310), .B2(n4309), .A(n4431), .ZN(n4314) );
  NAND2_X1 U4840 ( .A1(n4721), .A2(EAX_REG_8__SCAN_IN), .ZN(n4313) );
  INV_X1 U4841 ( .A(n4315), .ZN(n4311) );
  XNOR2_X1 U4842 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4311), .ZN(n5488) );
  AOI22_X1 U4843 ( .A1(n5203), .A2(n5488), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4312) );
  NAND3_X1 U4844 ( .A1(n4314), .A2(n4313), .A3(n4312), .ZN(n5196) );
  INV_X1 U4845 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5453) );
  XNOR2_X1 U4846 ( .A(n5453), .B(n4330), .ZN(n5747) );
  AOI22_X1 U4847 ( .A1(n4697), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U4848 ( .A1(n4485), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4318) );
  AOI22_X1 U4849 ( .A1(n3467), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U4850 ( .A1(n3468), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4316) );
  NAND4_X1 U4851 ( .A1(n4319), .A2(n4318), .A3(n4317), .A4(n4316), .ZN(n4325)
         );
  AOI22_X1 U4852 ( .A1(n3458), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U4853 ( .A1(n4698), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U4854 ( .A1(n3434), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U4855 ( .A1(n3776), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4320) );
  NAND4_X1 U4856 ( .A1(n4323), .A2(n4322), .A3(n4321), .A4(n4320), .ZN(n4324)
         );
  OR2_X1 U4857 ( .A1(n4325), .A2(n4324), .ZN(n4326) );
  AOI22_X1 U4858 ( .A1(n4431), .A2(n4326), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4329) );
  NAND2_X1 U4859 ( .A1(n4284), .A2(EAX_REG_9__SCAN_IN), .ZN(n4328) );
  OAI211_X1 U4860 ( .C1(n5747), .C2(n4689), .A(n4329), .B(n4328), .ZN(n5446)
         );
  INV_X1 U4861 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4331) );
  XNOR2_X1 U4862 ( .A(n4347), .B(n4331), .ZN(n5737) );
  AOI22_X1 U4863 ( .A1(n4697), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U4864 ( .A1(n3467), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4335) );
  AOI22_X1 U4865 ( .A1(n3434), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U4866 ( .A1(n3447), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4333) );
  NAND4_X1 U4867 ( .A1(n4336), .A2(n4335), .A3(n4334), .A4(n4333), .ZN(n4342)
         );
  AOI22_X1 U4868 ( .A1(n3465), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U4869 ( .A1(n3456), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U4870 ( .A1(n3469), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U4871 ( .A1(n4698), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4337) );
  NAND4_X1 U4872 ( .A1(n4340), .A2(n4339), .A3(n4338), .A4(n4337), .ZN(n4341)
         );
  OAI21_X1 U4873 ( .B1(n4342), .B2(n4341), .A(n4431), .ZN(n4345) );
  NAND2_X1 U4874 ( .A1(n4721), .A2(EAX_REG_10__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U4875 ( .A1(n4720), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4343)
         );
  NAND3_X1 U4876 ( .A1(n4345), .A2(n4344), .A3(n4343), .ZN(n4346) );
  AOI21_X1 U4877 ( .B1(n5737), .B2(n5203), .A(n4346), .ZN(n5493) );
  XNOR2_X1 U4878 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4363), .ZN(n6907)
         );
  AOI22_X1 U4879 ( .A1(n4697), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4351) );
  AOI22_X1 U4880 ( .A1(n3798), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U4881 ( .A1(n3458), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U4882 ( .A1(n4698), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4348) );
  NAND4_X1 U4883 ( .A1(n4351), .A2(n4350), .A3(n4349), .A4(n4348), .ZN(n4357)
         );
  AOI22_X1 U4884 ( .A1(n3465), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4355) );
  AOI22_X1 U4885 ( .A1(n3467), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U4886 ( .A1(n3468), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U4887 ( .A1(n3660), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4352) );
  NAND4_X1 U4888 ( .A1(n4355), .A2(n4354), .A3(n4353), .A4(n4352), .ZN(n4356)
         );
  OAI21_X1 U4889 ( .B1(n4357), .B2(n4356), .A(n4431), .ZN(n4360) );
  NAND2_X1 U4890 ( .A1(n4284), .A2(EAX_REG_11__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U4891 ( .A1(n4720), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4358)
         );
  NAND3_X1 U4892 ( .A1(n4360), .A2(n4359), .A3(n4358), .ZN(n4361) );
  AOI21_X1 U4893 ( .B1(n6907), .B2(n4716), .A(n4361), .ZN(n5673) );
  NOR2_X1 U4894 ( .A1(n5493), .A2(n5673), .ZN(n4393) );
  XNOR2_X1 U4895 ( .A(n4399), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5754)
         );
  NAND2_X1 U4896 ( .A1(n5754), .A2(n4716), .ZN(n4368) );
  INV_X1 U4897 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4366) );
  AOI21_X1 U4898 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5759), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4364) );
  INV_X1 U4899 ( .A(n4364), .ZN(n4365) );
  OAI21_X1 U4900 ( .B1(n4327), .B2(n4366), .A(n4365), .ZN(n4367) );
  NAND2_X1 U4901 ( .A1(n4368), .A2(n4367), .ZN(n4380) );
  AOI22_X1 U4902 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3467), .B1(n4696), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4372) );
  AOI22_X1 U4903 ( .A1(n4485), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4371) );
  AOI22_X1 U4904 ( .A1(n4697), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4370) );
  AOI22_X1 U4905 ( .A1(n4698), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4369) );
  NAND4_X1 U4906 ( .A1(n4372), .A2(n4371), .A3(n4370), .A4(n4369), .ZN(n4378)
         );
  AOI22_X1 U4907 ( .A1(n3798), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U4908 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3434), .B1(n3456), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U4909 ( .A1(n3458), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U4910 ( .A1(n3469), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4373) );
  NAND4_X1 U4911 ( .A1(n4376), .A2(n4375), .A3(n4374), .A4(n4373), .ZN(n4377)
         );
  OAI21_X1 U4912 ( .B1(n4378), .B2(n4377), .A(n4431), .ZN(n4379) );
  NAND2_X1 U4913 ( .A1(n4380), .A2(n4379), .ZN(n5749) );
  AOI22_X1 U4914 ( .A1(n4697), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4384) );
  AOI22_X1 U4915 ( .A1(n3465), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U4916 ( .A1(n3434), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4917 ( .A1(n4698), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4381) );
  NAND4_X1 U4918 ( .A1(n4384), .A2(n4383), .A3(n4382), .A4(n4381), .ZN(n4390)
         );
  AOI22_X1 U4919 ( .A1(n3798), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4388) );
  AOI22_X1 U4920 ( .A1(n4696), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U4921 ( .A1(n3468), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U4922 ( .A1(n3470), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4385) );
  NAND4_X1 U4923 ( .A1(n4388), .A2(n4387), .A3(n4386), .A4(n4385), .ZN(n4389)
         );
  OR2_X1 U4924 ( .A1(n4390), .A2(n4389), .ZN(n4391) );
  AND2_X1 U4925 ( .A1(n4431), .A2(n4391), .ZN(n4395) );
  AND2_X1 U4926 ( .A1(n5749), .A2(n4395), .ZN(n4392) );
  INV_X1 U4927 ( .A(n4395), .ZN(n4396) );
  NAND2_X1 U4928 ( .A1(n4397), .A2(n4396), .ZN(n4398) );
  OR2_X1 U4929 ( .A1(n4400), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4401)
         );
  NAND2_X1 U4930 ( .A1(n4401), .A2(n4421), .ZN(n6918) );
  NAND2_X1 U4931 ( .A1(n6918), .A2(n4716), .ZN(n4403) );
  AOI22_X1 U4932 ( .A1(n4721), .A2(EAX_REG_13__SCAN_IN), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U4933 ( .A1(n4403), .A2(n4402), .ZN(n5839) );
  NAND2_X1 U4934 ( .A1(n5836), .A2(n5839), .ZN(n5837) );
  AOI22_X1 U4935 ( .A1(n4485), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4408) );
  AOI22_X1 U4936 ( .A1(n3467), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U4937 ( .A1(n3434), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3458), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U4938 ( .A1(n3468), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4405) );
  NAND4_X1 U4939 ( .A1(n4408), .A2(n4407), .A3(n4406), .A4(n4405), .ZN(n4414)
         );
  AOI22_X1 U4940 ( .A1(n4696), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4412) );
  AOI22_X1 U4941 ( .A1(n3776), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U4942 ( .A1(n4698), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U4943 ( .A1(n4697), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4409) );
  NAND4_X1 U4944 ( .A1(n4412), .A2(n4411), .A3(n4410), .A4(n4409), .ZN(n4413)
         );
  NOR2_X1 U4945 ( .A1(n4414), .A2(n4413), .ZN(n4418) );
  XNOR2_X1 U4946 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4421), .ZN(n6933)
         );
  INV_X1 U4947 ( .A(n6933), .ZN(n4415) );
  AOI22_X1 U4948 ( .A1(n4720), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n5203), 
        .B2(n4415), .ZN(n4417) );
  NAND2_X1 U4949 ( .A1(n4284), .A2(EAX_REG_14__SCAN_IN), .ZN(n4416) );
  OAI211_X1 U4950 ( .C1(n4419), .C2(n4418), .A(n4417), .B(n4416), .ZN(n5870)
         );
  INV_X1 U4951 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4420) );
  INV_X1 U4952 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4422) );
  XNOR2_X1 U4953 ( .A(n4437), .B(n4422), .ZN(n6942) );
  OR2_X1 U4954 ( .A1(n6942), .A2(n4689), .ZN(n4436) );
  AOI22_X1 U4955 ( .A1(n4721), .A2(EAX_REG_15__SCAN_IN), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4435) );
  AOI22_X1 U4956 ( .A1(n4697), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4426) );
  AOI22_X1 U4957 ( .A1(n3457), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U4958 ( .A1(n4696), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3458), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4424) );
  AOI22_X1 U4959 ( .A1(n3470), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4423) );
  NAND4_X1 U4960 ( .A1(n4426), .A2(n4425), .A3(n4424), .A4(n4423), .ZN(n4433)
         );
  AOI22_X1 U4961 ( .A1(n4485), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U4962 ( .A1(n3434), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4429) );
  AOI22_X1 U4963 ( .A1(n3798), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U4964 ( .A1(n4698), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4427) );
  NAND4_X1 U4965 ( .A1(n4430), .A2(n4429), .A3(n4428), .A4(n4427), .ZN(n4432)
         );
  OAI21_X1 U4966 ( .B1(n4433), .B2(n4432), .A(n4431), .ZN(n4434) );
  XOR2_X1 U4967 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4452), .Z(n6955) );
  INV_X1 U4968 ( .A(n6955), .ZN(n4451) );
  NAND2_X1 U4969 ( .A1(n5969), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4671) );
  AOI22_X1 U4970 ( .A1(n3798), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4441) );
  AOI22_X1 U4971 ( .A1(n4485), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4440) );
  AOI22_X1 U4972 ( .A1(n3467), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4439) );
  AOI22_X1 U4973 ( .A1(n3470), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4438) );
  NAND4_X1 U4974 ( .A1(n4441), .A2(n4440), .A3(n4439), .A4(n4438), .ZN(n4447)
         );
  AOI22_X1 U4975 ( .A1(n4697), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U4976 ( .A1(n3458), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U4977 ( .A1(n4696), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4443) );
  AOI22_X1 U4978 ( .A1(n4698), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4442) );
  NAND4_X1 U4979 ( .A1(n4445), .A2(n4444), .A3(n4443), .A4(n4442), .ZN(n4446)
         );
  NOR2_X1 U4980 ( .A1(n4447), .A2(n4446), .ZN(n4449) );
  AOI22_X1 U4981 ( .A1(n4721), .A2(EAX_REG_16__SCAN_IN), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4448) );
  OAI21_X1 U4982 ( .B1(n4671), .B2(n4449), .A(n4448), .ZN(n4450) );
  AOI21_X1 U4983 ( .B1(n4451), .B2(n4716), .A(n4450), .ZN(n5925) );
  XNOR2_X1 U4984 ( .A(n4468), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6259)
         );
  AOI22_X1 U4985 ( .A1(n4698), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4456) );
  AOI22_X1 U4986 ( .A1(n3465), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4455) );
  AOI22_X1 U4987 ( .A1(n3467), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4454) );
  AOI22_X1 U4988 ( .A1(n3798), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4453) );
  NAND4_X1 U4989 ( .A1(n4456), .A2(n4455), .A3(n4454), .A4(n4453), .ZN(n4462)
         );
  AOI22_X1 U4990 ( .A1(n4697), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4460) );
  AOI22_X1 U4991 ( .A1(n3458), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4459) );
  AOI22_X1 U4992 ( .A1(n3470), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U4993 ( .A1(n3468), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4457) );
  NAND4_X1 U4994 ( .A1(n4460), .A2(n4459), .A3(n4458), .A4(n4457), .ZN(n4461)
         );
  OR2_X1 U4995 ( .A1(n4462), .A2(n4461), .ZN(n4466) );
  INV_X1 U4996 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U4997 ( .A1(n7076), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4463)
         );
  OAI211_X1 U4998 ( .C1(n4327), .C2(n4464), .A(n4689), .B(n4463), .ZN(n4465)
         );
  AOI21_X1 U4999 ( .B1(n4711), .B2(n4466), .A(n4465), .ZN(n4467) );
  AOI21_X1 U5000 ( .B1(n6259), .B2(n4716), .A(n4467), .ZN(n5920) );
  NAND2_X1 U5001 ( .A1(n5917), .A2(n5920), .ZN(n5918) );
  INV_X1 U5002 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5940) );
  OR2_X1 U5003 ( .A1(n4469), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4470)
         );
  NAND2_X1 U5004 ( .A1(n4470), .A2(n4501), .ZN(n6959) );
  AOI22_X1 U5005 ( .A1(n3464), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U5006 ( .A1(n4696), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U5007 ( .A1(n3458), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5008 ( .A1(n3469), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4471) );
  NAND4_X1 U5009 ( .A1(n4474), .A2(n4473), .A3(n4472), .A4(n4471), .ZN(n4480)
         );
  AOI22_X1 U5010 ( .A1(n3467), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4478) );
  AOI22_X1 U5011 ( .A1(n3776), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U5012 ( .A1(n4698), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4476) );
  AOI22_X1 U5013 ( .A1(n4697), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4475) );
  NAND4_X1 U5014 ( .A1(n4478), .A2(n4477), .A3(n4476), .A4(n4475), .ZN(n4479)
         );
  NOR2_X1 U5015 ( .A1(n4480), .A2(n4479), .ZN(n4483) );
  OAI21_X1 U5016 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6581), .A(n7076), 
        .ZN(n4482) );
  NAND2_X1 U5017 ( .A1(n4284), .A2(EAX_REG_18__SCAN_IN), .ZN(n4481) );
  OAI211_X1 U5018 ( .C1(n4671), .C2(n4483), .A(n4482), .B(n4481), .ZN(n4484)
         );
  OAI21_X1 U5019 ( .B1(n6959), .B2(n4689), .A(n4484), .ZN(n6149) );
  AOI22_X1 U5020 ( .A1(n3465), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U5021 ( .A1(n4696), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4488) );
  AOI22_X1 U5022 ( .A1(n3467), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4487) );
  AOI22_X1 U5023 ( .A1(n3700), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4486) );
  NAND4_X1 U5024 ( .A1(n4489), .A2(n4488), .A3(n4487), .A4(n4486), .ZN(n4495)
         );
  AOI22_X1 U5025 ( .A1(n4697), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4493) );
  AOI22_X1 U5026 ( .A1(n3776), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4492) );
  AOI22_X1 U5027 ( .A1(n4698), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U5028 ( .A1(n3447), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4490) );
  NAND4_X1 U5029 ( .A1(n4493), .A2(n4492), .A3(n4491), .A4(n4490), .ZN(n4494)
         );
  NOR2_X1 U5030 ( .A1(n4495), .A2(n4494), .ZN(n4498) );
  INV_X1 U5031 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6252) );
  AOI21_X1 U5032 ( .B1(n6252), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4496) );
  AOI21_X1 U5033 ( .B1(n4284), .B2(EAX_REG_19__SCAN_IN), .A(n4496), .ZN(n4497)
         );
  OAI21_X1 U5034 ( .B1(n4671), .B2(n4498), .A(n4497), .ZN(n4500) );
  XNOR2_X1 U5035 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4501), .ZN(n6971)
         );
  NAND2_X1 U5036 ( .A1(n6971), .A2(n4716), .ZN(n4499) );
  NAND2_X1 U5037 ( .A1(n4500), .A2(n4499), .ZN(n6250) );
  INV_X1 U5038 ( .A(n4534), .ZN(n4504) );
  OR2_X1 U5039 ( .A1(n4502), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4503)
         );
  NAND2_X1 U5040 ( .A1(n4504), .A2(n4503), .ZN(n6979) );
  AOI22_X1 U5041 ( .A1(n3798), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4508) );
  AOI22_X1 U5042 ( .A1(n3467), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4507) );
  AOI22_X1 U5043 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4698), .B1(n3660), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5044 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3469), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4505) );
  NAND4_X1 U5045 ( .A1(n4508), .A2(n4507), .A3(n4506), .A4(n4505), .ZN(n4514)
         );
  AOI22_X1 U5046 ( .A1(n4485), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4512) );
  AOI22_X1 U5047 ( .A1(n3700), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U5048 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3776), .B1(n3460), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U5049 ( .A1(n4697), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4509) );
  NAND4_X1 U5050 ( .A1(n4512), .A2(n4511), .A3(n4510), .A4(n4509), .ZN(n4513)
         );
  NOR2_X1 U5051 ( .A1(n4514), .A2(n4513), .ZN(n4517) );
  OAI21_X1 U5052 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6581), .A(n7076), 
        .ZN(n4516) );
  NAND2_X1 U5053 ( .A1(n4284), .A2(EAX_REG_20__SCAN_IN), .ZN(n4515) );
  OAI211_X1 U5054 ( .C1(n4671), .C2(n4517), .A(n4516), .B(n4515), .ZN(n4518)
         );
  INV_X1 U5055 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6241) );
  XNOR2_X1 U5056 ( .A(n4534), .B(n6241), .ZN(n6243) );
  AOI22_X1 U5057 ( .A1(n4698), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U5058 ( .A1(n4485), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5059 ( .A1(n3434), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U5060 ( .A1(n3776), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4520) );
  NAND4_X1 U5061 ( .A1(n4523), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(n4529)
         );
  AOI22_X1 U5062 ( .A1(n3798), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U5063 ( .A1(n3467), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5064 ( .A1(n3470), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U5065 ( .A1(n3468), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4524) );
  NAND4_X1 U5066 ( .A1(n4527), .A2(n4526), .A3(n4525), .A4(n4524), .ZN(n4528)
         );
  OR2_X1 U5067 ( .A1(n4529), .A2(n4528), .ZN(n4532) );
  NAND2_X1 U5068 ( .A1(n4284), .A2(EAX_REG_21__SCAN_IN), .ZN(n4530) );
  OAI211_X1 U5069 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6241), .A(n4530), .B(
        n4689), .ZN(n4531) );
  AOI21_X1 U5070 ( .B1(n4711), .B2(n4532), .A(n4531), .ZN(n4533) );
  AOI21_X1 U5071 ( .B1(n6243), .B2(n4716), .A(n4533), .ZN(n6103) );
  NAND2_X1 U5072 ( .A1(n6100), .A2(n6103), .ZN(n6101) );
  INV_X1 U5073 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4547) );
  AND2_X1 U5074 ( .A1(n4535), .A2(n4547), .ZN(n4536) );
  OR2_X1 U5075 ( .A1(n4536), .A2(n4578), .ZN(n7000) );
  AOI22_X1 U5076 ( .A1(n3464), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4540) );
  AOI22_X1 U5077 ( .A1(n3467), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5078 ( .A1(n3458), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5079 ( .A1(n3469), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4537) );
  NAND4_X1 U5080 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), .ZN(n4546)
         );
  AOI22_X1 U5081 ( .A1(n4696), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U5082 ( .A1(n3776), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U5083 ( .A1(n4697), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4542) );
  AOI22_X1 U5084 ( .A1(n4698), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4541) );
  NAND4_X1 U5085 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(n4545)
         );
  NOR2_X1 U5086 ( .A1(n4546), .A2(n4545), .ZN(n4550) );
  OAI21_X1 U5087 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4547), .A(n4689), .ZN(
        n4548) );
  AOI21_X1 U5088 ( .B1(n4284), .B2(EAX_REG_22__SCAN_IN), .A(n4548), .ZN(n4549)
         );
  OAI21_X1 U5089 ( .B1(n4671), .B2(n4550), .A(n4549), .ZN(n4551) );
  OAI21_X1 U5090 ( .B1(n7000), .B2(n4689), .A(n4551), .ZN(n6134) );
  NOR2_X2 U5091 ( .A1(n6101), .A2(n6134), .ZN(n6085) );
  INV_X1 U5092 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4552) );
  XNOR2_X1 U5093 ( .A(n4578), .B(n4552), .ZN(n6226) );
  AOI22_X1 U5094 ( .A1(n4697), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5095 ( .A1(n3467), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U5096 ( .A1(n3456), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5097 ( .A1(n3470), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4553) );
  NAND4_X1 U5098 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .ZN(n4562)
         );
  AOI22_X1 U5099 ( .A1(n3798), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5100 ( .A1(n3465), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U5101 ( .A1(n3458), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4558) );
  AOI22_X1 U5102 ( .A1(n4698), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4557) );
  NAND4_X1 U5103 ( .A1(n4560), .A2(n4559), .A3(n4558), .A4(n4557), .ZN(n4561)
         );
  NOR2_X1 U5104 ( .A1(n4562), .A2(n4561), .ZN(n4580) );
  AOI22_X1 U5105 ( .A1(n4485), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4566) );
  AOI22_X1 U5106 ( .A1(n4696), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5107 ( .A1(n4697), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4564) );
  AOI22_X1 U5108 ( .A1(n3469), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4563) );
  NAND4_X1 U5109 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .ZN(n4572)
         );
  AOI22_X1 U5110 ( .A1(n3467), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5111 ( .A1(n3700), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5112 ( .A1(n4698), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5113 ( .A1(n3776), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4567) );
  NAND4_X1 U5114 ( .A1(n4570), .A2(n4569), .A3(n4568), .A4(n4567), .ZN(n4571)
         );
  NOR2_X1 U5115 ( .A1(n4572), .A2(n4571), .ZN(n4579) );
  XOR2_X1 U5116 ( .A(n4580), .B(n4579), .Z(n4576) );
  INV_X1 U5117 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4574) );
  OAI21_X1 U5118 ( .B1(n6581), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n7076), 
        .ZN(n4573) );
  OAI21_X1 U5119 ( .B1(n4327), .B2(n4574), .A(n4573), .ZN(n4575) );
  AOI21_X1 U5120 ( .B1(n4711), .B2(n4576), .A(n4575), .ZN(n4577) );
  AOI21_X1 U5121 ( .B1(n6226), .B2(n4716), .A(n4577), .ZN(n6088) );
  NAND2_X1 U5122 ( .A1(n4578), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4609)
         );
  XNOR2_X1 U5123 ( .A(n4609), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n7018)
         );
  INV_X1 U5124 ( .A(n7018), .ZN(n6220) );
  OR2_X1 U5125 ( .A1(n4580), .A2(n4579), .ZN(n4605) );
  AOI22_X1 U5126 ( .A1(n4698), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U5127 ( .A1(n4697), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U5128 ( .A1(n3465), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4582) );
  AOI22_X1 U5129 ( .A1(n3469), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4581) );
  NAND4_X1 U5130 ( .A1(n4584), .A2(n4583), .A3(n4582), .A4(n4581), .ZN(n4590)
         );
  AOI22_X1 U5131 ( .A1(n3456), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U5132 ( .A1(n3467), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3458), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5133 ( .A1(n4679), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U5134 ( .A1(n3776), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4585) );
  NAND4_X1 U5135 ( .A1(n4588), .A2(n4587), .A3(n4586), .A4(n4585), .ZN(n4589)
         );
  NOR2_X1 U5136 ( .A1(n4590), .A2(n4589), .ZN(n4604) );
  XNOR2_X1 U5137 ( .A(n4605), .B(n4604), .ZN(n4592) );
  AOI22_X1 U5138 ( .A1(n4721), .A2(EAX_REG_24__SCAN_IN), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4591) );
  OAI21_X1 U5139 ( .B1(n4592), .B2(n4671), .A(n4591), .ZN(n4593) );
  AOI21_X1 U5140 ( .B1(n6220), .B2(n4716), .A(n4593), .ZN(n6218) );
  AOI22_X1 U5141 ( .A1(n4697), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4597) );
  AOI22_X1 U5142 ( .A1(n3798), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4596) );
  AOI22_X1 U5143 ( .A1(n3467), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3700), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U5144 ( .A1(n3470), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4594) );
  NAND4_X1 U5145 ( .A1(n4597), .A2(n4596), .A3(n4595), .A4(n4594), .ZN(n4603)
         );
  AOI22_X1 U5146 ( .A1(n3464), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3457), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5147 ( .A1(n3434), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4600) );
  AOI22_X1 U5148 ( .A1(n3468), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5149 ( .A1(n4698), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4598) );
  NAND4_X1 U5150 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(n4602)
         );
  NOR2_X1 U5151 ( .A1(n4603), .A2(n4602), .ZN(n4619) );
  OR2_X1 U5152 ( .A1(n4605), .A2(n4604), .ZN(n4618) );
  XOR2_X1 U5153 ( .A(n4619), .B(n4618), .Z(n4606) );
  NAND2_X1 U5154 ( .A1(n4606), .A2(n4711), .ZN(n4612) );
  INV_X1 U5155 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6076) );
  AOI21_X1 U5156 ( .B1(n6076), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4607) );
  AOI21_X1 U5157 ( .B1(n4284), .B2(EAX_REG_25__SCAN_IN), .A(n4607), .ZN(n4611)
         );
  INV_X1 U5158 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4608) );
  XNOR2_X1 U5159 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4613), .ZN(n6078)
         );
  AOI21_X1 U5160 ( .B1(n4612), .B2(n4611), .A(n4610), .ZN(n6068) );
  INV_X1 U5161 ( .A(n4615), .ZN(n4616) );
  INV_X1 U5162 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U5163 ( .A1(n4616), .A2(n6059), .ZN(n4617) );
  NAND2_X1 U5164 ( .A1(n4651), .A2(n4617), .ZN(n6201) );
  NOR2_X1 U5165 ( .A1(n4619), .A2(n4618), .ZN(n4645) );
  AOI22_X1 U5166 ( .A1(n3464), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5167 ( .A1(n4696), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4622) );
  AOI22_X1 U5168 ( .A1(n3467), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4621) );
  AOI22_X1 U5169 ( .A1(n3458), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4620) );
  NAND4_X1 U5170 ( .A1(n4623), .A2(n4622), .A3(n4621), .A4(n4620), .ZN(n4629)
         );
  AOI22_X1 U5171 ( .A1(n4697), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4627) );
  AOI22_X1 U5172 ( .A1(n3776), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4626) );
  AOI22_X1 U5173 ( .A1(n4698), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4625) );
  AOI22_X1 U5174 ( .A1(n3447), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4624) );
  NAND4_X1 U5175 ( .A1(n4627), .A2(n4626), .A3(n4625), .A4(n4624), .ZN(n4628)
         );
  OR2_X1 U5176 ( .A1(n4629), .A2(n4628), .ZN(n4644) );
  XNOR2_X1 U5177 ( .A(n4645), .B(n4644), .ZN(n4632) );
  AOI21_X1 U5178 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n7076), .A(n5203), 
        .ZN(n4631) );
  NAND2_X1 U5179 ( .A1(n4284), .A2(EAX_REG_26__SCAN_IN), .ZN(n4630) );
  OAI211_X1 U5180 ( .C1(n4632), .C2(n4671), .A(n4631), .B(n4630), .ZN(n4633)
         );
  OAI21_X1 U5181 ( .B1(n4689), .B2(n6201), .A(n4633), .ZN(n6058) );
  AOI22_X1 U5182 ( .A1(n3464), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4637) );
  AOI22_X1 U5183 ( .A1(n3467), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5184 ( .A1(n3434), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3458), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U5185 ( .A1(n3468), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4634) );
  NAND4_X1 U5186 ( .A1(n4637), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4643)
         );
  AOI22_X1 U5187 ( .A1(n4696), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4641) );
  AOI22_X1 U5188 ( .A1(n4698), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5189 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3798), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5190 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3776), .B1(n3447), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4638) );
  NAND4_X1 U5191 ( .A1(n4641), .A2(n4640), .A3(n4639), .A4(n4638), .ZN(n4642)
         );
  NOR2_X1 U5192 ( .A1(n4643), .A2(n4642), .ZN(n4657) );
  NAND2_X1 U5193 ( .A1(n4645), .A2(n4644), .ZN(n4656) );
  XOR2_X1 U5194 ( .A(n4657), .B(n4656), .Z(n4646) );
  NAND2_X1 U5195 ( .A1(n4646), .A2(n4711), .ZN(n4649) );
  INV_X1 U5196 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4650) );
  AOI21_X1 U5197 ( .B1(n4650), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4647) );
  AOI21_X1 U5198 ( .B1(n4284), .B2(EAX_REG_27__SCAN_IN), .A(n4647), .ZN(n4648)
         );
  XNOR2_X1 U5199 ( .A(n4651), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6050)
         );
  NAND2_X1 U5200 ( .A1(n4652), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4715)
         );
  INV_X1 U5201 ( .A(n4652), .ZN(n4654) );
  INV_X1 U5202 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U5203 ( .A1(n4654), .A2(n4653), .ZN(n4655) );
  NAND2_X1 U5204 ( .A1(n4715), .A2(n4655), .ZN(n6186) );
  NOR2_X1 U5205 ( .A1(n4657), .A2(n4656), .ZN(n4687) );
  AOI22_X1 U5206 ( .A1(n3465), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5207 ( .A1(n4696), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5208 ( .A1(n3467), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5209 ( .A1(n3458), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4659) );
  NAND4_X1 U5210 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4668)
         );
  AOI22_X1 U5211 ( .A1(n4697), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5212 ( .A1(n3776), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4665) );
  AOI22_X1 U5213 ( .A1(n4698), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U5214 ( .A1(n3447), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4663) );
  NAND4_X1 U5215 ( .A1(n4666), .A2(n4665), .A3(n4664), .A4(n4663), .ZN(n4667)
         );
  OR2_X1 U5216 ( .A1(n4668), .A2(n4667), .ZN(n4686) );
  XNOR2_X1 U5217 ( .A(n4687), .B(n4686), .ZN(n4672) );
  AOI21_X1 U5218 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n7076), .A(n5203), 
        .ZN(n4670) );
  NAND2_X1 U5219 ( .A1(n4721), .A2(EAX_REG_28__SCAN_IN), .ZN(n4669) );
  OAI211_X1 U5220 ( .C1(n4672), .C2(n4671), .A(n4670), .B(n4669), .ZN(n4673)
         );
  OAI21_X1 U5221 ( .B1(n4689), .B2(n6186), .A(n4673), .ZN(n6033) );
  XNOR2_X1 U5222 ( .A(n4715), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6021)
         );
  AOI22_X1 U5223 ( .A1(n4697), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5224 ( .A1(n3464), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4677) );
  AOI22_X1 U5225 ( .A1(n4696), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5226 ( .A1(n3660), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4675) );
  NAND4_X1 U5227 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4685)
         );
  AOI22_X1 U5228 ( .A1(n3467), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4683) );
  AOI22_X1 U5229 ( .A1(n3458), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4682) );
  AOI22_X1 U5230 ( .A1(n3776), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4681) );
  AOI22_X1 U5231 ( .A1(n4698), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4680) );
  NAND4_X1 U5232 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .ZN(n4684)
         );
  NOR2_X1 U5233 ( .A1(n4685), .A2(n4684), .ZN(n4695) );
  NAND2_X1 U5234 ( .A1(n4687), .A2(n4686), .ZN(n4694) );
  XOR2_X1 U5235 ( .A(n4695), .B(n4694), .Z(n4692) );
  INV_X1 U5236 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U5237 ( .A1(n7076), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4688)
         );
  OAI211_X1 U5238 ( .C1(n4327), .C2(n4690), .A(n4689), .B(n4688), .ZN(n4691)
         );
  AOI21_X1 U5239 ( .B1(n4692), .B2(n4711), .A(n4691), .ZN(n4693) );
  AOI21_X1 U5240 ( .B1(n4716), .B2(n6021), .A(n4693), .ZN(n4762) );
  NOR2_X1 U5241 ( .A1(n4695), .A2(n4694), .ZN(n4710) );
  AOI22_X1 U5242 ( .A1(n3465), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4696), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4702) );
  AOI22_X1 U5243 ( .A1(n3798), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5244 ( .A1(n4697), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4700) );
  AOI22_X1 U5245 ( .A1(n4698), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3681), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4699) );
  NAND4_X1 U5246 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4699), .ZN(n4708)
         );
  AOI22_X1 U5247 ( .A1(n3456), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U5248 ( .A1(n3467), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5249 ( .A1(n3700), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4679), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5250 ( .A1(n3468), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4703) );
  NAND4_X1 U5251 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .ZN(n4707)
         );
  NOR2_X1 U5252 ( .A1(n4708), .A2(n4707), .ZN(n4709) );
  XNOR2_X1 U5253 ( .A(n4710), .B(n4709), .ZN(n4712) );
  NAND2_X1 U5254 ( .A1(n4712), .A2(n4711), .ZN(n4719) );
  INV_X1 U5255 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4713) );
  AOI21_X1 U5256 ( .B1(n4713), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4714) );
  AOI21_X1 U5257 ( .B1(n4284), .B2(EAX_REG_30__SCAN_IN), .A(n4714), .ZN(n4718)
         );
  INV_X1 U5258 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6022) );
  XNOR2_X1 U5259 ( .A(n4729), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5977)
         );
  AND2_X1 U5260 ( .A1(n5977), .A2(n4716), .ZN(n4717) );
  AOI22_X1 U5261 ( .A1(n4721), .A2(EAX_REG_31__SCAN_IN), .B1(n4720), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4722) );
  INV_X1 U5262 ( .A(n4722), .ZN(n4723) );
  NOR2_X1 U5263 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7077), .ZN(n5202) );
  NAND2_X1 U5264 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5202), .ZN(n6767) );
  INV_X1 U5265 ( .A(n6767), .ZN(n4724) );
  NAND2_X1 U5266 ( .A1(n5764), .A2(n4724), .ZN(n6742) );
  OR2_X1 U5267 ( .A1(n4725), .A2(n5764), .ZN(n6770) );
  NAND2_X1 U5268 ( .A1(n6770), .A2(n7096), .ZN(n4726) );
  AND2_X2 U5269 ( .A1(n7033), .A2(n4726), .ZN(n6749) );
  NAND2_X1 U5270 ( .A1(n7096), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4728) );
  NAND2_X1 U5271 ( .A1(n6581), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4727) );
  AND2_X1 U5272 ( .A1(n4728), .A2(n4727), .ZN(n6709) );
  INV_X1 U5273 ( .A(n4729), .ZN(n4730) );
  NAND2_X1 U5274 ( .A1(n4730), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4731)
         );
  INV_X1 U5275 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6009) );
  XNOR2_X1 U5276 ( .A(n4731), .B(n6009), .ZN(n5227) );
  AOI21_X1 U5277 ( .B1(n6749), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4732), 
        .ZN(n4733) );
  OAI21_X1 U5278 ( .B1(n4736), .B2(n7033), .A(n4735), .ZN(U2955) );
  NAND2_X1 U5279 ( .A1(n3453), .A2(n6369), .ZN(n4737) );
  XNOR2_X1 U5280 ( .A(n4740), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5984)
         );
  INV_X1 U5281 ( .A(n4768), .ZN(n6029) );
  XNOR2_X2 U5282 ( .A(n4745), .B(n4744), .ZN(n5968) );
  INV_X1 U5283 ( .A(n5968), .ZN(n4751) );
  INV_X1 U5284 ( .A(n4746), .ZN(n6277) );
  AND2_X1 U5285 ( .A1(n6847), .A2(REIP_REG_30__SCAN_IN), .ZN(n5978) );
  NOR3_X1 U5286 ( .A1(n6292), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4747), 
        .ZN(n4748) );
  AOI211_X1 U5287 ( .C1(n6277), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5978), .B(n4748), .ZN(n4749) );
  OAI21_X1 U5288 ( .B1(n5984), .B2(n6878), .A(n4752), .ZN(U2988) );
  XNOR2_X1 U5289 ( .A(n4764), .B(n4754), .ZN(n5982) );
  INV_X1 U5290 ( .A(n5982), .ZN(n5954) );
  NAND2_X1 U5291 ( .A1(n7026), .A2(n4822), .ZN(n4804) );
  NOR2_X1 U5292 ( .A1(n3820), .A2(n4755), .ZN(n4756) );
  INV_X1 U5293 ( .A(n4868), .ZN(n6016) );
  NAND4_X1 U5294 ( .A1(n4756), .A2(n6016), .A3(n3720), .A4(n3718), .ZN(n4861)
         );
  INV_X1 U5295 ( .A(n4861), .ZN(n4757) );
  NAND3_X1 U5296 ( .A1(n4757), .A2(n4944), .A3(n4791), .ZN(n4758) );
  NAND2_X1 U5297 ( .A1(n4804), .A2(n4758), .ZN(n4759) );
  INV_X1 U5298 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5961) );
  OAI21_X1 U5299 ( .B1(n5954), .B2(n6156), .A(n4761), .ZN(U2829) );
  INV_X1 U5300 ( .A(n4762), .ZN(n4766) );
  INV_X1 U5301 ( .A(n4763), .ZN(n4765) );
  AOI21_X2 U5302 ( .B1(n4766), .B2(n4765), .A(n4764), .ZN(n6179) );
  INV_X1 U5303 ( .A(n6179), .ZN(n6160) );
  OAI21_X1 U5304 ( .B1(n4768), .B2(n4767), .A(n3471), .ZN(n6275) );
  NAND2_X1 U5305 ( .A1(n4769), .A2(EBX_REG_29__SCAN_IN), .ZN(n4770) );
  INV_X1 U5306 ( .A(n4774), .ZN(n6757) );
  INV_X1 U5307 ( .A(n7030), .ZN(n4775) );
  NOR2_X1 U5308 ( .A1(n4775), .A2(n7029), .ZN(n6756) );
  NAND2_X1 U5309 ( .A1(n6756), .A2(n7092), .ZN(n7118) );
  NAND2_X1 U5310 ( .A1(n6773), .A2(n5213), .ZN(n6772) );
  INV_X1 U5311 ( .A(n5212), .ZN(n4776) );
  NAND2_X1 U5312 ( .A1(n7122), .A2(n4776), .ZN(n7117) );
  INV_X1 U5313 ( .A(n7118), .ZN(n4777) );
  NOR3_X1 U5314 ( .A1(n7117), .A2(n4777), .A3(READREQUEST_REG_SCAN_IN), .ZN(
        n4778) );
  AOI21_X1 U5315 ( .B1(n6769), .B2(n6772), .A(n4778), .ZN(U3474) );
  INV_X1 U5316 ( .A(EAX_REG_21__SCAN_IN), .ZN(n7151) );
  INV_X1 U5317 ( .A(n7069), .ZN(n7120) );
  INV_X1 U5318 ( .A(n6771), .ZN(n4794) );
  OAI21_X1 U5319 ( .B1(n7120), .B2(n5010), .A(n4794), .ZN(n4779) );
  NAND2_X1 U5320 ( .A1(n6613), .A2(n4097), .ZN(n4844) );
  AND2_X2 U5321 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5202), .ZN(n6631) );
  AOI22_X1 U5322 ( .A1(n6631), .A2(UWORD_REG_5__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4781) );
  OAI21_X1 U5323 ( .B1(n7151), .B2(n4844), .A(n4781), .ZN(U2902) );
  INV_X1 U5324 ( .A(EAX_REG_22__SCAN_IN), .ZN(n7156) );
  AOI22_X1 U5325 ( .A1(n6631), .A2(UWORD_REG_6__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4782) );
  OAI21_X1 U5326 ( .B1(n7156), .B2(n4844), .A(n4782), .ZN(U2901) );
  INV_X1 U5327 ( .A(EAX_REG_25__SCAN_IN), .ZN(n7168) );
  AOI22_X1 U5328 ( .A1(n6631), .A2(UWORD_REG_9__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4783) );
  OAI21_X1 U5329 ( .B1(n7168), .B2(n4844), .A(n4783), .ZN(U2898) );
  INV_X1 U5330 ( .A(EAX_REG_24__SCAN_IN), .ZN(n7163) );
  AOI22_X1 U5331 ( .A1(n6631), .A2(UWORD_REG_8__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4784) );
  OAI21_X1 U5332 ( .B1(n7163), .B2(n4844), .A(n4784), .ZN(U2899) );
  INV_X1 U5333 ( .A(EAX_REG_20__SCAN_IN), .ZN(n7146) );
  AOI22_X1 U5334 ( .A1(n6631), .A2(UWORD_REG_4__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4785) );
  OAI21_X1 U5335 ( .B1(n7146), .B2(n4844), .A(n4785), .ZN(U2903) );
  AOI22_X1 U5336 ( .A1(n6631), .A2(UWORD_REG_7__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4786) );
  OAI21_X1 U5337 ( .B1(n4574), .B2(n4844), .A(n4786), .ZN(U2900) );
  INV_X1 U5338 ( .A(EAX_REG_26__SCAN_IN), .ZN(n7173) );
  AOI22_X1 U5339 ( .A1(n6631), .A2(UWORD_REG_10__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4787) );
  OAI21_X1 U5340 ( .B1(n7173), .B2(n4844), .A(n4787), .ZN(U2897) );
  NOR2_X1 U5341 ( .A1(n4789), .A2(n4788), .ZN(n4790) );
  OR2_X1 U5342 ( .A1(n4874), .A2(n4790), .ZN(n6714) );
  XNOR2_X1 U5343 ( .A(n6122), .B(n4791), .ZN(n4888) );
  AOI22_X1 U5344 ( .A1(n6702), .A2(n4888), .B1(EBX_REG_1__SCAN_IN), .B2(n4769), 
        .ZN(n4792) );
  OAI21_X1 U5345 ( .B1(n6156), .B2(n6714), .A(n4792), .ZN(U2858) );
  NAND2_X1 U5346 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7096), .ZN(n7082) );
  INV_X1 U5347 ( .A(n7082), .ZN(n4808) );
  INV_X1 U5348 ( .A(n4793), .ZN(n4797) );
  NAND2_X1 U5349 ( .A1(n5010), .A2(n4794), .ZN(n4795) );
  NAND2_X1 U5350 ( .A1(n4795), .A2(n4774), .ZN(n4796) );
  NAND2_X1 U5351 ( .A1(n4797), .A2(n4796), .ZN(n4807) );
  OR2_X1 U5352 ( .A1(n7026), .A2(n4823), .ZN(n4800) );
  NAND2_X1 U5353 ( .A1(n5024), .A2(n4798), .ZN(n4799) );
  NAND2_X1 U5354 ( .A1(n4800), .A2(n4799), .ZN(n4864) );
  INV_X1 U5355 ( .A(n4864), .ZN(n4806) );
  INV_X1 U5356 ( .A(n4801), .ZN(n4802) );
  AND3_X1 U5357 ( .A1(n4804), .A2(n4803), .A3(n4802), .ZN(n4805) );
  INV_X1 U5358 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7034) );
  NOR2_X1 U5359 ( .A1(n7076), .A2(n7077), .ZN(n5364) );
  NAND2_X1 U5360 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5364), .ZN(n7083) );
  OAI22_X1 U5361 ( .A1(n7047), .A2(n7073), .B1(n7034), .B2(n7083), .ZN(n7037)
         );
  NOR2_X1 U5362 ( .A1(n4808), .A2(n7037), .ZN(n5999) );
  NOR2_X1 U5363 ( .A1(n4809), .A2(n4810), .ZN(n4816) );
  AND3_X1 U5364 ( .A1(n4070), .A2(n4812), .A3(n4862), .ZN(n4813) );
  NAND2_X1 U5365 ( .A1(n4814), .A2(n4813), .ZN(n5971) );
  NAND2_X1 U5366 ( .A1(n4811), .A2(n5971), .ZN(n4815) );
  NAND2_X1 U5367 ( .A1(n5010), .A2(n3582), .ZN(n5003) );
  OAI211_X1 U5368 ( .C1(n4816), .C2(n3736), .A(n4815), .B(n5003), .ZN(n7042)
         );
  INV_X1 U5369 ( .A(n7075), .ZN(n6003) );
  AOI22_X1 U5370 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4015), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3835), .ZN(n4832) );
  NAND2_X1 U5371 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4831) );
  INV_X1 U5372 ( .A(n4831), .ZN(n4818) );
  INV_X1 U5373 ( .A(n4816), .ZN(n4817) );
  AOI222_X1 U5374 ( .A1(n7042), .A2(n6003), .B1(n4832), .B2(n4818), .C1(n4817), 
        .C2(n7087), .ZN(n4820) );
  NAND2_X1 U5375 ( .A1(n5999), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4819) );
  OAI21_X1 U5376 ( .B1(n5999), .B2(n4820), .A(n4819), .ZN(U3460) );
  INV_X1 U5377 ( .A(n4821), .ZN(n5007) );
  AOI21_X1 U5378 ( .B1(n7087), .B2(n5007), .A(n5999), .ZN(n6006) );
  NAND2_X1 U5379 ( .A1(n5010), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4826) );
  INV_X1 U5380 ( .A(n4822), .ZN(n7023) );
  NAND2_X1 U5381 ( .A1(n4823), .A2(n7023), .ZN(n5009) );
  INV_X1 U5382 ( .A(n5003), .ZN(n4824) );
  AOI21_X1 U5383 ( .B1(n5009), .B2(n4821), .A(n4824), .ZN(n4825) );
  MUX2_X1 U5384 ( .A(n4826), .B(n4825), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4828) );
  NOR2_X1 U5385 ( .A1(n4821), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4827)
         );
  NAND2_X1 U5386 ( .A1(n5009), .A2(n4827), .ZN(n5004) );
  NAND2_X1 U5387 ( .A1(n4828), .A2(n5004), .ZN(n4829) );
  AOI21_X1 U5388 ( .B1(n4975), .B2(n5971), .A(n4829), .ZN(n5000) );
  INV_X1 U5389 ( .A(n5000), .ZN(n4834) );
  NAND3_X1 U5390 ( .A1(n4821), .A2(n7087), .A3(n3509), .ZN(n4830) );
  OAI21_X1 U5391 ( .B1(n4832), .B2(n4831), .A(n4830), .ZN(n4833) );
  AOI21_X1 U5392 ( .B1(n4834), .B2(n6003), .A(n4833), .ZN(n4835) );
  OAI22_X1 U5393 ( .A1(n6006), .A2(n3509), .B1(n5999), .B2(n4835), .ZN(U3459)
         );
  INV_X1 U5394 ( .A(EAX_REG_18__SCAN_IN), .ZN(n7136) );
  AOI22_X1 U5395 ( .A1(n6631), .A2(UWORD_REG_2__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4836) );
  OAI21_X1 U5396 ( .B1(n7136), .B2(n4844), .A(n4836), .ZN(U2905) );
  INV_X1 U5397 ( .A(EAX_REG_30__SCAN_IN), .ZN(n7191) );
  AOI22_X1 U5398 ( .A1(n6631), .A2(UWORD_REG_14__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4837) );
  OAI21_X1 U5399 ( .B1(n7191), .B2(n4844), .A(n4837), .ZN(U2893) );
  INV_X1 U5400 ( .A(EAX_REG_16__SCAN_IN), .ZN(n7127) );
  AOI22_X1 U5401 ( .A1(n6631), .A2(UWORD_REG_0__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4838) );
  OAI21_X1 U5402 ( .B1(n7127), .B2(n4844), .A(n4838), .ZN(U2907) );
  AOI22_X1 U5403 ( .A1(n6631), .A2(UWORD_REG_1__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4839) );
  OAI21_X1 U5404 ( .B1(n4464), .B2(n4844), .A(n4839), .ZN(U2906) );
  INV_X1 U5405 ( .A(EAX_REG_19__SCAN_IN), .ZN(n7141) );
  AOI22_X1 U5406 ( .A1(n6631), .A2(UWORD_REG_3__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4840) );
  OAI21_X1 U5407 ( .B1(n7141), .B2(n4844), .A(n4840), .ZN(U2904) );
  INV_X1 U5408 ( .A(EAX_REG_27__SCAN_IN), .ZN(n7178) );
  AOI22_X1 U5409 ( .A1(n6631), .A2(UWORD_REG_11__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4841) );
  OAI21_X1 U5410 ( .B1(n7178), .B2(n4844), .A(n4841), .ZN(U2896) );
  INV_X1 U5411 ( .A(EAX_REG_28__SCAN_IN), .ZN(n7183) );
  AOI22_X1 U5412 ( .A1(n6631), .A2(UWORD_REG_12__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4842) );
  OAI21_X1 U5413 ( .B1(n7183), .B2(n4844), .A(n4842), .ZN(U2895) );
  AOI22_X1 U5414 ( .A1(n6631), .A2(UWORD_REG_13__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4843) );
  OAI21_X1 U5415 ( .B1(n4690), .B2(n4844), .A(n4843), .ZN(U2894) );
  OAI21_X1 U5416 ( .B1(n4845), .B2(n4848), .A(n4847), .ZN(n5655) );
  INV_X1 U5417 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4852) );
  AND2_X1 U5418 ( .A1(n4858), .A2(n4849), .ZN(n4851) );
  OR2_X1 U5419 ( .A1(n4851), .A2(n4850), .ZN(n5473) );
  OAI222_X1 U5420 ( .A1(n5655), .A2(n6156), .B1(n4852), .B2(n6706), .C1(n5473), 
        .C2(n6154), .ZN(U2854) );
  AOI21_X1 U5421 ( .B1(n4855), .B2(n4854), .A(n4845), .ZN(n5664) );
  INV_X1 U5422 ( .A(n5664), .ZN(n5234) );
  NAND2_X1 U5423 ( .A1(n4895), .A2(n4856), .ZN(n4857) );
  NAND2_X1 U5424 ( .A1(n4858), .A2(n4857), .ZN(n5223) );
  INV_X1 U5425 ( .A(n5223), .ZN(n4859) );
  AOI22_X1 U5426 ( .A1(n6702), .A2(n4859), .B1(EBX_REG_4__SCAN_IN), .B2(n4769), 
        .ZN(n4860) );
  OAI21_X1 U5427 ( .B1(n5234), .B2(n6156), .A(n4860), .ZN(U2855) );
  NOR2_X1 U5428 ( .A1(n4862), .A2(n4861), .ZN(n4863) );
  NOR2_X1 U5429 ( .A1(n4865), .A2(READY_N), .ZN(n4866) );
  NAND2_X1 U5430 ( .A1(n3747), .A2(n4868), .ZN(n4871) );
  NAND2_X2 U5431 ( .A1(n6015), .A2(n4871), .ZN(n7201) );
  XOR2_X1 U5432 ( .A(n4870), .B(n4869), .Z(n6711) );
  INV_X1 U5433 ( .A(n6711), .ZN(n4902) );
  INV_X1 U5434 ( .A(n4871), .ZN(n4872) );
  INV_X1 U5435 ( .A(DATAI_0_), .ZN(n6560) );
  INV_X1 U5436 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7130) );
  OAI222_X1 U5437 ( .A1(n7201), .A2(n4902), .B1(n5916), .B2(n6560), .C1(n6015), 
        .C2(n7130), .ZN(U2891) );
  INV_X1 U5438 ( .A(DATAI_4_), .ZN(n6448) );
  INV_X1 U5439 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7149) );
  OAI222_X1 U5440 ( .A1(n5234), .A2(n7201), .B1(n5916), .B2(n6448), .C1(n7149), 
        .C2(n6015), .ZN(U2887) );
  INV_X1 U5441 ( .A(DATAI_1_), .ZN(n6558) );
  INV_X1 U5442 ( .A(EAX_REG_1__SCAN_IN), .ZN(n7134) );
  OAI222_X1 U5443 ( .A1(n6714), .A2(n7201), .B1(n5916), .B2(n6558), .C1(n6015), 
        .C2(n7134), .ZN(U2890) );
  INV_X1 U5444 ( .A(n4874), .ZN(n4876) );
  NAND2_X1 U5445 ( .A1(n4876), .A2(n4875), .ZN(n4879) );
  NAND2_X1 U5446 ( .A1(n4878), .A2(n4877), .ZN(n4891) );
  OAI21_X1 U5447 ( .B1(n4873), .B2(n4879), .A(n4891), .ZN(n6722) );
  INV_X1 U5448 ( .A(DATAI_2_), .ZN(n6450) );
  INV_X1 U5449 ( .A(EAX_REG_2__SCAN_IN), .ZN(n7139) );
  OAI222_X1 U5450 ( .A1(n6722), .A2(n7201), .B1(n5916), .B2(n6450), .C1(n6015), 
        .C2(n7139), .ZN(U2889) );
  NAND2_X1 U5451 ( .A1(n4881), .A2(n4880), .ZN(n4882) );
  XNOR2_X1 U5452 ( .A(n4882), .B(n6707), .ZN(n6715) );
  NOR2_X1 U5453 ( .A1(n4884), .A2(n4883), .ZN(n4886) );
  INV_X1 U5454 ( .A(n6818), .ZN(n5138) );
  AOI21_X1 U5455 ( .B1(n6816), .B2(n6870), .A(n5138), .ZN(n6869) );
  INV_X1 U5456 ( .A(n6869), .ZN(n4885) );
  MUX2_X1 U5457 ( .A(n4886), .B(n4885), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4887) );
  INV_X1 U5458 ( .A(n4887), .ZN(n4890) );
  AOI22_X1 U5459 ( .A1(n6873), .A2(n4888), .B1(n6847), .B2(REIP_REG_1__SCAN_IN), .ZN(n4889) );
  OAI211_X1 U5460 ( .C1(n6878), .C2(n6715), .A(n4890), .B(n4889), .ZN(U3017)
         );
  INV_X1 U5461 ( .A(n4891), .ZN(n4893) );
  OAI21_X1 U5462 ( .B1(n4893), .B2(n4892), .A(n4854), .ZN(n5663) );
  INV_X1 U5463 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4897) );
  OAI21_X1 U5464 ( .B1(n4894), .B2(n4896), .A(n4895), .ZN(n5347) );
  OAI222_X1 U5465 ( .A1(n5663), .A2(n6156), .B1(n4897), .B2(n6706), .C1(n5347), 
        .C2(n6154), .ZN(U2856) );
  INV_X1 U5466 ( .A(n4898), .ZN(n4901) );
  INV_X1 U5467 ( .A(n4899), .ZN(n4900) );
  AOI21_X1 U5468 ( .B1(n4901), .B2(n6870), .A(n4900), .ZN(n6874) );
  INV_X1 U5469 ( .A(n6874), .ZN(n4903) );
  OAI222_X1 U5470 ( .A1(n4903), .A2(n6154), .B1(n5458), .B2(n6706), .C1(n6156), 
        .C2(n4902), .ZN(U2859) );
  XNOR2_X1 U5471 ( .A(n4847), .B(n4294), .ZN(n6885) );
  INV_X1 U5472 ( .A(n6885), .ZN(n4909) );
  INV_X1 U5473 ( .A(n4905), .ZN(n5102) );
  OAI21_X1 U5474 ( .B1(n4850), .B2(n4906), .A(n5102), .ZN(n6882) );
  INV_X1 U5475 ( .A(n6882), .ZN(n4907) );
  AOI22_X1 U5476 ( .A1(n6702), .A2(n4907), .B1(EBX_REG_6__SCAN_IN), .B2(n4769), 
        .ZN(n4908) );
  OAI21_X1 U5477 ( .B1(n4909), .B2(n6156), .A(n4908), .ZN(U2853) );
  INV_X1 U5478 ( .A(DATAI_6_), .ZN(n6507) );
  OAI222_X1 U5479 ( .A1(n7201), .A2(n4909), .B1(n5916), .B2(n6507), .C1(n6015), 
        .C2(n4291), .ZN(U2885) );
  NAND3_X1 U5480 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n7054), .A3(n5534), .ZN(n5499) );
  NOR2_X1 U5481 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5499), .ZN(n5378)
         );
  INV_X1 U5482 ( .A(n5378), .ZN(n4912) );
  INV_X1 U5483 ( .A(n4977), .ZN(n4910) );
  INV_X1 U5484 ( .A(n4960), .ZN(n4976) );
  NOR2_X1 U5485 ( .A1(n4910), .A2(n4976), .ZN(n5171) );
  NOR2_X1 U5486 ( .A1(n5171), .A2(n7076), .ZN(n5172) );
  NAND2_X1 U5487 ( .A1(n7076), .A2(n7077), .ZN(n6766) );
  INV_X1 U5488 ( .A(n5364), .ZN(n4911) );
  NAND2_X1 U5489 ( .A1(n4922), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U5490 ( .A1(n4966), .A2(n4959), .ZN(n5771) );
  AOI211_X1 U5491 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4912), .A(n5172), .B(
        n5771), .ZN(n4921) );
  INV_X1 U5492 ( .A(n5764), .ZN(n5687) );
  OR2_X1 U5493 ( .A1(n4975), .A2(n4811), .ZN(n4925) );
  NOR2_X1 U5494 ( .A1(n5538), .A2(n5687), .ZN(n4993) );
  NAND2_X1 U5495 ( .A1(n4267), .A2(n5106), .ZN(n5174) );
  INV_X1 U5496 ( .A(n5502), .ZN(n4916) );
  INV_X1 U5497 ( .A(n5594), .ZN(n4918) );
  INV_X1 U5498 ( .A(n5042), .ZN(n4962) );
  AND2_X1 U5499 ( .A1(n3462), .A2(n4962), .ZN(n4917) );
  AND2_X1 U5500 ( .A1(n3463), .A2(n4917), .ZN(n5304) );
  OAI21_X1 U5501 ( .B1(n4918), .B2(n5433), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4919) );
  OAI21_X1 U5502 ( .B1(n5302), .B2(n4993), .A(n4919), .ZN(n4920) );
  INV_X1 U5503 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4931) );
  INV_X1 U5504 ( .A(n5306), .ZN(n4926) );
  INV_X1 U5505 ( .A(n4922), .ZN(n4923) );
  NAND2_X1 U5506 ( .A1(n4923), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4965) );
  INV_X1 U5507 ( .A(n5171), .ZN(n4924) );
  OAI22_X1 U5508 ( .A1(n4926), .A2(n4925), .B1(n4965), .B2(n4924), .ZN(n5381)
         );
  NAND2_X1 U5509 ( .A1(n6254), .A2(DATAI_18_), .ZN(n5794) );
  NOR2_X1 U5510 ( .A1(n5119), .A2(n3720), .ZN(n5792) );
  NAND2_X1 U5511 ( .A1(n6254), .A2(DATAI_26_), .ZN(n5518) );
  INV_X1 U5512 ( .A(n5518), .ZN(n5796) );
  AOI22_X1 U5513 ( .A1(n5792), .A2(n5378), .B1(n5796), .B2(n5433), .ZN(n4928)
         );
  OAI21_X1 U5514 ( .B1(n5594), .B2(n5794), .A(n4928), .ZN(n4929) );
  AOI21_X1 U5515 ( .B1(n5715), .B2(n5381), .A(n4929), .ZN(n4930) );
  OAI21_X1 U5516 ( .B1(n5384), .B2(n4931), .A(n4930), .ZN(U3086) );
  INV_X1 U5517 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4935) );
  INV_X1 U5518 ( .A(DATAI_7_), .ZN(n6506) );
  NAND2_X1 U5519 ( .A1(n6254), .A2(DATAI_23_), .ZN(n5697) );
  NAND2_X1 U5520 ( .A1(n6254), .A2(DATAI_31_), .ZN(n5778) );
  INV_X1 U5521 ( .A(n5778), .ZN(n5682) );
  AOI22_X1 U5522 ( .A1(n5776), .A2(n5378), .B1(n5682), .B2(n5433), .ZN(n4932)
         );
  OAI21_X1 U5523 ( .B1(n5594), .B2(n5697), .A(n4932), .ZN(n4933) );
  AOI21_X1 U5524 ( .B1(n5694), .B2(n5381), .A(n4933), .ZN(n4934) );
  OAI21_X1 U5525 ( .B1(n5384), .B2(n4935), .A(n4934), .ZN(U3091) );
  INV_X1 U5526 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U5527 ( .A1(n6254), .A2(DATAI_16_), .ZN(n5831) );
  NOR2_X1 U5528 ( .A1(n5119), .A2(n3445), .ZN(n7221) );
  NAND2_X1 U5529 ( .A1(n6254), .A2(DATAI_24_), .ZN(n5555) );
  INV_X1 U5530 ( .A(n5555), .ZN(n7223) );
  AOI22_X1 U5531 ( .A1(n7221), .A2(n5378), .B1(n7223), .B2(n5433), .ZN(n4936)
         );
  OAI21_X1 U5532 ( .B1(n5594), .B2(n5831), .A(n4936), .ZN(n4937) );
  AOI21_X1 U5533 ( .B1(n5581), .B2(n5381), .A(n4937), .ZN(n4938) );
  OAI21_X1 U5534 ( .B1(n5384), .B2(n4939), .A(n4938), .ZN(U3084) );
  INV_X1 U5535 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U5536 ( .A1(n6254), .A2(DATAI_17_), .ZN(n5822) );
  NOR2_X1 U5537 ( .A1(n5119), .A2(n4034), .ZN(n5820) );
  NAND2_X1 U5538 ( .A1(n6254), .A2(DATAI_25_), .ZN(n5505) );
  INV_X1 U5539 ( .A(n5505), .ZN(n5824) );
  AOI22_X1 U5540 ( .A1(n5820), .A2(n5378), .B1(n5824), .B2(n5433), .ZN(n4940)
         );
  OAI21_X1 U5541 ( .B1(n5594), .B2(n5822), .A(n4940), .ZN(n4941) );
  AOI21_X1 U5542 ( .B1(n5720), .B2(n5381), .A(n4941), .ZN(n4942) );
  OAI21_X1 U5543 ( .B1(n5384), .B2(n4943), .A(n4942), .ZN(U3085) );
  INV_X1 U5544 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4948) );
  INV_X1 U5545 ( .A(DATAI_3_), .ZN(n6503) );
  NAND2_X1 U5546 ( .A1(n6254), .A2(DATAI_19_), .ZN(n5801) );
  NAND2_X1 U5547 ( .A1(n6254), .A2(DATAI_27_), .ZN(n5521) );
  INV_X1 U5548 ( .A(n5521), .ZN(n5803) );
  AOI22_X1 U5549 ( .A1(n5799), .A2(n5378), .B1(n5803), .B2(n5433), .ZN(n4945)
         );
  OAI21_X1 U5550 ( .B1(n5594), .B2(n5801), .A(n4945), .ZN(n4946) );
  AOI21_X1 U5551 ( .B1(n5710), .B2(n5381), .A(n4946), .ZN(n4947) );
  OAI21_X1 U5552 ( .B1(n5384), .B2(n4948), .A(n4947), .ZN(U3087) );
  INV_X1 U5553 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7060) );
  NAND2_X1 U5554 ( .A1(n4976), .A2(n7060), .ZN(n4953) );
  INV_X1 U5555 ( .A(n4953), .ZN(n5301) );
  INV_X1 U5556 ( .A(n4965), .ZN(n5768) );
  AOI22_X1 U5557 ( .A1(n5302), .A2(n3490), .B1(n5301), .B2(n5768), .ZN(n5169)
         );
  INV_X1 U5558 ( .A(n4267), .ZN(n4950) );
  NAND3_X1 U5559 ( .A1(n4950), .A2(n5106), .A3(n5173), .ZN(n5536) );
  NOR2_X1 U5560 ( .A1(n3463), .A2(n5173), .ZN(n4949) );
  NAND2_X1 U5561 ( .A1(n4950), .A2(n4949), .ZN(n5397) );
  NAND2_X1 U5562 ( .A1(n5764), .A2(n6581), .ZN(n5765) );
  OAI21_X1 U5563 ( .B1(n5583), .B2(n5441), .A(n5765), .ZN(n4952) );
  INV_X1 U5564 ( .A(n5387), .ZN(n5250) );
  NAND2_X1 U5565 ( .A1(n5250), .A2(n3490), .ZN(n4951) );
  AOI21_X1 U5566 ( .B1(n4952), .B2(n4951), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4955) );
  NOR2_X1 U5567 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U5568 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5535), .ZN(n5402) );
  NOR2_X1 U5569 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5402), .ZN(n5166)
         );
  NAND2_X1 U5570 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4953), .ZN(n5310) );
  INV_X1 U5571 ( .A(n5771), .ZN(n4954) );
  OAI211_X1 U5572 ( .C1(n4955), .C2(n5166), .A(n5310), .B(n4954), .ZN(n5162)
         );
  NAND2_X1 U5573 ( .A1(n5162), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4958) );
  INV_X1 U5574 ( .A(n5583), .ZN(n5164) );
  INV_X1 U5575 ( .A(n5441), .ZN(n5163) );
  OAI22_X1 U5576 ( .A1(n5164), .A2(n5555), .B1(n5163), .B2(n5831), .ZN(n4956)
         );
  AOI21_X1 U5577 ( .B1(n7221), .B2(n5166), .A(n4956), .ZN(n4957) );
  OAI211_X1 U5578 ( .C1(n5169), .C2(n7227), .A(n4958), .B(n4957), .ZN(U3036)
         );
  INV_X1 U5579 ( .A(n4975), .ZN(n5993) );
  INV_X1 U5580 ( .A(n4959), .ZN(n5300) );
  OR2_X1 U5581 ( .A1(n4960), .A2(n7060), .ZN(n4964) );
  INV_X1 U5582 ( .A(n4964), .ZN(n5767) );
  AOI22_X1 U5583 ( .A1(n5389), .A2(n5306), .B1(n5300), .B2(n5767), .ZN(n5135)
         );
  AND2_X1 U5584 ( .A1(n3462), .A2(n5042), .ZN(n4961) );
  AND2_X1 U5585 ( .A1(n3463), .A2(n4961), .ZN(n5280) );
  NAND2_X1 U5586 ( .A1(n5280), .A2(n4915), .ZN(n5358) );
  NOR2_X1 U5587 ( .A1(n3462), .A2(n4962), .ZN(n4963) );
  AOI21_X1 U5588 ( .B1(n5358), .B2(n7217), .A(n6581), .ZN(n4970) );
  NOR2_X1 U5589 ( .A1(n5389), .A2(n5687), .ZN(n5305) );
  NOR2_X1 U5590 ( .A1(n5305), .A2(n5302), .ZN(n4969) );
  NAND3_X1 U5591 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5281) );
  NOR2_X1 U5592 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5281), .ZN(n5132)
         );
  INV_X1 U5593 ( .A(n5132), .ZN(n4967) );
  AND2_X1 U5594 ( .A1(n4964), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U5595 ( .A1(n4966), .A2(n4965), .ZN(n5307) );
  AOI211_X1 U5596 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4967), .A(n5772), .B(
        n5307), .ZN(n4968) );
  OAI21_X1 U5597 ( .B1(n4970), .B2(n4969), .A(n4968), .ZN(n5130) );
  NAND2_X1 U5598 ( .A1(n5130), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4973)
         );
  OAI22_X1 U5599 ( .A1(n5555), .A2(n7217), .B1(n5358), .B2(n5831), .ZN(n4971)
         );
  AOI21_X1 U5600 ( .B1(n7221), .B2(n5132), .A(n4971), .ZN(n4972) );
  OAI211_X1 U5601 ( .C1(n5135), .C2(n7227), .A(n4973), .B(n4972), .ZN(U3132)
         );
  AND2_X1 U5602 ( .A1(n4975), .A2(n4974), .ZN(n5684) );
  NOR2_X1 U5603 ( .A1(n4977), .A2(n4976), .ZN(n4986) );
  AOI22_X1 U5604 ( .A1(n5302), .A2(n5684), .B1(n5300), .B2(n4986), .ZN(n5126)
         );
  NAND3_X1 U5605 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7060), .A3(n5534), .ZN(n5511) );
  NOR2_X1 U5606 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5511), .ZN(n5123)
         );
  INV_X1 U5607 ( .A(n5123), .ZN(n4978) );
  NOR2_X1 U5608 ( .A1(n4986), .A2(n7076), .ZN(n4988) );
  AOI211_X1 U5609 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4978), .A(n4988), .B(
        n5307), .ZN(n4982) );
  NOR2_X1 U5610 ( .A1(n5684), .A2(n5687), .ZN(n5178) );
  NOR2_X1 U5611 ( .A1(n3462), .A2(n5042), .ZN(n4979) );
  OAI21_X1 U5612 ( .B1(n5440), .B2(n5567), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4980) );
  OAI21_X1 U5613 ( .B1(n5306), .B2(n5178), .A(n4980), .ZN(n4981) );
  NAND2_X1 U5614 ( .A1(n4982), .A2(n4981), .ZN(n5118) );
  NAND2_X1 U5615 ( .A1(n5118), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4985) );
  INV_X1 U5616 ( .A(n5440), .ZN(n5121) );
  OAI22_X1 U5617 ( .A1(n5121), .A2(n5555), .B1(n5831), .B2(n5120), .ZN(n4983)
         );
  AOI21_X1 U5618 ( .B1(n7221), .B2(n5123), .A(n4983), .ZN(n4984) );
  OAI211_X1 U5619 ( .C1(n5126), .C2(n7227), .A(n4985), .B(n4984), .ZN(U3052)
         );
  AOI22_X1 U5620 ( .A1(n5302), .A2(n5538), .B1(n5768), .B2(n4986), .ZN(n5155)
         );
  INV_X1 U5621 ( .A(n5535), .ZN(n4987) );
  INV_X1 U5622 ( .A(n5152), .ZN(n4989) );
  AOI211_X1 U5623 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4989), .A(n4988), .B(
        n5771), .ZN(n4995) );
  INV_X1 U5624 ( .A(n5280), .ZN(n4990) );
  INV_X1 U5625 ( .A(n5357), .ZN(n4991) );
  OAI21_X1 U5626 ( .B1(n5584), .B2(n4991), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4992) );
  OAI21_X1 U5627 ( .B1(n4993), .B2(n5306), .A(n4992), .ZN(n4994) );
  NAND2_X1 U5628 ( .A1(n4995), .A2(n4994), .ZN(n5149) );
  NAND2_X1 U5629 ( .A1(n5149), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4998) );
  INV_X1 U5630 ( .A(n5584), .ZN(n5150) );
  OAI22_X1 U5631 ( .A1(n5150), .A2(n5831), .B1(n5555), .B2(n5357), .ZN(n4996)
         );
  AOI21_X1 U5632 ( .B1(n7221), .B2(n5152), .A(n4996), .ZN(n4997) );
  OAI211_X1 U5633 ( .C1(n5155), .C2(n7227), .A(n4998), .B(n4997), .ZN(U3020)
         );
  INV_X1 U5634 ( .A(n7047), .ZN(n4999) );
  AOI211_X1 U5635 ( .C1(n7077), .C2(n4999), .A(FLUSH_REG_SCAN_IN), .B(n7040), 
        .ZN(n5034) );
  INV_X1 U5636 ( .A(n5034), .ZN(n5031) );
  OR2_X1 U5637 ( .A1(n7047), .A2(n5000), .ZN(n5002) );
  NAND2_X1 U5638 ( .A1(n7047), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U5639 ( .A1(n5002), .A2(n5001), .ZN(n7055) );
  AND2_X1 U5640 ( .A1(n7055), .A2(n7077), .ZN(n5029) );
  NAND2_X1 U5641 ( .A1(n5387), .A2(n5971), .ZN(n5016) );
  INV_X1 U5642 ( .A(n5010), .ZN(n5974) );
  OAI211_X1 U5643 ( .C1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(n5974), .A(n5004), .B(n5003), .ZN(n5014) );
  INV_X1 U5644 ( .A(n5005), .ZN(n5006) );
  OAI21_X1 U5645 ( .B1(n5007), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n5006), 
        .ZN(n5008) );
  NAND2_X1 U5646 ( .A1(n5009), .A2(n5008), .ZN(n5012) );
  NAND3_X1 U5647 ( .A1(n5010), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n5005), .ZN(n5011) );
  NAND2_X1 U5648 ( .A1(n5012), .A2(n5011), .ZN(n5013) );
  AOI21_X1 U5649 ( .B1(n5014), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n5013), 
        .ZN(n5015) );
  NAND2_X1 U5650 ( .A1(n5016), .A2(n5015), .ZN(n6002) );
  OR2_X1 U5651 ( .A1(n7047), .A2(n6002), .ZN(n5018) );
  NAND2_X1 U5652 ( .A1(n7047), .A2(n3581), .ZN(n5017) );
  NAND2_X1 U5653 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7034), .ZN(n5027) );
  INV_X1 U5654 ( .A(n5019), .ZN(n5026) );
  INV_X1 U5655 ( .A(n5020), .ZN(n5021) );
  NOR2_X1 U5656 ( .A1(n5022), .A2(n5021), .ZN(n5023) );
  XNOR2_X1 U5657 ( .A(n5023), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5215)
         );
  NAND2_X1 U5658 ( .A1(n5024), .A2(n7077), .ZN(n5025) );
  OAI21_X1 U5659 ( .B1(n5027), .B2(n5026), .A(n7036), .ZN(n5028) );
  AOI21_X1 U5660 ( .B1(n5029), .B2(n7059), .A(n5028), .ZN(n5030) );
  NAND2_X1 U5661 ( .A1(n5031), .A2(n5030), .ZN(n7063) );
  INV_X1 U5662 ( .A(n5032), .ZN(n5033) );
  OR2_X1 U5663 ( .A1(n5034), .A2(n5033), .ZN(n5035) );
  NAND2_X1 U5664 ( .A1(n7063), .A2(n5035), .ZN(n5365) );
  NAND2_X1 U5665 ( .A1(n5365), .A2(n7034), .ZN(n5037) );
  INV_X1 U5666 ( .A(n7083), .ZN(n5036) );
  NAND2_X1 U5667 ( .A1(n5037), .A2(n5036), .ZN(n5038) );
  INV_X1 U5668 ( .A(n6399), .ZN(n5108) );
  NAND2_X1 U5669 ( .A1(n5108), .A2(n5764), .ZN(n5369) );
  NAND2_X1 U5670 ( .A1(n3462), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5105) );
  OAI21_X1 U5671 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3462), .A(n5105), .ZN(
        n5040) );
  AOI21_X1 U5672 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n7084), .A(n6399), .ZN(
        n5041) );
  AOI22_X1 U5673 ( .A1(n6399), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n4811), .B2(n5041), .ZN(n5039) );
  OAI21_X1 U5674 ( .B1(n5369), .B2(n5040), .A(n5039), .ZN(U3464) );
  INV_X1 U5675 ( .A(n5041), .ZN(n5366) );
  AND2_X1 U5676 ( .A1(n5176), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5683) );
  INV_X1 U5677 ( .A(n5683), .ZN(n5045) );
  NOR2_X1 U5678 ( .A1(n5105), .A2(n5042), .ZN(n5043) );
  AND2_X1 U5679 ( .A1(n3463), .A2(n5043), .ZN(n5385) );
  AOI21_X1 U5680 ( .B1(n4267), .B2(n6581), .A(n5385), .ZN(n5044) );
  AND3_X1 U5681 ( .A1(n5045), .A2(n5044), .A3(n5174), .ZN(n5046) );
  OAI222_X1 U5682 ( .A1(n5366), .A2(n5250), .B1(n5108), .B2(n7060), .C1(n5369), 
        .C2(n5046), .ZN(U3462) );
  NAND2_X1 U5683 ( .A1(n5149), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5049) );
  OAI22_X1 U5684 ( .A1(n5150), .A2(n5801), .B1(n5521), .B2(n5357), .ZN(n5047)
         );
  AOI21_X1 U5685 ( .B1(n5799), .B2(n5152), .A(n5047), .ZN(n5048) );
  OAI211_X1 U5686 ( .C1(n5155), .C2(n5805), .A(n5049), .B(n5048), .ZN(U3023)
         );
  NAND2_X1 U5687 ( .A1(n5118), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5052) );
  OAI22_X1 U5688 ( .A1(n5121), .A2(n5778), .B1(n5697), .B2(n5120), .ZN(n5050)
         );
  AOI21_X1 U5689 ( .B1(n5776), .B2(n5123), .A(n5050), .ZN(n5051) );
  OAI211_X1 U5690 ( .C1(n5126), .C2(n5784), .A(n5052), .B(n5051), .ZN(U3059)
         );
  NAND2_X1 U5691 ( .A1(n5130), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5055)
         );
  OAI22_X1 U5692 ( .A1(n5778), .A2(n7217), .B1(n5358), .B2(n5697), .ZN(n5053)
         );
  AOI21_X1 U5693 ( .B1(n5776), .B2(n5132), .A(n5053), .ZN(n5054) );
  OAI211_X1 U5694 ( .C1(n5135), .C2(n5784), .A(n5055), .B(n5054), .ZN(U3139)
         );
  NAND2_X1 U5695 ( .A1(n5149), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5058) );
  OAI22_X1 U5696 ( .A1(n5150), .A2(n5697), .B1(n5778), .B2(n5357), .ZN(n5056)
         );
  AOI21_X1 U5697 ( .B1(n5776), .B2(n5152), .A(n5056), .ZN(n5057) );
  OAI211_X1 U5698 ( .C1(n5155), .C2(n5784), .A(n5058), .B(n5057), .ZN(U3027)
         );
  NAND2_X1 U5699 ( .A1(n5130), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5061)
         );
  OAI22_X1 U5700 ( .A1(n5521), .A2(n7217), .B1(n5358), .B2(n5801), .ZN(n5059)
         );
  AOI21_X1 U5701 ( .B1(n5799), .B2(n5132), .A(n5059), .ZN(n5060) );
  OAI211_X1 U5702 ( .C1(n5135), .C2(n5805), .A(n5061), .B(n5060), .ZN(U3135)
         );
  NAND2_X1 U5703 ( .A1(n5118), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5064) );
  OAI22_X1 U5704 ( .A1(n5121), .A2(n5505), .B1(n5822), .B2(n5120), .ZN(n5062)
         );
  AOI21_X1 U5705 ( .B1(n5820), .B2(n5123), .A(n5062), .ZN(n5063) );
  OAI211_X1 U5706 ( .C1(n5126), .C2(n5826), .A(n5064), .B(n5063), .ZN(U3053)
         );
  NAND2_X1 U5707 ( .A1(n5162), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5067) );
  OAI22_X1 U5708 ( .A1(n5164), .A2(n5778), .B1(n5163), .B2(n5697), .ZN(n5065)
         );
  AOI21_X1 U5709 ( .B1(n5776), .B2(n5166), .A(n5065), .ZN(n5066) );
  OAI211_X1 U5710 ( .C1(n5169), .C2(n5784), .A(n5067), .B(n5066), .ZN(U3043)
         );
  NAND2_X1 U5711 ( .A1(n5162), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5070) );
  OAI22_X1 U5712 ( .A1(n5164), .A2(n5521), .B1(n5163), .B2(n5801), .ZN(n5068)
         );
  AOI21_X1 U5713 ( .B1(n5799), .B2(n5166), .A(n5068), .ZN(n5069) );
  OAI211_X1 U5714 ( .C1(n5169), .C2(n5805), .A(n5070), .B(n5069), .ZN(U3039)
         );
  NAND2_X1 U5715 ( .A1(n5149), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5073) );
  OAI22_X1 U5716 ( .A1(n5150), .A2(n5794), .B1(n5518), .B2(n5357), .ZN(n5071)
         );
  AOI21_X1 U5717 ( .B1(n5792), .B2(n5152), .A(n5071), .ZN(n5072) );
  OAI211_X1 U5718 ( .C1(n5155), .C2(n5798), .A(n5073), .B(n5072), .ZN(U3022)
         );
  NAND2_X1 U5719 ( .A1(n5162), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5076) );
  OAI22_X1 U5720 ( .A1(n5164), .A2(n5505), .B1(n5163), .B2(n5822), .ZN(n5074)
         );
  AOI21_X1 U5721 ( .B1(n5820), .B2(n5166), .A(n5074), .ZN(n5075) );
  OAI211_X1 U5722 ( .C1(n5169), .C2(n5826), .A(n5076), .B(n5075), .ZN(U3037)
         );
  NAND2_X1 U5723 ( .A1(n5118), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5079) );
  OAI22_X1 U5724 ( .A1(n5121), .A2(n5518), .B1(n5794), .B2(n5120), .ZN(n5077)
         );
  AOI21_X1 U5725 ( .B1(n5792), .B2(n5123), .A(n5077), .ZN(n5078) );
  OAI211_X1 U5726 ( .C1(n5126), .C2(n5798), .A(n5079), .B(n5078), .ZN(U3054)
         );
  NAND2_X1 U5727 ( .A1(n5130), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5082)
         );
  OAI22_X1 U5728 ( .A1(n5518), .A2(n7217), .B1(n5358), .B2(n5794), .ZN(n5080)
         );
  AOI21_X1 U5729 ( .B1(n5792), .B2(n5132), .A(n5080), .ZN(n5081) );
  OAI211_X1 U5730 ( .C1(n5135), .C2(n5798), .A(n5082), .B(n5081), .ZN(U3134)
         );
  NAND2_X1 U5731 ( .A1(n5130), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5085)
         );
  OAI22_X1 U5732 ( .A1(n5505), .A2(n7217), .B1(n5358), .B2(n5822), .ZN(n5083)
         );
  AOI21_X1 U5733 ( .B1(n5820), .B2(n5132), .A(n5083), .ZN(n5084) );
  OAI211_X1 U5734 ( .C1(n5135), .C2(n5826), .A(n5085), .B(n5084), .ZN(U3133)
         );
  NAND2_X1 U5735 ( .A1(n5149), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5088) );
  OAI22_X1 U5736 ( .A1(n5150), .A2(n5822), .B1(n5505), .B2(n5357), .ZN(n5086)
         );
  AOI21_X1 U5737 ( .B1(n5820), .B2(n5152), .A(n5086), .ZN(n5087) );
  OAI211_X1 U5738 ( .C1(n5155), .C2(n5826), .A(n5088), .B(n5087), .ZN(U3021)
         );
  NAND2_X1 U5739 ( .A1(n5162), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5091) );
  OAI22_X1 U5740 ( .A1(n5164), .A2(n5518), .B1(n5163), .B2(n5794), .ZN(n5089)
         );
  AOI21_X1 U5741 ( .B1(n5792), .B2(n5166), .A(n5089), .ZN(n5090) );
  OAI211_X1 U5742 ( .C1(n5169), .C2(n5798), .A(n5091), .B(n5090), .ZN(U3038)
         );
  NAND2_X1 U5743 ( .A1(n5118), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5094) );
  OAI22_X1 U5744 ( .A1(n5121), .A2(n5521), .B1(n5801), .B2(n5120), .ZN(n5092)
         );
  AOI21_X1 U5745 ( .B1(n5799), .B2(n5123), .A(n5092), .ZN(n5093) );
  OAI211_X1 U5746 ( .C1(n5126), .C2(n5805), .A(n5094), .B(n5093), .ZN(U3055)
         );
  AOI21_X1 U5747 ( .B1(n5095), .B2(n5098), .A(n5097), .ZN(n6896) );
  INV_X1 U5748 ( .A(n6896), .ZN(n5170) );
  INV_X1 U5749 ( .A(n5099), .ZN(n5103) );
  INV_X1 U5750 ( .A(n5100), .ZN(n5101) );
  AOI21_X1 U5751 ( .B1(n5103), .B2(n5102), .A(n5101), .ZN(n6890) );
  AOI22_X1 U5752 ( .A1(n6702), .A2(n6890), .B1(EBX_REG_7__SCAN_IN), .B2(n4769), 
        .ZN(n5104) );
  OAI21_X1 U5753 ( .B1(n5170), .B2(n6156), .A(n5104), .ZN(U2852) );
  XNOR2_X1 U5754 ( .A(n5106), .B(n5105), .ZN(n5107) );
  OAI222_X1 U5755 ( .A1(n5108), .A2(n7054), .B1(n5366), .B2(n5993), .C1(n5369), 
        .C2(n5107), .ZN(U3463) );
  NAND2_X1 U5756 ( .A1(n5130), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5111)
         );
  NOR2_X1 U5757 ( .A1(n5119), .A2(n3746), .ZN(n5785) );
  NAND2_X1 U5758 ( .A1(n6254), .A2(DATAI_30_), .ZN(n5617) );
  NAND2_X1 U5759 ( .A1(n6254), .A2(DATAI_22_), .ZN(n5787) );
  OAI22_X1 U5760 ( .A1(n5617), .A2(n7217), .B1(n5358), .B2(n5787), .ZN(n5109)
         );
  AOI21_X1 U5761 ( .B1(n5785), .B2(n5132), .A(n5109), .ZN(n5110) );
  OAI211_X1 U5762 ( .C1(n5135), .C2(n5791), .A(n5111), .B(n5110), .ZN(U3138)
         );
  NAND2_X1 U5763 ( .A1(n5118), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5114) );
  OAI22_X1 U5764 ( .A1(n5121), .A2(n5617), .B1(n5787), .B2(n5120), .ZN(n5112)
         );
  AOI21_X1 U5765 ( .B1(n5785), .B2(n5123), .A(n5112), .ZN(n5113) );
  OAI211_X1 U5766 ( .C1(n5126), .C2(n5791), .A(n5114), .B(n5113), .ZN(U3058)
         );
  NAND2_X1 U5767 ( .A1(n5118), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U5768 ( .A1(n6254), .A2(DATAI_28_), .ZN(n5628) );
  NAND2_X1 U5769 ( .A1(n6254), .A2(DATAI_20_), .ZN(n5808) );
  OAI22_X1 U5770 ( .A1(n5121), .A2(n5628), .B1(n5808), .B2(n5120), .ZN(n5115)
         );
  AOI21_X1 U5771 ( .B1(n5806), .B2(n5123), .A(n5115), .ZN(n5116) );
  OAI211_X1 U5772 ( .C1(n5126), .C2(n5812), .A(n5117), .B(n5116), .ZN(U3056)
         );
  INV_X1 U5773 ( .A(DATAI_5_), .ZN(n6504) );
  NAND2_X1 U5774 ( .A1(n5118), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5125) );
  NOR2_X1 U5775 ( .A1(n5119), .A2(n3724), .ZN(n5813) );
  NAND2_X1 U5776 ( .A1(n6254), .A2(DATAI_29_), .ZN(n5622) );
  NAND2_X1 U5777 ( .A1(n6254), .A2(DATAI_21_), .ZN(n5815) );
  OAI22_X1 U5778 ( .A1(n5121), .A2(n5622), .B1(n5815), .B2(n5120), .ZN(n5122)
         );
  AOI21_X1 U5779 ( .B1(n5813), .B2(n5123), .A(n5122), .ZN(n5124) );
  OAI211_X1 U5780 ( .C1(n5126), .C2(n5819), .A(n5125), .B(n5124), .ZN(U3057)
         );
  NAND2_X1 U5781 ( .A1(n5130), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5129)
         );
  OAI22_X1 U5782 ( .A1(n5628), .A2(n7217), .B1(n5358), .B2(n5808), .ZN(n5127)
         );
  AOI21_X1 U5783 ( .B1(n5806), .B2(n5132), .A(n5127), .ZN(n5128) );
  OAI211_X1 U5784 ( .C1(n5135), .C2(n5812), .A(n5129), .B(n5128), .ZN(U3136)
         );
  NAND2_X1 U5785 ( .A1(n5130), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5134)
         );
  OAI22_X1 U5786 ( .A1(n5622), .A2(n7217), .B1(n5358), .B2(n5815), .ZN(n5131)
         );
  AOI21_X1 U5787 ( .B1(n5813), .B2(n5132), .A(n5131), .ZN(n5133) );
  OAI211_X1 U5788 ( .C1(n5135), .C2(n5819), .A(n5134), .B(n5133), .ZN(U3137)
         );
  XNOR2_X1 U5789 ( .A(n5136), .B(n5137), .ZN(n5671) );
  INV_X1 U5790 ( .A(n5857), .ZN(n6814) );
  NAND2_X1 U5791 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6779) );
  AOI21_X1 U5792 ( .B1(n6814), .B2(n6779), .A(n5138), .ZN(n6787) );
  OAI21_X1 U5793 ( .B1(n5878), .B2(n6778), .A(n6787), .ZN(n6791) );
  INV_X1 U5794 ( .A(n6847), .ZN(n6860) );
  INV_X1 U5795 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6639) );
  NOR2_X1 U5796 ( .A1(n6860), .A2(n6639), .ZN(n5667) );
  NOR2_X1 U5797 ( .A1(n6794), .A2(n5223), .ZN(n5139) );
  AOI211_X1 U5798 ( .C1(n6791), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5667), 
        .B(n5139), .ZN(n5142) );
  INV_X1 U5799 ( .A(n6778), .ZN(n5468) );
  NAND2_X1 U5800 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6378), .ZN(n6788)
         );
  OAI22_X1 U5801 ( .A1(n5468), .A2(n5878), .B1(n3872), .B2(n6788), .ZN(n6808)
         );
  NAND2_X1 U5802 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5140) );
  OAI211_X1 U5803 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6808), .B(n5140), .ZN(n5141) );
  OAI211_X1 U5804 ( .C1(n5671), .C2(n6878), .A(n5142), .B(n5141), .ZN(U3014)
         );
  NAND2_X1 U5805 ( .A1(n5149), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5145) );
  OAI22_X1 U5806 ( .A1(n5150), .A2(n5808), .B1(n5628), .B2(n5357), .ZN(n5143)
         );
  AOI21_X1 U5807 ( .B1(n5806), .B2(n5152), .A(n5143), .ZN(n5144) );
  OAI211_X1 U5808 ( .C1(n5155), .C2(n5812), .A(n5145), .B(n5144), .ZN(U3024)
         );
  NAND2_X1 U5809 ( .A1(n5149), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5148) );
  OAI22_X1 U5810 ( .A1(n5150), .A2(n5787), .B1(n5617), .B2(n5357), .ZN(n5146)
         );
  AOI21_X1 U5811 ( .B1(n5785), .B2(n5152), .A(n5146), .ZN(n5147) );
  OAI211_X1 U5812 ( .C1(n5155), .C2(n5791), .A(n5148), .B(n5147), .ZN(U3026)
         );
  NAND2_X1 U5813 ( .A1(n5149), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5154) );
  OAI22_X1 U5814 ( .A1(n5150), .A2(n5815), .B1(n5622), .B2(n5357), .ZN(n5151)
         );
  AOI21_X1 U5815 ( .B1(n5813), .B2(n5152), .A(n5151), .ZN(n5153) );
  OAI211_X1 U5816 ( .C1(n5155), .C2(n5819), .A(n5154), .B(n5153), .ZN(U3025)
         );
  NAND2_X1 U5817 ( .A1(n5162), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5158) );
  OAI22_X1 U5818 ( .A1(n5164), .A2(n5628), .B1(n5163), .B2(n5808), .ZN(n5156)
         );
  AOI21_X1 U5819 ( .B1(n5806), .B2(n5166), .A(n5156), .ZN(n5157) );
  OAI211_X1 U5820 ( .C1(n5169), .C2(n5812), .A(n5158), .B(n5157), .ZN(U3040)
         );
  NAND2_X1 U5821 ( .A1(n5162), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5161) );
  OAI22_X1 U5822 ( .A1(n5164), .A2(n5617), .B1(n5163), .B2(n5787), .ZN(n5159)
         );
  AOI21_X1 U5823 ( .B1(n5785), .B2(n5166), .A(n5159), .ZN(n5160) );
  OAI211_X1 U5824 ( .C1(n5169), .C2(n5791), .A(n5161), .B(n5160), .ZN(U3042)
         );
  NAND2_X1 U5825 ( .A1(n5162), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5168) );
  OAI22_X1 U5826 ( .A1(n5164), .A2(n5622), .B1(n5163), .B2(n5815), .ZN(n5165)
         );
  AOI21_X1 U5827 ( .B1(n5813), .B2(n5166), .A(n5165), .ZN(n5167) );
  OAI211_X1 U5828 ( .C1(n5169), .C2(n5819), .A(n5168), .B(n5167), .ZN(U3041)
         );
  INV_X1 U5829 ( .A(EAX_REG_5__SCAN_IN), .ZN(n7154) );
  OAI222_X1 U5830 ( .A1(n5655), .A2(n7201), .B1(n5916), .B2(n6504), .C1(n6015), 
        .C2(n7154), .ZN(U2886) );
  INV_X1 U5831 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7144) );
  OAI222_X1 U5832 ( .A1(n5663), .A2(n7201), .B1(n5916), .B2(n6503), .C1(n6015), 
        .C2(n7144), .ZN(U2888) );
  OAI222_X1 U5833 ( .A1(n5170), .A2(n7201), .B1(n5916), .B2(n6506), .C1(n6015), 
        .C2(n4298), .ZN(U2884) );
  AOI22_X1 U5834 ( .A1(n5306), .A2(n5684), .B1(n5300), .B2(n5171), .ZN(n5648)
         );
  NOR3_X1 U5835 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7054), .A3(n7060), 
        .ZN(n5693) );
  INV_X1 U5836 ( .A(n5693), .ZN(n5686) );
  OR2_X1 U5837 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5686), .ZN(n5643)
         );
  AOI211_X1 U5838 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5643), .A(n5172), .B(
        n5307), .ZN(n5180) );
  INV_X1 U5839 ( .A(n5261), .ZN(n5175) );
  NOR2_X2 U5840 ( .A1(n5175), .A2(n4915), .ZN(n5645) );
  OAI21_X1 U5841 ( .B1(n5645), .B2(n7222), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5177) );
  OAI21_X1 U5842 ( .B1(n5302), .B2(n5178), .A(n5177), .ZN(n5179) );
  NAND2_X1 U5843 ( .A1(n5180), .A2(n5179), .ZN(n5641) );
  NAND2_X1 U5844 ( .A1(n5641), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5183)
         );
  OAI22_X1 U5845 ( .A1(n5560), .A2(n5643), .B1(n5697), .B2(n5642), .ZN(n5181)
         );
  AOI21_X1 U5846 ( .B1(n5682), .B2(n5645), .A(n5181), .ZN(n5182) );
  OAI211_X1 U5847 ( .C1(n5648), .C2(n5784), .A(n5183), .B(n5182), .ZN(U3123)
         );
  NAND2_X1 U5848 ( .A1(n5641), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5186)
         );
  OAI22_X1 U5849 ( .A1(n5714), .A2(n5643), .B1(n5801), .B2(n5642), .ZN(n5184)
         );
  AOI21_X1 U5850 ( .B1(n5803), .B2(n5645), .A(n5184), .ZN(n5185) );
  OAI211_X1 U5851 ( .C1(n5648), .C2(n5805), .A(n5186), .B(n5185), .ZN(U3119)
         );
  NAND2_X1 U5852 ( .A1(n5641), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5189)
         );
  INV_X1 U5853 ( .A(n5820), .ZN(n5724) );
  OAI22_X1 U5854 ( .A1(n5724), .A2(n5643), .B1(n5822), .B2(n5642), .ZN(n5187)
         );
  AOI21_X1 U5855 ( .B1(n5824), .B2(n5645), .A(n5187), .ZN(n5188) );
  OAI211_X1 U5856 ( .C1(n5648), .C2(n5826), .A(n5189), .B(n5188), .ZN(U3117)
         );
  NAND2_X1 U5857 ( .A1(n5641), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5192)
         );
  INV_X1 U5858 ( .A(n7221), .ZN(n5588) );
  OAI22_X1 U5859 ( .A1(n5588), .A2(n5643), .B1(n5831), .B2(n5642), .ZN(n5190)
         );
  AOI21_X1 U5860 ( .B1(n7223), .B2(n5645), .A(n5190), .ZN(n5191) );
  OAI211_X1 U5861 ( .C1(n5648), .C2(n7227), .A(n5192), .B(n5191), .ZN(U3116)
         );
  NAND2_X1 U5862 ( .A1(n5641), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5195)
         );
  INV_X1 U5863 ( .A(n5792), .ZN(n5719) );
  OAI22_X1 U5864 ( .A1(n5719), .A2(n5643), .B1(n5794), .B2(n5642), .ZN(n5193)
         );
  AOI21_X1 U5865 ( .B1(n5796), .B2(n5645), .A(n5193), .ZN(n5194) );
  OAI211_X1 U5866 ( .C1(n5648), .C2(n5798), .A(n5195), .B(n5194), .ZN(U3118)
         );
  NOR2_X1 U5867 ( .A1(n5097), .A2(n5196), .ZN(n5197) );
  OR2_X1 U5868 ( .A1(n3485), .A2(n5197), .ZN(n5486) );
  NAND2_X1 U5869 ( .A1(n5100), .A2(n5198), .ZN(n5199) );
  NAND2_X1 U5870 ( .A1(n5447), .A2(n5199), .ZN(n6795) );
  INV_X1 U5871 ( .A(n6795), .ZN(n5200) );
  AOI22_X1 U5872 ( .A1(n6702), .A2(n5200), .B1(EBX_REG_8__SCAN_IN), .B2(n4769), 
        .ZN(n5201) );
  OAI21_X1 U5873 ( .B1(n5486), .B2(n6156), .A(n5201), .ZN(U2851) );
  NOR3_X1 U5874 ( .A1(n7096), .A2(n7084), .A3(n6766), .ZN(n7090) );
  NAND2_X1 U5875 ( .A1(n5203), .A2(n5202), .ZN(n7080) );
  INV_X1 U5876 ( .A(n7080), .ZN(n5204) );
  OR2_X1 U5877 ( .A1(n6847), .A2(n5204), .ZN(n5205) );
  OR2_X1 U5878 ( .A1(n7090), .A2(n5205), .ZN(n5206) );
  NOR2_X1 U5879 ( .A1(n5227), .A2(n7077), .ZN(n5207) );
  NAND2_X1 U5880 ( .A1(n6007), .A2(n4035), .ZN(n5208) );
  NAND2_X1 U5881 ( .A1(n7124), .A2(n6581), .ZN(n5219) );
  INV_X1 U5882 ( .A(n5219), .ZN(n5209) );
  AND3_X1 U5883 ( .A1(n5210), .A2(n5209), .A3(n4097), .ZN(n5211) );
  INV_X1 U5884 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6690) );
  INV_X1 U5885 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6780) );
  OR2_X1 U5886 ( .A1(n6690), .A2(n6780), .ZN(n5989) );
  INV_X1 U5887 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U5888 ( .A1(n5989), .A2(n6637), .ZN(n5235) );
  OAI21_X1 U5889 ( .B1(n7010), .B2(n5235), .A(n6107), .ZN(n5253) );
  NAND3_X1 U5890 ( .A1(n6994), .A2(n5235), .A3(n6639), .ZN(n5231) );
  INV_X1 U5891 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5665) );
  INV_X1 U5892 ( .A(n5213), .ZN(n5214) );
  NAND2_X1 U5893 ( .A1(n6007), .A2(n5214), .ZN(n5992) );
  OAI22_X1 U5894 ( .A1(n5665), .A2(n6980), .B1(n5215), .B2(n5992), .ZN(n5226)
         );
  OR2_X1 U5895 ( .A1(n6771), .A2(n5219), .ZN(n7068) );
  NAND2_X1 U5896 ( .A1(n3821), .A2(n7068), .ZN(n5217) );
  INV_X1 U5897 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6127) );
  NAND3_X1 U5898 ( .A1(n4097), .A2(n6127), .A3(n5219), .ZN(n5216) );
  NAND2_X1 U5899 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  NAND2_X1 U5900 ( .A1(n5219), .A2(EBX_REG_31__SCAN_IN), .ZN(n5220) );
  NOR2_X1 U5901 ( .A1(n5221), .A2(n5220), .ZN(n5222) );
  OAI22_X1 U5902 ( .A1(n5224), .A2(n6998), .B1(n7006), .B2(n5223), .ZN(n5225)
         );
  NOR3_X1 U5903 ( .A1(n6974), .A2(n5226), .A3(n5225), .ZN(n5230) );
  AND2_X1 U5904 ( .A1(n5227), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U5905 ( .A1(n7017), .A2(n5668), .ZN(n5229) );
  NAND3_X1 U5906 ( .A1(n5231), .A2(n5230), .A3(n5229), .ZN(n5232) );
  AOI21_X1 U5907 ( .B1(n5253), .B2(REIP_REG_4__SCAN_IN), .A(n5232), .ZN(n5233)
         );
  OAI21_X1 U5908 ( .B1(n5234), .B2(n6120), .A(n5233), .ZN(U2823) );
  INV_X1 U5909 ( .A(n5488), .ZN(n5239) );
  NAND2_X1 U5910 ( .A1(n5235), .A2(REIP_REG_4__SCAN_IN), .ZN(n5478) );
  INV_X1 U5911 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6641) );
  NOR2_X1 U5912 ( .A1(n5478), .A2(n6641), .ZN(n5472) );
  NAND2_X1 U5913 ( .A1(n5472), .A2(REIP_REG_6__SCAN_IN), .ZN(n6889) );
  INV_X1 U5914 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6643) );
  NOR2_X1 U5915 ( .A1(n6889), .A2(n6643), .ZN(n5236) );
  INV_X1 U5916 ( .A(n5236), .ZN(n5237) );
  NAND2_X1 U5917 ( .A1(n5236), .A2(REIP_REG_8__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U5918 ( .A1(n6994), .A2(n5751), .ZN(n5240) );
  OAI22_X1 U5919 ( .A1(n7006), .A2(n6795), .B1(n5237), .B2(n5240), .ZN(n5238)
         );
  AOI21_X1 U5920 ( .B1(n7017), .B2(n5239), .A(n5238), .ZN(n5245) );
  NAND2_X1 U5921 ( .A1(n6107), .A2(n5240), .ZN(n5597) );
  OAI22_X1 U5922 ( .A1(n5242), .A2(n6980), .B1(n5241), .B2(n6998), .ZN(n5243)
         );
  AOI211_X1 U5923 ( .C1(REIP_REG_8__SCAN_IN), .C2(n5597), .A(n6974), .B(n5243), 
        .ZN(n5244) );
  OAI211_X1 U5924 ( .C1(n7001), .C2(n5486), .A(n5245), .B(n5244), .ZN(U2819)
         );
  INV_X1 U5925 ( .A(n6107), .ZN(n6116) );
  OAI21_X1 U5926 ( .B1(n6116), .B2(n5989), .A(n6637), .ZN(n5252) );
  INV_X1 U5927 ( .A(n5347), .ZN(n5246) );
  AOI22_X1 U5928 ( .A1(n7015), .A2(n5246), .B1(n7008), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5249) );
  INV_X1 U5929 ( .A(n5247), .ZN(n5660) );
  AOI22_X1 U5930 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n7009), .B1(n7017), 
        .B2(n5660), .ZN(n5248) );
  OAI211_X1 U5931 ( .C1(n5250), .C2(n5992), .A(n5249), .B(n5248), .ZN(n5251)
         );
  AOI21_X1 U5932 ( .B1(n5253), .B2(n5252), .A(n5251), .ZN(n5254) );
  OAI21_X1 U5933 ( .B1(n6120), .B2(n5663), .A(n5254), .ZN(U2824) );
  OAI21_X1 U5934 ( .B1(n5261), .B2(n5687), .A(n5765), .ZN(n5259) );
  NAND2_X1 U5935 ( .A1(n3490), .A2(n5387), .ZN(n5774) );
  INV_X1 U5936 ( .A(n5972), .ZN(n5386) );
  NAND3_X1 U5937 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7054), .ZN(n5770) );
  OR2_X1 U5938 ( .A1(n7043), .A2(n5770), .ZN(n5629) );
  OAI21_X1 U5939 ( .B1(n5774), .B2(n5386), .A(n5629), .ZN(n5257) );
  INV_X1 U5940 ( .A(n5770), .ZN(n5255) );
  AOI22_X1 U5941 ( .A1(n5259), .A2(n5257), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5255), .ZN(n5634) );
  INV_X1 U5942 ( .A(n5257), .ZN(n5258) );
  AOI22_X1 U5943 ( .A1(n5259), .A2(n5258), .B1(n5770), .B2(n5687), .ZN(n5260)
         );
  NAND2_X1 U5944 ( .A1(n5689), .A2(n5260), .ZN(n5627) );
  NAND2_X1 U5945 ( .A1(n5627), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5264)
         );
  INV_X1 U5946 ( .A(n5697), .ZN(n5782) );
  OAI22_X1 U5947 ( .A1(n5560), .A2(n5629), .B1(n5778), .B2(n5830), .ZN(n5262)
         );
  AOI21_X1 U5948 ( .B1(n5782), .B2(n5645), .A(n5262), .ZN(n5263) );
  OAI211_X1 U5949 ( .C1(n5634), .C2(n5784), .A(n5264), .B(n5263), .ZN(U3115)
         );
  NAND2_X1 U5950 ( .A1(n5627), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n5267)
         );
  INV_X1 U5951 ( .A(n5831), .ZN(n7219) );
  OAI22_X1 U5952 ( .A1(n5588), .A2(n5629), .B1(n5555), .B2(n5830), .ZN(n5265)
         );
  AOI21_X1 U5953 ( .B1(n7219), .B2(n5645), .A(n5265), .ZN(n5266) );
  OAI211_X1 U5954 ( .C1(n5634), .C2(n7227), .A(n5267), .B(n5266), .ZN(U3108)
         );
  INV_X1 U5955 ( .A(DATAI_8_), .ZN(n6552) );
  INV_X1 U5956 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7166) );
  OAI222_X1 U5957 ( .A1(n5486), .A2(n7201), .B1(n5916), .B2(n6552), .C1(n6015), 
        .C2(n7166), .ZN(U2883) );
  NAND2_X1 U5958 ( .A1(n5627), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5270)
         );
  INV_X1 U5959 ( .A(n5801), .ZN(n5550) );
  OAI22_X1 U5960 ( .A1(n5714), .A2(n5629), .B1(n5521), .B2(n5830), .ZN(n5268)
         );
  AOI21_X1 U5961 ( .B1(n5550), .B2(n5645), .A(n5268), .ZN(n5269) );
  OAI211_X1 U5962 ( .C1(n5634), .C2(n5805), .A(n5270), .B(n5269), .ZN(U3111)
         );
  NAND2_X1 U5963 ( .A1(n5627), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5273)
         );
  INV_X1 U5964 ( .A(n5794), .ZN(n5575) );
  OAI22_X1 U5965 ( .A1(n5719), .A2(n5629), .B1(n5518), .B2(n5830), .ZN(n5271)
         );
  AOI21_X1 U5966 ( .B1(n5575), .B2(n5645), .A(n5271), .ZN(n5272) );
  OAI211_X1 U5967 ( .C1(n5634), .C2(n5798), .A(n5273), .B(n5272), .ZN(U3110)
         );
  NAND2_X1 U5968 ( .A1(n5627), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n5276)
         );
  INV_X1 U5969 ( .A(n5822), .ZN(n5568) );
  OAI22_X1 U5970 ( .A1(n5724), .A2(n5629), .B1(n5505), .B2(n5830), .ZN(n5274)
         );
  AOI21_X1 U5971 ( .B1(n5568), .B2(n5645), .A(n5274), .ZN(n5275) );
  OAI211_X1 U5972 ( .C1(n5634), .C2(n5826), .A(n5276), .B(n5275), .ZN(U3109)
         );
  AND2_X1 U5973 ( .A1(n5387), .A2(n5972), .ZN(n5685) );
  NOR2_X1 U5974 ( .A1(n5277), .A2(n7060), .ZN(n5360) );
  AOI21_X1 U5975 ( .B1(n5389), .B2(n5685), .A(n5360), .ZN(n5283) );
  INV_X1 U5976 ( .A(n5283), .ZN(n5279) );
  INV_X1 U5977 ( .A(n5281), .ZN(n5278) );
  AOI22_X1 U5978 ( .A1(n5279), .A2(n5764), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5278), .ZN(n5363) );
  OAI21_X1 U5979 ( .B1(n5280), .B2(n6742), .A(n5765), .ZN(n5282) );
  AOI22_X1 U5980 ( .A1(n5283), .A2(n5282), .B1(n5687), .B2(n5281), .ZN(n5284)
         );
  NAND2_X1 U5981 ( .A1(n5689), .A2(n5284), .ZN(n5356) );
  NAND2_X1 U5982 ( .A1(n5356), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5287)
         );
  OAI22_X1 U5983 ( .A1(n5518), .A2(n5358), .B1(n5357), .B2(n5794), .ZN(n5285)
         );
  AOI21_X1 U5984 ( .B1(n5792), .B2(n5360), .A(n5285), .ZN(n5286) );
  OAI211_X1 U5985 ( .C1(n5363), .C2(n5798), .A(n5287), .B(n5286), .ZN(U3142)
         );
  NAND2_X1 U5986 ( .A1(n5356), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5290)
         );
  OAI22_X1 U5987 ( .A1(n5555), .A2(n5358), .B1(n5357), .B2(n5831), .ZN(n5288)
         );
  AOI21_X1 U5988 ( .B1(n7221), .B2(n5360), .A(n5288), .ZN(n5289) );
  OAI211_X1 U5989 ( .C1(n5363), .C2(n7227), .A(n5290), .B(n5289), .ZN(U3140)
         );
  NAND2_X1 U5990 ( .A1(n5356), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5293)
         );
  OAI22_X1 U5991 ( .A1(n5521), .A2(n5358), .B1(n5357), .B2(n5801), .ZN(n5291)
         );
  AOI21_X1 U5992 ( .B1(n5799), .B2(n5360), .A(n5291), .ZN(n5292) );
  OAI211_X1 U5993 ( .C1(n5363), .C2(n5805), .A(n5293), .B(n5292), .ZN(U3143)
         );
  NAND2_X1 U5994 ( .A1(n5356), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5296)
         );
  OAI22_X1 U5995 ( .A1(n5505), .A2(n5358), .B1(n5357), .B2(n5822), .ZN(n5294)
         );
  AOI21_X1 U5996 ( .B1(n5820), .B2(n5360), .A(n5294), .ZN(n5295) );
  OAI211_X1 U5997 ( .C1(n5363), .C2(n5826), .A(n5296), .B(n5295), .ZN(U3141)
         );
  NAND2_X1 U5998 ( .A1(n5356), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5299)
         );
  OAI22_X1 U5999 ( .A1(n5778), .A2(n5358), .B1(n5357), .B2(n5697), .ZN(n5297)
         );
  AOI21_X1 U6000 ( .B1(n5776), .B2(n5360), .A(n5297), .ZN(n5298) );
  OAI211_X1 U6001 ( .C1(n5363), .C2(n5784), .A(n5299), .B(n5298), .ZN(U3147)
         );
  AOI22_X1 U6002 ( .A1(n5302), .A2(n5389), .B1(n5301), .B2(n5300), .ZN(n5340)
         );
  NAND3_X1 U6003 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7060), .ZN(n5392) );
  NOR2_X1 U6004 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5392), .ZN(n5337)
         );
  NAND2_X1 U6005 ( .A1(n5507), .A2(n5303), .ZN(n5335) );
  NAND2_X1 U6006 ( .A1(n5304), .A2(n4915), .ZN(n5334) );
  NOR2_X1 U6007 ( .A1(n5569), .A2(n5434), .ZN(n5309) );
  OR2_X1 U6008 ( .A1(n5306), .A2(n5305), .ZN(n5308) );
  AOI221_X1 U6009 ( .B1(n5309), .B2(n5308), .C1(n6581), .C2(n5308), .A(n5307), 
        .ZN(n5311) );
  OAI211_X1 U6010 ( .C1(n5337), .C2(n7084), .A(n5311), .B(n5310), .ZN(n5333)
         );
  NAND2_X1 U6011 ( .A1(n5333), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5314) );
  OAI22_X1 U6012 ( .A1(n5628), .A2(n5335), .B1(n5334), .B2(n5808), .ZN(n5312)
         );
  AOI21_X1 U6013 ( .B1(n5806), .B2(n5337), .A(n5312), .ZN(n5313) );
  OAI211_X1 U6014 ( .C1(n5340), .C2(n5812), .A(n5314), .B(n5313), .ZN(U3072)
         );
  NAND2_X1 U6015 ( .A1(n5333), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5317) );
  OAI22_X1 U6016 ( .A1(n5617), .A2(n5335), .B1(n5334), .B2(n5787), .ZN(n5315)
         );
  AOI21_X1 U6017 ( .B1(n5785), .B2(n5337), .A(n5315), .ZN(n5316) );
  OAI211_X1 U6018 ( .C1(n5340), .C2(n5791), .A(n5317), .B(n5316), .ZN(U3074)
         );
  NAND2_X1 U6019 ( .A1(n5333), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5320) );
  OAI22_X1 U6020 ( .A1(n5505), .A2(n5335), .B1(n5334), .B2(n5822), .ZN(n5318)
         );
  AOI21_X1 U6021 ( .B1(n5820), .B2(n5337), .A(n5318), .ZN(n5319) );
  OAI211_X1 U6022 ( .C1(n5340), .C2(n5826), .A(n5320), .B(n5319), .ZN(U3069)
         );
  NAND2_X1 U6023 ( .A1(n5333), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5323) );
  OAI22_X1 U6024 ( .A1(n5521), .A2(n5335), .B1(n5334), .B2(n5801), .ZN(n5321)
         );
  AOI21_X1 U6025 ( .B1(n5799), .B2(n5337), .A(n5321), .ZN(n5322) );
  OAI211_X1 U6026 ( .C1(n5340), .C2(n5805), .A(n5323), .B(n5322), .ZN(U3071)
         );
  NAND2_X1 U6027 ( .A1(n5333), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5326) );
  OAI22_X1 U6028 ( .A1(n5555), .A2(n5335), .B1(n5334), .B2(n5831), .ZN(n5324)
         );
  AOI21_X1 U6029 ( .B1(n7221), .B2(n5337), .A(n5324), .ZN(n5325) );
  OAI211_X1 U6030 ( .C1(n5340), .C2(n7227), .A(n5326), .B(n5325), .ZN(U3068)
         );
  NAND2_X1 U6031 ( .A1(n5333), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5329) );
  OAI22_X1 U6032 ( .A1(n5622), .A2(n5335), .B1(n5334), .B2(n5815), .ZN(n5327)
         );
  AOI21_X1 U6033 ( .B1(n5813), .B2(n5337), .A(n5327), .ZN(n5328) );
  OAI211_X1 U6034 ( .C1(n5340), .C2(n5819), .A(n5329), .B(n5328), .ZN(U3073)
         );
  NAND2_X1 U6035 ( .A1(n5333), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5332) );
  OAI22_X1 U6036 ( .A1(n5778), .A2(n5335), .B1(n5334), .B2(n5697), .ZN(n5330)
         );
  AOI21_X1 U6037 ( .B1(n5776), .B2(n5337), .A(n5330), .ZN(n5331) );
  OAI211_X1 U6038 ( .C1(n5340), .C2(n5784), .A(n5332), .B(n5331), .ZN(U3075)
         );
  NAND2_X1 U6039 ( .A1(n5333), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5339) );
  OAI22_X1 U6040 ( .A1(n5518), .A2(n5335), .B1(n5334), .B2(n5794), .ZN(n5336)
         );
  AOI21_X1 U6041 ( .B1(n5792), .B2(n5337), .A(n5336), .ZN(n5338) );
  OAI211_X1 U6042 ( .C1(n5340), .C2(n5798), .A(n5339), .B(n5338), .ZN(U3070)
         );
  NAND2_X1 U6043 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  XOR2_X1 U6044 ( .A(n5344), .B(n5343), .Z(n5656) );
  INV_X1 U6045 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5345) );
  AOI22_X1 U6046 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n6791), .B1(n6808), 
        .B2(n5345), .ZN(n5346) );
  NAND2_X1 U6047 ( .A1(n6847), .A2(REIP_REG_3__SCAN_IN), .ZN(n5657) );
  OAI211_X1 U6048 ( .C1(n6794), .C2(n5347), .A(n5346), .B(n5657), .ZN(n5348)
         );
  AOI21_X1 U6049 ( .B1(n5656), .B2(n6857), .A(n5348), .ZN(n5349) );
  INV_X1 U6050 ( .A(n5349), .ZN(U3015) );
  NAND2_X1 U6051 ( .A1(n5356), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5352)
         );
  OAI22_X1 U6052 ( .A1(n5628), .A2(n5358), .B1(n5357), .B2(n5808), .ZN(n5350)
         );
  AOI21_X1 U6053 ( .B1(n5806), .B2(n5360), .A(n5350), .ZN(n5351) );
  OAI211_X1 U6054 ( .C1(n5363), .C2(n5812), .A(n5352), .B(n5351), .ZN(U3144)
         );
  NAND2_X1 U6055 ( .A1(n5356), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5355)
         );
  OAI22_X1 U6056 ( .A1(n5617), .A2(n5358), .B1(n5357), .B2(n5787), .ZN(n5353)
         );
  AOI21_X1 U6057 ( .B1(n5785), .B2(n5360), .A(n5353), .ZN(n5354) );
  OAI211_X1 U6058 ( .C1(n5363), .C2(n5791), .A(n5355), .B(n5354), .ZN(U3146)
         );
  NAND2_X1 U6059 ( .A1(n5356), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5362)
         );
  OAI22_X1 U6060 ( .A1(n5622), .A2(n5358), .B1(n5357), .B2(n5815), .ZN(n5359)
         );
  AOI21_X1 U6061 ( .B1(n5813), .B2(n5360), .A(n5359), .ZN(n5361) );
  OAI211_X1 U6062 ( .C1(n5363), .C2(n5819), .A(n5362), .B(n5361), .ZN(U3145)
         );
  NAND2_X1 U6063 ( .A1(n5365), .A2(n5364), .ZN(n7095) );
  OAI22_X1 U6064 ( .A1(n6399), .A2(n7095), .B1(n5386), .B2(n5366), .ZN(n5367)
         );
  AOI21_X1 U6065 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6399), .A(n5367), 
        .ZN(n5368) );
  OAI21_X1 U6066 ( .B1(n4915), .B2(n5369), .A(n5368), .ZN(U3465) );
  INV_X1 U6067 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5373) );
  INV_X1 U6068 ( .A(n5628), .ZN(n5810) );
  AOI22_X1 U6069 ( .A1(n5806), .A2(n5378), .B1(n5810), .B2(n5433), .ZN(n5370)
         );
  OAI21_X1 U6070 ( .B1(n5594), .B2(n5808), .A(n5370), .ZN(n5371) );
  AOI21_X1 U6071 ( .B1(n5700), .B2(n5381), .A(n5371), .ZN(n5372) );
  OAI21_X1 U6072 ( .B1(n5384), .B2(n5373), .A(n5372), .ZN(U3088) );
  INV_X1 U6073 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5377) );
  INV_X1 U6074 ( .A(n5617), .ZN(n5789) );
  AOI22_X1 U6075 ( .A1(n5785), .A2(n5378), .B1(n5789), .B2(n5433), .ZN(n5374)
         );
  OAI21_X1 U6076 ( .B1(n5594), .B2(n5787), .A(n5374), .ZN(n5375) );
  AOI21_X1 U6077 ( .B1(n5726), .B2(n5381), .A(n5375), .ZN(n5376) );
  OAI21_X1 U6078 ( .B1(n5384), .B2(n5377), .A(n5376), .ZN(U3090) );
  INV_X1 U6079 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5383) );
  INV_X1 U6080 ( .A(n5622), .ZN(n5817) );
  AOI22_X1 U6081 ( .A1(n5813), .A2(n5378), .B1(n5817), .B2(n5433), .ZN(n5379)
         );
  OAI21_X1 U6082 ( .B1(n5594), .B2(n5815), .A(n5379), .ZN(n5380) );
  AOI21_X1 U6083 ( .B1(n5705), .B2(n5381), .A(n5380), .ZN(n5382) );
  OAI21_X1 U6084 ( .B1(n5384), .B2(n5383), .A(n5382), .ZN(U3089) );
  NOR2_X1 U6085 ( .A1(n5385), .A2(n5687), .ZN(n5391) );
  NOR2_X1 U6086 ( .A1(n5387), .A2(n5386), .ZN(n5539) );
  INV_X1 U6087 ( .A(n5437), .ZN(n5388) );
  AOI21_X1 U6088 ( .B1(n5539), .B2(n5389), .A(n5388), .ZN(n5394) );
  AOI22_X1 U6089 ( .A1(n5391), .A2(n5394), .B1(n5687), .B2(n5392), .ZN(n5390)
         );
  NAND2_X1 U6090 ( .A1(n5689), .A2(n5390), .ZN(n5432) );
  INV_X1 U6091 ( .A(n5391), .ZN(n5393) );
  OAI22_X1 U6092 ( .A1(n5394), .A2(n5393), .B1(n7076), .B2(n5392), .ZN(n5431)
         );
  AOI22_X1 U6093 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5432), .B1(n5694), 
        .B2(n5431), .ZN(n5396) );
  AOI22_X1 U6094 ( .A1(n5434), .A2(n5682), .B1(n5433), .B2(n5782), .ZN(n5395)
         );
  OAI211_X1 U6095 ( .C1(n5437), .C2(n5560), .A(n5396), .B(n5395), .ZN(U3083)
         );
  NAND2_X1 U6096 ( .A1(n7050), .A2(n5535), .ZN(n5444) );
  OR2_X1 U6097 ( .A1(n5397), .A2(n6581), .ZN(n5398) );
  INV_X1 U6098 ( .A(n5444), .ZN(n5399) );
  AOI21_X1 U6099 ( .B1(n5539), .B2(n3490), .A(n5399), .ZN(n5404) );
  AOI22_X1 U6100 ( .A1(n5401), .A2(n5404), .B1(n5687), .B2(n5402), .ZN(n5400)
         );
  NAND2_X1 U6101 ( .A1(n5689), .A2(n5400), .ZN(n5439) );
  INV_X1 U6102 ( .A(n5401), .ZN(n5403) );
  OAI22_X1 U6103 ( .A1(n5404), .A2(n5403), .B1(n7076), .B2(n5402), .ZN(n5438)
         );
  AOI22_X1 U6104 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5439), .B1(n5715), 
        .B2(n5438), .ZN(n5406) );
  AOI22_X1 U6105 ( .A1(n5796), .A2(n5441), .B1(n5440), .B2(n5575), .ZN(n5405)
         );
  OAI211_X1 U6106 ( .C1(n5719), .C2(n5444), .A(n5406), .B(n5405), .ZN(U3046)
         );
  AOI22_X1 U6107 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5439), .B1(n5710), 
        .B2(n5438), .ZN(n5408) );
  AOI22_X1 U6108 ( .A1(n5803), .A2(n5441), .B1(n5440), .B2(n5550), .ZN(n5407)
         );
  OAI211_X1 U6109 ( .C1(n5714), .C2(n5444), .A(n5408), .B(n5407), .ZN(U3047)
         );
  AOI22_X1 U6110 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5439), .B1(n5581), 
        .B2(n5438), .ZN(n5410) );
  AOI22_X1 U6111 ( .A1(n7223), .A2(n5441), .B1(n5440), .B2(n7219), .ZN(n5409)
         );
  OAI211_X1 U6112 ( .C1(n5588), .C2(n5444), .A(n5410), .B(n5409), .ZN(U3044)
         );
  AOI22_X1 U6113 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5432), .B1(n5705), 
        .B2(n5431), .ZN(n5412) );
  INV_X1 U6114 ( .A(n5815), .ZN(n5624) );
  AOI22_X1 U6115 ( .A1(n5434), .A2(n5817), .B1(n5433), .B2(n5624), .ZN(n5411)
         );
  OAI211_X1 U6116 ( .C1(n5437), .C2(n5709), .A(n5412), .B(n5411), .ZN(U3081)
         );
  AOI22_X1 U6117 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5432), .B1(n5700), 
        .B2(n5431), .ZN(n5414) );
  INV_X1 U6118 ( .A(n5808), .ZN(n5631) );
  AOI22_X1 U6119 ( .A1(n5434), .A2(n5810), .B1(n5433), .B2(n5631), .ZN(n5413)
         );
  OAI211_X1 U6120 ( .C1(n5437), .C2(n5704), .A(n5414), .B(n5413), .ZN(U3080)
         );
  AOI22_X1 U6121 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5432), .B1(n5710), 
        .B2(n5431), .ZN(n5416) );
  AOI22_X1 U6122 ( .A1(n5434), .A2(n5803), .B1(n5433), .B2(n5550), .ZN(n5415)
         );
  OAI211_X1 U6123 ( .C1(n5437), .C2(n5714), .A(n5416), .B(n5415), .ZN(U3079)
         );
  INV_X1 U6124 ( .A(n5785), .ZN(n5731) );
  AOI22_X1 U6125 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5432), .B1(n5726), 
        .B2(n5431), .ZN(n5418) );
  INV_X1 U6126 ( .A(n5787), .ZN(n5619) );
  AOI22_X1 U6127 ( .A1(n5434), .A2(n5789), .B1(n5433), .B2(n5619), .ZN(n5417)
         );
  OAI211_X1 U6128 ( .C1(n5437), .C2(n5731), .A(n5418), .B(n5417), .ZN(U3082)
         );
  AOI22_X1 U6129 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5432), .B1(n5720), 
        .B2(n5431), .ZN(n5420) );
  AOI22_X1 U6130 ( .A1(n5434), .A2(n5824), .B1(n5433), .B2(n5568), .ZN(n5419)
         );
  OAI211_X1 U6131 ( .C1(n5437), .C2(n5724), .A(n5420), .B(n5419), .ZN(U3077)
         );
  AOI22_X1 U6132 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5432), .B1(n5581), 
        .B2(n5431), .ZN(n5422) );
  AOI22_X1 U6133 ( .A1(n5434), .A2(n7223), .B1(n5433), .B2(n7219), .ZN(n5421)
         );
  OAI211_X1 U6134 ( .C1(n5437), .C2(n5588), .A(n5422), .B(n5421), .ZN(U3076)
         );
  AOI22_X1 U6135 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5439), .B1(n5694), 
        .B2(n5438), .ZN(n5424) );
  AOI22_X1 U6136 ( .A1(n5682), .A2(n5441), .B1(n5440), .B2(n5782), .ZN(n5423)
         );
  OAI211_X1 U6137 ( .C1(n5560), .C2(n5444), .A(n5424), .B(n5423), .ZN(U3051)
         );
  AOI22_X1 U6138 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5439), .B1(n5700), 
        .B2(n5438), .ZN(n5426) );
  AOI22_X1 U6139 ( .A1(n5810), .A2(n5441), .B1(n5440), .B2(n5631), .ZN(n5425)
         );
  OAI211_X1 U6140 ( .C1(n5704), .C2(n5444), .A(n5426), .B(n5425), .ZN(U3048)
         );
  AOI22_X1 U6141 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5439), .B1(n5720), 
        .B2(n5438), .ZN(n5428) );
  AOI22_X1 U6142 ( .A1(n5824), .A2(n5441), .B1(n5440), .B2(n5568), .ZN(n5427)
         );
  OAI211_X1 U6143 ( .C1(n5724), .C2(n5444), .A(n5428), .B(n5427), .ZN(U3045)
         );
  AOI22_X1 U6144 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5439), .B1(n5726), 
        .B2(n5438), .ZN(n5430) );
  AOI22_X1 U6145 ( .A1(n5789), .A2(n5441), .B1(n5440), .B2(n5619), .ZN(n5429)
         );
  OAI211_X1 U6146 ( .C1(n5731), .C2(n5444), .A(n5430), .B(n5429), .ZN(U3050)
         );
  AOI22_X1 U6147 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5432), .B1(n5715), 
        .B2(n5431), .ZN(n5436) );
  AOI22_X1 U6148 ( .A1(n5434), .A2(n5796), .B1(n5433), .B2(n5575), .ZN(n5435)
         );
  OAI211_X1 U6149 ( .C1(n5437), .C2(n5719), .A(n5436), .B(n5435), .ZN(U3078)
         );
  AOI22_X1 U6150 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5439), .B1(n5705), 
        .B2(n5438), .ZN(n5443) );
  AOI22_X1 U6151 ( .A1(n5817), .A2(n5441), .B1(n5440), .B2(n5624), .ZN(n5442)
         );
  OAI211_X1 U6152 ( .C1(n5709), .C2(n5444), .A(n5443), .B(n5442), .ZN(U3049)
         );
  OAI21_X1 U6153 ( .B1(n3485), .B2(n5446), .A(n5445), .ZN(n5744) );
  NOR2_X1 U6154 ( .A1(n7010), .A2(n5751), .ZN(n6902) );
  INV_X1 U6155 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6647) );
  INV_X1 U6156 ( .A(n5447), .ZN(n5450) );
  INV_X1 U6157 ( .A(n5448), .ZN(n5449) );
  OAI21_X1 U6158 ( .B1(n5450), .B2(n5449), .A(n5676), .ZN(n6823) );
  AOI21_X1 U6159 ( .B1(n5747), .B2(n7017), .A(n6974), .ZN(n5451) );
  OAI21_X1 U6160 ( .B1(n7006), .B2(n6823), .A(n5451), .ZN(n5455) );
  AOI22_X1 U6161 ( .A1(EBX_REG_9__SCAN_IN), .A2(n7008), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5597), .ZN(n5452) );
  OAI21_X1 U6162 ( .B1(n5453), .B2(n6980), .A(n5452), .ZN(n5454) );
  AOI211_X1 U6163 ( .C1(n6902), .C2(n6647), .A(n5455), .B(n5454), .ZN(n5456)
         );
  OAI21_X1 U6164 ( .B1(n7001), .B2(n5744), .A(n5456), .ZN(U2818) );
  NOR2_X1 U6165 ( .A1(n6994), .A2(n6116), .ZN(n6929) );
  INV_X1 U6166 ( .A(REIP_REG_0__SCAN_IN), .ZN(n5463) );
  INV_X1 U6167 ( .A(n6120), .ZN(n5460) );
  OAI21_X1 U6168 ( .B1(n7009), .B2(n7017), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5457) );
  OAI21_X1 U6169 ( .B1(n6998), .B2(n5458), .A(n5457), .ZN(n5459) );
  AOI21_X1 U6170 ( .B1(n5460), .B2(n6711), .A(n5459), .ZN(n5462) );
  INV_X1 U6171 ( .A(n5992), .ZN(n6123) );
  AOI22_X1 U6172 ( .A1(n6123), .A2(n5972), .B1(n7015), .B2(n6874), .ZN(n5461)
         );
  OAI211_X1 U6173 ( .C1(n6929), .C2(n5463), .A(n5462), .B(n5461), .ZN(U2827)
         );
  INV_X1 U6174 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5464) );
  OAI222_X1 U6175 ( .A1(n5744), .A2(n6156), .B1(n5464), .B2(n6706), .C1(n6154), 
        .C2(n6823), .ZN(U2850) );
  INV_X1 U6176 ( .A(DATAI_9_), .ZN(n6550) );
  INV_X1 U6177 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7171) );
  OAI222_X1 U6178 ( .A1(n5744), .A2(n7201), .B1(n5916), .B2(n6550), .C1(n6015), 
        .C2(n7171), .ZN(U2882) );
  XOR2_X1 U6179 ( .A(n5465), .B(n5466), .Z(n5649) );
  OAI22_X1 U6180 ( .A1(n6794), .A2(n5473), .B1(n6641), .B2(n6860), .ZN(n5470)
         );
  NAND3_X1 U6181 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6808), .ZN(n5609) );
  NAND3_X1 U6182 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n5467) );
  INV_X1 U6183 ( .A(n6787), .ZN(n6789) );
  AOI221_X1 U6184 ( .B1(n5468), .B2(n6790), .C1(n5467), .C2(n6790), .A(n6789), 
        .ZN(n5611) );
  AOI21_X1 U6185 ( .B1(n5610), .B2(n5609), .A(n5611), .ZN(n5469) );
  AOI211_X1 U6186 ( .C1(n5649), .C2(n6857), .A(n5470), .B(n5469), .ZN(n5471)
         );
  INV_X1 U6187 ( .A(n5471), .ZN(U3013) );
  INV_X1 U6188 ( .A(n5472), .ZN(n6879) );
  NAND2_X1 U6189 ( .A1(n6994), .A2(n6879), .ZN(n5479) );
  NAND2_X1 U6190 ( .A1(n5479), .A2(n6107), .ZN(n6897) );
  INV_X1 U6191 ( .A(n5652), .ZN(n5477) );
  NAND2_X1 U6192 ( .A1(n7008), .A2(EBX_REG_5__SCAN_IN), .ZN(n5476) );
  OAI22_X1 U6193 ( .A1(n5650), .A2(n6980), .B1(n7006), .B2(n5473), .ZN(n5474)
         );
  NOR2_X1 U6194 ( .A1(n6974), .A2(n5474), .ZN(n5475) );
  OAI211_X1 U6195 ( .C1(n6999), .C2(n5477), .A(n5476), .B(n5475), .ZN(n5481)
         );
  NOR2_X1 U6196 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  AOI211_X1 U6197 ( .C1(REIP_REG_5__SCAN_IN), .C2(n6897), .A(n5481), .B(n5480), 
        .ZN(n5482) );
  OAI21_X1 U6198 ( .B1(n6120), .B2(n5655), .A(n5482), .ZN(U2822) );
  OAI21_X1 U6199 ( .B1(n5485), .B2(n5484), .A(n5483), .ZN(n6792) );
  INV_X1 U6200 ( .A(n5486), .ZN(n5490) );
  AOI22_X1 U6201 ( .A1(n6749), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6847), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5487) );
  OAI21_X1 U6202 ( .B1(n6755), .B2(n5488), .A(n5487), .ZN(n5489) );
  AOI21_X1 U6203 ( .B1(n5490), .B2(n6254), .A(n5489), .ZN(n5491) );
  OAI21_X1 U6204 ( .B1(n6792), .B2(n7033), .A(n5491), .ZN(U2978) );
  INV_X1 U6205 ( .A(n5493), .ZN(n5494) );
  OR2_X1 U6206 ( .A1(n5445), .A2(n5493), .ZN(n5674) );
  OAI21_X1 U6207 ( .B1(n5492), .B2(n5494), .A(n5674), .ZN(n5741) );
  INV_X1 U6208 ( .A(n5678), .ZN(n5495) );
  XNOR2_X1 U6209 ( .A(n5676), .B(n5495), .ZN(n5600) );
  INV_X1 U6210 ( .A(n5600), .ZN(n6812) );
  AOI22_X1 U6211 ( .A1(n6702), .A2(n6812), .B1(EBX_REG_10__SCAN_IN), .B2(n4769), .ZN(n5496) );
  OAI21_X1 U6212 ( .B1(n5741), .B2(n6156), .A(n5496), .ZN(U2849) );
  OAI21_X1 U6213 ( .B1(n5502), .B2(n6581), .A(n5764), .ZN(n5501) );
  NOR2_X1 U6214 ( .A1(n7043), .A2(n5499), .ZN(n5591) );
  AOI21_X1 U6215 ( .B1(n5685), .B2(n5538), .A(n5591), .ZN(n5500) );
  INV_X1 U6216 ( .A(n5500), .ZN(n5498) );
  NAND2_X1 U6217 ( .A1(n5687), .A2(n5499), .ZN(n5497) );
  OAI211_X1 U6218 ( .C1(n5501), .C2(n5498), .A(n5689), .B(n5497), .ZN(n5590)
         );
  OAI22_X1 U6219 ( .A1(n5501), .A2(n5500), .B1(n7076), .B2(n5499), .ZN(n5589)
         );
  AOI22_X1 U6220 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5590), .B1(n5720), 
        .B2(n5589), .ZN(n5504) );
  AOI22_X1 U6221 ( .A1(n5833), .A2(n5568), .B1(n5820), .B2(n5591), .ZN(n5503)
         );
  OAI211_X1 U6222 ( .C1(n5594), .C2(n5505), .A(n5504), .B(n5503), .ZN(U3093)
         );
  NOR2_X1 U6223 ( .A1(n7043), .A2(n5511), .ZN(n5506) );
  INV_X1 U6224 ( .A(n5506), .ZN(n5572) );
  AOI21_X1 U6225 ( .B1(n5539), .B2(n5684), .A(n5506), .ZN(n5513) );
  INV_X1 U6226 ( .A(n5513), .ZN(n5510) );
  INV_X1 U6227 ( .A(n5507), .ZN(n5508) );
  OAI21_X1 U6228 ( .B1(n5508), .B2(n6581), .A(n5764), .ZN(n5512) );
  NAND2_X1 U6229 ( .A1(n5687), .A2(n5511), .ZN(n5509) );
  OAI211_X1 U6230 ( .C1(n5510), .C2(n5512), .A(n5689), .B(n5509), .ZN(n5566)
         );
  OAI22_X1 U6231 ( .A1(n5513), .A2(n5512), .B1(n7076), .B2(n5511), .ZN(n5565)
         );
  AOI22_X1 U6232 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5566), .B1(n5581), 
        .B2(n5565), .ZN(n5515) );
  AOI22_X1 U6233 ( .A1(n5569), .A2(n7219), .B1(n5567), .B2(n7223), .ZN(n5514)
         );
  OAI211_X1 U6234 ( .C1(n5588), .C2(n5572), .A(n5515), .B(n5514), .ZN(U3060)
         );
  AOI22_X1 U6235 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5590), .B1(n5715), 
        .B2(n5589), .ZN(n5517) );
  AOI22_X1 U6236 ( .A1(n5833), .A2(n5575), .B1(n5792), .B2(n5591), .ZN(n5516)
         );
  OAI211_X1 U6237 ( .C1(n5594), .C2(n5518), .A(n5517), .B(n5516), .ZN(U3094)
         );
  AOI22_X1 U6238 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5590), .B1(n5710), 
        .B2(n5589), .ZN(n5520) );
  AOI22_X1 U6239 ( .A1(n5833), .A2(n5550), .B1(n5799), .B2(n5591), .ZN(n5519)
         );
  OAI211_X1 U6240 ( .C1(n5594), .C2(n5521), .A(n5520), .B(n5519), .ZN(U3095)
         );
  AOI22_X1 U6241 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5566), .B1(n5710), 
        .B2(n5565), .ZN(n5523) );
  AOI22_X1 U6242 ( .A1(n5569), .A2(n5550), .B1(n5567), .B2(n5803), .ZN(n5522)
         );
  OAI211_X1 U6243 ( .C1(n5714), .C2(n5572), .A(n5523), .B(n5522), .ZN(U3063)
         );
  AOI22_X1 U6244 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5566), .B1(n5700), 
        .B2(n5565), .ZN(n5525) );
  AOI22_X1 U6245 ( .A1(n5569), .A2(n5631), .B1(n5567), .B2(n5810), .ZN(n5524)
         );
  OAI211_X1 U6246 ( .C1(n5704), .C2(n5572), .A(n5525), .B(n5524), .ZN(U3064)
         );
  AOI22_X1 U6247 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5566), .B1(n5715), 
        .B2(n5565), .ZN(n5527) );
  AOI22_X1 U6248 ( .A1(n5569), .A2(n5575), .B1(n5567), .B2(n5796), .ZN(n5526)
         );
  OAI211_X1 U6249 ( .C1(n5719), .C2(n5572), .A(n5527), .B(n5526), .ZN(U3062)
         );
  AOI22_X1 U6250 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5566), .B1(n5726), 
        .B2(n5565), .ZN(n5529) );
  AOI22_X1 U6251 ( .A1(n5569), .A2(n5619), .B1(n5567), .B2(n5789), .ZN(n5528)
         );
  OAI211_X1 U6252 ( .C1(n5731), .C2(n5572), .A(n5529), .B(n5528), .ZN(U3066)
         );
  AOI22_X1 U6253 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5566), .B1(n5694), 
        .B2(n5565), .ZN(n5531) );
  AOI22_X1 U6254 ( .A1(n5569), .A2(n5782), .B1(n5567), .B2(n5682), .ZN(n5530)
         );
  OAI211_X1 U6255 ( .C1(n5560), .C2(n5572), .A(n5531), .B(n5530), .ZN(U3067)
         );
  AOI22_X1 U6256 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5566), .B1(n5705), 
        .B2(n5565), .ZN(n5533) );
  AOI22_X1 U6257 ( .A1(n5569), .A2(n5624), .B1(n5567), .B2(n5817), .ZN(n5532)
         );
  OAI211_X1 U6258 ( .C1(n5709), .C2(n5572), .A(n5533), .B(n5532), .ZN(U3065)
         );
  NAND2_X1 U6259 ( .A1(n5535), .A2(n5534), .ZN(n5543) );
  NOR2_X1 U6260 ( .A1(n7043), .A2(n5543), .ZN(n5537) );
  INV_X1 U6261 ( .A(n5537), .ZN(n5587) );
  INV_X1 U6262 ( .A(n5543), .ZN(n5542) );
  OAI21_X1 U6263 ( .B1(n5536), .B2(n6581), .A(n5764), .ZN(n5544) );
  INV_X1 U6264 ( .A(n5544), .ZN(n5540) );
  AOI21_X1 U6265 ( .B1(n5539), .B2(n5538), .A(n5537), .ZN(n5545) );
  NAND2_X1 U6266 ( .A1(n5540), .A2(n5545), .ZN(n5541) );
  OAI211_X1 U6267 ( .C1(n5764), .C2(n5542), .A(n5689), .B(n5541), .ZN(n5582)
         );
  OAI22_X1 U6268 ( .A1(n5545), .A2(n5544), .B1(n7076), .B2(n5543), .ZN(n5580)
         );
  AOI22_X1 U6269 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5582), .B1(n5705), 
        .B2(n5580), .ZN(n5547) );
  AOI22_X1 U6270 ( .A1(n5817), .A2(n5584), .B1(n5583), .B2(n5624), .ZN(n5546)
         );
  OAI211_X1 U6271 ( .C1(n5709), .C2(n5587), .A(n5547), .B(n5546), .ZN(U3033)
         );
  AOI22_X1 U6272 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5582), .B1(n5700), 
        .B2(n5580), .ZN(n5549) );
  AOI22_X1 U6273 ( .A1(n5810), .A2(n5584), .B1(n5583), .B2(n5631), .ZN(n5548)
         );
  OAI211_X1 U6274 ( .C1(n5704), .C2(n5587), .A(n5549), .B(n5548), .ZN(U3032)
         );
  AOI22_X1 U6275 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5582), .B1(n5710), 
        .B2(n5580), .ZN(n5552) );
  AOI22_X1 U6276 ( .A1(n5803), .A2(n5584), .B1(n5583), .B2(n5550), .ZN(n5551)
         );
  OAI211_X1 U6277 ( .C1(n5714), .C2(n5587), .A(n5552), .B(n5551), .ZN(U3031)
         );
  AOI22_X1 U6278 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5590), .B1(n5581), 
        .B2(n5589), .ZN(n5554) );
  AOI22_X1 U6279 ( .A1(n7219), .A2(n5833), .B1(n7221), .B2(n5591), .ZN(n5553)
         );
  OAI211_X1 U6280 ( .C1(n5594), .C2(n5555), .A(n5554), .B(n5553), .ZN(U3092)
         );
  AOI22_X1 U6281 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5582), .B1(n5720), 
        .B2(n5580), .ZN(n5557) );
  AOI22_X1 U6282 ( .A1(n5824), .A2(n5584), .B1(n5583), .B2(n5568), .ZN(n5556)
         );
  OAI211_X1 U6283 ( .C1(n5724), .C2(n5587), .A(n5557), .B(n5556), .ZN(U3029)
         );
  AOI22_X1 U6284 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5582), .B1(n5694), 
        .B2(n5580), .ZN(n5559) );
  AOI22_X1 U6285 ( .A1(n5682), .A2(n5584), .B1(n5583), .B2(n5782), .ZN(n5558)
         );
  OAI211_X1 U6286 ( .C1(n5560), .C2(n5587), .A(n5559), .B(n5558), .ZN(U3035)
         );
  AOI22_X1 U6287 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5582), .B1(n5726), 
        .B2(n5580), .ZN(n5562) );
  AOI22_X1 U6288 ( .A1(n5789), .A2(n5584), .B1(n5583), .B2(n5619), .ZN(n5561)
         );
  OAI211_X1 U6289 ( .C1(n5731), .C2(n5587), .A(n5562), .B(n5561), .ZN(U3034)
         );
  AOI22_X1 U6290 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5590), .B1(n5694), 
        .B2(n5589), .ZN(n5564) );
  AOI22_X1 U6291 ( .A1(n5833), .A2(n5782), .B1(n5776), .B2(n5591), .ZN(n5563)
         );
  OAI211_X1 U6292 ( .C1(n5594), .C2(n5778), .A(n5564), .B(n5563), .ZN(U3099)
         );
  AOI22_X1 U6293 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5566), .B1(n5720), 
        .B2(n5565), .ZN(n5571) );
  AOI22_X1 U6294 ( .A1(n5569), .A2(n5568), .B1(n5567), .B2(n5824), .ZN(n5570)
         );
  OAI211_X1 U6295 ( .C1(n5724), .C2(n5572), .A(n5571), .B(n5570), .ZN(U3061)
         );
  AOI22_X1 U6296 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5590), .B1(n5705), 
        .B2(n5589), .ZN(n5574) );
  AOI22_X1 U6297 ( .A1(n5833), .A2(n5624), .B1(n5813), .B2(n5591), .ZN(n5573)
         );
  OAI211_X1 U6298 ( .C1(n5594), .C2(n5622), .A(n5574), .B(n5573), .ZN(U3097)
         );
  AOI22_X1 U6299 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5582), .B1(n5715), 
        .B2(n5580), .ZN(n5577) );
  AOI22_X1 U6300 ( .A1(n5796), .A2(n5584), .B1(n5583), .B2(n5575), .ZN(n5576)
         );
  OAI211_X1 U6301 ( .C1(n5719), .C2(n5587), .A(n5577), .B(n5576), .ZN(U3030)
         );
  AOI22_X1 U6302 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5590), .B1(n5700), 
        .B2(n5589), .ZN(n5579) );
  AOI22_X1 U6303 ( .A1(n5833), .A2(n5631), .B1(n5806), .B2(n5591), .ZN(n5578)
         );
  OAI211_X1 U6304 ( .C1(n5594), .C2(n5628), .A(n5579), .B(n5578), .ZN(U3096)
         );
  AOI22_X1 U6305 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5582), .B1(n5581), 
        .B2(n5580), .ZN(n5586) );
  AOI22_X1 U6306 ( .A1(n7223), .A2(n5584), .B1(n5583), .B2(n7219), .ZN(n5585)
         );
  OAI211_X1 U6307 ( .C1(n5588), .C2(n5587), .A(n5586), .B(n5585), .ZN(U3028)
         );
  AOI22_X1 U6308 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5590), .B1(n5726), 
        .B2(n5589), .ZN(n5593) );
  AOI22_X1 U6309 ( .A1(n5833), .A2(n5619), .B1(n5785), .B2(n5591), .ZN(n5592)
         );
  OAI211_X1 U6310 ( .C1(n5594), .C2(n5617), .A(n5593), .B(n5592), .ZN(U3098)
         );
  INV_X1 U6311 ( .A(n5737), .ZN(n5602) );
  OAI22_X1 U6312 ( .A1(n4331), .A2(n6980), .B1(n5595), .B2(n6998), .ZN(n5596)
         );
  AOI211_X1 U6313 ( .C1(REIP_REG_10__SCAN_IN), .C2(n5597), .A(n6974), .B(n5596), .ZN(n5599) );
  NAND2_X1 U6314 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n6903) );
  OAI211_X1 U6315 ( .C1(REIP_REG_9__SCAN_IN), .C2(REIP_REG_10__SCAN_IN), .A(
        n6902), .B(n6903), .ZN(n5598) );
  OAI211_X1 U6316 ( .C1(n5600), .C2(n7006), .A(n5599), .B(n5598), .ZN(n5601)
         );
  AOI21_X1 U6317 ( .B1(n7017), .B2(n5602), .A(n5601), .ZN(n5603) );
  OAI21_X1 U6318 ( .B1(n7001), .B2(n5741), .A(n5603), .ZN(U2817) );
  NAND2_X1 U6319 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  XNOR2_X1 U6320 ( .A(n5604), .B(n5607), .ZN(n6728) );
  INV_X1 U6321 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5608) );
  OAI22_X1 U6322 ( .A1(n6794), .A2(n6882), .B1(n6860), .B2(n5608), .ZN(n5615)
         );
  NOR2_X1 U6323 ( .A1(n5610), .A2(n5609), .ZN(n5613) );
  INV_X1 U6324 ( .A(n5611), .ZN(n5612) );
  MUX2_X1 U6325 ( .A(n5613), .B(n5612), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n5614) );
  AOI211_X1 U6326 ( .C1(n6857), .C2(n6728), .A(n5615), .B(n5614), .ZN(n5616)
         );
  INV_X1 U6327 ( .A(n5616), .ZN(U3012) );
  NAND2_X1 U6328 ( .A1(n5627), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5621)
         );
  OAI22_X1 U6329 ( .A1(n5731), .A2(n5629), .B1(n5617), .B2(n5830), .ZN(n5618)
         );
  AOI21_X1 U6330 ( .B1(n5619), .B2(n5645), .A(n5618), .ZN(n5620) );
  OAI211_X1 U6331 ( .C1(n5634), .C2(n5791), .A(n5621), .B(n5620), .ZN(U3114)
         );
  NAND2_X1 U6332 ( .A1(n5627), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5626)
         );
  OAI22_X1 U6333 ( .A1(n5709), .A2(n5629), .B1(n5622), .B2(n5830), .ZN(n5623)
         );
  AOI21_X1 U6334 ( .B1(n5624), .B2(n5645), .A(n5623), .ZN(n5625) );
  OAI211_X1 U6335 ( .C1(n5634), .C2(n5819), .A(n5626), .B(n5625), .ZN(U3113)
         );
  NAND2_X1 U6336 ( .A1(n5627), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5633)
         );
  OAI22_X1 U6337 ( .A1(n5704), .A2(n5629), .B1(n5628), .B2(n5830), .ZN(n5630)
         );
  AOI21_X1 U6338 ( .B1(n5631), .B2(n5645), .A(n5630), .ZN(n5632) );
  OAI211_X1 U6339 ( .C1(n5634), .C2(n5812), .A(n5633), .B(n5632), .ZN(U3112)
         );
  NAND2_X1 U6340 ( .A1(n5641), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5637)
         );
  OAI22_X1 U6341 ( .A1(n5709), .A2(n5643), .B1(n5815), .B2(n5642), .ZN(n5635)
         );
  AOI21_X1 U6342 ( .B1(n5817), .B2(n5645), .A(n5635), .ZN(n5636) );
  OAI211_X1 U6343 ( .C1(n5648), .C2(n5819), .A(n5637), .B(n5636), .ZN(U3121)
         );
  NAND2_X1 U6344 ( .A1(n5641), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5640)
         );
  OAI22_X1 U6345 ( .A1(n5704), .A2(n5643), .B1(n5808), .B2(n5642), .ZN(n5638)
         );
  AOI21_X1 U6346 ( .B1(n5810), .B2(n5645), .A(n5638), .ZN(n5639) );
  OAI211_X1 U6347 ( .C1(n5648), .C2(n5812), .A(n5640), .B(n5639), .ZN(U3120)
         );
  NAND2_X1 U6348 ( .A1(n5641), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5647)
         );
  OAI22_X1 U6349 ( .A1(n5731), .A2(n5643), .B1(n5787), .B2(n5642), .ZN(n5644)
         );
  AOI21_X1 U6350 ( .B1(n5789), .B2(n5645), .A(n5644), .ZN(n5646) );
  OAI211_X1 U6351 ( .C1(n5648), .C2(n5791), .A(n5647), .B(n5646), .ZN(U3122)
         );
  NAND2_X1 U6352 ( .A1(n5649), .A2(n6751), .ZN(n5654) );
  INV_X1 U6353 ( .A(n6749), .ZN(n6710) );
  OAI22_X1 U6354 ( .A1(n6710), .A2(n5650), .B1(n6860), .B2(n6641), .ZN(n5651)
         );
  AOI21_X1 U6355 ( .B1(n5652), .B2(n6269), .A(n5651), .ZN(n5653) );
  OAI211_X1 U6356 ( .C1(n6742), .C2(n5655), .A(n5654), .B(n5653), .ZN(U2981)
         );
  NAND2_X1 U6357 ( .A1(n5656), .A2(n6751), .ZN(n5662) );
  INV_X1 U6358 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5658) );
  OAI21_X1 U6359 ( .B1(n6710), .B2(n5658), .A(n5657), .ZN(n5659) );
  AOI21_X1 U6360 ( .B1(n5660), .B2(n6269), .A(n5659), .ZN(n5661) );
  OAI211_X1 U6361 ( .C1(n6742), .C2(n5663), .A(n5662), .B(n5661), .ZN(U2983)
         );
  INV_X1 U6362 ( .A(DATAI_10_), .ZN(n6546) );
  INV_X1 U6363 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7176) );
  OAI222_X1 U6364 ( .A1(n5741), .A2(n7201), .B1(n5916), .B2(n6546), .C1(n6015), 
        .C2(n7176), .ZN(U2881) );
  NAND2_X1 U6365 ( .A1(n5664), .A2(n6254), .ZN(n5670) );
  NOR2_X1 U6366 ( .A1(n6710), .A2(n5665), .ZN(n5666) );
  AOI211_X1 U6367 ( .C1(n6269), .C2(n5668), .A(n5667), .B(n5666), .ZN(n5669)
         );
  OAI211_X1 U6368 ( .C1(n5671), .C2(n7033), .A(n5670), .B(n5669), .ZN(U2982)
         );
  INV_X1 U6369 ( .A(n5672), .ZN(n5750) );
  NAND2_X1 U6370 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND2_X1 U6371 ( .A1(n5750), .A2(n5675), .ZN(n6908) );
  INV_X1 U6372 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5681) );
  INV_X1 U6373 ( .A(n5676), .ZN(n5679) );
  AOI21_X1 U6374 ( .B1(n5679), .B2(n5678), .A(n5677), .ZN(n5680) );
  OR2_X1 U6375 ( .A1(n5680), .A2(n3475), .ZN(n6833) );
  OAI222_X1 U6376 ( .A1(n6908), .A2(n6156), .B1(n5681), .B2(n6706), .C1(n6154), 
        .C2(n6833), .ZN(U2848) );
  INV_X1 U6377 ( .A(DATAI_11_), .ZN(n6544) );
  INV_X1 U6378 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7181) );
  OAI222_X1 U6379 ( .A1(n6908), .A2(n7201), .B1(n5916), .B2(n6544), .C1(n6015), 
        .C2(n7181), .ZN(U2880) );
  NOR2_X1 U6380 ( .A1(n7043), .A2(n5686), .ZN(n7220) );
  NAND2_X1 U6381 ( .A1(n7222), .A2(n5682), .ZN(n5696) );
  NOR2_X1 U6382 ( .A1(n5683), .A2(n5687), .ZN(n5692) );
  AOI21_X1 U6383 ( .B1(n5685), .B2(n5684), .A(n7220), .ZN(n5690) );
  AOI22_X1 U6384 ( .A1(n5692), .A2(n5690), .B1(n5687), .B2(n5686), .ZN(n5688)
         );
  NAND2_X1 U6385 ( .A1(n5689), .A2(n5688), .ZN(n7224) );
  INV_X1 U6386 ( .A(n5690), .ZN(n5691) );
  AOI22_X1 U6387 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5693), .B1(n5692), .B2(
        n5691), .ZN(n7228) );
  INV_X1 U6388 ( .A(n7228), .ZN(n5725) );
  AOI22_X1 U6389 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n7224), .B1(n5694), 
        .B2(n5725), .ZN(n5695) );
  OAI211_X1 U6390 ( .C1(n7217), .C2(n5697), .A(n5696), .B(n5695), .ZN(n5698)
         );
  AOI21_X1 U6391 ( .B1(n5776), .B2(n7220), .A(n5698), .ZN(n5699) );
  INV_X1 U6392 ( .A(n5699), .ZN(U3131) );
  INV_X1 U6393 ( .A(n7220), .ZN(n5730) );
  AOI22_X1 U6394 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n7224), .B1(n5700), 
        .B2(n5725), .ZN(n5701) );
  OAI21_X1 U6395 ( .B1(n7217), .B2(n5808), .A(n5701), .ZN(n5702) );
  AOI21_X1 U6396 ( .B1(n5810), .B2(n7222), .A(n5702), .ZN(n5703) );
  OAI21_X1 U6397 ( .B1(n5704), .B2(n5730), .A(n5703), .ZN(U3128) );
  AOI22_X1 U6398 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n7224), .B1(n5705), 
        .B2(n5725), .ZN(n5706) );
  OAI21_X1 U6399 ( .B1(n7217), .B2(n5815), .A(n5706), .ZN(n5707) );
  AOI21_X1 U6400 ( .B1(n5817), .B2(n7222), .A(n5707), .ZN(n5708) );
  OAI21_X1 U6401 ( .B1(n5709), .B2(n5730), .A(n5708), .ZN(U3129) );
  AOI22_X1 U6402 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n7224), .B1(n5710), 
        .B2(n5725), .ZN(n5711) );
  OAI21_X1 U6403 ( .B1(n7217), .B2(n5801), .A(n5711), .ZN(n5712) );
  AOI21_X1 U6404 ( .B1(n5803), .B2(n7222), .A(n5712), .ZN(n5713) );
  OAI21_X1 U6405 ( .B1(n5714), .B2(n5730), .A(n5713), .ZN(U3127) );
  AOI22_X1 U6406 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n7224), .B1(n5715), 
        .B2(n5725), .ZN(n5716) );
  OAI21_X1 U6407 ( .B1(n7217), .B2(n5794), .A(n5716), .ZN(n5717) );
  AOI21_X1 U6408 ( .B1(n5796), .B2(n7222), .A(n5717), .ZN(n5718) );
  OAI21_X1 U6409 ( .B1(n5719), .B2(n5730), .A(n5718), .ZN(U3126) );
  AOI22_X1 U6410 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n7224), .B1(n5720), 
        .B2(n5725), .ZN(n5721) );
  OAI21_X1 U6411 ( .B1(n7217), .B2(n5822), .A(n5721), .ZN(n5722) );
  AOI21_X1 U6412 ( .B1(n5824), .B2(n7222), .A(n5722), .ZN(n5723) );
  OAI21_X1 U6413 ( .B1(n5724), .B2(n5730), .A(n5723), .ZN(U3125) );
  AOI22_X1 U6414 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n7224), .B1(n5726), 
        .B2(n5725), .ZN(n5727) );
  OAI21_X1 U6415 ( .B1(n7217), .B2(n5787), .A(n5727), .ZN(n5728) );
  AOI21_X1 U6416 ( .B1(n5789), .B2(n7222), .A(n5728), .ZN(n5729) );
  OAI21_X1 U6417 ( .B1(n5731), .B2(n5730), .A(n5729), .ZN(U3130) );
  NAND2_X1 U6418 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  XNOR2_X1 U6419 ( .A(n5732), .B(n5735), .ZN(n6819) );
  NAND2_X1 U6420 ( .A1(n6819), .A2(n6751), .ZN(n5740) );
  INV_X1 U6421 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5736) );
  NOR2_X1 U6422 ( .A1(n6860), .A2(n5736), .ZN(n6811) );
  NOR2_X1 U6423 ( .A1(n6755), .A2(n5737), .ZN(n5738) );
  AOI211_X1 U6424 ( .C1(n6749), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6811), 
        .B(n5738), .ZN(n5739) );
  OAI211_X1 U6425 ( .C1(n6742), .C2(n5741), .A(n5740), .B(n5739), .ZN(U2976)
         );
  NAND2_X1 U6426 ( .A1(n6847), .A2(REIP_REG_9__SCAN_IN), .ZN(n6824) );
  OAI21_X1 U6427 ( .B1(n6710), .B2(n5453), .A(n6824), .ZN(n5746) );
  NOR2_X1 U6428 ( .A1(n5744), .A2(n6742), .ZN(n5745) );
  AOI211_X1 U6429 ( .C1(n6269), .C2(n5747), .A(n5746), .B(n5745), .ZN(n5748)
         );
  OAI21_X1 U6430 ( .B1(n7033), .B2(n6827), .A(n5748), .ZN(U2977) );
  XNOR2_X1 U6431 ( .A(n5750), .B(n5749), .ZN(n5851) );
  INV_X1 U6432 ( .A(n5851), .ZN(n5763) );
  INV_X1 U6433 ( .A(DATAI_12_), .ZN(n6509) );
  OAI222_X1 U6434 ( .A1(n7201), .A2(n5763), .B1(n5916), .B2(n6509), .C1(n6015), 
        .C2(n4366), .ZN(U2879) );
  INV_X1 U6435 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6650) );
  NOR3_X1 U6436 ( .A1(n5751), .A2(n6903), .A3(n6650), .ZN(n5937) );
  OAI21_X1 U6437 ( .B1(n7010), .B2(n5937), .A(n6107), .ZN(n6921) );
  INV_X1 U6438 ( .A(n5937), .ZN(n5752) );
  NOR2_X1 U6439 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5752), .ZN(n5753) );
  AND2_X1 U6440 ( .A1(n6994), .A2(n5753), .ZN(n6922) );
  INV_X1 U6441 ( .A(n5754), .ZN(n5849) );
  NOR2_X1 U6442 ( .A1(n6999), .A2(n5849), .ZN(n5756) );
  NOR2_X1 U6443 ( .A1(n4147), .A2(n6998), .ZN(n5755) );
  OR4_X1 U6444 ( .A1(n6922), .A2(n5756), .A3(n5755), .A4(n6974), .ZN(n5761) );
  OR2_X1 U6445 ( .A1(n3475), .A2(n5757), .ZN(n5758) );
  NAND2_X1 U6446 ( .A1(n5841), .A2(n5758), .ZN(n5853) );
  OAI22_X1 U6447 ( .A1(n5759), .A2(n6980), .B1(n7006), .B2(n5853), .ZN(n5760)
         );
  AOI211_X1 U6448 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6921), .A(n5761), .B(n5760), .ZN(n5762) );
  OAI21_X1 U6449 ( .B1(n5763), .B2(n7001), .A(n5762), .ZN(U2815) );
  OAI222_X1 U6450 ( .A1(n6154), .A2(n5853), .B1(n6706), .B2(n4147), .C1(n6156), 
        .C2(n5763), .ZN(U2847) );
  INV_X1 U6451 ( .A(n5833), .ZN(n5779) );
  NAND3_X1 U6452 ( .A1(n5779), .A2(n5764), .A3(n5830), .ZN(n5766) );
  NAND2_X1 U6453 ( .A1(n5766), .A2(n5765), .ZN(n5773) );
  INV_X1 U6454 ( .A(n5774), .ZN(n5769) );
  INV_X1 U6455 ( .A(n5830), .ZN(n5781) );
  NOR2_X1 U6456 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5770), .ZN(n5828)
         );
  AOI211_X1 U6457 ( .C1(n5774), .C2(n5773), .A(n5772), .B(n5771), .ZN(n5775)
         );
  AOI22_X1 U6458 ( .A1(n5776), .A2(n5828), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5827), .ZN(n5777) );
  OAI21_X1 U6459 ( .B1(n5779), .B2(n5778), .A(n5777), .ZN(n5780) );
  AOI21_X1 U6460 ( .B1(n5782), .B2(n5781), .A(n5780), .ZN(n5783) );
  OAI21_X1 U6461 ( .B1(n5835), .B2(n5784), .A(n5783), .ZN(U3107) );
  AOI22_X1 U6462 ( .A1(n5785), .A2(n5828), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5827), .ZN(n5786) );
  OAI21_X1 U6463 ( .B1(n5787), .B2(n5830), .A(n5786), .ZN(n5788) );
  AOI21_X1 U6464 ( .B1(n5833), .B2(n5789), .A(n5788), .ZN(n5790) );
  OAI21_X1 U6465 ( .B1(n5835), .B2(n5791), .A(n5790), .ZN(U3106) );
  AOI22_X1 U6466 ( .A1(n5792), .A2(n5828), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5827), .ZN(n5793) );
  OAI21_X1 U6467 ( .B1(n5794), .B2(n5830), .A(n5793), .ZN(n5795) );
  AOI21_X1 U6468 ( .B1(n5833), .B2(n5796), .A(n5795), .ZN(n5797) );
  OAI21_X1 U6469 ( .B1(n5835), .B2(n5798), .A(n5797), .ZN(U3102) );
  AOI22_X1 U6470 ( .A1(n5799), .A2(n5828), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5827), .ZN(n5800) );
  OAI21_X1 U6471 ( .B1(n5801), .B2(n5830), .A(n5800), .ZN(n5802) );
  AOI21_X1 U6472 ( .B1(n5833), .B2(n5803), .A(n5802), .ZN(n5804) );
  OAI21_X1 U6473 ( .B1(n5835), .B2(n5805), .A(n5804), .ZN(U3103) );
  AOI22_X1 U6474 ( .A1(n5806), .A2(n5828), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5827), .ZN(n5807) );
  OAI21_X1 U6475 ( .B1(n5808), .B2(n5830), .A(n5807), .ZN(n5809) );
  AOI21_X1 U6476 ( .B1(n5833), .B2(n5810), .A(n5809), .ZN(n5811) );
  OAI21_X1 U6477 ( .B1(n5835), .B2(n5812), .A(n5811), .ZN(U3104) );
  AOI22_X1 U6478 ( .A1(n5813), .A2(n5828), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5827), .ZN(n5814) );
  OAI21_X1 U6479 ( .B1(n5815), .B2(n5830), .A(n5814), .ZN(n5816) );
  AOI21_X1 U6480 ( .B1(n5833), .B2(n5817), .A(n5816), .ZN(n5818) );
  OAI21_X1 U6481 ( .B1(n5835), .B2(n5819), .A(n5818), .ZN(U3105) );
  AOI22_X1 U6482 ( .A1(n5820), .A2(n5828), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5827), .ZN(n5821) );
  OAI21_X1 U6483 ( .B1(n5822), .B2(n5830), .A(n5821), .ZN(n5823) );
  AOI21_X1 U6484 ( .B1(n5833), .B2(n5824), .A(n5823), .ZN(n5825) );
  OAI21_X1 U6485 ( .B1(n5835), .B2(n5826), .A(n5825), .ZN(U3101) );
  AOI22_X1 U6486 ( .A1(n7221), .A2(n5828), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5827), .ZN(n5829) );
  OAI21_X1 U6487 ( .B1(n5831), .B2(n5830), .A(n5829), .ZN(n5832) );
  AOI21_X1 U6488 ( .B1(n7223), .B2(n5833), .A(n5832), .ZN(n5834) );
  OAI21_X1 U6489 ( .B1(n5835), .B2(n7227), .A(n5834), .ZN(U3100) );
  OAI21_X1 U6490 ( .B1(n5836), .B2(n5839), .A(n5838), .ZN(n6917) );
  INV_X1 U6491 ( .A(n5872), .ZN(n5840) );
  AOI21_X1 U6492 ( .B1(n5842), .B2(n5841), .A(n5840), .ZN(n6914) );
  AOI22_X1 U6493 ( .A1(n6914), .A2(n6702), .B1(EBX_REG_13__SCAN_IN), .B2(n4769), .ZN(n5843) );
  OAI21_X1 U6494 ( .B1(n6917), .B2(n6156), .A(n5843), .ZN(U2846) );
  NAND2_X1 U6495 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  XNOR2_X1 U6496 ( .A(n5847), .B(n5846), .ZN(n5867) );
  AND2_X1 U6497 ( .A1(n6847), .A2(REIP_REG_12__SCAN_IN), .ZN(n5864) );
  AOI21_X1 U6498 ( .B1(n6749), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5864), 
        .ZN(n5848) );
  OAI21_X1 U6499 ( .B1(n6755), .B2(n5849), .A(n5848), .ZN(n5850) );
  AOI21_X1 U6500 ( .B1(n5851), .B2(n6254), .A(n5850), .ZN(n5852) );
  OAI21_X1 U6501 ( .B1(n5867), .B2(n7033), .A(n5852), .ZN(U2974) );
  INV_X1 U6502 ( .A(n5853), .ZN(n5865) );
  NAND2_X1 U6503 ( .A1(n6378), .A2(n5856), .ZN(n5855) );
  INV_X1 U6504 ( .A(n5859), .ZN(n5854) );
  OR2_X1 U6505 ( .A1(n5878), .A2(n5854), .ZN(n5905) );
  NAND2_X1 U6506 ( .A1(n5855), .A2(n5905), .ZN(n6835) );
  NOR2_X1 U6507 ( .A1(n6350), .A2(n6834), .ZN(n5862) );
  OR2_X1 U6508 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  OAI211_X1 U6509 ( .C1(n5859), .C2(n5878), .A(n6818), .B(n5858), .ZN(n6836)
         );
  AOI221_X1 U6510 ( .B1(n6816), .B2(n6834), .C1(n6378), .C2(n6834), .A(n6836), 
        .ZN(n5860) );
  INV_X1 U6511 ( .A(n5860), .ZN(n5861) );
  MUX2_X1 U6512 ( .A(n5862), .B(n5861), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n5863) );
  AOI211_X1 U6513 ( .C1(n6873), .C2(n5865), .A(n5864), .B(n5863), .ZN(n5866)
         );
  OAI21_X1 U6514 ( .B1(n5867), .B2(n6878), .A(n5866), .ZN(U3006) );
  OAI21_X1 U6515 ( .B1(n5868), .B2(n5870), .A(n5869), .ZN(n5912) );
  AND2_X1 U6516 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  OR2_X1 U6517 ( .A1(n5873), .A2(n5894), .ZN(n6930) );
  INV_X1 U6518 ( .A(n6930), .ZN(n5903) );
  AOI22_X1 U6519 ( .A1(n5903), .A2(n6702), .B1(EBX_REG_14__SCAN_IN), .B2(n4769), .ZN(n5874) );
  OAI21_X1 U6520 ( .B1(n5912), .B2(n6156), .A(n5874), .ZN(U2845) );
  INV_X1 U6521 ( .A(DATAI_13_), .ZN(n5875) );
  INV_X1 U6522 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7189) );
  OAI222_X1 U6523 ( .A1(n6917), .A2(n7201), .B1(n5916), .B2(n5875), .C1(n6015), 
        .C2(n7189), .ZN(U2878) );
  INV_X1 U6524 ( .A(DATAI_14_), .ZN(n6540) );
  INV_X1 U6525 ( .A(EAX_REG_14__SCAN_IN), .ZN(n7195) );
  OAI222_X1 U6526 ( .A1(n5912), .A2(n7201), .B1(n5916), .B2(n6540), .C1(n6015), 
        .C2(n7195), .ZN(U2877) );
  OAI21_X1 U6527 ( .B1(n3444), .B2(n5877), .A(n5876), .ZN(n5886) );
  INV_X1 U6528 ( .A(n5886), .ZN(n5885) );
  NAND2_X1 U6529 ( .A1(n5878), .A2(n5904), .ZN(n6867) );
  AOI21_X1 U6530 ( .B1(n5880), .B2(n6867), .A(n6836), .ZN(n5879) );
  OAI21_X1 U6531 ( .B1(n5900), .B2(n6868), .A(n5879), .ZN(n5907) );
  NOR2_X1 U6532 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5880), .ZN(n5881)
         );
  AOI22_X1 U6533 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5907), .B1(n5881), .B2(n6835), .ZN(n5884) );
  INV_X1 U6534 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5882) );
  NOR2_X1 U6535 ( .A1(n6860), .A2(n5882), .ZN(n5888) );
  AOI21_X1 U6536 ( .B1(n6873), .B2(n6914), .A(n5888), .ZN(n5883) );
  OAI211_X1 U6537 ( .C1(n5885), .C2(n6878), .A(n5884), .B(n5883), .ZN(U3005)
         );
  NAND2_X1 U6538 ( .A1(n5886), .A2(n6751), .ZN(n5890) );
  NOR2_X1 U6539 ( .A1(n6755), .A2(n6918), .ZN(n5887) );
  AOI211_X1 U6540 ( .C1(n6749), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5888), 
        .B(n5887), .ZN(n5889) );
  OAI211_X1 U6541 ( .C1(n6742), .C2(n6917), .A(n5890), .B(n5889), .ZN(U2973)
         );
  INV_X1 U6542 ( .A(n5869), .ZN(n5893) );
  BUF_X1 U6543 ( .A(n5891), .Z(n5892) );
  OAI21_X1 U6544 ( .B1(n5893), .B2(n3493), .A(n5892), .ZN(n6939) );
  AOI21_X1 U6545 ( .B1(n3492), .B2(n3517), .A(n5928), .ZN(n6940) );
  AOI22_X1 U6546 ( .A1(n6940), .A2(n6702), .B1(EBX_REG_15__SCAN_IN), .B2(n4769), .ZN(n5895) );
  OAI21_X1 U6547 ( .B1(n6939), .B2(n6156), .A(n5895), .ZN(U2844) );
  XNOR2_X1 U6548 ( .A(n6369), .B(n5899), .ZN(n5897) );
  XNOR2_X1 U6549 ( .A(n5896), .B(n5897), .ZN(n5915) );
  INV_X1 U6550 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5898) );
  NOR2_X1 U6551 ( .A1(n6860), .A2(n5898), .ZN(n5911) );
  NAND2_X1 U6552 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  NOR2_X1 U6553 ( .A1(n6350), .A2(n5901), .ZN(n5902) );
  AOI211_X1 U6554 ( .C1(n6873), .C2(n5903), .A(n5911), .B(n5902), .ZN(n5909)
         );
  AOI21_X1 U6555 ( .B1(n5905), .B2(n5904), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5906) );
  OAI21_X1 U6556 ( .B1(n5907), .B2(n5906), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5908) );
  OAI211_X1 U6557 ( .C1(n5915), .C2(n6878), .A(n5909), .B(n5908), .ZN(U3004)
         );
  AND2_X1 U6558 ( .A1(n6749), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5910)
         );
  AOI211_X1 U6559 ( .C1(n6933), .C2(n6269), .A(n5911), .B(n5910), .ZN(n5914)
         );
  INV_X1 U6560 ( .A(n5912), .ZN(n6934) );
  NAND2_X1 U6561 ( .A1(n6934), .A2(n6254), .ZN(n5913) );
  OAI211_X1 U6562 ( .C1(n5915), .C2(n7033), .A(n5914), .B(n5913), .ZN(U2972)
         );
  INV_X1 U6563 ( .A(DATAI_15_), .ZN(n6409) );
  INV_X1 U6564 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7200) );
  OAI222_X1 U6565 ( .A1(n6939), .A2(n7201), .B1(n5916), .B2(n6409), .C1(n6015), 
        .C2(n7200), .ZN(U2876) );
  OAI21_X1 U6567 ( .B1(n5917), .B2(n5920), .A(n5919), .ZN(n6262) );
  NAND2_X1 U6568 ( .A1(n5930), .A2(n5921), .ZN(n5922) );
  AND2_X1 U6569 ( .A1(n6152), .A2(n5922), .ZN(n6849) );
  INV_X1 U6570 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5939) );
  NOR2_X1 U6571 ( .A1(n6706), .A2(n5939), .ZN(n5923) );
  AOI21_X1 U6572 ( .B1(n6849), .B2(n6702), .A(n5923), .ZN(n5924) );
  OAI21_X1 U6573 ( .B1(n6262), .B2(n6156), .A(n5924), .ZN(U2842) );
  AND2_X1 U6574 ( .A1(n5892), .A2(n5925), .ZN(n5926) );
  OR2_X1 U6575 ( .A1(n5926), .A2(n5917), .ZN(n6266) );
  INV_X1 U6576 ( .A(n6156), .ZN(n6703) );
  OR2_X1 U6577 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U6578 ( .A1(n5930), .A2(n5929), .ZN(n6958) );
  OAI22_X1 U6579 ( .A1(n6958), .A2(n6154), .B1(n6953), .B2(n6706), .ZN(n5931)
         );
  AOI21_X1 U6580 ( .B1(n7202), .B2(n6703), .A(n5931), .ZN(n5932) );
  INV_X1 U6581 ( .A(n5932), .ZN(U2843) );
  NOR2_X2 U6582 ( .A1(n7235), .A2(n5933), .ZN(n7232) );
  AOI22_X1 U6583 ( .A1(n7232), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n7235), .ZN(n5936) );
  NOR2_X1 U6584 ( .A1(n6016), .A2(n3820), .ZN(n5934) );
  NAND2_X1 U6585 ( .A1(n7236), .A2(DATAI_1_), .ZN(n5935) );
  OAI211_X1 U6586 ( .C1(n6262), .C2(n7201), .A(n5936), .B(n5935), .ZN(U2874)
         );
  NAND3_X1 U6587 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .ZN(n5955) );
  INV_X1 U6588 ( .A(n5955), .ZN(n5938) );
  NAND2_X1 U6589 ( .A1(n5937), .A2(REIP_REG_12__SCAN_IN), .ZN(n6915) );
  NOR2_X1 U6590 ( .A1(n6915), .A2(n5882), .ZN(n6927) );
  NAND2_X1 U6591 ( .A1(n6927), .A2(REIP_REG_14__SCAN_IN), .ZN(n5956) );
  NOR2_X1 U6592 ( .A1(n6116), .A2(n5956), .ZN(n6928) );
  AOI21_X1 U6593 ( .B1(n5938), .B2(n6928), .A(n6929), .ZN(n6968) );
  INV_X1 U6594 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6963) );
  NOR2_X1 U6595 ( .A1(n7010), .A2(n5956), .ZN(n6950) );
  NAND3_X1 U6596 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        n6950), .ZN(n6962) );
  NAND2_X1 U6597 ( .A1(n6963), .A2(n6962), .ZN(n5942) );
  OAI22_X1 U6598 ( .A1(n5940), .A2(n6980), .B1(n5939), .B2(n6998), .ZN(n5941)
         );
  AOI211_X1 U6599 ( .C1(n6968), .C2(n5942), .A(n6974), .B(n5941), .ZN(n5944)
         );
  AOI22_X1 U6600 ( .A1(n7015), .A2(n6849), .B1(n7017), .B2(n6259), .ZN(n5943)
         );
  OAI211_X1 U6601 ( .C1(n6262), .C2(n7001), .A(n5944), .B(n5943), .ZN(U2810)
         );
  XNOR2_X1 U6602 ( .A(n3461), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5946)
         );
  XNOR2_X1 U6603 ( .A(n5945), .B(n5946), .ZN(n6842) );
  NAND2_X1 U6604 ( .A1(n6842), .A2(n6751), .ZN(n5951) );
  INV_X1 U6605 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5947) );
  NOR2_X1 U6606 ( .A1(n6860), .A2(n5947), .ZN(n6840) );
  INV_X1 U6607 ( .A(n6942), .ZN(n5948) );
  NOR2_X1 U6608 ( .A1(n6755), .A2(n5948), .ZN(n5949) );
  AOI211_X1 U6609 ( .C1(n6749), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6840), 
        .B(n5949), .ZN(n5950) );
  OAI211_X1 U6610 ( .C1(n6742), .C2(n6939), .A(n5951), .B(n5950), .ZN(U2971)
         );
  AOI22_X1 U6611 ( .A1(n7232), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n7235), .ZN(n5953) );
  NAND2_X1 U6612 ( .A1(n7236), .A2(DATAI_14_), .ZN(n5952) );
  OAI211_X1 U6613 ( .C1(n5954), .C2(n7201), .A(n5953), .B(n5952), .ZN(U2861)
         );
  NAND2_X1 U6614 ( .A1(n5982), .A2(n7016), .ZN(n5967) );
  INV_X1 U6615 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6678) );
  INV_X1 U6616 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6674) );
  NOR2_X1 U6617 ( .A1(n6678), .A2(n6674), .ZN(n5959) );
  NAND2_X1 U6618 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5958) );
  INV_X1 U6619 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6491) );
  INV_X1 U6620 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6859) );
  INV_X1 U6621 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6605) );
  INV_X1 U6622 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6969) );
  NOR3_X1 U6623 ( .A1(n6969), .A2(n5956), .A3(n5955), .ZN(n5957) );
  NAND3_X1 U6624 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n5957), .ZN(n6109) );
  NOR2_X1 U6625 ( .A1(n6605), .A2(n6109), .ZN(n6993) );
  NAND2_X1 U6626 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6993), .ZN(n6092) );
  NOR2_X1 U6627 ( .A1(n6859), .A2(n6092), .ZN(n7012) );
  NAND2_X1 U6628 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7012), .ZN(n6079) );
  NOR2_X1 U6629 ( .A1(n6491), .A2(n6079), .ZN(n6060) );
  AND2_X1 U6630 ( .A1(n6060), .A2(REIP_REG_26__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U6631 ( .A1(n6107), .A2(n5962), .ZN(n6046) );
  INV_X1 U6632 ( .A(n6929), .ZN(n6047) );
  OAI21_X1 U6633 ( .B1(n5958), .B2(n6046), .A(n6047), .ZN(n6020) );
  OAI21_X1 U6634 ( .B1(n5959), .B2(n7010), .A(n6020), .ZN(n6012) );
  AOI22_X1 U6635 ( .A1(n5977), .A2(n7017), .B1(n7009), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5960) );
  OAI21_X1 U6636 ( .B1(n6998), .B2(n5961), .A(n5960), .ZN(n5965) );
  NAND2_X1 U6637 ( .A1(n6994), .A2(n5962), .ZN(n6049) );
  INV_X1 U6638 ( .A(n6049), .ZN(n5963) );
  NAND3_X1 U6639 ( .A1(n5963), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n6025) );
  NOR3_X1 U6640 ( .A1(n6025), .A2(REIP_REG_30__SCAN_IN), .A3(n6674), .ZN(n5964) );
  AOI211_X1 U6641 ( .C1(REIP_REG_30__SCAN_IN), .C2(n6012), .A(n5965), .B(n5964), .ZN(n5966) );
  OAI211_X1 U6642 ( .C1(n5968), .C2(n7006), .A(n5967), .B(n5966), .ZN(U2797)
         );
  INV_X1 U6643 ( .A(n5999), .ZN(n7041) );
  AND2_X1 U6644 ( .A1(n5969), .A2(n3510), .ZN(n5970) );
  AOI21_X1 U6645 ( .B1(n5972), .B2(n5971), .A(n5970), .ZN(n7051) );
  AOI22_X1 U6646 ( .A1(n3510), .A2(n7087), .B1(n6870), .B2(
        STATE2_REG_1__SCAN_IN), .ZN(n5973) );
  OAI21_X1 U6647 ( .B1(n7051), .B2(n7075), .A(n5973), .ZN(n5975) );
  NOR2_X1 U6648 ( .A1(n5974), .A2(n3510), .ZN(n7048) );
  AOI22_X1 U6649 ( .A1(n7041), .A2(n5975), .B1(n6003), .B2(n7048), .ZN(n5976)
         );
  OAI21_X1 U6650 ( .B1(n3510), .B2(n7041), .A(n5976), .ZN(U3461) );
  INV_X1 U6651 ( .A(n5977), .ZN(n5980) );
  AOI21_X1 U6652 ( .B1(n6749), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5978), 
        .ZN(n5979) );
  OAI21_X1 U6653 ( .B1(n6755), .B2(n5980), .A(n5979), .ZN(n5981) );
  AOI21_X1 U6654 ( .B1(n5982), .B2(n6254), .A(n5981), .ZN(n5983) );
  OAI21_X1 U6655 ( .B1(n5984), .B2(n7033), .A(n5983), .ZN(U2956) );
  NOR2_X1 U6656 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  OR2_X1 U6657 ( .A1(n4894), .A2(n5987), .ZN(n6781) );
  INV_X1 U6658 ( .A(n6781), .ZN(n5997) );
  AOI22_X1 U6659 ( .A1(n6702), .A2(n5997), .B1(EBX_REG_2__SCAN_IN), .B2(n4769), 
        .ZN(n5988) );
  OAI21_X1 U6660 ( .B1(n6722), .B2(n6156), .A(n5988), .ZN(U2857) );
  OAI211_X1 U6661 ( .C1(REIP_REG_1__SCAN_IN), .C2(REIP_REG_2__SCAN_IN), .A(
        n6994), .B(n5989), .ZN(n5991) );
  AOI22_X1 U6662 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7009), .B1(n6116), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n5990) );
  OAI211_X1 U6663 ( .C1(n6727), .C2(n6999), .A(n5991), .B(n5990), .ZN(n5996)
         );
  OAI22_X1 U6664 ( .A1(n6998), .A2(n5994), .B1(n5993), .B2(n5992), .ZN(n5995)
         );
  AOI211_X1 U6665 ( .C1(n7015), .C2(n5997), .A(n5996), .B(n5995), .ZN(n5998)
         );
  OAI21_X1 U6666 ( .B1(n6120), .B2(n6722), .A(n5998), .ZN(U2825) );
  NOR2_X1 U6667 ( .A1(n5999), .A2(n3885), .ZN(n6001) );
  OAI21_X1 U6668 ( .B1(n6001), .B2(n6000), .A(n7087), .ZN(n6005) );
  NAND3_X1 U6669 ( .A1(n7041), .A2(n6003), .A3(n6002), .ZN(n6004) );
  OAI211_X1 U6670 ( .C1(n6006), .C2(n3581), .A(n6005), .B(n6004), .ZN(U3456)
         );
  NAND2_X1 U6671 ( .A1(n6017), .A2(n7016), .ZN(n6014) );
  NAND4_X1 U6672 ( .A1(n6007), .A2(n3821), .A3(EBX_REG_31__SCAN_IN), .A4(n7068), .ZN(n6008) );
  OAI21_X1 U6673 ( .B1(n6980), .B2(n6009), .A(n6008), .ZN(n6011) );
  NOR4_X1 U6674 ( .A1(n6025), .A2(REIP_REG_31__SCAN_IN), .A3(n6678), .A4(n6674), .ZN(n6010) );
  AOI211_X1 U6675 ( .C1(REIP_REG_31__SCAN_IN), .C2(n6012), .A(n6011), .B(n6010), .ZN(n6013) );
  OAI211_X1 U6676 ( .C1(n6128), .C2(n7006), .A(n6014), .B(n6013), .ZN(U2796)
         );
  NAND3_X1 U6677 ( .A1(n6017), .A2(n6016), .A3(n6015), .ZN(n6019) );
  AOI22_X1 U6678 ( .A1(n7232), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7235), .ZN(n6018) );
  NAND2_X1 U6679 ( .A1(n6019), .A2(n6018), .ZN(U2860) );
  NAND2_X1 U6680 ( .A1(n6179), .A2(n7016), .ZN(n6028) );
  INV_X1 U6681 ( .A(n6020), .ZN(n6038) );
  INV_X1 U6682 ( .A(n6021), .ZN(n6177) );
  OAI22_X1 U6683 ( .A1(n6022), .A2(n6980), .B1(n6999), .B2(n6177), .ZN(n6023)
         );
  AOI21_X1 U6684 ( .B1(n7008), .B2(EBX_REG_29__SCAN_IN), .A(n6023), .ZN(n6024)
         );
  OAI21_X1 U6685 ( .B1(n6025), .B2(REIP_REG_29__SCAN_IN), .A(n6024), .ZN(n6026) );
  AOI21_X1 U6686 ( .B1(n6038), .B2(REIP_REG_29__SCAN_IN), .A(n6026), .ZN(n6027) );
  OAI211_X1 U6687 ( .C1(n7006), .C2(n6275), .A(n6028), .B(n6027), .ZN(U2798)
         );
  OAI21_X1 U6688 ( .B1(n6044), .B2(n6030), .A(n6029), .ZN(n6281) );
  AOI21_X1 U6690 ( .B1(n6033), .B2(n6032), .A(n4763), .ZN(n6188) );
  NAND2_X1 U6691 ( .A1(n6188), .A2(n7016), .ZN(n6040) );
  INV_X1 U6692 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6669) );
  NOR3_X1 U6693 ( .A1(n6049), .A2(REIP_REG_28__SCAN_IN), .A3(n6669), .ZN(n6037) );
  INV_X1 U6694 ( .A(n6186), .ZN(n6034) );
  AOI22_X1 U6695 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n7009), .B1(n7017), 
        .B2(n6034), .ZN(n6035) );
  OAI21_X1 U6696 ( .B1(n6998), .B2(n6129), .A(n6035), .ZN(n6036) );
  AOI211_X1 U6697 ( .C1(n6038), .C2(REIP_REG_28__SCAN_IN), .A(n6037), .B(n6036), .ZN(n6039) );
  OAI211_X1 U6698 ( .C1(n7006), .C2(n6281), .A(n6040), .B(n6039), .ZN(U2799)
         );
  BUF_X1 U6699 ( .A(n6041), .Z(n6042) );
  OAI21_X1 U6700 ( .B1(n6042), .B2(n6043), .A(n6032), .ZN(n6192) );
  AOI21_X1 U6701 ( .B1(n6045), .B2(n6056), .A(n6044), .ZN(n6290) );
  NAND2_X1 U6702 ( .A1(n6047), .A2(n6046), .ZN(n6062) );
  AOI22_X1 U6703 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n7009), .B1(
        EBX_REG_27__SCAN_IN), .B2(n7008), .ZN(n6048) );
  OAI221_X1 U6704 ( .B1(REIP_REG_27__SCAN_IN), .B2(n6049), .C1(n6669), .C2(
        n6062), .A(n6048), .ZN(n6052) );
  INV_X1 U6705 ( .A(n6050), .ZN(n6194) );
  NOR2_X1 U6706 ( .A1(n6999), .A2(n6194), .ZN(n6051) );
  AOI211_X1 U6707 ( .C1(n6290), .C2(n7015), .A(n6052), .B(n6051), .ZN(n6053)
         );
  OAI21_X1 U6708 ( .B1(n6192), .B2(n7001), .A(n6053), .ZN(U2800) );
  NAND2_X1 U6709 ( .A1(n6072), .A2(n6054), .ZN(n6055) );
  NAND2_X1 U6710 ( .A1(n6056), .A2(n6055), .ZN(n6297) );
  AOI21_X1 U6711 ( .B1(n6058), .B2(n6057), .A(n6042), .ZN(n6203) );
  NAND2_X1 U6712 ( .A1(n6203), .A2(n7016), .ZN(n6066) );
  OAI22_X1 U6713 ( .A1(n6059), .A2(n6980), .B1(n6999), .B2(n6201), .ZN(n6064)
         );
  AOI21_X1 U6714 ( .B1(n6994), .B2(n6060), .A(REIP_REG_26__SCAN_IN), .ZN(n6061) );
  NOR2_X1 U6715 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  AOI211_X1 U6716 ( .C1(EBX_REG_26__SCAN_IN), .C2(n7008), .A(n6064), .B(n6063), 
        .ZN(n6065) );
  OAI211_X1 U6717 ( .C1(n7006), .C2(n6297), .A(n6066), .B(n6065), .ZN(U2801)
         );
  XOR2_X1 U6718 ( .A(n6068), .B(n6067), .Z(n7234) );
  INV_X1 U6719 ( .A(n7234), .ZN(n6133) );
  INV_X1 U6720 ( .A(n6315), .ZN(n6069) );
  NAND2_X1 U6721 ( .A1(n6316), .A2(n6069), .ZN(n6071) );
  NAND2_X1 U6722 ( .A1(n6071), .A2(n6070), .ZN(n6073) );
  AND2_X1 U6723 ( .A1(n6073), .A2(n6072), .ZN(n6307) );
  INV_X1 U6724 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6664) );
  INV_X1 U6725 ( .A(n7012), .ZN(n6074) );
  NAND2_X1 U6726 ( .A1(n6994), .A2(n6074), .ZN(n6075) );
  NAND2_X1 U6727 ( .A1(n6075), .A2(n6107), .ZN(n7013) );
  AOI21_X1 U6728 ( .B1(n6994), .B2(n6664), .A(n7013), .ZN(n6077) );
  OAI22_X1 U6729 ( .A1(n6077), .A2(n6491), .B1(n6076), .B2(n6980), .ZN(n6083)
         );
  INV_X1 U6730 ( .A(n6078), .ZN(n6208) );
  OR3_X1 U6731 ( .A1(n7010), .A2(REIP_REG_25__SCAN_IN), .A3(n6079), .ZN(n6081)
         );
  NAND2_X1 U6732 ( .A1(n7008), .A2(EBX_REG_25__SCAN_IN), .ZN(n6080) );
  OAI211_X1 U6733 ( .C1(n6208), .C2(n6999), .A(n6081), .B(n6080), .ZN(n6082)
         );
  AOI211_X1 U6734 ( .C1(n6307), .C2(n7015), .A(n6083), .B(n6082), .ZN(n6084)
         );
  OAI21_X1 U6735 ( .B1(n6133), .B2(n7001), .A(n6084), .ZN(U2802) );
  BUF_X1 U6736 ( .A(n6085), .Z(n6086) );
  OAI21_X1 U6737 ( .B1(n6086), .B2(n6088), .A(n6087), .ZN(n6171) );
  INV_X1 U6738 ( .A(n6171), .ZN(n6230) );
  INV_X1 U6739 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6089) );
  OAI22_X1 U6740 ( .A1(n4552), .A2(n6980), .B1(n6089), .B2(n6998), .ZN(n6098)
         );
  NOR2_X1 U6741 ( .A1(n6137), .A2(n6090), .ZN(n6091) );
  OR2_X1 U6742 ( .A1(n6316), .A2(n6091), .ZN(n6855) );
  INV_X1 U6743 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U6744 ( .A1(n6994), .A2(n6093), .ZN(n6094) );
  NAND2_X1 U6745 ( .A1(n6094), .A2(n6859), .ZN(n6095) );
  AOI22_X1 U6746 ( .A1(n7013), .A2(n6095), .B1(n6226), .B2(n7017), .ZN(n6096)
         );
  OAI21_X1 U6747 ( .B1(n6855), .B2(n7006), .A(n6096), .ZN(n6097) );
  AOI211_X1 U6748 ( .C1(n6230), .C2(n7016), .A(n6098), .B(n6097), .ZN(n6099)
         );
  INV_X1 U6749 ( .A(n6099), .ZN(U2804) );
  OAI21_X1 U6751 ( .B1(n6100), .B2(n6103), .A(n6102), .ZN(n6246) );
  NAND2_X1 U6752 ( .A1(n6104), .A2(n6105), .ZN(n6106) );
  AND2_X1 U6753 ( .A1(n6136), .A2(n6106), .ZN(n6336) );
  INV_X1 U6754 ( .A(n6109), .ZN(n6108) );
  OAI21_X1 U6755 ( .B1(n7010), .B2(n6108), .A(n6107), .ZN(n6990) );
  INV_X1 U6756 ( .A(n6990), .ZN(n6113) );
  INV_X1 U6757 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6141) );
  OAI22_X1 U6758 ( .A1(n6241), .A2(n6980), .B1(n6141), .B2(n6998), .ZN(n6111)
         );
  NOR2_X1 U6759 ( .A1(n6109), .A2(REIP_REG_21__SCAN_IN), .ZN(n6110) );
  AND2_X1 U6760 ( .A1(n6994), .A2(n6110), .ZN(n6991) );
  AOI211_X1 U6761 ( .C1(n7017), .C2(n6243), .A(n6111), .B(n6991), .ZN(n6112)
         );
  OAI21_X1 U6762 ( .B1(n6113), .B2(n6605), .A(n6112), .ZN(n6114) );
  AOI21_X1 U6763 ( .B1(n7015), .B2(n6336), .A(n6114), .ZN(n6115) );
  OAI21_X1 U6764 ( .B1(n6246), .B2(n7001), .A(n6115), .ZN(U2806) );
  INV_X1 U6765 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6117) );
  AOI22_X1 U6766 ( .A1(n7017), .A2(n6117), .B1(n6116), .B2(REIP_REG_1__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U6767 ( .A1(n7009), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6118)
         );
  OAI211_X1 U6768 ( .C1(n6120), .C2(n6714), .A(n6119), .B(n6118), .ZN(n6121)
         );
  INV_X1 U6769 ( .A(n6121), .ZN(n6126) );
  AOI22_X1 U6770 ( .A1(n7008), .A2(EBX_REG_1__SCAN_IN), .B1(n6994), .B2(n6690), 
        .ZN(n6125) );
  AOI22_X1 U6771 ( .A1(n6123), .A2(n4811), .B1(n7015), .B2(n6122), .ZN(n6124)
         );
  NAND3_X1 U6772 ( .A1(n6126), .A2(n6125), .A3(n6124), .ZN(U2826) );
  OAI22_X1 U6773 ( .A1(n6128), .A2(n6154), .B1(n6706), .B2(n6127), .ZN(U2828)
         );
  INV_X1 U6774 ( .A(n6188), .ZN(n6163) );
  OAI222_X1 U6775 ( .A1(n6156), .A2(n6163), .B1(n6129), .B2(n6706), .C1(n6281), 
        .C2(n6154), .ZN(U2831) );
  AOI22_X1 U6776 ( .A1(n6290), .A2(n6702), .B1(EBX_REG_27__SCAN_IN), .B2(n4769), .ZN(n6130) );
  OAI21_X1 U6777 ( .B1(n6192), .B2(n6156), .A(n6130), .ZN(U2832) );
  INV_X1 U6778 ( .A(n6203), .ZN(n6168) );
  OAI222_X1 U6779 ( .A1(n6156), .A2(n6168), .B1(n6131), .B2(n6706), .C1(n6297), 
        .C2(n6154), .ZN(U2833) );
  AOI22_X1 U6780 ( .A1(n6307), .A2(n6702), .B1(EBX_REG_25__SCAN_IN), .B2(n4769), .ZN(n6132) );
  OAI21_X1 U6781 ( .B1(n6133), .B2(n6156), .A(n6132), .ZN(U2834) );
  OAI222_X1 U6782 ( .A1(n6156), .A2(n6171), .B1(n6089), .B2(n6706), .C1(n6855), 
        .C2(n6154), .ZN(U2836) );
  AND2_X1 U6783 ( .A1(n6136), .A2(n6135), .ZN(n6138) );
  OR2_X1 U6784 ( .A1(n6138), .A2(n6137), .ZN(n7007) );
  OAI22_X1 U6785 ( .A1(n7007), .A2(n6154), .B1(n6997), .B2(n6706), .ZN(n6139)
         );
  AOI21_X1 U6786 ( .B1(n7214), .B2(n6703), .A(n6139), .ZN(n6140) );
  INV_X1 U6787 ( .A(n6140), .ZN(U2837) );
  NOR2_X1 U6788 ( .A1(n6706), .A2(n6141), .ZN(n6142) );
  AOI21_X1 U6789 ( .B1(n6336), .B2(n6702), .A(n6142), .ZN(n6143) );
  OAI21_X1 U6790 ( .B1(n6246), .B2(n6156), .A(n6143), .ZN(U2838) );
  NOR2_X1 U6791 ( .A1(n3477), .A2(n6144), .ZN(n6145) );
  OR2_X1 U6792 ( .A1(n6100), .A2(n6145), .ZN(n6750) );
  OAI21_X1 U6793 ( .B1(n6357), .B2(n6146), .A(n6104), .ZN(n6989) );
  OAI222_X1 U6794 ( .A1(n6750), .A2(n6156), .B1(n6147), .B2(n6706), .C1(n6154), 
        .C2(n6989), .ZN(U2839) );
  NAND2_X1 U6795 ( .A1(n5919), .A2(n6149), .ZN(n6150) );
  AND2_X1 U6796 ( .A1(n6148), .A2(n6150), .ZN(n7205) );
  INV_X1 U6797 ( .A(n7205), .ZN(n6157) );
  NAND2_X1 U6798 ( .A1(n6152), .A2(n6151), .ZN(n6153) );
  NAND2_X1 U6799 ( .A1(n6358), .A2(n6153), .ZN(n6960) );
  OAI222_X1 U6800 ( .A1(n6157), .A2(n6156), .B1(n6155), .B2(n6706), .C1(n6154), 
        .C2(n6960), .ZN(U2841) );
  AOI22_X1 U6801 ( .A1(n7232), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n7235), .ZN(n6159) );
  NAND2_X1 U6802 ( .A1(n7236), .A2(DATAI_13_), .ZN(n6158) );
  OAI211_X1 U6803 ( .C1(n6160), .C2(n7201), .A(n6159), .B(n6158), .ZN(U2862)
         );
  AOI22_X1 U6804 ( .A1(n7232), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n7235), .ZN(n6162) );
  NAND2_X1 U6805 ( .A1(n7236), .A2(DATAI_12_), .ZN(n6161) );
  OAI211_X1 U6806 ( .C1(n6163), .C2(n7201), .A(n6162), .B(n6161), .ZN(U2863)
         );
  AOI22_X1 U6807 ( .A1(n7232), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n7235), .ZN(n6165) );
  NAND2_X1 U6808 ( .A1(n7236), .A2(DATAI_11_), .ZN(n6164) );
  OAI211_X1 U6809 ( .C1(n6192), .C2(n7201), .A(n6165), .B(n6164), .ZN(U2864)
         );
  AOI22_X1 U6810 ( .A1(n7232), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n7235), .ZN(n6167) );
  NAND2_X1 U6811 ( .A1(n7236), .A2(DATAI_10_), .ZN(n6166) );
  OAI211_X1 U6812 ( .C1(n6168), .C2(n7201), .A(n6167), .B(n6166), .ZN(U2865)
         );
  AOI22_X1 U6813 ( .A1(n7232), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n7235), .ZN(n6170) );
  NAND2_X1 U6814 ( .A1(n7236), .A2(DATAI_7_), .ZN(n6169) );
  OAI211_X1 U6815 ( .C1(n6171), .C2(n7201), .A(n6170), .B(n6169), .ZN(U2868)
         );
  AOI22_X1 U6816 ( .A1(n7232), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n7235), .ZN(n6173) );
  NAND2_X1 U6817 ( .A1(n7236), .A2(DATAI_5_), .ZN(n6172) );
  OAI211_X1 U6818 ( .C1(n6246), .C2(n7201), .A(n6173), .B(n6172), .ZN(U2870)
         );
  AND2_X1 U6819 ( .A1(n6847), .A2(REIP_REG_29__SCAN_IN), .ZN(n6271) );
  AOI21_X1 U6820 ( .B1(n6749), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6271), 
        .ZN(n6176) );
  OAI21_X1 U6821 ( .B1(n6755), .B2(n6177), .A(n6176), .ZN(n6178) );
  AOI21_X1 U6822 ( .B1(n6179), .B2(n6254), .A(n6178), .ZN(n6180) );
  NAND2_X1 U6823 ( .A1(n6182), .A2(n6181), .ZN(n6184) );
  XNOR2_X1 U6824 ( .A(n3461), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6183)
         );
  XNOR2_X1 U6825 ( .A(n6184), .B(n6183), .ZN(n6288) );
  AND2_X1 U6826 ( .A1(n6847), .A2(REIP_REG_28__SCAN_IN), .ZN(n6283) );
  AOI21_X1 U6827 ( .B1(n6749), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6283), 
        .ZN(n6185) );
  OAI21_X1 U6828 ( .B1(n6755), .B2(n6186), .A(n6185), .ZN(n6187) );
  AOI21_X1 U6829 ( .B1(n6188), .B2(n6254), .A(n6187), .ZN(n6189) );
  OAI21_X1 U6830 ( .B1(n6288), .B2(n7033), .A(n6189), .ZN(U2958) );
  NOR2_X1 U6831 ( .A1(n6369), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6190)
         );
  MUX2_X1 U6832 ( .A(n6369), .B(n6190), .S(n3440), .Z(n6191) );
  XNOR2_X1 U6833 ( .A(n6191), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6296)
         );
  INV_X1 U6834 ( .A(n6192), .ZN(n6196) );
  AND2_X1 U6835 ( .A1(n6847), .A2(REIP_REG_27__SCAN_IN), .ZN(n6289) );
  AOI21_X1 U6836 ( .B1(n6749), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6289), 
        .ZN(n6193) );
  OAI21_X1 U6837 ( .B1(n6755), .B2(n6194), .A(n6193), .ZN(n6195) );
  AOI21_X1 U6838 ( .B1(n6196), .B2(n6254), .A(n6195), .ZN(n6197) );
  OAI21_X1 U6839 ( .B1(n6296), .B2(n7033), .A(n6197), .ZN(U2959) );
  XNOR2_X1 U6840 ( .A(n3461), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6199)
         );
  XNOR2_X1 U6841 ( .A(n6198), .B(n6199), .ZN(n6306) );
  AND2_X1 U6842 ( .A1(n6847), .A2(REIP_REG_26__SCAN_IN), .ZN(n6302) );
  AOI21_X1 U6843 ( .B1(n6749), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6302), 
        .ZN(n6200) );
  OAI21_X1 U6844 ( .B1(n6755), .B2(n6201), .A(n6200), .ZN(n6202) );
  AOI21_X1 U6845 ( .B1(n6203), .B2(n6254), .A(n6202), .ZN(n6204) );
  OAI21_X1 U6846 ( .B1(n6306), .B2(n7033), .A(n6204), .ZN(U2960) );
  XNOR2_X1 U6847 ( .A(n6205), .B(n6206), .ZN(n6314) );
  AOI22_X1 U6848 ( .A1(n6749), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n6847), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n6207) );
  OAI21_X1 U6849 ( .B1(n6755), .B2(n6208), .A(n6207), .ZN(n6209) );
  AOI21_X1 U6850 ( .B1(n7234), .B2(n6254), .A(n6209), .ZN(n6210) );
  OAI21_X1 U6851 ( .B1(n6314), .B2(n7033), .A(n6210), .ZN(U2961) );
  NOR2_X1 U6852 ( .A1(n6368), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6340)
         );
  AOI21_X1 U6853 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n6368), .A(n6340), 
        .ZN(n6247) );
  NAND2_X1 U6854 ( .A1(n6211), .A2(n6247), .ZN(n6214) );
  NOR2_X1 U6855 ( .A1(n3461), .A2(n6346), .ZN(n6213) );
  XNOR2_X1 U6856 ( .A(n3461), .B(n6332), .ZN(n6240) );
  NOR2_X1 U6857 ( .A1(n6239), .A2(n6240), .ZN(n6238) );
  AOI21_X1 U6858 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n6368), .A(n6238), 
        .ZN(n6232) );
  NAND3_X1 U6859 ( .A1(n3461), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6216) );
  INV_X1 U6860 ( .A(n6214), .ZN(n6341) );
  NOR4_X1 U6861 ( .A1(n6369), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A4(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n6215) );
  NAND2_X1 U6862 ( .A1(n6341), .A2(n6215), .ZN(n6223) );
  OAI22_X1 U6863 ( .A1(n6232), .A2(n6216), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6223), .ZN(n6217) );
  XNOR2_X1 U6864 ( .A(n6217), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6322)
         );
  AOI21_X1 U6865 ( .B1(n6218), .B2(n6087), .A(n6067), .ZN(n7229) );
  NOR2_X1 U6866 ( .A1(n6860), .A2(n6664), .ZN(n6320) );
  AOI21_X1 U6867 ( .B1(n6749), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6320), 
        .ZN(n6219) );
  OAI21_X1 U6868 ( .B1(n6755), .B2(n6220), .A(n6219), .ZN(n6221) );
  AOI21_X1 U6869 ( .B1(n7229), .B2(n6254), .A(n6221), .ZN(n6222) );
  OAI21_X1 U6870 ( .B1(n6322), .B2(n7033), .A(n6222), .ZN(U2962) );
  OAI21_X1 U6871 ( .B1(n6368), .B2(n6224), .A(n6223), .ZN(n6225) );
  XNOR2_X1 U6872 ( .A(n6225), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6854)
         );
  INV_X1 U6873 ( .A(n6226), .ZN(n6228) );
  AOI22_X1 U6874 ( .A1(n6749), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .B1(n6847), 
        .B2(REIP_REG_23__SCAN_IN), .ZN(n6227) );
  OAI21_X1 U6875 ( .B1(n6755), .B2(n6228), .A(n6227), .ZN(n6229) );
  AOI21_X1 U6876 ( .B1(n6230), .B2(n6254), .A(n6229), .ZN(n6231) );
  OAI21_X1 U6877 ( .B1(n6854), .B2(n7033), .A(n6231), .ZN(U2963) );
  XNOR2_X1 U6878 ( .A(n3461), .B(n6233), .ZN(n6234) );
  XNOR2_X1 U6879 ( .A(n6232), .B(n6234), .ZN(n6329) );
  NAND2_X1 U6880 ( .A1(n6847), .A2(REIP_REG_22__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U6881 ( .A1(n6749), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6235)
         );
  OAI211_X1 U6882 ( .C1(n6755), .C2(n7000), .A(n6325), .B(n6235), .ZN(n6236)
         );
  AOI21_X1 U6883 ( .B1(n7214), .B2(n6254), .A(n6236), .ZN(n6237) );
  OAI21_X1 U6884 ( .B1(n6329), .B2(n7033), .A(n6237), .ZN(U2964) );
  INV_X1 U6885 ( .A(n6238), .ZN(n6331) );
  NAND2_X1 U6886 ( .A1(n6239), .A2(n6240), .ZN(n6330) );
  NAND3_X1 U6887 ( .A1(n6331), .A2(n6751), .A3(n6330), .ZN(n6245) );
  AND2_X1 U6888 ( .A1(n6847), .A2(REIP_REG_21__SCAN_IN), .ZN(n6335) );
  NOR2_X1 U6889 ( .A1(n6710), .A2(n6241), .ZN(n6242) );
  AOI211_X1 U6890 ( .C1(n6269), .C2(n6243), .A(n6335), .B(n6242), .ZN(n6244)
         );
  OAI211_X1 U6891 ( .C1(n6742), .C2(n6246), .A(n6245), .B(n6244), .ZN(U2965)
         );
  INV_X1 U6892 ( .A(n6211), .ZN(n6249) );
  INV_X1 U6893 ( .A(n6247), .ZN(n6248) );
  AOI21_X1 U6894 ( .B1(n6249), .B2(n6248), .A(n6341), .ZN(n6367) );
  XOR2_X1 U6895 ( .A(n6250), .B(n6148), .Z(n7208) );
  NAND2_X1 U6896 ( .A1(n6269), .A2(n6971), .ZN(n6251) );
  NAND2_X1 U6897 ( .A1(n6847), .A2(REIP_REG_19__SCAN_IN), .ZN(n6360) );
  OAI211_X1 U6898 ( .C1(n6710), .C2(n6252), .A(n6251), .B(n6360), .ZN(n6253)
         );
  AOI21_X1 U6899 ( .B1(n7208), .B2(n6254), .A(n6253), .ZN(n6255) );
  OAI21_X1 U6900 ( .B1(n6367), .B2(n7033), .A(n6255), .ZN(U2967) );
  OAI21_X1 U6901 ( .B1(n4157), .B2(n3461), .A(n6256), .ZN(n6372) );
  XNOR2_X1 U6902 ( .A(n6369), .B(n6377), .ZN(n6257) );
  XNOR2_X1 U6903 ( .A(n6372), .B(n6257), .ZN(n6850) );
  NAND2_X1 U6904 ( .A1(n6850), .A2(n6751), .ZN(n6261) );
  OAI22_X1 U6905 ( .A1(n6710), .A2(n5940), .B1(n6860), .B2(n6963), .ZN(n6258)
         );
  AOI21_X1 U6906 ( .B1(n6269), .B2(n6259), .A(n6258), .ZN(n6260) );
  OAI211_X1 U6907 ( .C1(n6742), .C2(n6262), .A(n6261), .B(n6260), .ZN(U2969)
         );
  MUX2_X1 U6908 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n4157), .S(n6369), 
        .Z(n6264) );
  XOR2_X1 U6909 ( .A(n6264), .B(n6263), .Z(n6395) );
  INV_X1 U6910 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U6911 ( .A1(n6847), .A2(REIP_REG_16__SCAN_IN), .ZN(n6391) );
  OAI21_X1 U6912 ( .B1(n6710), .B2(n6265), .A(n6391), .ZN(n6268) );
  NOR2_X1 U6913 ( .A1(n6266), .A2(n6742), .ZN(n6267) );
  AOI211_X1 U6914 ( .C1(n6269), .C2(n6955), .A(n6268), .B(n6267), .ZN(n6270)
         );
  OAI21_X1 U6915 ( .B1(n6395), .B2(n7033), .A(n6270), .ZN(U2970) );
  INV_X1 U6916 ( .A(n6271), .ZN(n6274) );
  INV_X1 U6917 ( .A(n6292), .ZN(n6284) );
  NAND3_X1 U6918 ( .A1(n6284), .A2(n6272), .A3(n4010), .ZN(n6273) );
  OAI211_X1 U6919 ( .C1(n6275), .C2(n6794), .A(n6274), .B(n6273), .ZN(n6276)
         );
  AOI21_X1 U6920 ( .B1(n6277), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n6276), 
        .ZN(n6278) );
  OAI21_X1 U6921 ( .B1(n6279), .B2(n6878), .A(n6278), .ZN(U2989) );
  XNOR2_X1 U6922 ( .A(n6280), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6285)
         );
  NOR2_X1 U6923 ( .A1(n6281), .A2(n6794), .ZN(n6282) );
  AOI211_X1 U6924 ( .C1(n6285), .C2(n6284), .A(n6283), .B(n6282), .ZN(n6287)
         );
  NAND2_X1 U6925 ( .A1(n6294), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6286) );
  OAI211_X1 U6926 ( .C1(n6288), .C2(n6878), .A(n6287), .B(n6286), .ZN(U2990)
         );
  AOI21_X1 U6927 ( .B1(n6290), .B2(n6873), .A(n6289), .ZN(n6291) );
  OAI21_X1 U6928 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6292), .A(n6291), 
        .ZN(n6293) );
  AOI21_X1 U6929 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6294), .A(n6293), 
        .ZN(n6295) );
  OAI21_X1 U6930 ( .B1(n6296), .B2(n6878), .A(n6295), .ZN(U2991) );
  INV_X1 U6931 ( .A(n6297), .ZN(n6303) );
  AOI211_X1 U6932 ( .C1(n6300), .C2(n6299), .A(n6298), .B(n6310), .ZN(n6301)
         );
  AOI211_X1 U6933 ( .C1(n6303), .C2(n6873), .A(n6302), .B(n6301), .ZN(n6305)
         );
  NAND2_X1 U6934 ( .A1(n6312), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6304) );
  OAI211_X1 U6935 ( .C1(n6306), .C2(n6878), .A(n6305), .B(n6304), .ZN(U2992)
         );
  NAND2_X1 U6936 ( .A1(n6307), .A2(n6873), .ZN(n6309) );
  NAND2_X1 U6937 ( .A1(n6847), .A2(REIP_REG_25__SCAN_IN), .ZN(n6308) );
  OAI211_X1 U6938 ( .C1(n6310), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6309), .B(n6308), .ZN(n6311) );
  AOI21_X1 U6939 ( .B1(n6312), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6311), 
        .ZN(n6313) );
  OAI21_X1 U6940 ( .B1(n6314), .B2(n6878), .A(n6313), .ZN(U2993) );
  XNOR2_X1 U6941 ( .A(n6316), .B(n6315), .ZN(n7014) );
  AOI21_X1 U6942 ( .B1(n6864), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6317) );
  NOR2_X1 U6943 ( .A1(n6318), .A2(n6317), .ZN(n6319) );
  AOI211_X1 U6944 ( .C1(n6873), .C2(n7014), .A(n6320), .B(n6319), .ZN(n6321)
         );
  OAI21_X1 U6945 ( .B1(n6322), .B2(n6878), .A(n6321), .ZN(U2994) );
  INV_X1 U6946 ( .A(n6339), .ZN(n6324) );
  NAND3_X1 U6947 ( .A1(n6324), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n6323), .ZN(n6326) );
  OAI211_X1 U6948 ( .C1(n6794), .C2(n7007), .A(n6326), .B(n6325), .ZN(n6327)
         );
  AOI21_X1 U6949 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6862), .A(n6327), 
        .ZN(n6328) );
  OAI21_X1 U6950 ( .B1(n6329), .B2(n6878), .A(n6328), .ZN(U2996) );
  NAND3_X1 U6951 ( .A1(n6331), .A2(n6857), .A3(n6330), .ZN(n6338) );
  NOR2_X1 U6952 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  AOI211_X1 U6953 ( .C1(n6873), .C2(n6336), .A(n6335), .B(n6334), .ZN(n6337)
         );
  OAI211_X1 U6954 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n6339), .A(n6338), .B(n6337), .ZN(U2997) );
  NOR2_X1 U6955 ( .A1(n6341), .A2(n6340), .ZN(n6343) );
  XNOR2_X1 U6956 ( .A(n6369), .B(n6346), .ZN(n6342) );
  XNOR2_X1 U6957 ( .A(n6343), .B(n6342), .ZN(n6752) );
  INV_X1 U6958 ( .A(n6752), .ZN(n6356) );
  INV_X1 U6959 ( .A(n6989), .ZN(n6348) );
  NOR2_X1 U6960 ( .A1(n6345), .A2(n6344), .ZN(n6362) );
  INV_X1 U6961 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6983) );
  OAI22_X1 U6962 ( .A1(n6362), .A2(n6346), .B1(n6860), .B2(n6983), .ZN(n6347)
         );
  AOI21_X1 U6963 ( .B1(n6873), .B2(n6348), .A(n6347), .ZN(n6355) );
  INV_X1 U6964 ( .A(n6349), .ZN(n6388) );
  NOR2_X1 U6965 ( .A1(n6350), .A2(n6386), .ZN(n6841) );
  NAND2_X1 U6966 ( .A1(n6388), .A2(n6841), .ZN(n6853) );
  NOR2_X1 U6967 ( .A1(n6853), .A2(n6351), .ZN(n6365) );
  NAND3_X1 U6968 ( .A1(n6365), .A2(n6353), .A3(n6352), .ZN(n6354) );
  OAI211_X1 U6969 ( .C1(n6356), .C2(n6878), .A(n6355), .B(n6354), .ZN(U2998)
         );
  AOI21_X1 U6970 ( .B1(n6359), .B2(n6358), .A(n6357), .ZN(n6975) );
  NAND2_X1 U6971 ( .A1(n6975), .A2(n6873), .ZN(n6361) );
  OAI211_X1 U6972 ( .C1(n6362), .C2(n6364), .A(n6361), .B(n6360), .ZN(n6363)
         );
  AOI21_X1 U6973 ( .B1(n6365), .B2(n6364), .A(n6363), .ZN(n6366) );
  OAI21_X1 U6974 ( .B1(n6367), .B2(n6878), .A(n6366), .ZN(U2999) );
  NAND2_X1 U6975 ( .A1(n6368), .A2(n6377), .ZN(n6371) );
  NAND2_X1 U6976 ( .A1(n3461), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6370) );
  OAI22_X1 U6977 ( .A1(n6372), .A2(n6371), .B1(n6256), .B2(n6370), .ZN(n6373)
         );
  XNOR2_X1 U6978 ( .A(n6373), .B(n6379), .ZN(n6746) );
  INV_X1 U6979 ( .A(n6746), .ZN(n6385) );
  INV_X1 U6980 ( .A(n6960), .ZN(n6383) );
  NOR3_X1 U6981 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6377), .A3(n6853), 
        .ZN(n6382) );
  AOI22_X1 U6982 ( .A1(n6816), .A2(n6375), .B1(n6814), .B2(n6374), .ZN(n6376)
         );
  NAND2_X1 U6983 ( .A1(n6818), .A2(n6376), .ZN(n6848) );
  AOI21_X1 U6984 ( .B1(n6378), .B2(n6377), .A(n6848), .ZN(n6380) );
  OAI22_X1 U6985 ( .A1(n6380), .A2(n6379), .B1(n6860), .B2(n6969), .ZN(n6381)
         );
  AOI211_X1 U6986 ( .C1(n6873), .C2(n6383), .A(n6382), .B(n6381), .ZN(n6384)
         );
  OAI21_X1 U6987 ( .B1(n6385), .B2(n6878), .A(n6384), .ZN(U3000) );
  AND2_X1 U6988 ( .A1(n6790), .A2(n6386), .ZN(n6387) );
  NOR2_X1 U6989 ( .A1(n6836), .A2(n6387), .ZN(n6846) );
  INV_X1 U6990 ( .A(n6846), .ZN(n6393) );
  AOI21_X1 U6991 ( .B1(n4157), .B2(n6845), .A(n6388), .ZN(n6389) );
  NAND2_X1 U6992 ( .A1(n6389), .A2(n6841), .ZN(n6390) );
  OAI211_X1 U6993 ( .C1(n6958), .C2(n6794), .A(n6391), .B(n6390), .ZN(n6392)
         );
  AOI21_X1 U6994 ( .B1(n6393), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6392), 
        .ZN(n6394) );
  OAI21_X1 U6995 ( .B1(n6395), .B2(n6878), .A(n6394), .ZN(U3002) );
  INV_X1 U6996 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6396) );
  AOI21_X1 U6997 ( .B1(n6396), .B2(STATE_REG_1__SCAN_IN), .A(n7105), .ZN(n6401) );
  INV_X1 U6998 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6397) );
  INV_X1 U6999 ( .A(BS16_N), .ZN(n6569) );
  NAND2_X1 U7000 ( .A1(n6396), .A2(n7105), .ZN(n6762) );
  AOI21_X1 U7001 ( .B1(n6569), .B2(n6762), .A(n6398), .ZN(n7098) );
  AOI21_X1 U7002 ( .B1(n6398), .B2(n6397), .A(n7098), .ZN(U3451) );
  AND2_X1 U7003 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6398), .ZN(U3180) );
  AND2_X1 U7004 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6398), .ZN(U3179) );
  AND2_X1 U7005 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6398), .ZN(U3178) );
  AND2_X1 U7006 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6398), .ZN(U3177) );
  AND2_X1 U7007 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6398), .ZN(U3176) );
  AND2_X1 U7008 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6398), .ZN(U3175) );
  AND2_X1 U7009 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6398), .ZN(U3174) );
  AND2_X1 U7010 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6398), .ZN(U3173) );
  AND2_X1 U7011 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6398), .ZN(U3172) );
  AND2_X1 U7012 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6398), .ZN(U3170) );
  AND2_X1 U7013 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6398), .ZN(U3169) );
  AND2_X1 U7014 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6398), .ZN(U3168) );
  AND2_X1 U7015 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6398), .ZN(U3167) );
  AND2_X1 U7016 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6398), .ZN(U3166) );
  AND2_X1 U7017 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6398), .ZN(U3165) );
  AND2_X1 U7018 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6398), .ZN(U3164) );
  AND2_X1 U7019 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6398), .ZN(U3163) );
  AND2_X1 U7020 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6398), .ZN(U3162) );
  AND2_X1 U7021 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6398), .ZN(U3161) );
  AND2_X1 U7022 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6398), .ZN(U3160) );
  AND2_X1 U7023 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6398), .ZN(U3159) );
  AND2_X1 U7024 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6398), .ZN(U3158) );
  AND2_X1 U7025 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6398), .ZN(U3157) );
  AND2_X1 U7026 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6398), .ZN(U3156) );
  AND2_X1 U7027 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6398), .ZN(U3155) );
  AND2_X1 U7028 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6398), .ZN(U3154) );
  AND2_X1 U7029 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6398), .ZN(U3153) );
  AND2_X1 U7030 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6398), .ZN(U3152) );
  AND2_X1 U7031 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6398), .ZN(U3151) );
  AND2_X1 U7032 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6399), .ZN(U3019)
         );
  AND2_X1 U7033 ( .A1(n6620), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7034 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6400) );
  AOI21_X1 U7035 ( .B1(n6401), .B2(n6400), .A(n7116), .ZN(U2789) );
  NAND2_X1 U7036 ( .A1(n6398), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6612) );
  OAI22_X1 U7037 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput_126), .B1(
        keyinput_127), .B2(REIP_REG_19__SCAN_IN), .ZN(n6402) );
  AOI221_X1 U7038 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_126), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput_127), .A(n6402), .ZN(n6610) );
  INV_X1 U7039 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6992) );
  OAI22_X1 U7040 ( .A1(n6992), .A2(keyinput_124), .B1(keyinput_123), .B2(
        REIP_REG_23__SCAN_IN), .ZN(n6403) );
  AOI221_X1 U7041 ( .B1(n6992), .B2(keyinput_124), .C1(REIP_REG_23__SCAN_IN), 
        .C2(keyinput_123), .A(n6403), .ZN(n6493) );
  OAI22_X1 U7042 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_116), .B1(
        keyinput_117), .B2(REIP_REG_29__SCAN_IN), .ZN(n6404) );
  AOI221_X1 U7043 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_116), .C1(
        REIP_REG_29__SCAN_IN), .C2(keyinput_117), .A(n6404), .ZN(n6486) );
  XNOR2_X1 U7044 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_104), .ZN(n6468) );
  INV_X1 U7045 ( .A(keyinput_103), .ZN(n6466) );
  INV_X1 U7046 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6577) );
  OAI22_X1 U7047 ( .A1(HOLD), .A2(keyinput_100), .B1(keyinput_101), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n6405) );
  AOI221_X1 U7048 ( .B1(HOLD), .B2(keyinput_100), .C1(READREQUEST_REG_SCAN_IN), 
        .C2(keyinput_101), .A(n6405), .ZN(n6463) );
  INV_X1 U7049 ( .A(keyinput_99), .ZN(n6461) );
  INV_X1 U7050 ( .A(keyinput_98), .ZN(n6459) );
  INV_X1 U7051 ( .A(NA_N), .ZN(n7107) );
  INV_X1 U7052 ( .A(keyinput_97), .ZN(n6457) );
  AOI22_X1 U7053 ( .A1(n6507), .A2(keyinput_89), .B1(n6506), .B2(keyinput_88), 
        .ZN(n6406) );
  OAI221_X1 U7054 ( .B1(n6507), .B2(keyinput_89), .C1(n6506), .C2(keyinput_88), 
        .A(n6406), .ZN(n6446) );
  INV_X1 U7055 ( .A(keyinput_87), .ZN(n6443) );
  INV_X1 U7056 ( .A(keyinput_86), .ZN(n6441) );
  INV_X1 U7057 ( .A(keyinput_85), .ZN(n6439) );
  OAI22_X1 U7058 ( .A1(n6509), .A2(keyinput_83), .B1(DATAI_13_), .B2(
        keyinput_82), .ZN(n6407) );
  AOI221_X1 U7059 ( .B1(n6509), .B2(keyinput_83), .C1(keyinput_82), .C2(
        DATAI_13_), .A(n6407), .ZN(n6436) );
  INV_X1 U7060 ( .A(DATAI_16_), .ZN(n6410) );
  AOI22_X1 U7061 ( .A1(n6410), .A2(keyinput_79), .B1(keyinput_80), .B2(n6409), 
        .ZN(n6408) );
  OAI221_X1 U7062 ( .B1(n6410), .B2(keyinput_79), .C1(n6409), .C2(keyinput_80), 
        .A(n6408), .ZN(n6434) );
  INV_X1 U7063 ( .A(keyinput_78), .ZN(n6431) );
  INV_X1 U7064 ( .A(DATAI_17_), .ZN(n6535) );
  INV_X1 U7065 ( .A(DATAI_18_), .ZN(n6529) );
  OAI22_X1 U7066 ( .A1(n6529), .A2(keyinput_77), .B1(keyinput_75), .B2(
        DATAI_20_), .ZN(n6411) );
  AOI221_X1 U7067 ( .B1(n6529), .B2(keyinput_77), .C1(DATAI_20_), .C2(
        keyinput_75), .A(n6411), .ZN(n6428) );
  INV_X1 U7068 ( .A(DATAI_27_), .ZN(n6417) );
  INV_X1 U7069 ( .A(DATAI_29_), .ZN(n6514) );
  INV_X1 U7070 ( .A(DATAI_28_), .ZN(n6515) );
  AOI22_X1 U7071 ( .A1(n6514), .A2(keyinput_66), .B1(keyinput_67), .B2(n6515), 
        .ZN(n6412) );
  OAI221_X1 U7072 ( .B1(n6514), .B2(keyinput_66), .C1(n6515), .C2(keyinput_67), 
        .A(n6412), .ZN(n6415) );
  OAI22_X1 U7073 ( .A1(DATAI_31_), .A2(keyinput_64), .B1(DATAI_30_), .B2(
        keyinput_65), .ZN(n6413) );
  AOI221_X1 U7074 ( .B1(DATAI_31_), .B2(keyinput_64), .C1(keyinput_65), .C2(
        DATAI_30_), .A(n6413), .ZN(n6414) );
  OAI22_X1 U7075 ( .A1(keyinput_68), .A2(n6417), .B1(n6415), .B2(n6414), .ZN(
        n6416) );
  AOI21_X1 U7076 ( .B1(keyinput_68), .B2(n6417), .A(n6416), .ZN(n6426) );
  INV_X1 U7077 ( .A(DATAI_25_), .ZN(n6419) );
  INV_X1 U7078 ( .A(DATAI_26_), .ZN(n6512) );
  AOI22_X1 U7079 ( .A1(n6419), .A2(keyinput_70), .B1(n6512), .B2(keyinput_69), 
        .ZN(n6418) );
  OAI221_X1 U7080 ( .B1(n6419), .B2(keyinput_70), .C1(n6512), .C2(keyinput_69), 
        .A(n6418), .ZN(n6425) );
  INV_X1 U7081 ( .A(DATAI_24_), .ZN(n6521) );
  INV_X1 U7082 ( .A(DATAI_22_), .ZN(n6522) );
  OAI22_X1 U7083 ( .A1(n6521), .A2(keyinput_71), .B1(n6522), .B2(keyinput_73), 
        .ZN(n6420) );
  AOI221_X1 U7084 ( .B1(n6521), .B2(keyinput_71), .C1(keyinput_73), .C2(n6522), 
        .A(n6420), .ZN(n6424) );
  INV_X1 U7085 ( .A(DATAI_23_), .ZN(n6422) );
  OAI22_X1 U7086 ( .A1(n6422), .A2(keyinput_72), .B1(DATAI_21_), .B2(
        keyinput_74), .ZN(n6421) );
  AOI221_X1 U7087 ( .B1(n6422), .B2(keyinput_72), .C1(keyinput_74), .C2(
        DATAI_21_), .A(n6421), .ZN(n6423) );
  OAI211_X1 U7088 ( .C1(n6426), .C2(n6425), .A(n6424), .B(n6423), .ZN(n6427)
         );
  OAI211_X1 U7089 ( .C1(DATAI_19_), .C2(keyinput_76), .A(n6428), .B(n6427), 
        .ZN(n6429) );
  AOI21_X1 U7090 ( .B1(DATAI_19_), .B2(keyinput_76), .A(n6429), .ZN(n6430) );
  AOI221_X1 U7091 ( .B1(DATAI_17_), .B2(n6431), .C1(n6535), .C2(keyinput_78), 
        .A(n6430), .ZN(n6433) );
  NAND2_X1 U7092 ( .A1(n6540), .A2(keyinput_81), .ZN(n6432) );
  OAI221_X1 U7093 ( .B1(n6434), .B2(n6433), .C1(n6540), .C2(keyinput_81), .A(
        n6432), .ZN(n6435) );
  OAI211_X1 U7094 ( .C1(n6544), .C2(keyinput_84), .A(n6436), .B(n6435), .ZN(
        n6437) );
  AOI21_X1 U7095 ( .B1(n6544), .B2(keyinput_84), .A(n6437), .ZN(n6438) );
  AOI221_X1 U7096 ( .B1(DATAI_10_), .B2(n6439), .C1(n6546), .C2(keyinput_85), 
        .A(n6438), .ZN(n6440) );
  AOI221_X1 U7097 ( .B1(DATAI_9_), .B2(keyinput_86), .C1(n6550), .C2(n6441), 
        .A(n6440), .ZN(n6442) );
  AOI221_X1 U7098 ( .B1(DATAI_8_), .B2(keyinput_87), .C1(n6552), .C2(n6443), 
        .A(n6442), .ZN(n6445) );
  NAND2_X1 U7099 ( .A1(keyinput_90), .A2(DATAI_5_), .ZN(n6444) );
  OAI221_X1 U7100 ( .B1(n6446), .B2(n6445), .C1(keyinput_90), .C2(DATAI_5_), 
        .A(n6444), .ZN(n6455) );
  AOI22_X1 U7101 ( .A1(DATAI_3_), .A2(keyinput_92), .B1(n6448), .B2(
        keyinput_91), .ZN(n6447) );
  OAI221_X1 U7102 ( .B1(DATAI_3_), .B2(keyinput_92), .C1(n6448), .C2(
        keyinput_91), .A(n6447), .ZN(n6454) );
  OAI22_X1 U7103 ( .A1(n6450), .A2(keyinput_93), .B1(n6558), .B2(keyinput_94), 
        .ZN(n6449) );
  AOI221_X1 U7104 ( .B1(n6450), .B2(keyinput_93), .C1(keyinput_94), .C2(n6558), 
        .A(n6449), .ZN(n6453) );
  OAI22_X1 U7105 ( .A1(DATAI_0_), .A2(keyinput_95), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_96), .ZN(n6451) );
  AOI221_X1 U7106 ( .B1(DATAI_0_), .B2(keyinput_95), .C1(keyinput_96), .C2(
        MEMORYFETCH_REG_SCAN_IN), .A(n6451), .ZN(n6452) );
  OAI211_X1 U7107 ( .C1(n6455), .C2(n6454), .A(n6453), .B(n6452), .ZN(n6456)
         );
  OAI221_X1 U7108 ( .B1(NA_N), .B2(keyinput_97), .C1(n7107), .C2(n6457), .A(
        n6456), .ZN(n6458) );
  OAI221_X1 U7109 ( .B1(BS16_N), .B2(n6459), .C1(n6569), .C2(keyinput_98), .A(
        n6458), .ZN(n6460) );
  OAI221_X1 U7110 ( .B1(READY_N), .B2(n6461), .C1(n7124), .C2(keyinput_99), 
        .A(n6460), .ZN(n6462) );
  AOI22_X1 U7111 ( .A1(n6463), .A2(n6462), .B1(keyinput_102), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n6464) );
  OAI21_X1 U7112 ( .B1(keyinput_102), .B2(ADS_N_REG_SCAN_IN), .A(n6464), .ZN(
        n6465) );
  OAI221_X1 U7113 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6466), .C1(n6577), .C2(
        keyinput_103), .A(n6465), .ZN(n6467) );
  AOI22_X1 U7114 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_105), .B1(n6468), .B2(
        n6467), .ZN(n6471) );
  INV_X1 U7115 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6764) );
  AOI22_X1 U7116 ( .A1(n6764), .A2(keyinput_106), .B1(n6581), .B2(keyinput_107), .ZN(n6469) );
  OAI221_X1 U7117 ( .B1(n6764), .B2(keyinput_106), .C1(n6581), .C2(
        keyinput_107), .A(n6469), .ZN(n6470) );
  AOI221_X1 U7118 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6471), .C1(keyinput_105), 
        .C2(n6471), .A(n6470), .ZN(n6477) );
  OAI22_X1 U7119 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_109), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_108), .ZN(n6472) );
  AOI221_X1 U7120 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_109), .C1(
        keyinput_108), .C2(MORE_REG_SCAN_IN), .A(n6472), .ZN(n6476) );
  XOR2_X1 U7121 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_110), .Z(n6475) );
  AOI22_X1 U7122 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_111), .B1(
        BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_112), .ZN(n6473) );
  OAI221_X1 U7123 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_111), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_112), .A(n6473), .ZN(n6474)
         );
  AOI211_X1 U7124 ( .C1(n6477), .C2(n6476), .A(n6475), .B(n6474), .ZN(n6480)
         );
  INV_X1 U7125 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6498) );
  AOI22_X1 U7126 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_113), .B1(
        n6498), .B2(keyinput_114), .ZN(n6478) );
  OAI221_X1 U7127 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_113), .C1(
        n6498), .C2(keyinput_114), .A(n6478), .ZN(n6479) );
  AOI211_X1 U7128 ( .C1(REIP_REG_31__SCAN_IN), .C2(keyinput_115), .A(n6480), 
        .B(n6479), .ZN(n6481) );
  OAI21_X1 U7129 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_115), .A(n6481), 
        .ZN(n6485) );
  INV_X1 U7130 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6483) );
  AOI22_X1 U7131 ( .A1(n6483), .A2(keyinput_118), .B1(keyinput_119), .B2(n6669), .ZN(n6482) );
  OAI221_X1 U7132 ( .B1(n6483), .B2(keyinput_118), .C1(n6669), .C2(
        keyinput_119), .A(n6482), .ZN(n6484) );
  AOI21_X1 U7133 ( .B1(n6486), .B2(n6485), .A(n6484), .ZN(n6489) );
  INV_X1 U7134 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6667) );
  AOI22_X1 U7135 ( .A1(n6667), .A2(keyinput_120), .B1(n6664), .B2(keyinput_122), .ZN(n6487) );
  OAI221_X1 U7136 ( .B1(n6667), .B2(keyinput_120), .C1(n6664), .C2(
        keyinput_122), .A(n6487), .ZN(n6488) );
  AOI211_X1 U7137 ( .C1(n6491), .C2(keyinput_121), .A(n6489), .B(n6488), .ZN(
        n6490) );
  OAI21_X1 U7138 ( .B1(n6491), .B2(keyinput_121), .A(n6490), .ZN(n6492) );
  AOI22_X1 U7139 ( .A1(n6493), .A2(n6492), .B1(keyinput_125), .B2(
        REIP_REG_21__SCAN_IN), .ZN(n6494) );
  OAI21_X1 U7140 ( .B1(keyinput_125), .B2(REIP_REG_21__SCAN_IN), .A(n6494), 
        .ZN(n6609) );
  AOI22_X1 U7141 ( .A1(n6859), .A2(keyinput_59), .B1(n6992), .B2(keyinput_60), 
        .ZN(n6495) );
  OAI221_X1 U7142 ( .B1(n6859), .B2(keyinput_59), .C1(n6992), .C2(keyinput_60), 
        .A(n6495), .ZN(n6603) );
  OAI22_X1 U7143 ( .A1(n6667), .A2(keyinput_56), .B1(keyinput_57), .B2(
        REIP_REG_25__SCAN_IN), .ZN(n6496) );
  AOI221_X1 U7144 ( .B1(n6667), .B2(keyinput_56), .C1(REIP_REG_25__SCAN_IN), 
        .C2(keyinput_57), .A(n6496), .ZN(n6600) );
  INV_X1 U7145 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6693) );
  INV_X1 U7146 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6499) );
  OAI22_X1 U7147 ( .A1(n6499), .A2(keyinput_51), .B1(n6498), .B2(keyinput_50), 
        .ZN(n6497) );
  AOI221_X1 U7148 ( .B1(n6499), .B2(keyinput_51), .C1(keyinput_50), .C2(n6498), 
        .A(n6497), .ZN(n6592) );
  XOR2_X1 U7149 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_41), .Z(n6586) );
  INV_X1 U7150 ( .A(keyinput_40), .ZN(n6579) );
  INV_X1 U7151 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7114) );
  INV_X1 U7152 ( .A(keyinput_39), .ZN(n6576) );
  INV_X1 U7153 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6501) );
  OAI22_X1 U7154 ( .A1(n6501), .A2(keyinput_37), .B1(HOLD), .B2(keyinput_36), 
        .ZN(n6500) );
  AOI221_X1 U7155 ( .B1(n6501), .B2(keyinput_37), .C1(keyinput_36), .C2(HOLD), 
        .A(n6500), .ZN(n6573) );
  INV_X1 U7156 ( .A(keyinput_35), .ZN(n6571) );
  INV_X1 U7157 ( .A(keyinput_34), .ZN(n6568) );
  INV_X1 U7158 ( .A(keyinput_33), .ZN(n6566) );
  AOI22_X1 U7159 ( .A1(n6504), .A2(keyinput_26), .B1(keyinput_28), .B2(n6503), 
        .ZN(n6502) );
  OAI221_X1 U7160 ( .B1(n6504), .B2(keyinput_26), .C1(n6503), .C2(keyinput_28), 
        .A(n6502), .ZN(n6564) );
  AOI22_X1 U7161 ( .A1(n6507), .A2(keyinput_25), .B1(n6506), .B2(keyinput_24), 
        .ZN(n6505) );
  OAI221_X1 U7162 ( .B1(n6507), .B2(keyinput_25), .C1(n6506), .C2(keyinput_24), 
        .A(n6505), .ZN(n6556) );
  INV_X1 U7163 ( .A(keyinput_23), .ZN(n6553) );
  INV_X1 U7164 ( .A(keyinput_22), .ZN(n6549) );
  INV_X1 U7165 ( .A(keyinput_21), .ZN(n6547) );
  OAI22_X1 U7166 ( .A1(n6509), .A2(keyinput_19), .B1(DATAI_13_), .B2(
        keyinput_18), .ZN(n6508) );
  AOI221_X1 U7167 ( .B1(n6509), .B2(keyinput_19), .C1(keyinput_18), .C2(
        DATAI_13_), .A(n6508), .ZN(n6542) );
  OAI22_X1 U7168 ( .A1(DATAI_16_), .A2(keyinput_15), .B1(DATAI_15_), .B2(
        keyinput_16), .ZN(n6510) );
  AOI221_X1 U7169 ( .B1(DATAI_16_), .B2(keyinput_15), .C1(keyinput_16), .C2(
        DATAI_15_), .A(n6510), .ZN(n6538) );
  INV_X1 U7170 ( .A(keyinput_14), .ZN(n6536) );
  OAI22_X1 U7171 ( .A1(n6512), .A2(keyinput_5), .B1(keyinput_6), .B2(DATAI_25_), .ZN(n6511) );
  AOI221_X1 U7172 ( .B1(n6512), .B2(keyinput_5), .C1(DATAI_25_), .C2(
        keyinput_6), .A(n6511), .ZN(n6527) );
  AOI22_X1 U7173 ( .A1(n6515), .A2(keyinput_3), .B1(n6514), .B2(keyinput_2), 
        .ZN(n6513) );
  OAI221_X1 U7174 ( .B1(n6515), .B2(keyinput_3), .C1(n6514), .C2(keyinput_2), 
        .A(n6513), .ZN(n6519) );
  OAI22_X1 U7175 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(DATAI_30_), .B2(
        keyinput_1), .ZN(n6516) );
  AOI221_X1 U7176 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(keyinput_1), .C2(
        DATAI_30_), .A(n6516), .ZN(n6518) );
  NAND2_X1 U7177 ( .A1(DATAI_27_), .A2(keyinput_4), .ZN(n6517) );
  OAI221_X1 U7178 ( .B1(n6519), .B2(n6518), .C1(DATAI_27_), .C2(keyinput_4), 
        .A(n6517), .ZN(n6526) );
  AOI22_X1 U7179 ( .A1(n6522), .A2(keyinput_9), .B1(n6521), .B2(keyinput_7), 
        .ZN(n6520) );
  OAI221_X1 U7180 ( .B1(n6522), .B2(keyinput_9), .C1(n6521), .C2(keyinput_7), 
        .A(n6520), .ZN(n6525) );
  AOI22_X1 U7181 ( .A1(DATAI_21_), .A2(keyinput_10), .B1(DATAI_23_), .B2(
        keyinput_8), .ZN(n6523) );
  OAI221_X1 U7182 ( .B1(DATAI_21_), .B2(keyinput_10), .C1(DATAI_23_), .C2(
        keyinput_8), .A(n6523), .ZN(n6524) );
  AOI211_X1 U7183 ( .C1(n6527), .C2(n6526), .A(n6525), .B(n6524), .ZN(n6532)
         );
  INV_X1 U7184 ( .A(DATAI_19_), .ZN(n6530) );
  AOI22_X1 U7185 ( .A1(n6530), .A2(keyinput_12), .B1(keyinput_13), .B2(n6529), 
        .ZN(n6528) );
  OAI221_X1 U7186 ( .B1(n6530), .B2(keyinput_12), .C1(n6529), .C2(keyinput_13), 
        .A(n6528), .ZN(n6531) );
  AOI211_X1 U7187 ( .C1(DATAI_20_), .C2(keyinput_11), .A(n6532), .B(n6531), 
        .ZN(n6533) );
  OAI21_X1 U7188 ( .B1(DATAI_20_), .B2(keyinput_11), .A(n6533), .ZN(n6534) );
  OAI221_X1 U7189 ( .B1(DATAI_17_), .B2(n6536), .C1(n6535), .C2(keyinput_14), 
        .A(n6534), .ZN(n6537) );
  AOI22_X1 U7190 ( .A1(keyinput_17), .A2(n6540), .B1(n6538), .B2(n6537), .ZN(
        n6539) );
  OAI21_X1 U7191 ( .B1(n6540), .B2(keyinput_17), .A(n6539), .ZN(n6541) );
  OAI211_X1 U7192 ( .C1(n6544), .C2(keyinput_20), .A(n6542), .B(n6541), .ZN(
        n6543) );
  AOI21_X1 U7193 ( .B1(n6544), .B2(keyinput_20), .A(n6543), .ZN(n6545) );
  AOI221_X1 U7194 ( .B1(DATAI_10_), .B2(n6547), .C1(n6546), .C2(keyinput_21), 
        .A(n6545), .ZN(n6548) );
  AOI221_X1 U7195 ( .B1(DATAI_9_), .B2(keyinput_22), .C1(n6550), .C2(n6549), 
        .A(n6548), .ZN(n6551) );
  AOI221_X1 U7196 ( .B1(DATAI_8_), .B2(n6553), .C1(n6552), .C2(keyinput_23), 
        .A(n6551), .ZN(n6555) );
  NAND2_X1 U7197 ( .A1(keyinput_27), .A2(DATAI_4_), .ZN(n6554) );
  OAI221_X1 U7198 ( .B1(n6556), .B2(n6555), .C1(keyinput_27), .C2(DATAI_4_), 
        .A(n6554), .ZN(n6563) );
  INV_X1 U7199 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7115) );
  OAI22_X1 U7200 ( .A1(n6558), .A2(keyinput_30), .B1(n7115), .B2(keyinput_32), 
        .ZN(n6557) );
  AOI221_X1 U7201 ( .B1(n6558), .B2(keyinput_30), .C1(keyinput_32), .C2(n7115), 
        .A(n6557), .ZN(n6562) );
  OAI22_X1 U7202 ( .A1(n6560), .A2(keyinput_31), .B1(DATAI_2_), .B2(
        keyinput_29), .ZN(n6559) );
  AOI221_X1 U7203 ( .B1(n6560), .B2(keyinput_31), .C1(keyinput_29), .C2(
        DATAI_2_), .A(n6559), .ZN(n6561) );
  OAI211_X1 U7204 ( .C1(n6564), .C2(n6563), .A(n6562), .B(n6561), .ZN(n6565)
         );
  OAI221_X1 U7205 ( .B1(NA_N), .B2(keyinput_33), .C1(n7107), .C2(n6566), .A(
        n6565), .ZN(n6567) );
  OAI221_X1 U7206 ( .B1(BS16_N), .B2(keyinput_34), .C1(n6569), .C2(n6568), .A(
        n6567), .ZN(n6570) );
  OAI221_X1 U7207 ( .B1(READY_N), .B2(keyinput_35), .C1(n7124), .C2(n6571), 
        .A(n6570), .ZN(n6572) );
  AOI22_X1 U7208 ( .A1(n6573), .A2(n6572), .B1(ADS_N_REG_SCAN_IN), .B2(
        keyinput_38), .ZN(n6574) );
  OAI21_X1 U7209 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput_38), .A(n6574), .ZN(
        n6575) );
  OAI221_X1 U7210 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_39), .C1(n6577), 
        .C2(n6576), .A(n6575), .ZN(n6578) );
  OAI221_X1 U7211 ( .B1(M_IO_N_REG_SCAN_IN), .B2(n6579), .C1(n7114), .C2(
        keyinput_40), .A(n6578), .ZN(n6585) );
  AOI22_X1 U7212 ( .A1(n6581), .A2(keyinput_43), .B1(keyinput_45), .B2(n7034), 
        .ZN(n6580) );
  OAI221_X1 U7213 ( .B1(n6581), .B2(keyinput_43), .C1(n7034), .C2(keyinput_45), 
        .A(n6580), .ZN(n6584) );
  AOI22_X1 U7214 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_44), .B1(n6764), .B2(
        keyinput_42), .ZN(n6582) );
  OAI221_X1 U7215 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_44), .C1(n6764), .C2(
        keyinput_42), .A(n6582), .ZN(n6583) );
  AOI211_X1 U7216 ( .C1(n6586), .C2(n6585), .A(n6584), .B(n6583), .ZN(n6589)
         );
  INV_X1 U7217 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6698) );
  AOI22_X1 U7218 ( .A1(keyinput_46), .A2(W_R_N_REG_SCAN_IN), .B1(n6698), .B2(
        keyinput_47), .ZN(n6587) );
  OAI221_X1 U7219 ( .B1(keyinput_46), .B2(W_R_N_REG_SCAN_IN), .C1(n6698), .C2(
        keyinput_47), .A(n6587), .ZN(n6588) );
  AOI211_X1 U7220 ( .C1(BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_48), .A(n6589), .B(n6588), .ZN(n6590) );
  OAI21_X1 U7221 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_48), .A(n6590), 
        .ZN(n6591) );
  OAI211_X1 U7222 ( .C1(n6693), .C2(keyinput_49), .A(n6592), .B(n6591), .ZN(
        n6593) );
  AOI21_X1 U7223 ( .B1(n6693), .B2(keyinput_49), .A(n6593), .ZN(n6598) );
  AOI22_X1 U7224 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_53), .B1(n6678), 
        .B2(keyinput_52), .ZN(n6594) );
  OAI221_X1 U7225 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_53), .C1(n6678), 
        .C2(keyinput_52), .A(n6594), .ZN(n6597) );
  OAI22_X1 U7226 ( .A1(n6669), .A2(keyinput_55), .B1(keyinput_54), .B2(
        REIP_REG_28__SCAN_IN), .ZN(n6595) );
  AOI221_X1 U7227 ( .B1(n6669), .B2(keyinput_55), .C1(REIP_REG_28__SCAN_IN), 
        .C2(keyinput_54), .A(n6595), .ZN(n6596) );
  OAI21_X1 U7228 ( .B1(n6598), .B2(n6597), .A(n6596), .ZN(n6599) );
  OAI211_X1 U7229 ( .C1(REIP_REG_24__SCAN_IN), .C2(keyinput_58), .A(n6600), 
        .B(n6599), .ZN(n6601) );
  AOI21_X1 U7230 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_58), .A(n6601), 
        .ZN(n6602) );
  OAI22_X1 U7231 ( .A1(keyinput_61), .A2(n6605), .B1(n6603), .B2(n6602), .ZN(
        n6604) );
  AOI21_X1 U7232 ( .B1(keyinput_61), .B2(n6605), .A(n6604), .ZN(n6608) );
  INV_X1 U7233 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U7234 ( .A1(n6985), .A2(keyinput_63), .B1(n6983), .B2(keyinput_62), 
        .ZN(n6606) );
  OAI221_X1 U7235 ( .B1(n6985), .B2(keyinput_63), .C1(n6983), .C2(keyinput_62), 
        .A(n6606), .ZN(n6607) );
  AOI211_X1 U7236 ( .C1(n6610), .C2(n6609), .A(n6608), .B(n6607), .ZN(n6611)
         );
  XNOR2_X1 U7237 ( .A(n6612), .B(n6611), .ZN(U3171) );
  AOI22_X1 U7238 ( .A1(n6631), .A2(LWORD_REG_0__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6614) );
  OAI21_X1 U7239 ( .B1(n7130), .B2(n6633), .A(n6614), .ZN(U2923) );
  AOI22_X1 U7240 ( .A1(n6631), .A2(LWORD_REG_1__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6615) );
  OAI21_X1 U7241 ( .B1(n7134), .B2(n6633), .A(n6615), .ZN(U2922) );
  AOI22_X1 U7242 ( .A1(n6631), .A2(LWORD_REG_2__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6616) );
  OAI21_X1 U7243 ( .B1(n7139), .B2(n6633), .A(n6616), .ZN(U2921) );
  AOI22_X1 U7244 ( .A1(n6631), .A2(LWORD_REG_3__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6617) );
  OAI21_X1 U7245 ( .B1(n7144), .B2(n6633), .A(n6617), .ZN(U2920) );
  AOI22_X1 U7246 ( .A1(n6631), .A2(LWORD_REG_4__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6618) );
  OAI21_X1 U7247 ( .B1(n7149), .B2(n6633), .A(n6618), .ZN(U2919) );
  AOI22_X1 U7248 ( .A1(n6631), .A2(LWORD_REG_5__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6619) );
  OAI21_X1 U7249 ( .B1(n7154), .B2(n6633), .A(n6619), .ZN(U2918) );
  AOI22_X1 U7250 ( .A1(n6631), .A2(LWORD_REG_6__SCAN_IN), .B1(n6620), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6621) );
  OAI21_X1 U7251 ( .B1(n4291), .B2(n6633), .A(n6621), .ZN(U2917) );
  AOI22_X1 U7252 ( .A1(n6631), .A2(LWORD_REG_7__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6622) );
  OAI21_X1 U7253 ( .B1(n4298), .B2(n6633), .A(n6622), .ZN(U2916) );
  AOI22_X1 U7254 ( .A1(n6631), .A2(LWORD_REG_8__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6623) );
  OAI21_X1 U7255 ( .B1(n7166), .B2(n6633), .A(n6623), .ZN(U2915) );
  AOI22_X1 U7256 ( .A1(n6631), .A2(LWORD_REG_9__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6624) );
  OAI21_X1 U7257 ( .B1(n7171), .B2(n6633), .A(n6624), .ZN(U2914) );
  AOI22_X1 U7258 ( .A1(n6631), .A2(LWORD_REG_10__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6625) );
  OAI21_X1 U7259 ( .B1(n7176), .B2(n6633), .A(n6625), .ZN(U2913) );
  AOI22_X1 U7260 ( .A1(n6631), .A2(LWORD_REG_11__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6626) );
  OAI21_X1 U7261 ( .B1(n7181), .B2(n6633), .A(n6626), .ZN(U2912) );
  AOI22_X1 U7262 ( .A1(n6631), .A2(LWORD_REG_12__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6627) );
  OAI21_X1 U7263 ( .B1(n4366), .B2(n6633), .A(n6627), .ZN(U2911) );
  AOI22_X1 U7264 ( .A1(n6631), .A2(LWORD_REG_13__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6628) );
  OAI21_X1 U7265 ( .B1(n7189), .B2(n6633), .A(n6628), .ZN(U2910) );
  AOI22_X1 U7266 ( .A1(n6631), .A2(LWORD_REG_14__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6629) );
  OAI21_X1 U7267 ( .B1(n7195), .B2(n6633), .A(n6629), .ZN(U2909) );
  AOI22_X1 U7268 ( .A1(n6631), .A2(LWORD_REG_15__SCAN_IN), .B1(n6630), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6632) );
  OAI21_X1 U7269 ( .B1(n7200), .B2(n6633), .A(n6632), .ZN(U2908) );
  NAND2_X1 U7270 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7116), .ZN(n6677) );
  INV_X2 U7271 ( .A(n7116), .ZN(n7113) );
  NOR2_X2 U7272 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7113), .ZN(n6675) );
  AOI22_X1 U7273 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n7113), .ZN(n6634) );
  OAI21_X1 U7274 ( .B1(n6690), .B2(n6677), .A(n6634), .ZN(U3184) );
  AOI22_X1 U7275 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n7113), .ZN(n6635) );
  OAI21_X1 U7276 ( .B1(n6780), .B2(n6677), .A(n6635), .ZN(U3185) );
  AOI22_X1 U7277 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n7113), .ZN(n6636) );
  OAI21_X1 U7278 ( .B1(n6637), .B2(n6677), .A(n6636), .ZN(U3186) );
  AOI22_X1 U7279 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n7113), .ZN(n6638) );
  OAI21_X1 U7280 ( .B1(n6639), .B2(n6677), .A(n6638), .ZN(U3187) );
  AOI22_X1 U7281 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n7113), .ZN(n6640) );
  OAI21_X1 U7282 ( .B1(n6641), .B2(n6677), .A(n6640), .ZN(U3188) );
  INV_X1 U7283 ( .A(n6675), .ZN(n6672) );
  INV_X1 U7284 ( .A(n6677), .ZN(n6670) );
  AOI22_X1 U7285 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n7113), .ZN(n6642) );
  OAI21_X1 U7286 ( .B1(n6643), .B2(n6672), .A(n6642), .ZN(U3189) );
  INV_X1 U7287 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6793) );
  AOI22_X1 U7288 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n7113), .ZN(n6644) );
  OAI21_X1 U7289 ( .B1(n6793), .B2(n6672), .A(n6644), .ZN(U3190) );
  AOI22_X1 U7290 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n7113), .ZN(n6645) );
  OAI21_X1 U7291 ( .B1(n6793), .B2(n6677), .A(n6645), .ZN(U3191) );
  AOI22_X1 U7292 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n7113), .ZN(n6646) );
  OAI21_X1 U7293 ( .B1(n6647), .B2(n6677), .A(n6646), .ZN(U3192) );
  AOI22_X1 U7294 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n7113), .ZN(n6648) );
  OAI21_X1 U7295 ( .B1(n6650), .B2(n6672), .A(n6648), .ZN(U3193) );
  AOI22_X1 U7296 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n7113), .ZN(n6649) );
  OAI21_X1 U7297 ( .B1(n6650), .B2(n6677), .A(n6649), .ZN(U3194) );
  AOI22_X1 U7298 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n7113), .ZN(n6651) );
  OAI21_X1 U7299 ( .B1(n5882), .B2(n6672), .A(n6651), .ZN(U3195) );
  AOI22_X1 U7300 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n7113), .ZN(n6652) );
  OAI21_X1 U7301 ( .B1(n5882), .B2(n6677), .A(n6652), .ZN(U3196) );
  AOI22_X1 U7302 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n7113), .ZN(n6653) );
  OAI21_X1 U7303 ( .B1(n5947), .B2(n6672), .A(n6653), .ZN(U3197) );
  INV_X1 U7304 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6949) );
  AOI22_X1 U7305 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n7113), .ZN(n6654) );
  OAI21_X1 U7306 ( .B1(n6949), .B2(n6672), .A(n6654), .ZN(U3198) );
  AOI22_X1 U7307 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n7113), .ZN(n6655) );
  OAI21_X1 U7308 ( .B1(n6963), .B2(n6672), .A(n6655), .ZN(U3199) );
  AOI22_X1 U7309 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n7113), .ZN(n6656) );
  OAI21_X1 U7310 ( .B1(n6969), .B2(n6672), .A(n6656), .ZN(U3200) );
  AOI22_X1 U7311 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n7113), .ZN(n6657) );
  OAI21_X1 U7312 ( .B1(n6969), .B2(n6677), .A(n6657), .ZN(U3201) );
  AOI22_X1 U7313 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n7113), .ZN(n6658) );
  OAI21_X1 U7314 ( .B1(n6983), .B2(n6672), .A(n6658), .ZN(U3202) );
  AOI22_X1 U7315 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n7113), .ZN(n6659) );
  OAI21_X1 U7316 ( .B1(n6983), .B2(n6677), .A(n6659), .ZN(U3203) );
  AOI22_X1 U7317 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n7113), .ZN(n6660) );
  OAI21_X1 U7318 ( .B1(n6992), .B2(n6672), .A(n6660), .ZN(U3204) );
  AOI22_X1 U7319 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n7113), .ZN(n6661) );
  OAI21_X1 U7320 ( .B1(n6859), .B2(n6672), .A(n6661), .ZN(U3205) );
  AOI22_X1 U7321 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n7113), .ZN(n6662) );
  OAI21_X1 U7322 ( .B1(n6664), .B2(n6672), .A(n6662), .ZN(U3206) );
  AOI22_X1 U7323 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n7113), .ZN(n6663) );
  OAI21_X1 U7324 ( .B1(n6664), .B2(n6677), .A(n6663), .ZN(U3207) );
  AOI22_X1 U7325 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n7113), .ZN(n6665) );
  OAI21_X1 U7326 ( .B1(n6667), .B2(n6672), .A(n6665), .ZN(U3208) );
  AOI22_X1 U7327 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n7113), .ZN(n6666) );
  OAI21_X1 U7328 ( .B1(n6667), .B2(n6677), .A(n6666), .ZN(U3209) );
  AOI22_X1 U7329 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n7113), .ZN(n6668) );
  OAI21_X1 U7330 ( .B1(n6669), .B2(n6677), .A(n6668), .ZN(U3210) );
  AOI22_X1 U7331 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6670), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n7113), .ZN(n6671) );
  OAI21_X1 U7332 ( .B1(n6674), .B2(n6672), .A(n6671), .ZN(U3211) );
  AOI22_X1 U7333 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n7113), .ZN(n6673) );
  OAI21_X1 U7334 ( .B1(n6674), .B2(n6677), .A(n6673), .ZN(U3212) );
  AOI22_X1 U7335 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6675), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n7113), .ZN(n6676) );
  OAI21_X1 U7336 ( .B1(n6678), .B2(n6677), .A(n6676), .ZN(U3213) );
  MUX2_X1 U7337 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n7116), .Z(U3445) );
  AOI221_X1 U7338 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6689) );
  NOR4_X1 U7339 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6682) );
  NOR4_X1 U7340 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6681) );
  NOR4_X1 U7341 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6680) );
  NOR4_X1 U7342 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6679) );
  NAND4_X1 U7343 ( .A1(n6682), .A2(n6681), .A3(n6680), .A4(n6679), .ZN(n6688)
         );
  NOR4_X1 U7344 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6686) );
  AOI211_X1 U7345 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_11__SCAN_IN), .B(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6685) );
  NOR4_X1 U7346 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6684) );
  NOR4_X1 U7347 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6683) );
  NAND4_X1 U7348 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n6687)
         );
  NOR2_X1 U7349 ( .A1(n6688), .A2(n6687), .ZN(n6699) );
  MUX2_X1 U7350 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n6689), .S(n6699), .Z(
        U2795) );
  MUX2_X1 U7351 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n7116), .Z(U3446) );
  AOI21_X1 U7352 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6691) );
  OAI221_X1 U7353 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6691), .C1(n6690), .C2(
        REIP_REG_0__SCAN_IN), .A(n6699), .ZN(n6692) );
  OAI21_X1 U7354 ( .B1(n6699), .B2(n6693), .A(n6692), .ZN(U3468) );
  MUX2_X1 U7355 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n7116), .Z(U3447) );
  INV_X1 U7356 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6696) );
  NOR3_X1 U7357 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6694) );
  OAI21_X1 U7358 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6694), .A(n6699), .ZN(n6695)
         );
  OAI21_X1 U7359 ( .B1(n6699), .B2(n6696), .A(n6695), .ZN(U2794) );
  MUX2_X1 U7360 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n7116), .Z(U3448) );
  OAI21_X1 U7361 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6699), .ZN(n6697) );
  OAI21_X1 U7362 ( .B1(n6699), .B2(n6698), .A(n6697), .ZN(U3469) );
  INV_X1 U7363 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6701) );
  AOI22_X1 U7364 ( .A1(n7208), .A2(n6703), .B1(n6702), .B2(n6975), .ZN(n6700)
         );
  OAI21_X1 U7365 ( .B1(n6706), .B2(n6701), .A(n6700), .ZN(U2840) );
  AOI22_X1 U7366 ( .A1(n7229), .A2(n6703), .B1(n6702), .B2(n7014), .ZN(n6704)
         );
  OAI21_X1 U7367 ( .B1(n6706), .B2(n6705), .A(n6704), .ZN(U2835) );
  OAI21_X1 U7368 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6708), .A(n6707), 
        .ZN(n6877) );
  NAND2_X1 U7369 ( .A1(n6710), .A2(n6709), .ZN(n6712) );
  AOI22_X1 U7370 ( .A1(n6712), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6254), 
        .B2(n6711), .ZN(n6713) );
  NAND2_X1 U7371 ( .A1(n6847), .A2(REIP_REG_0__SCAN_IN), .ZN(n6875) );
  OAI211_X1 U7372 ( .C1(n7033), .C2(n6877), .A(n6713), .B(n6875), .ZN(U2986)
         );
  AOI22_X1 U7373 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6749), .B1(n6847), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6718) );
  OAI22_X1 U7374 ( .A1(n6715), .A2(n7033), .B1(n6742), .B2(n6714), .ZN(n6716)
         );
  INV_X1 U7375 ( .A(n6716), .ZN(n6717) );
  OAI211_X1 U7376 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6755), .A(n6718), 
        .B(n6717), .ZN(U2985) );
  AOI22_X1 U7377 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6749), .B1(n6847), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6726) );
  XNOR2_X1 U7378 ( .A(n6719), .B(n3872), .ZN(n6721) );
  XNOR2_X1 U7379 ( .A(n6721), .B(n6720), .ZN(n6782) );
  INV_X1 U7380 ( .A(n6782), .ZN(n6724) );
  INV_X1 U7381 ( .A(n6722), .ZN(n6723) );
  AOI22_X1 U7382 ( .A1(n6724), .A2(n6751), .B1(n6254), .B2(n6723), .ZN(n6725)
         );
  OAI211_X1 U7383 ( .C1(n6755), .C2(n6727), .A(n6726), .B(n6725), .ZN(U2984)
         );
  AOI22_X1 U7384 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6749), .B1(n6847), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6730) );
  AOI22_X1 U7385 ( .A1(n6728), .A2(n6751), .B1(n6254), .B2(n6885), .ZN(n6729)
         );
  OAI211_X1 U7386 ( .C1(n6755), .C2(n6888), .A(n6730), .B(n6729), .ZN(U2980)
         );
  AOI22_X1 U7387 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6749), .B1(n6847), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6736) );
  OAI21_X1 U7388 ( .B1(n6733), .B2(n6732), .A(n6731), .ZN(n6734) );
  INV_X1 U7389 ( .A(n6734), .ZN(n6802) );
  AOI22_X1 U7390 ( .A1(n6802), .A2(n6751), .B1(n6254), .B2(n6896), .ZN(n6735)
         );
  OAI211_X1 U7391 ( .C1(n6755), .C2(n6901), .A(n6736), .B(n6735), .ZN(U2979)
         );
  INV_X1 U7392 ( .A(n6738), .ZN(n6739) );
  NOR2_X1 U7393 ( .A1(n6740), .A2(n6739), .ZN(n6741) );
  XNOR2_X1 U7394 ( .A(n6737), .B(n6741), .ZN(n6839) );
  AOI22_X1 U7395 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6749), .B1(n6847), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n6745) );
  OAI22_X1 U7396 ( .A1(n6908), .A2(n6742), .B1(n6755), .B2(n6907), .ZN(n6743)
         );
  INV_X1 U7397 ( .A(n6743), .ZN(n6744) );
  OAI211_X1 U7398 ( .C1(n6839), .C2(n7033), .A(n6745), .B(n6744), .ZN(U2975)
         );
  AOI22_X1 U7399 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6749), .B1(n6847), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n6748) );
  AOI22_X1 U7400 ( .A1(n6746), .A2(n6751), .B1(n6254), .B2(n7205), .ZN(n6747)
         );
  OAI211_X1 U7401 ( .C1(n6755), .C2(n6959), .A(n6748), .B(n6747), .ZN(U2968)
         );
  AOI22_X1 U7402 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6749), .B1(n6847), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n6754) );
  AOI22_X1 U7403 ( .A1(n6752), .A2(n6751), .B1(n6254), .B2(n7211), .ZN(n6753)
         );
  OAI211_X1 U7404 ( .C1(n6755), .C2(n6979), .A(n6754), .B(n6753), .ZN(U2966)
         );
  INV_X1 U7405 ( .A(n6766), .ZN(n7088) );
  NAND2_X1 U7406 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7088), .ZN(n6760) );
  INV_X1 U7407 ( .A(n7026), .ZN(n6758) );
  OAI22_X1 U7408 ( .A1(n6758), .A2(n4035), .B1(n6757), .B2(n6756), .ZN(n7032)
         );
  OAI21_X1 U7409 ( .B1(n7032), .B2(n7073), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6759) );
  OAI21_X1 U7410 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6760), .A(n6759), .ZN(
        U2790) );
  NOR2_X1 U7411 ( .A1(n7116), .A2(D_C_N_REG_SCAN_IN), .ZN(n6761) );
  AOI22_X1 U7412 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7116), .B1(n6762), .B2(
        n6761), .ZN(U2791) );
  INV_X1 U7413 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6763) );
  AOI22_X1 U7414 ( .A1(n7116), .A2(READREQUEST_REG_SCAN_IN), .B1(n6763), .B2(
        n7113), .ZN(U3470) );
  AND2_X1 U7415 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n7100) );
  NOR2_X1 U7416 ( .A1(n7105), .A2(n6764), .ZN(n7108) );
  AOI21_X1 U7417 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7108), .ZN(n6765)
         );
  NAND2_X1 U7418 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7109) );
  OAI211_X1 U7419 ( .C1(n7100), .C2(n6765), .A(n6771), .B(n7109), .ZN(U3182)
         );
  NAND2_X1 U7420 ( .A1(n6766), .A2(n7083), .ZN(n6768) );
  NAND2_X1 U7421 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7124), .ZN(n7074) );
  OAI221_X1 U7422 ( .B1(n6768), .B2(n7076), .C1(n6768), .C2(n7074), .A(n6767), 
        .ZN(U3150) );
  AOI211_X1 U7423 ( .C1(n6631), .C2(n7124), .A(n6770), .B(n6769), .ZN(n6777)
         );
  AOI21_X1 U7424 ( .B1(n6772), .B2(n6771), .A(READY_N), .ZN(n7031) );
  OAI211_X1 U7425 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6773), .A(n7031), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6774) );
  AOI21_X1 U7426 ( .B1(n6774), .B2(STATE2_REG_0__SCAN_IN), .A(n7088), .ZN(
        n6776) );
  NAND2_X1 U7427 ( .A1(n6777), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6775) );
  OAI21_X1 U7428 ( .B1(n6777), .B2(n6776), .A(n6775), .ZN(U3472) );
  OAI21_X1 U7429 ( .B1(n6779), .B2(n6870), .A(n6778), .ZN(n6785) );
  OAI22_X1 U7430 ( .A1(n6794), .A2(n6781), .B1(n6780), .B2(n6860), .ZN(n6784)
         );
  NOR2_X1 U7431 ( .A1(n6782), .A2(n6878), .ZN(n6783) );
  AOI211_X1 U7432 ( .C1(n6816), .C2(n6785), .A(n6784), .B(n6783), .ZN(n6786)
         );
  OAI221_X1 U7433 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6788), .C1(n3872), .C2(n6787), .A(n6786), .ZN(U3016) );
  OAI22_X1 U7434 ( .A1(n6797), .A2(n6791), .B1(n6790), .B2(n6789), .ZN(n6806)
         );
  OAI222_X1 U7435 ( .A1(n6795), .A2(n6794), .B1(n6860), .B2(n6793), .C1(n6878), 
        .C2(n6792), .ZN(n6796) );
  INV_X1 U7436 ( .A(n6796), .ZN(n6800) );
  INV_X1 U7437 ( .A(n6808), .ZN(n6798) );
  NOR2_X1 U7438 ( .A1(n6798), .A2(n6797), .ZN(n6803) );
  OAI221_X1 U7439 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n6801), .C2(n6807), .A(n6803), 
        .ZN(n6799) );
  OAI211_X1 U7440 ( .C1(n6806), .C2(n6801), .A(n6800), .B(n6799), .ZN(U3010)
         );
  AOI22_X1 U7441 ( .A1(n6873), .A2(n6890), .B1(n6847), .B2(REIP_REG_7__SCAN_IN), .ZN(n6805) );
  AOI22_X1 U7442 ( .A1(n6803), .A2(n6807), .B1(n6802), .B2(n6857), .ZN(n6804)
         );
  OAI211_X1 U7443 ( .C1(n6807), .C2(n6806), .A(n6805), .B(n6804), .ZN(U3011)
         );
  NAND2_X1 U7444 ( .A1(n6809), .A2(n6808), .ZN(n6832) );
  OAI21_X1 U7445 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6810), .ZN(n6822) );
  AOI21_X1 U7446 ( .B1(n6873), .B2(n6812), .A(n6811), .ZN(n6821) );
  AOI22_X1 U7447 ( .A1(n6816), .A2(n6815), .B1(n6814), .B2(n6813), .ZN(n6817)
         );
  NAND2_X1 U7448 ( .A1(n6818), .A2(n6817), .ZN(n6828) );
  AOI22_X1 U7449 ( .A1(n6819), .A2(n6857), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6828), .ZN(n6820) );
  OAI211_X1 U7450 ( .C1(n6832), .C2(n6822), .A(n6821), .B(n6820), .ZN(U3008)
         );
  INV_X1 U7451 ( .A(n6823), .ZN(n6826) );
  INV_X1 U7452 ( .A(n6824), .ZN(n6825) );
  AOI21_X1 U7453 ( .B1(n6873), .B2(n6826), .A(n6825), .ZN(n6831) );
  INV_X1 U7454 ( .A(n6827), .ZN(n6829) );
  AOI22_X1 U7455 ( .A1(n6829), .A2(n6857), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6828), .ZN(n6830) );
  OAI211_X1 U7456 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6832), .A(n6831), 
        .B(n6830), .ZN(U3009) );
  INV_X1 U7457 ( .A(n6833), .ZN(n6906) );
  AOI22_X1 U7458 ( .A1(n6873), .A2(n6906), .B1(n6847), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7459 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6836), .B1(n6835), .B2(n6834), .ZN(n6837) );
  OAI211_X1 U7460 ( .C1(n6839), .C2(n6878), .A(n6838), .B(n6837), .ZN(U3007)
         );
  AOI21_X1 U7461 ( .B1(n6940), .B2(n6873), .A(n6840), .ZN(n6844) );
  AOI22_X1 U7462 ( .A1(n6842), .A2(n6857), .B1(n6841), .B2(n6845), .ZN(n6843)
         );
  OAI211_X1 U7463 ( .C1(n6846), .C2(n6845), .A(n6844), .B(n6843), .ZN(U3003)
         );
  AOI22_X1 U7464 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6848), .B1(n6847), .B2(REIP_REG_17__SCAN_IN), .ZN(n6852) );
  AOI22_X1 U7465 ( .A1(n6850), .A2(n6857), .B1(n6873), .B2(n6849), .ZN(n6851)
         );
  OAI211_X1 U7466 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n6853), .A(n6852), .B(n6851), .ZN(U3001) );
  INV_X1 U7467 ( .A(n6854), .ZN(n6858) );
  INV_X1 U7468 ( .A(n6855), .ZN(n6856) );
  AOI22_X1 U7469 ( .A1(n6858), .A2(n6857), .B1(n6873), .B2(n6856), .ZN(n6866)
         );
  NOR2_X1 U7470 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  AOI221_X1 U7471 ( .B1(n6864), .B2(n6863), .C1(n6862), .C2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A(n6861), .ZN(n6865) );
  NAND2_X1 U7472 ( .A1(n6866), .A2(n6865), .ZN(U2995) );
  INV_X1 U7473 ( .A(n6867), .ZN(n6871) );
  AOI22_X1 U7474 ( .A1(n6871), .A2(n6870), .B1(n6869), .B2(n6868), .ZN(n6872)
         );
  AOI21_X1 U7475 ( .B1(n6874), .B2(n6873), .A(n6872), .ZN(n6876) );
  OAI211_X1 U7476 ( .C1(n6878), .C2(n6877), .A(n6876), .B(n6875), .ZN(U3018)
         );
  NOR3_X1 U7477 ( .A1(n7010), .A2(REIP_REG_6__SCAN_IN), .A3(n6879), .ZN(n6898)
         );
  NOR2_X1 U7478 ( .A1(n6880), .A2(n6998), .ZN(n6881) );
  AOI211_X1 U7479 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6897), .A(n6898), .B(n6881), 
        .ZN(n6887) );
  INV_X1 U7480 ( .A(n6974), .ZN(n6891) );
  OAI21_X1 U7481 ( .B1(n6980), .B2(n4286), .A(n6891), .ZN(n6884) );
  NOR2_X1 U7482 ( .A1(n7006), .A2(n6882), .ZN(n6883) );
  AOI211_X1 U7483 ( .C1(n7016), .C2(n6885), .A(n6884), .B(n6883), .ZN(n6886)
         );
  OAI211_X1 U7484 ( .C1(n6888), .C2(n6999), .A(n6887), .B(n6886), .ZN(U2821)
         );
  NOR3_X1 U7485 ( .A1(n7010), .A2(REIP_REG_7__SCAN_IN), .A3(n6889), .ZN(n6895)
         );
  INV_X1 U7486 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6893) );
  AOI22_X1 U7487 ( .A1(EBX_REG_7__SCAN_IN), .A2(n7008), .B1(n7015), .B2(n6890), 
        .ZN(n6892) );
  OAI211_X1 U7488 ( .C1(n6980), .C2(n6893), .A(n6892), .B(n6891), .ZN(n6894)
         );
  AOI211_X1 U7489 ( .C1(n6896), .C2(n7016), .A(n6895), .B(n6894), .ZN(n6900)
         );
  OAI21_X1 U7490 ( .B1(n6898), .B2(n6897), .A(REIP_REG_7__SCAN_IN), .ZN(n6899)
         );
  OAI211_X1 U7491 ( .C1(n6999), .C2(n6901), .A(n6900), .B(n6899), .ZN(U2820)
         );
  INV_X1 U7492 ( .A(n6902), .ZN(n6904) );
  NOR3_X1 U7493 ( .A1(n6904), .A2(REIP_REG_11__SCAN_IN), .A3(n6903), .ZN(n6905) );
  AOI21_X1 U7494 ( .B1(n6906), .B2(n7015), .A(n6905), .ZN(n6913) );
  AOI22_X1 U7495 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n7009), .B1(
        EBX_REG_11__SCAN_IN), .B2(n7008), .ZN(n6912) );
  AOI21_X1 U7496 ( .B1(REIP_REG_11__SCAN_IN), .B2(n6921), .A(n6974), .ZN(n6911) );
  OAI22_X1 U7497 ( .A1(n6908), .A2(n7001), .B1(n6999), .B2(n6907), .ZN(n6909)
         );
  INV_X1 U7498 ( .A(n6909), .ZN(n6910) );
  NAND4_X1 U7499 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(U2816)
         );
  AOI22_X1 U7500 ( .A1(EBX_REG_13__SCAN_IN), .A2(n7008), .B1(n7015), .B2(n6914), .ZN(n6926) );
  NOR3_X1 U7501 ( .A1(n7010), .A2(REIP_REG_13__SCAN_IN), .A3(n6915), .ZN(n6916) );
  AOI211_X1 U7502 ( .C1(n7009), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6974), 
        .B(n6916), .ZN(n6925) );
  INV_X1 U7503 ( .A(n6917), .ZN(n6920) );
  INV_X1 U7504 ( .A(n6918), .ZN(n6919) );
  AOI22_X1 U7505 ( .A1(n6920), .A2(n7016), .B1(n6919), .B2(n7017), .ZN(n6924)
         );
  OAI21_X1 U7506 ( .B1(n6922), .B2(n6921), .A(REIP_REG_13__SCAN_IN), .ZN(n6923) );
  NAND4_X1 U7507 ( .A1(n6926), .A2(n6925), .A3(n6924), .A4(n6923), .ZN(U2814)
         );
  AOI21_X1 U7508 ( .B1(n6994), .B2(n6927), .A(REIP_REG_14__SCAN_IN), .ZN(n6938) );
  NOR2_X1 U7509 ( .A1(n6929), .A2(n6928), .ZN(n6947) );
  INV_X1 U7510 ( .A(n6947), .ZN(n6937) );
  OAI22_X1 U7511 ( .A1(n6931), .A2(n6998), .B1(n7006), .B2(n6930), .ZN(n6932)
         );
  AOI211_X1 U7512 ( .C1(n7009), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6974), 
        .B(n6932), .ZN(n6936) );
  AOI22_X1 U7513 ( .A1(n6934), .A2(n7016), .B1(n7017), .B2(n6933), .ZN(n6935)
         );
  OAI211_X1 U7514 ( .C1(n6938), .C2(n6937), .A(n6936), .B(n6935), .ZN(U2813)
         );
  AOI22_X1 U7515 ( .A1(EBX_REG_15__SCAN_IN), .A2(n7008), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6947), .ZN(n6946) );
  AND2_X1 U7516 ( .A1(n5947), .A2(n6950), .ZN(n6948) );
  AOI211_X1 U7517 ( .C1(n7009), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6974), 
        .B(n6948), .ZN(n6945) );
  INV_X1 U7518 ( .A(n6939), .ZN(n6941) );
  AOI22_X1 U7519 ( .A1(n6941), .A2(n7016), .B1(n7015), .B2(n6940), .ZN(n6944)
         );
  NAND2_X1 U7520 ( .A1(n6942), .A2(n7017), .ZN(n6943) );
  NAND4_X1 U7521 ( .A1(n6946), .A2(n6945), .A3(n6944), .A4(n6943), .ZN(U2812)
         );
  OAI21_X1 U7522 ( .B1(n6948), .B2(n6947), .A(REIP_REG_16__SCAN_IN), .ZN(n6952) );
  NAND3_X1 U7523 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6950), .A3(n6949), .ZN(
        n6951) );
  OAI211_X1 U7524 ( .C1(n6998), .C2(n6953), .A(n6952), .B(n6951), .ZN(n6954)
         );
  AOI211_X1 U7525 ( .C1(n7009), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6974), 
        .B(n6954), .ZN(n6957) );
  AOI22_X1 U7526 ( .A1(n7202), .A2(n7016), .B1(n7017), .B2(n6955), .ZN(n6956)
         );
  OAI211_X1 U7527 ( .C1(n7006), .C2(n6958), .A(n6957), .B(n6956), .ZN(U2811)
         );
  AOI21_X1 U7528 ( .B1(n7009), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6974), 
        .ZN(n6967) );
  AOI22_X1 U7529 ( .A1(EBX_REG_18__SCAN_IN), .A2(n7008), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6968), .ZN(n6966) );
  OAI22_X1 U7530 ( .A1(n7006), .A2(n6960), .B1(n6959), .B2(n6999), .ZN(n6961)
         );
  AOI21_X1 U7531 ( .B1(n7205), .B2(n7016), .A(n6961), .ZN(n6965) );
  NOR2_X1 U7532 ( .A1(n6963), .A2(n6962), .ZN(n6970) );
  NAND2_X1 U7533 ( .A1(n6970), .A2(n6969), .ZN(n6964) );
  NAND4_X1 U7534 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(U2809)
         );
  AOI21_X1 U7535 ( .B1(n6970), .B2(n6969), .A(n6968), .ZN(n6978) );
  NAND2_X1 U7536 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6970), .ZN(n6984) );
  AOI22_X1 U7537 ( .A1(n6971), .A2(n7017), .B1(EBX_REG_19__SCAN_IN), .B2(n7008), .ZN(n6972) );
  OAI21_X1 U7538 ( .B1(REIP_REG_19__SCAN_IN), .B2(n6984), .A(n6972), .ZN(n6973) );
  AOI211_X1 U7539 ( .C1(n7009), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6974), 
        .B(n6973), .ZN(n6977) );
  AOI22_X1 U7540 ( .A1(n7208), .A2(n7016), .B1(n7015), .B2(n6975), .ZN(n6976)
         );
  OAI211_X1 U7541 ( .C1(n6978), .C2(n6985), .A(n6977), .B(n6976), .ZN(U2808)
         );
  INV_X1 U7542 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6981) );
  OAI22_X1 U7543 ( .A1(n6981), .A2(n6980), .B1(n6979), .B2(n6999), .ZN(n6982)
         );
  AOI21_X1 U7544 ( .B1(EBX_REG_20__SCAN_IN), .B2(n7008), .A(n6982), .ZN(n6988)
         );
  OAI21_X1 U7545 ( .B1(n6985), .B2(n6984), .A(n6983), .ZN(n6986) );
  AOI22_X1 U7546 ( .A1(n7211), .A2(n7016), .B1(n6986), .B2(n6990), .ZN(n6987)
         );
  OAI211_X1 U7547 ( .C1(n6989), .C2(n7006), .A(n6988), .B(n6987), .ZN(U2807)
         );
  OAI21_X1 U7548 ( .B1(n6991), .B2(n6990), .A(REIP_REG_22__SCAN_IN), .ZN(n6996) );
  NAND3_X1 U7549 ( .A1(n6994), .A2(n6993), .A3(n6992), .ZN(n6995) );
  OAI211_X1 U7550 ( .C1(n6998), .C2(n6997), .A(n6996), .B(n6995), .ZN(n7004)
         );
  INV_X1 U7551 ( .A(n7214), .ZN(n7002) );
  OAI22_X1 U7552 ( .A1(n7002), .A2(n7001), .B1(n7000), .B2(n6999), .ZN(n7003)
         );
  AOI211_X1 U7553 ( .C1(PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n7009), .A(n7004), 
        .B(n7003), .ZN(n7005) );
  OAI21_X1 U7554 ( .B1(n7007), .B2(n7006), .A(n7005), .ZN(U2805) );
  AOI22_X1 U7555 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n7009), .B1(
        EBX_REG_24__SCAN_IN), .B2(n7008), .ZN(n7022) );
  NOR2_X1 U7556 ( .A1(n7010), .A2(REIP_REG_24__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U7557 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7013), .B1(n7012), .B2(
        n7011), .ZN(n7021) );
  AOI22_X1 U7558 ( .A1(n7229), .A2(n7016), .B1(n7015), .B2(n7014), .ZN(n7020)
         );
  NAND2_X1 U7559 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  NAND4_X1 U7560 ( .A1(n7022), .A2(n7021), .A3(n7020), .A4(n7019), .ZN(U2803)
         );
  OR2_X1 U7561 ( .A1(n7026), .A2(n7023), .ZN(n7028) );
  NAND2_X1 U7562 ( .A1(n7024), .A2(n4774), .ZN(n7025) );
  NAND2_X1 U7563 ( .A1(n7026), .A2(n7025), .ZN(n7027) );
  OAI211_X1 U7564 ( .C1(n7030), .C2(n7029), .A(n7028), .B(n7027), .ZN(n7061)
         );
  NOR2_X1 U7565 ( .A1(n7032), .A2(n7031), .ZN(n7064) );
  NOR2_X1 U7566 ( .A1(n7064), .A2(n7073), .ZN(n7035) );
  MUX2_X1 U7567 ( .A(MORE_REG_SCAN_IN), .B(n7061), .S(n7035), .Z(U3471) );
  OAI21_X1 U7568 ( .B1(n7035), .B2(n7034), .A(n7033), .ZN(U2793) );
  INV_X1 U7569 ( .A(n7036), .ZN(n7038) );
  NAND3_X1 U7570 ( .A1(n7038), .A2(n7084), .A3(n7037), .ZN(n7039) );
  OAI21_X1 U7571 ( .B1(n7041), .B2(n7040), .A(n7039), .ZN(U3455) );
  INV_X1 U7572 ( .A(n7055), .ZN(n7057) );
  INV_X1 U7573 ( .A(n7042), .ZN(n7046) );
  INV_X1 U7574 ( .A(n7051), .ZN(n7044) );
  NOR3_X1 U7575 ( .A1(n7044), .A2(n7048), .A3(n7043), .ZN(n7045) );
  OAI22_X1 U7576 ( .A1(n7047), .A2(n7046), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n7045), .ZN(n7053) );
  INV_X1 U7577 ( .A(n7048), .ZN(n7049) );
  NAND3_X1 U7578 ( .A1(n7051), .A2(n7050), .A3(n7049), .ZN(n7052) );
  OAI211_X1 U7579 ( .C1(n7055), .C2(n7054), .A(n7053), .B(n7052), .ZN(n7056)
         );
  OAI21_X1 U7580 ( .B1(n7057), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n7056), 
        .ZN(n7058) );
  AOI222_X1 U7581 ( .A1(n7060), .A2(n7059), .B1(n7060), .B2(n7058), .C1(n7059), 
        .C2(n7058), .ZN(n7067) );
  NOR3_X1 U7582 ( .A1(n7063), .A2(n7062), .A3(n7061), .ZN(n7066) );
  OAI21_X1 U7583 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n7064), 
        .ZN(n7065) );
  OAI211_X1 U7584 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n7067), .A(n7066), .B(n7065), .ZN(n7091) );
  OR2_X1 U7585 ( .A1(n7091), .A2(n7073), .ZN(n7072) );
  NAND2_X1 U7586 ( .A1(READY_N), .A2(n6631), .ZN(n7071) );
  NOR2_X1 U7587 ( .A1(n7069), .A2(n7068), .ZN(n7070) );
  AOI21_X1 U7588 ( .B1(n7072), .B2(n7071), .A(n7070), .ZN(n7086) );
  INV_X1 U7589 ( .A(n7086), .ZN(n7085) );
  OAI21_X1 U7590 ( .B1(n7075), .B2(n7074), .A(n7073), .ZN(n7079) );
  OAI221_X1 U7591 ( .B1(n7086), .B2(READY_N), .C1(n7086), .C2(n7076), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n7093) );
  AOI21_X1 U7592 ( .B1(n7093), .B2(n7085), .A(n7077), .ZN(n7078) );
  AOI21_X1 U7593 ( .B1(n7085), .B2(n7079), .A(n7078), .ZN(n7081) );
  NAND2_X1 U7594 ( .A1(n7081), .A2(n7080), .ZN(U3149) );
  OAI211_X1 U7595 ( .C1(n7085), .C2(n7084), .A(n7083), .B(n7082), .ZN(U3453)
         );
  AOI211_X1 U7596 ( .C1(n7088), .C2(n7087), .A(STATE2_REG_0__SCAN_IN), .B(
        n7086), .ZN(n7089) );
  AOI211_X1 U7597 ( .C1(n7092), .C2(n7091), .A(n7090), .B(n7089), .ZN(n7094)
         );
  OAI211_X1 U7598 ( .C1(n7096), .C2(n7095), .A(n7094), .B(n7093), .ZN(U3148)
         );
  AOI21_X1 U7599 ( .B1(n6398), .B2(STATEBS16_REG_SCAN_IN), .A(n7098), .ZN(
        n7097) );
  INV_X1 U7600 ( .A(n7097), .ZN(U2792) );
  AOI21_X1 U7601 ( .B1(n6398), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(n7098), .ZN(
        n7099) );
  INV_X1 U7602 ( .A(n7099), .ZN(U3452) );
  NAND2_X1 U7603 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n7104) );
  INV_X1 U7604 ( .A(n7109), .ZN(n7102) );
  AOI221_X1 U7605 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7107), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7111) );
  AOI221_X1 U7606 ( .B1(n7102), .B2(n7101), .C1(n7100), .C2(n7101), .A(n7111), 
        .ZN(n7103) );
  OAI221_X1 U7607 ( .B1(n7116), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7116), 
        .C2(n7104), .A(n7103), .ZN(U3181) );
  AOI221_X1 U7608 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7124), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7106) );
  AOI221_X1 U7609 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7106), .C2(HOLD), .A(n7105), .ZN(n7112) );
  AOI21_X1 U7610 ( .B1(n7108), .B2(n7107), .A(STATE_REG_2__SCAN_IN), .ZN(n7110) );
  OAI22_X1 U7611 ( .A1(n7112), .A2(n7111), .B1(n7110), .B2(n7109), .ZN(U3183)
         );
  AOI22_X1 U7612 ( .A1(n7116), .A2(n7115), .B1(n7114), .B2(n7113), .ZN(U3473)
         );
  AOI21_X1 U7613 ( .B1(n7118), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n7117), .ZN(
        n7119) );
  INV_X1 U7614 ( .A(n7119), .ZN(U2788) );
  NAND2_X2 U7615 ( .A1(n7121), .A2(n7120), .ZN(n7199) );
  INV_X1 U7616 ( .A(n7122), .ZN(n7123) );
  OAI21_X1 U7617 ( .B1(n3821), .B2(n7124), .A(n7123), .ZN(n7193) );
  AND2_X1 U7618 ( .A1(n7196), .A2(DATAI_0_), .ZN(n7128) );
  AOI21_X1 U7619 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n7197), .A(n7128), .ZN(n7126) );
  OAI21_X1 U7620 ( .B1(n7127), .B2(n7199), .A(n7126), .ZN(U2924) );
  AOI21_X1 U7621 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n7197), .A(n7128), .ZN(n7129) );
  OAI21_X1 U7622 ( .B1(n7130), .B2(n7199), .A(n7129), .ZN(U2939) );
  AND2_X1 U7623 ( .A1(n7196), .A2(DATAI_1_), .ZN(n7132) );
  AOI21_X1 U7624 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n7197), .A(n7132), .ZN(n7131) );
  OAI21_X1 U7625 ( .B1(n4464), .B2(n7199), .A(n7131), .ZN(U2925) );
  AOI21_X1 U7626 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n7197), .A(n7132), .ZN(n7133) );
  OAI21_X1 U7627 ( .B1(n7134), .B2(n7199), .A(n7133), .ZN(U2940) );
  AND2_X1 U7628 ( .A1(n7196), .A2(DATAI_2_), .ZN(n7137) );
  AOI21_X1 U7629 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n7197), .A(n7137), .ZN(n7135) );
  OAI21_X1 U7630 ( .B1(n7136), .B2(n7199), .A(n7135), .ZN(U2926) );
  AOI21_X1 U7631 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n7197), .A(n7137), .ZN(n7138) );
  OAI21_X1 U7632 ( .B1(n7139), .B2(n7199), .A(n7138), .ZN(U2941) );
  AND2_X1 U7633 ( .A1(n7196), .A2(DATAI_3_), .ZN(n7142) );
  AOI21_X1 U7634 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n7197), .A(n7142), .ZN(n7140) );
  OAI21_X1 U7635 ( .B1(n7141), .B2(n7199), .A(n7140), .ZN(U2927) );
  AOI21_X1 U7636 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n7197), .A(n7142), .ZN(n7143) );
  OAI21_X1 U7637 ( .B1(n7144), .B2(n7199), .A(n7143), .ZN(U2942) );
  AND2_X1 U7638 ( .A1(n7196), .A2(DATAI_4_), .ZN(n7147) );
  AOI21_X1 U7639 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n7197), .A(n7147), .ZN(n7145) );
  OAI21_X1 U7640 ( .B1(n7146), .B2(n7199), .A(n7145), .ZN(U2928) );
  AOI21_X1 U7641 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n7197), .A(n7147), .ZN(n7148) );
  OAI21_X1 U7642 ( .B1(n7149), .B2(n7199), .A(n7148), .ZN(U2943) );
  AND2_X1 U7643 ( .A1(n7196), .A2(DATAI_5_), .ZN(n7152) );
  AOI21_X1 U7644 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n7197), .A(n7152), .ZN(n7150) );
  OAI21_X1 U7645 ( .B1(n7151), .B2(n7199), .A(n7150), .ZN(U2929) );
  AOI21_X1 U7646 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n7197), .A(n7152), .ZN(n7153) );
  OAI21_X1 U7647 ( .B1(n7154), .B2(n7199), .A(n7153), .ZN(U2944) );
  AND2_X1 U7648 ( .A1(n7196), .A2(DATAI_6_), .ZN(n7157) );
  AOI21_X1 U7649 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n7197), .A(n7157), .ZN(n7155) );
  OAI21_X1 U7650 ( .B1(n7156), .B2(n7199), .A(n7155), .ZN(U2930) );
  AOI21_X1 U7651 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n7197), .A(n7157), .ZN(n7158) );
  OAI21_X1 U7652 ( .B1(n4291), .B2(n7199), .A(n7158), .ZN(U2945) );
  AND2_X1 U7653 ( .A1(n7196), .A2(DATAI_7_), .ZN(n7160) );
  AOI21_X1 U7654 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n7197), .A(n7160), .ZN(n7159) );
  OAI21_X1 U7655 ( .B1(n4574), .B2(n7199), .A(n7159), .ZN(U2931) );
  AOI21_X1 U7656 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n7197), .A(n7160), .ZN(n7161) );
  OAI21_X1 U7657 ( .B1(n4298), .B2(n7199), .A(n7161), .ZN(U2946) );
  AND2_X1 U7658 ( .A1(n7196), .A2(DATAI_8_), .ZN(n7164) );
  AOI21_X1 U7659 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n7197), .A(n7164), .ZN(n7162) );
  OAI21_X1 U7660 ( .B1(n7163), .B2(n7199), .A(n7162), .ZN(U2932) );
  AOI21_X1 U7661 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n7197), .A(n7164), .ZN(n7165) );
  OAI21_X1 U7662 ( .B1(n7166), .B2(n7199), .A(n7165), .ZN(U2947) );
  AND2_X1 U7663 ( .A1(n7196), .A2(DATAI_9_), .ZN(n7169) );
  AOI21_X1 U7664 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n7197), .A(n7169), .ZN(n7167) );
  OAI21_X1 U7665 ( .B1(n7168), .B2(n7199), .A(n7167), .ZN(U2933) );
  AOI21_X1 U7666 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n7197), .A(n7169), .ZN(n7170) );
  OAI21_X1 U7667 ( .B1(n7171), .B2(n7199), .A(n7170), .ZN(U2948) );
  AND2_X1 U7668 ( .A1(n7196), .A2(DATAI_10_), .ZN(n7174) );
  AOI21_X1 U7669 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n7197), .A(n7174), .ZN(
        n7172) );
  OAI21_X1 U7670 ( .B1(n7173), .B2(n7199), .A(n7172), .ZN(U2934) );
  AOI21_X1 U7671 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n7197), .A(n7174), .ZN(
        n7175) );
  OAI21_X1 U7672 ( .B1(n7176), .B2(n7199), .A(n7175), .ZN(U2949) );
  AND2_X1 U7673 ( .A1(n7196), .A2(DATAI_11_), .ZN(n7179) );
  AOI21_X1 U7674 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n7197), .A(n7179), .ZN(
        n7177) );
  OAI21_X1 U7675 ( .B1(n7178), .B2(n7199), .A(n7177), .ZN(U2935) );
  AOI21_X1 U7676 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n7197), .A(n7179), .ZN(
        n7180) );
  OAI21_X1 U7677 ( .B1(n7181), .B2(n7199), .A(n7180), .ZN(U2950) );
  AND2_X1 U7678 ( .A1(n7196), .A2(DATAI_12_), .ZN(n7184) );
  AOI21_X1 U7679 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n7197), .A(n7184), .ZN(
        n7182) );
  OAI21_X1 U7680 ( .B1(n7183), .B2(n7199), .A(n7182), .ZN(U2936) );
  AOI21_X1 U7681 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n7193), .A(n7184), .ZN(
        n7185) );
  OAI21_X1 U7682 ( .B1(n4366), .B2(n7199), .A(n7185), .ZN(U2951) );
  AND2_X1 U7683 ( .A1(n7196), .A2(DATAI_13_), .ZN(n7187) );
  AOI21_X1 U7684 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n7193), .A(n7187), .ZN(
        n7186) );
  OAI21_X1 U7685 ( .B1(n4690), .B2(n7199), .A(n7186), .ZN(U2937) );
  AOI21_X1 U7686 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n7193), .A(n7187), .ZN(
        n7188) );
  OAI21_X1 U7687 ( .B1(n7189), .B2(n7199), .A(n7188), .ZN(U2952) );
  AND2_X1 U7688 ( .A1(n7196), .A2(DATAI_14_), .ZN(n7192) );
  AOI21_X1 U7689 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n7193), .A(n7192), .ZN(
        n7190) );
  OAI21_X1 U7690 ( .B1(n7191), .B2(n7199), .A(n7190), .ZN(U2938) );
  AOI21_X1 U7691 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n7193), .A(n7192), .ZN(
        n7194) );
  OAI21_X1 U7692 ( .B1(n7195), .B2(n7199), .A(n7194), .ZN(U2953) );
  AOI22_X1 U7693 ( .A1(n7197), .A2(LWORD_REG_15__SCAN_IN), .B1(n7196), .B2(
        DATAI_15_), .ZN(n7198) );
  OAI21_X1 U7694 ( .B1(n7200), .B2(n7199), .A(n7198), .ZN(U2954) );
  INV_X1 U7695 ( .A(n7201), .ZN(n7233) );
  AOI22_X1 U7696 ( .A1(n7202), .A2(n7233), .B1(n7232), .B2(DATAI_16_), .ZN(
        n7204) );
  AOI22_X1 U7697 ( .A1(n7236), .A2(DATAI_0_), .B1(n7235), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n7203) );
  NAND2_X1 U7698 ( .A1(n7204), .A2(n7203), .ZN(U2875) );
  AOI22_X1 U7699 ( .A1(n7205), .A2(n7233), .B1(n7232), .B2(DATAI_18_), .ZN(
        n7207) );
  AOI22_X1 U7700 ( .A1(n7236), .A2(DATAI_2_), .B1(n7235), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n7206) );
  NAND2_X1 U7701 ( .A1(n7207), .A2(n7206), .ZN(U2873) );
  AOI22_X1 U7702 ( .A1(n7208), .A2(n7233), .B1(n7232), .B2(DATAI_19_), .ZN(
        n7210) );
  AOI22_X1 U7703 ( .A1(n7236), .A2(DATAI_3_), .B1(n7235), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U7704 ( .A1(n7210), .A2(n7209), .ZN(U2872) );
  AOI22_X1 U7705 ( .A1(n7211), .A2(n7233), .B1(n7232), .B2(DATAI_20_), .ZN(
        n7213) );
  AOI22_X1 U7706 ( .A1(n7236), .A2(DATAI_4_), .B1(n7235), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n7212) );
  NAND2_X1 U7707 ( .A1(n7213), .A2(n7212), .ZN(U2871) );
  AOI22_X1 U7708 ( .A1(n7214), .A2(n7233), .B1(n7232), .B2(DATAI_22_), .ZN(
        n7216) );
  AOI22_X1 U7709 ( .A1(n7236), .A2(DATAI_6_), .B1(n7235), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n7215) );
  NAND2_X1 U7710 ( .A1(n7216), .A2(n7215), .ZN(U2869) );
  INV_X1 U7711 ( .A(n7217), .ZN(n7218) );
  AOI22_X1 U7712 ( .A1(n7221), .A2(n7220), .B1(n7219), .B2(n7218), .ZN(n7226)
         );
  AOI22_X1 U7713 ( .A1(n7224), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n7223), 
        .B2(n7222), .ZN(n7225) );
  OAI211_X1 U7714 ( .C1(n7228), .C2(n7227), .A(n7226), .B(n7225), .ZN(U3124)
         );
  AOI22_X1 U7715 ( .A1(n7229), .A2(n7233), .B1(n7232), .B2(DATAI_24_), .ZN(
        n7231) );
  AOI22_X1 U7716 ( .A1(n7236), .A2(DATAI_8_), .B1(n7235), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n7230) );
  NAND2_X1 U7717 ( .A1(n7231), .A2(n7230), .ZN(U2867) );
  AOI22_X1 U7718 ( .A1(n7234), .A2(n7233), .B1(n7232), .B2(DATAI_25_), .ZN(
        n7238) );
  AOI22_X1 U7719 ( .A1(n7236), .A2(DATAI_9_), .B1(n7235), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U7720 ( .A1(n7238), .A2(n7237), .ZN(U2866) );
  NAND2_X1 U3635 ( .A1(n3751), .A2(n3750), .ZN(n4070) );
  AND2_X1 U3902 ( .A1(n6000), .A2(n4821), .ZN(n3855) );
  AND2_X1 U4194 ( .A1(n3749), .A2(n3748), .ZN(n3751) );
  CLKBUF_X1 U3496 ( .A(n3699), .Z(n3466) );
  AND4_X1 U3504 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .ZN(n3593)
         );
  CLKBUF_X1 U3507 ( .A(n3838), .Z(n3446) );
  CLKBUF_X1 U3537 ( .A(n3511), .Z(n3445) );
  CLKBUF_X1 U3615 ( .A(n6031), .Z(n6032) );
  CLKBUF_X1 U6566 ( .A(n6620), .Z(n6630) );
  CLKBUF_X1 U6689 ( .A(n6101), .Z(n6102) );
  CLKBUF_X1 U6750 ( .A(n5918), .Z(n5919) );
endmodule

