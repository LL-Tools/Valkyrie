

module b15_C_AntiSAT_k_128_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819;

  CLKBUF_X2 U3458 ( .A(n3249), .Z(n4218) );
  CLKBUF_X2 U34590 ( .A(n3390), .Z(n4257) );
  CLKBUF_X2 U34600 ( .A(n3247), .Z(n4224) );
  AND2_X1 U34610 ( .A1(n3567), .A2(n3233), .ZN(n3589) );
  AND2_X1 U34620 ( .A1(n3609), .A2(n3331), .ZN(n3326) );
  INV_X1 U34630 ( .A(n3717), .ZN(n3725) );
  NAND2_X1 U34640 ( .A1(n4421), .A2(n3265), .ZN(n4353) );
  INV_X1 U34650 ( .A(n3839), .ZN(n4273) );
  INV_X1 U3466 ( .A(n3272), .ZN(n3612) );
  INV_X1 U3467 ( .A(n3237), .ZN(n3790) );
  INV_X1 U34690 ( .A(n6062), .ZN(n6101) );
  NAND2_X2 U34710 ( .A1(n3081), .A2(n4370), .ZN(n3459) );
  BUF_X8 U34720 ( .A(n3316), .Z(n4255) );
  XNOR2_X2 U34730 ( .A(n3349), .B(n3347), .ZN(n3417) );
  NOR2_X2 U34740 ( .A1(n5644), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5643) );
  NAND2_X2 U3475 ( .A1(n3076), .A2(n3075), .ZN(n5644) );
  NOR2_X4 U3476 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4588) );
  AOI22_X2 U3477 ( .A1(n6195), .A2(n3437), .B1(n3436), .B2(n3435), .ZN(n4540)
         );
  OR2_X2 U3478 ( .A1(n5631), .A2(n5632), .ZN(n5608) );
  NAND2_X1 U3479 ( .A1(n5234), .A2(n3528), .ZN(n5248) );
  OAI21_X1 U3481 ( .B1(n3791), .B2(STATE2_REG_0__SCAN_IN), .A(n3424), .ZN(
        n3309) );
  AND2_X1 U3482 ( .A1(n3334), .A2(n5032), .ZN(n4449) );
  BUF_X1 U3483 ( .A(n3680), .Z(n3026) );
  BUF_X2 U3484 ( .A(n3273), .Z(n3022) );
  NAND2_X1 U3485 ( .A1(n3325), .A2(n3237), .ZN(n3255) );
  INV_X1 U3486 ( .A(n3233), .ZN(n4564) );
  OR2_X2 U3487 ( .A1(n3230), .A2(n3229), .ZN(n3335) );
  CLKBUF_X2 U3488 ( .A(n3200), .Z(n3273) );
  BUF_X2 U3489 ( .A(n3366), .Z(n4249) );
  OR2_X1 U3491 ( .A1(n5408), .A2(n6224), .ZN(n3045) );
  CLKBUF_X1 U3492 ( .A(n3548), .Z(n3549) );
  AND2_X1 U3493 ( .A1(n5436), .A2(n4290), .ZN(n4291) );
  OR2_X1 U3494 ( .A1(n5451), .A2(n5450), .ZN(n5804) );
  XNOR2_X1 U3495 ( .A(n4276), .B(n4275), .ZN(n4344) );
  AND2_X2 U3496 ( .A1(n5466), .A2(n5468), .ZN(n5460) );
  AND2_X1 U3497 ( .A1(n3079), .A2(n3077), .ZN(n3033) );
  OR2_X1 U3498 ( .A1(n5663), .A2(n3539), .ZN(n3079) );
  NAND2_X1 U3499 ( .A1(n5248), .A2(n5249), .ZN(n3529) );
  OAI22_X1 U3500 ( .A1(n5401), .A2(n5536), .B1(n5538), .B2(n5431), .ZN(n4365)
         );
  AND2_X1 U3501 ( .A1(n3069), .A2(n3068), .ZN(n3067) );
  NOR2_X1 U3502 ( .A1(n5292), .A2(n3065), .ZN(n3064) );
  AND2_X1 U3503 ( .A1(n3533), .A2(n3070), .ZN(n3069) );
  OR2_X1 U3504 ( .A1(n3074), .A2(n3534), .ZN(n3073) );
  OR2_X2 U3505 ( .A1(n5533), .A2(n5532), .ZN(n5535) );
  NAND2_X1 U3506 ( .A1(n3398), .A2(n3397), .ZN(n4370) );
  AND2_X1 U3507 ( .A1(n4433), .A2(n4434), .ZN(n4436) );
  CLKBUF_X1 U3508 ( .A(n4369), .Z(n5778) );
  XNOR2_X1 U3509 ( .A(n4503), .B(n4970), .ZN(n4372) );
  NAND2_X1 U3510 ( .A1(n3379), .A2(n3378), .ZN(n4503) );
  INV_X2 U3511 ( .A(n5350), .ZN(n3010) );
  OAI21_X1 U3512 ( .B1(n4873), .B2(n3581), .A(n3430), .ZN(n4440) );
  AOI21_X1 U3513 ( .B1(n4375), .B2(n6506), .A(n3346), .ZN(n3416) );
  NAND2_X1 U3514 ( .A1(n3062), .A2(n3310), .ZN(n3349) );
  NAND2_X1 U3515 ( .A1(n3309), .A2(n3423), .ZN(n3062) );
  INV_X1 U3516 ( .A(n3015), .ZN(n3351) );
  NAND2_X1 U3517 ( .A1(n3383), .A2(n3382), .ZN(n4970) );
  NAND2_X1 U3518 ( .A1(n3279), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3355) );
  AND2_X1 U3519 ( .A1(n3654), .A2(n3653), .ZN(n4628) );
  INV_X1 U3520 ( .A(n3018), .ZN(n4292) );
  NAND2_X1 U3521 ( .A1(n4449), .A2(n4345), .ZN(n3732) );
  OR2_X1 U3522 ( .A1(n3680), .A2(n4353), .ZN(n3717) );
  CLKBUF_X3 U3523 ( .A(n4353), .Z(n3027) );
  INV_X1 U3524 ( .A(n3330), .ZN(n3636) );
  CLKBUF_X1 U3525 ( .A(n3402), .Z(n4424) );
  NAND2_X1 U3526 ( .A1(n3716), .A2(n3026), .ZN(n4428) );
  OAI211_X1 U3527 ( .C1(n3263), .C2(n3233), .A(n3335), .B(n3255), .ZN(n3269)
         );
  AND2_X1 U3528 ( .A1(n3265), .A2(n3612), .ZN(n3402) );
  BUF_X2 U3529 ( .A(n3272), .Z(n4421) );
  OR2_X1 U3530 ( .A1(n3305), .A2(n3304), .ZN(n3428) );
  NAND2_X1 U3531 ( .A1(n3197), .A2(n3196), .ZN(n3331) );
  NOR2_X2 U3532 ( .A1(n3237), .A2(n4378), .ZN(n3778) );
  OR2_X1 U3533 ( .A1(n3293), .A2(n3292), .ZN(n3522) );
  NAND4_X1 U3534 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n3200)
         );
  AND4_X1 U3535 ( .A1(n3191), .A2(n3190), .A3(n3189), .A4(n3188), .ZN(n3197)
         );
  AND4_X1 U3536 ( .A1(n3140), .A2(n3139), .A3(n3138), .A4(n3137), .ZN(n3156)
         );
  AND2_X1 U3537 ( .A1(n3125), .A2(n3124), .ZN(n3135) );
  NAND2_X2 U3538 ( .A1(n3166), .A2(n3165), .ZN(n3237) );
  AND4_X1 U3539 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3217)
         );
  AND4_X1 U3540 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3166)
         );
  AND4_X1 U3541 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3219)
         );
  AND4_X1 U3542 ( .A1(n3204), .A2(n3203), .A3(n3202), .A4(n3201), .ZN(n3220)
         );
  AND4_X1 U3543 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3165)
         );
  AND4_X1 U3544 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3218)
         );
  AND4_X1 U3545 ( .A1(n3179), .A2(n3178), .A3(n3177), .A4(n3176), .ZN(n3185)
         );
  AND4_X1 U3546 ( .A1(n3119), .A2(n3118), .A3(n3117), .A4(n3116), .ZN(n3125)
         );
  AND4_X1 U3547 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3124)
         );
  AND4_X1 U3548 ( .A1(n3195), .A2(n3194), .A3(n3193), .A4(n3192), .ZN(n3196)
         );
  AND4_X1 U3549 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3153)
         );
  AND4_X1 U3550 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .ZN(n3186)
         );
  AND4_X1 U3551 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3154)
         );
  AND4_X1 U3552 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3187)
         );
  AND4_X1 U3553 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3155)
         );
  AND4_X1 U3554 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3184)
         );
  AND4_X1 U3555 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3134)
         );
  BUF_X2 U3556 ( .A(n4121), .Z(n4099) );
  BUF_X2 U3557 ( .A(n3242), .Z(n4223) );
  BUF_X2 U3558 ( .A(n3240), .Z(n4226) );
  BUF_X2 U3559 ( .A(n3241), .Z(n4248) );
  BUF_X2 U3560 ( .A(n3175), .Z(n4157) );
  BUF_X2 U3561 ( .A(n3248), .Z(n4181) );
  AND2_X2 U3562 ( .A1(n4606), .A2(n3127), .ZN(n4121) );
  BUF_X2 U3563 ( .A(n3251), .Z(n4225) );
  AND2_X2 U3564 ( .A1(n3129), .A2(n4446), .ZN(n3366) );
  AND2_X2 U3565 ( .A1(n3127), .A2(n4446), .ZN(n3247) );
  AND2_X2 U3566 ( .A1(n3128), .A2(n3129), .ZN(n3240) );
  BUF_X2 U3567 ( .A(n3250), .Z(n4250) );
  AND2_X2 U3568 ( .A1(n4606), .A2(n4588), .ZN(n3390) );
  AND2_X2 U3569 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4446) );
  CLKBUF_X1 U3570 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n6598) );
  AND2_X2 U3571 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4603) );
  NAND2_X1 U3572 ( .A1(n3066), .A2(n3014), .ZN(n3011) );
  AND2_X2 U3573 ( .A1(n3011), .A2(n3012), .ZN(n5359) );
  OR2_X1 U3574 ( .A1(n3013), .A2(n5353), .ZN(n3012) );
  INV_X1 U3575 ( .A(n3535), .ZN(n3013) );
  AND2_X1 U3576 ( .A1(n3063), .A2(n3535), .ZN(n3014) );
  AND2_X2 U3577 ( .A1(n3353), .A2(n3343), .ZN(n3015) );
  NAND2_X1 U3578 ( .A1(n3282), .A2(n3283), .ZN(n3016) );
  NAND2_X1 U3579 ( .A1(n3282), .A2(n3283), .ZN(n3352) );
  OR2_X1 U3580 ( .A1(n3406), .A2(n3405), .ZN(n3408) );
  NAND2_X4 U3581 ( .A1(n3512), .A2(n3523), .ZN(n5650) );
  NOR2_X2 U3582 ( .A1(n3333), .A2(n3332), .ZN(n3619) );
  NAND2_X1 U3583 ( .A1(n4372), .A2(n6506), .ZN(n3398) );
  AND2_X1 U3584 ( .A1(n3329), .A2(n3265), .ZN(n3017) );
  NAND2_X1 U3585 ( .A1(n3020), .A2(n3265), .ZN(n3018) );
  CLKBUF_X1 U3586 ( .A(n5001), .Z(n3019) );
  NOR2_X1 U3587 ( .A1(n3616), .A2(n3327), .ZN(n3020) );
  AOI21_X1 U3588 ( .B1(n4368), .B2(n3563), .A(n3415), .ZN(n3021) );
  INV_X4 U3589 ( .A(n3614), .ZN(n3265) );
  NAND2_X1 U3590 ( .A1(n3231), .A2(n3335), .ZN(n3616) );
  NOR2_X1 U3591 ( .A1(n3616), .A2(n3327), .ZN(n3605) );
  AOI21_X1 U3592 ( .B1(n4368), .B2(n3563), .A(n3415), .ZN(n6195) );
  NAND2_X1 U3593 ( .A1(n3080), .A2(n3404), .ZN(n3438) );
  OAI21_X1 U3594 ( .B1(n3409), .B2(n3793), .A(n4131), .ZN(n3805) );
  NOR2_X4 U3595 ( .A1(n5535), .A2(n3694), .ZN(n5529) );
  OR2_X1 U3596 ( .A1(n3355), .A2(n3088), .ZN(n3361) );
  XNOR2_X1 U3597 ( .A(n3417), .B(n3416), .ZN(n4369) );
  AND2_X2 U3598 ( .A1(n5381), .A2(n5386), .ZN(n5385) );
  NOR2_X2 U3599 ( .A1(n5329), .A2(n5382), .ZN(n5381) );
  AOI211_X1 U3600 ( .C1(n4375), .C2(n5789), .A(n5788), .B(n5787), .ZN(n6464)
         );
  AOI21_X1 U3601 ( .B1(n3417), .B2(n3416), .A(n3350), .ZN(n3405) );
  OAI22_X2 U3602 ( .A1(n5615), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5625), .B2(n5609), .ZN(n5610) );
  NOR2_X2 U3603 ( .A1(n4509), .A2(n4625), .ZN(n4624) );
  NOR2_X4 U3604 ( .A1(n4754), .A2(n4755), .ZN(n4753) );
  BUF_X1 U3606 ( .A(n3316), .Z(n3025) );
  OAI21_X2 U3607 ( .B1(n5460), .B2(n5461), .A(n5435), .ZN(n5811) );
  NAND2_X1 U3608 ( .A1(n3272), .A2(n3331), .ZN(n3680) );
  NOR2_X4 U3609 ( .A1(n5500), .A2(n5501), .ZN(n5492) );
  NAND2_X2 U3610 ( .A1(n5385), .A2(n3097), .ZN(n5500) );
  INV_X1 U3611 ( .A(n3410), .ZN(n3400) );
  INV_X1 U3612 ( .A(n5292), .ZN(n3068) );
  NOR2_X1 U3613 ( .A1(n4862), .A2(n3093), .ZN(n3092) );
  INV_X1 U3614 ( .A(n4710), .ZN(n3095) );
  INV_X1 U3615 ( .A(n5260), .ZN(n3074) );
  OR2_X1 U3616 ( .A1(n4473), .A2(n6501), .ZN(n3775) );
  NAND2_X1 U3617 ( .A1(n5012), .A2(n4292), .ZN(n4422) );
  AND2_X1 U3618 ( .A1(n5273), .A2(n3934), .ZN(n3096) );
  OR2_X1 U3619 ( .A1(n3495), .A2(n3494), .ZN(n3514) );
  OR2_X1 U3620 ( .A1(n3322), .A2(n3321), .ZN(n3418) );
  AND2_X1 U3621 ( .A1(n3614), .A2(n3331), .ZN(n3413) );
  OAI211_X1 U3622 ( .C1(n3355), .C2(n4454), .A(n3339), .B(n3340), .ZN(n3353)
         );
  AOI21_X1 U3623 ( .B1(n3260), .B2(n3259), .A(n4334), .ZN(n3261) );
  INV_X1 U3624 ( .A(n3331), .ZN(n3640) );
  NAND2_X1 U3625 ( .A1(n3614), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3385) );
  OR2_X1 U3626 ( .A1(n3233), .A2(n6506), .ZN(n3384) );
  NOR2_X1 U3627 ( .A1(n5437), .A2(n3099), .ZN(n3098) );
  INV_X1 U3628 ( .A(n5461), .ZN(n3099) );
  NOR2_X1 U3629 ( .A1(n5786), .A2(n6506), .ZN(n4266) );
  INV_X1 U3630 ( .A(n4266), .ZN(n4238) );
  INV_X1 U3631 ( .A(n3073), .ZN(n3065) );
  NAND2_X1 U3632 ( .A1(n4378), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4131) );
  NOR2_X1 U3633 ( .A1(n3078), .A2(n3032), .ZN(n3077) );
  INV_X1 U3634 ( .A(n3538), .ZN(n3078) );
  NAND2_X1 U3635 ( .A1(n3675), .A2(n3050), .ZN(n3052) );
  NOR2_X1 U3636 ( .A1(n5268), .A2(n5245), .ZN(n3050) );
  NAND2_X1 U3637 ( .A1(n3044), .A2(n3027), .ZN(n3708) );
  OR2_X1 U3638 ( .A1(n3372), .A2(n3371), .ZN(n3410) );
  NOR2_X1 U3639 ( .A1(n3613), .A2(n3615), .ZN(n3637) );
  INV_X1 U3640 ( .A(n3738), .ZN(n3267) );
  AND3_X1 U3641 ( .A1(n3236), .A2(n3276), .A3(n3235), .ZN(n3268) );
  INV_X1 U3642 ( .A(n3589), .ZN(n3374) );
  OAI21_X1 U3643 ( .B1(n6614), .B2(n4620), .A(n6592), .ZN(n4383) );
  AOI22_X1 U3644 ( .A1(n3249), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3061) );
  AND2_X1 U3645 ( .A1(n3238), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U3646 ( .A1(n3385), .A2(n3384), .ZN(n3597) );
  AND2_X1 U3647 ( .A1(n3596), .A2(n3595), .ZN(n3627) );
  OR2_X1 U3648 ( .A1(n3594), .A2(n3593), .ZN(n3596) );
  NAND2_X1 U3649 ( .A1(n3589), .A2(n3563), .ZN(n3601) );
  OR2_X1 U3650 ( .A1(n6594), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4277) );
  INV_X1 U3651 ( .A(n6079), .ZN(n5163) );
  OR2_X1 U3652 ( .A1(n6609), .A2(n4297), .ZN(n6080) );
  OR2_X1 U3653 ( .A1(n6273), .A2(n4295), .ZN(n4296) );
  AND2_X1 U3654 ( .A1(n3700), .A2(n3699), .ZN(n5512) );
  INV_X1 U3655 ( .A(n4131), .ZN(n4272) );
  NOR2_X1 U3656 ( .A1(n4213), .A2(n5576), .ZN(n4240) );
  AND2_X1 U3657 ( .A1(n5460), .A2(n3038), .ZN(n3101) );
  AND2_X1 U3658 ( .A1(n4034), .A2(n3037), .ZN(n3097) );
  NAND2_X1 U3659 ( .A1(n3997), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4029)
         );
  NAND2_X1 U3660 ( .A1(n3952), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3953)
         );
  OR2_X1 U3661 ( .A1(n5650), .A2(n5360), .ZN(n3536) );
  INV_X1 U3662 ( .A(n5331), .ZN(n3950) );
  NAND2_X1 U3663 ( .A1(n6179), .A2(n3510), .ZN(n5003) );
  NAND2_X1 U3664 ( .A1(n3060), .A2(n3458), .ZN(n4965) );
  NAND2_X1 U3665 ( .A1(n4965), .A2(n4964), .ZN(n4963) );
  INV_X1 U3666 ( .A(n3775), .ZN(n5012) );
  NOR2_X1 U3667 ( .A1(n3086), .A2(n5591), .ZN(n3085) );
  INV_X1 U3668 ( .A(n3109), .ZN(n3086) );
  AOI21_X1 U3669 ( .B1(n5644), .B2(n3107), .A(n5645), .ZN(n3545) );
  OR2_X1 U3670 ( .A1(n5336), .A2(n5335), .ZN(n5533) );
  NAND2_X1 U3671 ( .A1(n5317), .A2(n5316), .ZN(n5336) );
  NAND2_X1 U3672 ( .A1(n3072), .A2(n3071), .ZN(n3070) );
  NAND2_X1 U3673 ( .A1(n3675), .A2(n3674), .ZN(n5269) );
  NAND2_X1 U3674 ( .A1(n5650), .A2(n6238), .ZN(n5249) );
  INV_X1 U3675 ( .A(n6301), .ZN(n6279) );
  NAND2_X1 U3676 ( .A1(n5363), .A2(n3751), .ZN(n6257) );
  OAI21_X1 U3677 ( .B1(n3775), .B2(n3633), .A(n3632), .ZN(n3753) );
  NAND2_X1 U3678 ( .A1(n3408), .A2(n3407), .ZN(n3409) );
  CLKBUF_X1 U3679 ( .A(n3619), .Z(n3620) );
  INV_X1 U3680 ( .A(n5119), .ZN(n5111) );
  AND2_X1 U3681 ( .A1(n4839), .A2(n3023), .ZN(n5187) );
  AND2_X1 U3682 ( .A1(n4374), .A2(n6090), .ZN(n5068) );
  AND2_X1 U3683 ( .A1(n5778), .A2(n4873), .ZN(n4973) );
  AND2_X1 U3684 ( .A1(n4605), .A2(n4604), .ZN(n6488) );
  INV_X1 U3685 ( .A(n6082), .ZN(n5875) );
  AND2_X1 U3686 ( .A1(n6609), .A2(n4302), .ZN(n6067) );
  NAND2_X1 U3687 ( .A1(n5403), .A2(n5402), .ZN(n3049) );
  AND2_X1 U3688 ( .A1(n5400), .A2(n5405), .ZN(n3048) );
  AOI21_X1 U3689 ( .B1(n4359), .B2(n3059), .A(n4358), .ZN(n4364) );
  INV_X1 U3690 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6632) );
  NOR2_X2 U3691 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6367) );
  INV_X1 U3692 ( .A(n3023), .ZN(n5171) );
  INV_X1 U3693 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6479) );
  AND2_X2 U3694 ( .A1(n3088), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3129)
         );
  AND2_X2 U3695 ( .A1(n3111), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3128)
         );
  NAND2_X1 U3696 ( .A1(n3556), .A2(n3555), .ZN(n3586) );
  INV_X1 U3697 ( .A(n5029), .ZN(n3093) );
  NAND2_X1 U3698 ( .A1(n3461), .A2(n3460), .ZN(n3485) );
  OR2_X1 U3699 ( .A1(n3472), .A2(n3471), .ZN(n3502) );
  OR2_X1 U3700 ( .A1(n3449), .A2(n3448), .ZN(n3503) );
  NAND2_X1 U3701 ( .A1(n3255), .A2(n4564), .ZN(n3260) );
  NOR2_X1 U3702 ( .A1(n3324), .A2(n3323), .ZN(n3347) );
  AND2_X1 U3703 ( .A1(n3413), .A2(n3263), .ZN(n3264) );
  NOR2_X1 U3704 ( .A1(n3272), .A2(n3271), .ZN(n3328) );
  NAND2_X1 U3705 ( .A1(n4256), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3114)
         );
  AND2_X1 U3706 ( .A1(n3265), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U3707 ( .A1(n3241), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3240), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U3708 ( .A1(n3366), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3163) );
  AND2_X2 U3709 ( .A1(n3087), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3127)
         );
  OR3_X1 U3710 ( .A1(n3594), .A2(n6479), .A3(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n3622) );
  INV_X1 U3711 ( .A(n3604), .ZN(n4335) );
  INV_X1 U3712 ( .A(n4290), .ZN(n4217) );
  AND2_X1 U3713 ( .A1(n5492), .A2(n3039), .ZN(n5466) );
  NOR2_X1 U3714 ( .A1(n5480), .A2(n3091), .ZN(n3089) );
  INV_X1 U3715 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3779) );
  NOR2_X1 U3716 ( .A1(n5250), .A2(n3074), .ZN(n3071) );
  INV_X1 U3717 ( .A(n3534), .ZN(n3072) );
  NAND2_X1 U3718 ( .A1(n5650), .A2(n3526), .ZN(n3527) );
  NAND2_X1 U3719 ( .A1(n3055), .A2(n4513), .ZN(n3054) );
  INV_X1 U3720 ( .A(n4531), .ZN(n3055) );
  NAND2_X1 U3721 ( .A1(n3027), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3043)
         );
  INV_X1 U3722 ( .A(n3384), .ZN(n4337) );
  AOI21_X1 U3723 ( .B1(n4373), .B2(n6506), .A(n3373), .ZN(n3376) );
  INV_X1 U3724 ( .A(n5778), .ZN(n4810) );
  OR2_X1 U3725 ( .A1(n3396), .A2(n3395), .ZN(n3452) );
  AND2_X1 U3726 ( .A1(n3023), .A2(n4841), .ZN(n4812) );
  INV_X1 U3727 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6474) );
  AND2_X1 U3728 ( .A1(n3996), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3997)
         );
  AND2_X1 U3729 ( .A1(n3857), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3874)
         );
  AND2_X1 U3730 ( .A1(n3999), .A2(n3998), .ZN(n5524) );
  OR2_X1 U3731 ( .A1(n5818), .A2(n3818), .ZN(n4153) );
  INV_X1 U3732 ( .A(n4449), .ZN(n4343) );
  INV_X1 U3733 ( .A(n6168), .ZN(n4494) );
  OR2_X1 U3734 ( .A1(n4281), .A2(n5424), .ZN(n4282) );
  AND2_X1 U3735 ( .A1(n4245), .A2(n4244), .ZN(n5449) );
  OR2_X1 U3736 ( .A1(n5587), .A2(n3818), .ZN(n4195) );
  AND2_X1 U3737 ( .A1(n5808), .A2(n4242), .ZN(n4172) );
  AND2_X1 U3738 ( .A1(n4150), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4151)
         );
  NAND2_X1 U3739 ( .A1(n4151), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4193)
         );
  AND2_X1 U3740 ( .A1(n4084), .A2(n4083), .ZN(n5487) );
  NOR2_X1 U3741 ( .A1(n4065), .A2(n5640), .ZN(n4066) );
  NAND2_X1 U3742 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4110)
         );
  AND2_X1 U3743 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4030), .ZN(n4031)
         );
  INV_X1 U3744 ( .A(n4029), .ZN(n4030) );
  NAND2_X1 U3745 ( .A1(n4031), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4065)
         );
  AND2_X1 U3746 ( .A1(n4014), .A2(n4013), .ZN(n5518) );
  INV_X1 U3747 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6666) );
  AND2_X1 U3748 ( .A1(n3968), .A2(n3967), .ZN(n5382) );
  AND2_X1 U3749 ( .A1(n3935), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3952)
         );
  AOI21_X1 U3750 ( .B1(n3069), .B2(n3064), .A(n3042), .ZN(n3063) );
  NAND2_X1 U3751 ( .A1(n3529), .A2(n3067), .ZN(n3066) );
  NAND2_X1 U3752 ( .A1(n3903), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3919)
         );
  AND2_X1 U3753 ( .A1(n3889), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3903)
         );
  AND2_X1 U3754 ( .A1(n3874), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3889)
         );
  CLKBUF_X1 U3755 ( .A(n5241), .Z(n5242) );
  INV_X1 U3756 ( .A(n5102), .ZN(n3872) );
  AND2_X1 U3757 ( .A1(n3852), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3857)
         );
  CLKBUF_X1 U3758 ( .A(n5027), .Z(n5028) );
  NAND2_X1 U3759 ( .A1(n3826), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3827)
         );
  INV_X1 U3760 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3829) );
  NOR2_X1 U3761 ( .A1(n3827), .A2(n3829), .ZN(n3852) );
  INV_X1 U3762 ( .A(n4359), .ZN(n4360) );
  NAND2_X1 U3763 ( .A1(n3059), .A2(n3058), .ZN(n4359) );
  INV_X1 U3764 ( .A(n5454), .ZN(n3058) );
  NOR2_X1 U3765 ( .A1(n5562), .A2(n5672), .ZN(n5396) );
  NAND2_X1 U3766 ( .A1(n3548), .A2(n3082), .ZN(n5562) );
  NOR2_X1 U3767 ( .A1(n3084), .A2(n3083), .ZN(n3082) );
  INV_X1 U3768 ( .A(n3085), .ZN(n3084) );
  OR2_X1 U3769 ( .A1(n5464), .A2(n5438), .ZN(n5440) );
  NAND2_X1 U3770 ( .A1(n5472), .A2(n5462), .ZN(n5464) );
  NOR2_X2 U3771 ( .A1(n5485), .A2(n5475), .ZN(n5476) );
  XNOR2_X1 U3772 ( .A(n5650), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5599)
         );
  NAND2_X1 U3773 ( .A1(n5529), .A2(n3056), .ZN(n5496) );
  NOR2_X1 U3774 ( .A1(n3703), .A2(n3057), .ZN(n3056) );
  AOI21_X1 U3775 ( .B1(n3539), .B2(n3077), .A(n3035), .ZN(n3075) );
  AND2_X1 U3776 ( .A1(n3686), .A2(n3685), .ZN(n5335) );
  AND2_X1 U3777 ( .A1(n3683), .A2(n3682), .ZN(n5316) );
  NOR2_X2 U3778 ( .A1(n3052), .A2(n3051), .ZN(n5317) );
  NAND2_X1 U3779 ( .A1(n4963), .A2(n3482), .ZN(n6181) );
  NAND2_X1 U3780 ( .A1(n6181), .A2(n6180), .ZN(n6179) );
  AND2_X1 U3781 ( .A1(n3662), .A2(n3661), .ZN(n4950) );
  OR2_X1 U3782 ( .A1(n4530), .A2(n3054), .ZN(n4629) );
  NOR2_X1 U3783 ( .A1(n3746), .A2(n3744), .ZN(n4466) );
  CLKBUF_X1 U3784 ( .A(n4373), .Z(n4374) );
  OR2_X1 U3785 ( .A1(n3263), .A2(n3611), .ZN(n5786) );
  INV_X1 U3786 ( .A(n3016), .ZN(n3344) );
  NOR2_X1 U3787 ( .A1(n4977), .A2(n5778), .ZN(n4874) );
  INV_X1 U3788 ( .A(n4977), .ZN(n4974) );
  NAND2_X1 U3789 ( .A1(n4847), .A2(n4810), .ZN(n4817) );
  NOR2_X1 U3790 ( .A1(n3777), .A2(n4368), .ZN(n4847) );
  OR2_X1 U3791 ( .A1(n3355), .A2(n3087), .ZN(n3383) );
  INV_X1 U3792 ( .A(n4983), .ZN(n4843) );
  INV_X1 U3793 ( .A(n4763), .ZN(n4633) );
  AOI21_X1 U3794 ( .B1(n3175), .B2(INSTQUEUE_REG_1__2__SCAN_IN), .A(n3239), 
        .ZN(n3246) );
  INV_X1 U3795 ( .A(n4873), .ZN(n4872) );
  INV_X1 U3796 ( .A(n4565), .ZN(n4578) );
  AOI21_X1 U3797 ( .B1(n6632), .B2(STATE2_REG_3__SCAN_IN), .A(n4910), .ZN(
        n4983) );
  AND2_X1 U3798 ( .A1(n4368), .A2(n4371), .ZN(n4547) );
  AND2_X1 U3799 ( .A1(n3603), .A2(n3602), .ZN(n4473) );
  AND2_X1 U3800 ( .A1(n6784), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3604) );
  NOR2_X1 U3801 ( .A1(n6784), .A2(n4378), .ZN(n4620) );
  AND2_X1 U3802 ( .A1(n6367), .A2(n6784), .ZN(n5947) );
  INV_X1 U3803 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6365) );
  NOR2_X1 U3804 ( .A1(n5831), .A2(n4312), .ZN(n5816) );
  AND2_X1 U3805 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5869), .ZN(n5862) );
  NOR2_X1 U3806 ( .A1(n5989), .A2(n4308), .ZN(n5882) );
  INV_X1 U3807 ( .A(n6087), .ZN(n6075) );
  AND2_X1 U3808 ( .A1(n6080), .A2(n4306), .ZN(n6062) );
  AND2_X1 U3809 ( .A1(n4305), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4306) );
  AND2_X1 U3810 ( .A1(n6609), .A2(n4317), .ZN(n6054) );
  AND2_X1 U3811 ( .A1(n5033), .A2(n6024), .ZN(n5415) );
  NAND2_X1 U3812 ( .A1(n6609), .A2(n4304), .ZN(n6079) );
  INV_X1 U3813 ( .A(n5415), .ZN(n6098) );
  INV_X1 U3814 ( .A(n5433), .ZN(n5401) );
  NAND2_X1 U3815 ( .A1(n5529), .A2(n5514), .ZN(n5503) );
  NAND2_X2 U3816 ( .A1(n5538), .A2(n4334), .ZN(n5536) );
  INV_X1 U3817 ( .A(n5422), .ZN(n5544) );
  INV_X1 U3818 ( .A(n5886), .ZN(n6623) );
  INV_X1 U3819 ( .A(n5541), .ZN(n6620) );
  NAND2_X2 U3820 ( .A1(n5541), .A2(n4553), .ZN(n5886) );
  INV_X1 U3821 ( .A(n5383), .ZN(n5290) );
  AND2_X1 U3822 ( .A1(n5015), .A2(n5014), .ZN(n6131) );
  NAND2_X1 U3823 ( .A1(n6144), .A2(n5013), .ZN(n5015) );
  CLKBUF_X1 U3824 ( .A(n5060), .Z(n6612) );
  INV_X2 U3825 ( .A(n6111), .ZN(n6139) );
  NAND2_X1 U3826 ( .A1(n5012), .A2(n4339), .ZN(n6168) );
  AND2_X1 U3827 ( .A1(n3020), .A2(n4338), .ZN(n4339) );
  XNOR2_X1 U3828 ( .A(n5451), .B(n4349), .ZN(n5422) );
  INV_X1 U3829 ( .A(n4348), .ZN(n4349) );
  INV_X1 U3830 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5576) );
  INV_X1 U3831 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5626) );
  INV_X1 U3832 ( .A(n5899), .ZN(n6102) );
  CLKBUF_X1 U3833 ( .A(n5312), .Z(n5313) );
  OR2_X1 U3834 ( .A1(n6511), .A2(n6316), .ZN(n6211) );
  INV_X1 U3835 ( .A(n5903), .ZN(n6208) );
  AND2_X1 U3836 ( .A1(n3549), .A2(n3085), .ZN(n5584) );
  OR2_X1 U3837 ( .A1(n5721), .A2(n3765), .ZN(n5705) );
  NOR2_X1 U3838 ( .A1(n5724), .A2(n3767), .ZN(n5712) );
  OR2_X1 U3839 ( .A1(n5916), .A2(n3758), .ZN(n5904) );
  NOR2_X1 U3840 ( .A1(n5364), .A2(n5932), .ZN(n5916) );
  OAI21_X1 U3841 ( .B1(n3529), .B2(n3073), .A(n3069), .ZN(n5294) );
  NAND2_X1 U3842 ( .A1(n5261), .A2(n5260), .ZN(n6170) );
  CLKBUF_X1 U3843 ( .A(n5105), .Z(n5246) );
  OR2_X1 U3844 ( .A1(n6257), .A2(n6279), .ZN(n6260) );
  INV_X1 U3845 ( .A(n4375), .ZN(n6090) );
  AND2_X1 U3846 ( .A1(n5778), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5781) );
  INV_X1 U3847 ( .A(n6367), .ZN(n6316) );
  OAI21_X1 U3848 ( .B1(n4613), .B2(n6589), .A(n4910), .ZN(n6312) );
  INV_X1 U3849 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6463) );
  INV_X1 U3850 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6784) );
  AND2_X1 U3851 ( .A1(n4386), .A2(n4385), .ZN(n4734) );
  OAI21_X1 U3852 ( .B1(n6322), .B2(n6338), .A(n6321), .ZN(n6340) );
  OAI21_X1 U3853 ( .B1(n5075), .B2(n6591), .A(n5067), .ZN(n5094) );
  OAI211_X1 U3854 ( .C1(n5188), .C2(n5187), .A(n6321), .B(n5186), .ZN(n5225)
         );
  AOI22_X1 U3855 ( .A1(n5182), .A2(n5187), .B1(n6360), .B2(n5181), .ZN(n5233)
         );
  NAND2_X1 U3856 ( .A1(n4847), .A2(n4973), .ZN(n6458) );
  NOR2_X1 U3857 ( .A1(n6151), .A2(n4910), .ZN(n6433) );
  INV_X1 U3858 ( .A(n5220), .ZN(n6432) );
  NOR2_X1 U3859 ( .A1(n6153), .A2(n4910), .ZN(n6418) );
  INV_X1 U3860 ( .A(n5215), .ZN(n6417) );
  NOR2_X1 U3861 ( .A1(n6155), .A2(n4910), .ZN(n6382) );
  INV_X1 U3862 ( .A(n5210), .ZN(n6383) );
  NOR2_X1 U3863 ( .A1(n4502), .A2(n4910), .ZN(n6439) );
  INV_X1 U3864 ( .A(n5227), .ZN(n6438) );
  NOR2_X1 U3865 ( .A1(n6158), .A2(n4910), .ZN(n6445) );
  NOR2_X1 U3866 ( .A1(n6160), .A2(n4910), .ZN(n6396) );
  NOR2_X1 U3867 ( .A1(n6162), .A2(n4910), .ZN(n6454) );
  INV_X1 U3868 ( .A(n5195), .ZN(n6452) );
  NOR2_X1 U3869 ( .A1(n6164), .A2(n4910), .ZN(n6407) );
  INV_X1 U3870 ( .A(n5200), .ZN(n6409) );
  INV_X1 U3871 ( .A(n6433), .ZN(n5224) );
  INV_X1 U3872 ( .A(n6418), .ZN(n5219) );
  INV_X1 U3873 ( .A(n6439), .ZN(n5232) );
  AND2_X1 U3874 ( .A1(n4547), .A2(n4872), .ZN(n4737) );
  INV_X1 U3875 ( .A(n6396), .ZN(n5209) );
  INV_X1 U3876 ( .A(n6407), .ZN(n5204) );
  INV_X1 U3877 ( .A(n4677), .ZN(n4660) );
  INV_X1 U3878 ( .A(n6503), .ZN(n6501) );
  AND3_X1 U3879 ( .A1(n6489), .A2(n6488), .A3(n6487), .ZN(n6502) );
  OR2_X1 U3880 ( .A1(n6591), .A2(n4473), .ZN(n6592) );
  INV_X1 U3881 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6506) );
  AND2_X1 U3882 ( .A1(n3604), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6503) );
  NOR2_X1 U3883 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6614) );
  INV_X1 U3884 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6591) );
  INV_X1 U3885 ( .A(n6510), .ZN(n6590) );
  OR2_X1 U3886 ( .A1(n5683), .A2(n6093), .ZN(n4322) );
  AOI211_X1 U3887 ( .C1(n6173), .C2(n5580), .A(n5579), .B(n5578), .ZN(n5581)
         );
  NAND2_X1 U3888 ( .A1(n3046), .A2(n3045), .ZN(U2988) );
  AOI21_X1 U3889 ( .B1(n5433), .B2(n6290), .A(n3047), .ZN(n3046) );
  NAND2_X1 U3890 ( .A1(n3049), .A2(n3048), .ZN(n3047) );
  INV_X1 U3891 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U3892 ( .A1(n5385), .A2(n3037), .ZN(n5509) );
  NAND2_X1 U3893 ( .A1(n5492), .A2(n3090), .ZN(n5479) );
  NAND2_X1 U3894 ( .A1(n5256), .A2(n5273), .ZN(n5272) );
  AND4_X1 U3895 ( .A1(n3243), .A2(n3252), .A3(n3244), .A4(n3253), .ZN(n3028)
         );
  NAND2_X1 U3896 ( .A1(n3079), .A2(n3538), .ZN(n5651) );
  NAND2_X1 U3897 ( .A1(n5492), .A2(n3089), .ZN(n3029) );
  INV_X1 U3898 ( .A(n3059), .ZN(n5453) );
  NOR2_X1 U3899 ( .A1(n5440), .A2(n4299), .ZN(n3059) );
  NAND2_X1 U3900 ( .A1(n3361), .A2(n3360), .ZN(n3378) );
  NAND2_X1 U3901 ( .A1(n3640), .A2(n3265), .ZN(n3716) );
  INV_X1 U3902 ( .A(n3716), .ZN(n3044) );
  AND2_X1 U3903 ( .A1(n5492), .A2(n5493), .ZN(n3030) );
  AND2_X1 U3904 ( .A1(n5385), .A2(n5524), .ZN(n3031) );
  OR2_X1 U3905 ( .A1(n4291), .A2(n3101), .ZN(n5577) );
  AND2_X2 U3906 ( .A1(n4446), .A2(n4603), .ZN(n3238) );
  AND2_X1 U3907 ( .A1(n5650), .A2(n3540), .ZN(n3032) );
  INV_X1 U3908 ( .A(n3200), .ZN(n3325) );
  NAND2_X1 U3909 ( .A1(n5570), .A2(n5599), .ZN(n3548) );
  INV_X1 U3910 ( .A(n5245), .ZN(n3674) );
  AND2_X1 U3911 ( .A1(n3708), .A2(n3043), .ZN(n3034) );
  NOR2_X1 U3912 ( .A1(n5650), .A2(n3541), .ZN(n3035) );
  AND3_X1 U3913 ( .A1(n3245), .A2(n3254), .A3(n3061), .ZN(n3036) );
  NAND2_X1 U3914 ( .A1(n3612), .A2(n3614), .ZN(n3561) );
  NAND2_X1 U3915 ( .A1(n3459), .A2(n3399), .ZN(n3777) );
  OR2_X1 U3916 ( .A1(n4710), .A2(n4862), .ZN(n4861) );
  NAND2_X1 U3917 ( .A1(n3529), .A2(n5250), .ZN(n5261) );
  AND2_X1 U3918 ( .A1(n5518), .A2(n5524), .ZN(n3037) );
  NAND2_X1 U3919 ( .A1(n3066), .A2(n3063), .ZN(n5352) );
  AND2_X1 U3920 ( .A1(n5241), .A2(n5257), .ZN(n5256) );
  AND2_X1 U3921 ( .A1(n4217), .A2(n3098), .ZN(n3038) );
  INV_X1 U3922 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3087) );
  NOR2_X1 U3923 ( .A1(n4861), .A2(n4948), .ZN(n5026) );
  INV_X1 U3924 ( .A(n3091), .ZN(n3090) );
  NAND2_X1 U3925 ( .A1(n5487), .A2(n5493), .ZN(n3091) );
  AND2_X1 U3926 ( .A1(n3022), .A2(n4421), .ZN(n3563) );
  INV_X1 U3927 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3088) );
  AND2_X1 U3928 ( .A1(n4134), .A2(n3089), .ZN(n3039) );
  AND2_X1 U3929 ( .A1(n3038), .A2(n5449), .ZN(n3040) );
  AND2_X1 U3930 ( .A1(n3753), .A2(n3733), .ZN(n6290) );
  NOR2_X1 U3931 ( .A1(n4530), .A2(n4531), .ZN(n3041) );
  AND2_X1 U3932 ( .A1(n5650), .A2(n5304), .ZN(n3042) );
  INV_X1 U3933 ( .A(n3259), .ZN(n3609) );
  INV_X1 U3934 ( .A(n5514), .ZN(n3057) );
  NAND2_X1 U3935 ( .A1(n3105), .A2(n3640), .ZN(n4352) );
  INV_X1 U3936 ( .A(n3335), .ZN(n4334) );
  INV_X1 U3937 ( .A(n5673), .ZN(n3083) );
  INV_X2 U3938 ( .A(n3027), .ZN(n4438) );
  INV_X1 U3939 ( .A(n3052), .ZN(n5276) );
  INV_X1 U3940 ( .A(n5275), .ZN(n3051) );
  OR2_X2 U3941 ( .A1(n4530), .A2(n3053), .ZN(n4754) );
  OR2_X2 U3942 ( .A1(n3054), .A2(n4628), .ZN(n3053) );
  NOR2_X2 U3943 ( .A1(n5496), .A2(n5495), .ZN(n5489) );
  OAI21_X1 U3944 ( .B1(n6189), .B2(n6188), .A(n3060), .ZN(n6190) );
  NAND2_X1 U3945 ( .A1(n6189), .A2(n6188), .ZN(n3060) );
  NAND2_X1 U3946 ( .A1(n5003), .A2(n5002), .ZN(n5001) );
  NAND3_X1 U3947 ( .A1(n3246), .A2(n3028), .A3(n3036), .ZN(n3259) );
  NAND2_X1 U3948 ( .A1(n3062), .A2(n3426), .ZN(n4873) );
  NAND2_X1 U3949 ( .A1(n5663), .A2(n3077), .ZN(n3076) );
  NAND3_X1 U3950 ( .A1(n3459), .A2(n3563), .A3(n3399), .ZN(n3080) );
  INV_X1 U3951 ( .A(n3407), .ZN(n3081) );
  NAND2_X1 U3952 ( .A1(n3548), .A2(n3109), .ZN(n5392) );
  AND3_X4 U3953 ( .A1(n3136), .A2(n3134), .A3(n3135), .ZN(n3614) );
  INV_X2 U3954 ( .A(n3409), .ZN(n4368) );
  INV_X1 U3955 ( .A(n4948), .ZN(n3094) );
  NAND3_X1 U3956 ( .A1(n3095), .A2(n3094), .A3(n3092), .ZN(n5027) );
  NAND2_X1 U3957 ( .A1(n5256), .A2(n3096), .ZN(n5312) );
  INV_X1 U3958 ( .A(n5312), .ZN(n3951) );
  AND2_X1 U3959 ( .A1(n5460), .A2(n3098), .ZN(n4289) );
  NAND2_X1 U3960 ( .A1(n5460), .A2(n5461), .ZN(n5435) );
  AND2_X1 U3961 ( .A1(n5460), .A2(n3040), .ZN(n5451) );
  OAI21_X2 U3962 ( .B1(n5359), .B2(n3537), .A(n3536), .ZN(n5663) );
  NAND2_X1 U3963 ( .A1(n3311), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U3964 ( .A1(n3311), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3158) );
  INV_X1 U3965 ( .A(n4289), .ZN(n5436) );
  AND2_X1 U3966 ( .A1(n4334), .A2(n5541), .ZN(n3100) );
  INV_X1 U3967 ( .A(READY_N), .ZN(n6611) );
  INV_X2 U3968 ( .A(n6211), .ZN(n6184) );
  INV_X1 U3969 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4507) );
  NOR2_X1 U3970 ( .A1(n6360), .A2(n4377), .ZN(n3102) );
  AND3_X1 U3971 ( .A1(n5713), .A2(n5728), .A3(n5607), .ZN(n3103) );
  OR2_X1 U3972 ( .A1(n3341), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3104)
         );
  AND2_X1 U3973 ( .A1(n3325), .A2(n3609), .ZN(n3105) );
  AND3_X1 U3974 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5445), .A3(n6673), .ZN(n3106) );
  AND3_X1 U3975 ( .A1(n3544), .A2(n3543), .A3(n3542), .ZN(n3107) );
  INV_X1 U3976 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3435) );
  INV_X1 U3977 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5618) );
  AND2_X1 U3978 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n3027), .ZN(n3108)
         );
  INV_X1 U3979 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4192) );
  OR2_X1 U3980 ( .A1(n5645), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3109)
         );
  NAND2_X2 U3981 ( .A1(n5012), .A2(n4408), .ZN(n6178) );
  INV_X1 U3982 ( .A(n6178), .ZN(n6206) );
  INV_X1 U3983 ( .A(n4478), .ZN(n6143) );
  INV_X1 U3984 ( .A(n6143), .ZN(n4498) );
  NOR2_X1 U3985 ( .A1(n3335), .A2(n4378), .ZN(n3794) );
  INV_X1 U3986 ( .A(n6024), .ZN(n4331) );
  INV_X1 U3987 ( .A(n5744), .ZN(n3543) );
  AND2_X1 U3988 ( .A1(n5329), .A2(n5382), .ZN(n3110) );
  NAND2_X2 U3989 ( .A1(n4357), .A2(n4356), .ZN(n5538) );
  AND2_X1 U3990 ( .A1(n5538), .A2(n3335), .ZN(n5350) );
  INV_X1 U3991 ( .A(n3765), .ZN(n3542) );
  AND2_X1 U3992 ( .A1(n6632), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3564)
         );
  INV_X1 U3993 ( .A(n4277), .ZN(n3359) );
  AND2_X1 U3994 ( .A1(n6479), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3593)
         );
  INV_X1 U3995 ( .A(n5511), .ZN(n4034) );
  INV_X1 U3996 ( .A(n3418), .ZN(n3345) );
  INV_X1 U3997 ( .A(n3280), .ZN(n3281) );
  INV_X1 U3998 ( .A(n3459), .ZN(n3461) );
  AOI22_X1 U3999 ( .A1(n3175), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3251), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3160) );
  OR2_X1 U4000 ( .A1(n4127), .A2(n4126), .ZN(n4145) );
  INV_X1 U4001 ( .A(n5314), .ZN(n3934) );
  NOR2_X2 U4002 ( .A1(n3485), .A2(n3484), .ZN(n3498) );
  OR2_X1 U4003 ( .A1(n3627), .A2(n3626), .ZN(n4406) );
  INV_X1 U4004 ( .A(n5474), .ZN(n4134) );
  OR2_X1 U4005 ( .A1(n4110), .A2(n5626), .ZN(n4111) );
  NOR2_X1 U4006 ( .A1(n3953), .A2(n6666), .ZN(n3996) );
  INV_X1 U4007 ( .A(n3794), .ZN(n3839) );
  XNOR2_X1 U4008 ( .A(n3459), .B(n3460), .ZN(n3821) );
  NAND2_X1 U4009 ( .A1(n3498), .A2(n3499), .ZN(n3512) );
  NAND2_X1 U4010 ( .A1(n4538), .A2(n4540), .ZN(n4539) );
  MUX2_X1 U4011 ( .A(n3716), .B(n3717), .S(n6095), .Z(n3641) );
  NAND2_X1 U4012 ( .A1(n4438), .A2(n3026), .ZN(n3720) );
  OR2_X1 U4013 ( .A1(n5860), .A2(n3818), .ZN(n4068) );
  OR3_X1 U4014 ( .A1(n4193), .A2(n5595), .A3(n4192), .ZN(n4213) );
  NOR2_X1 U4015 ( .A1(n4111), .A2(n5618), .ZN(n4150) );
  INV_X1 U4016 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3918) );
  INV_X1 U4017 ( .A(n3818), .ZN(n4242) );
  NOR2_X1 U4018 ( .A1(n3798), .A2(n3779), .ZN(n3810) );
  AND3_X1 U4019 ( .A1(n4337), .A2(n3563), .A3(n3522), .ZN(n3523) );
  OR2_X1 U4020 ( .A1(n5650), .A2(n3531), .ZN(n3532) );
  OR2_X1 U4021 ( .A1(n4374), .A2(n4375), .ZN(n5119) );
  OR2_X1 U4022 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  NAND2_X1 U4023 ( .A1(n4359), .A2(n3026), .ZN(n4363) );
  NAND2_X1 U4024 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5986), .ZN(n5989) );
  NOR2_X1 U4025 ( .A1(n3919), .A2(n3918), .ZN(n3935) );
  OR2_X1 U4026 ( .A1(n6496), .A2(n4296), .ZN(n4297) );
  INV_X1 U4027 ( .A(n3561), .ZN(n5032) );
  AND2_X1 U4028 ( .A1(n4069), .A2(n4068), .ZN(n5493) );
  AND2_X1 U4029 ( .A1(n4154), .A2(n4153), .ZN(n5468) );
  XNOR2_X1 U4030 ( .A(n4282), .B(n4328), .ZN(n4305) );
  INV_X1 U4031 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5595) );
  INV_X1 U4032 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5640) );
  AND2_X1 U4033 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3810), .ZN(n3826)
         );
  AND2_X1 U4034 ( .A1(n5392), .A2(n5394), .ZN(n5395) );
  OR2_X1 U4035 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5592)
         );
  AND2_X1 U4036 ( .A1(n6169), .A2(n3532), .ZN(n3533) );
  INV_X1 U4037 ( .A(n6282), .ZN(n6302) );
  AND2_X1 U4038 ( .A1(n4787), .A2(n6343), .ZN(n4788) );
  NAND2_X1 U4039 ( .A1(n3425), .A2(n3424), .ZN(n3426) );
  NAND2_X1 U4040 ( .A1(n4368), .A2(n4614), .ZN(n4977) );
  INV_X1 U4041 ( .A(n6424), .ZN(n5155) );
  INV_X1 U4042 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6467) );
  OR2_X1 U4043 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3818) );
  OR2_X1 U4044 ( .A1(n4402), .A2(n6501), .ZN(n4416) );
  NAND2_X1 U4045 ( .A1(n4422), .A2(n4416), .ZN(n6609) );
  NOR2_X1 U4046 ( .A1(n3106), .A2(n4320), .ZN(n4321) );
  NOR2_X1 U4047 ( .A1(n6568), .A2(n5840), .ZN(n5836) );
  NOR3_X1 U4048 ( .A1(n6562), .A2(n5972), .A3(n6560), .ZN(n5869) );
  AND2_X1 U4049 ( .A1(n5163), .A2(n4307), .ZN(n5986) );
  OR2_X1 U4050 ( .A1(n6086), .A2(n4949), .ZN(n6018) );
  NOR2_X1 U4051 ( .A1(n4305), .A2(n6784), .ZN(n4298) );
  AND2_X1 U4052 ( .A1(n6080), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U4053 ( .A1(n6079), .A2(n6080), .ZN(n6082) );
  INV_X1 U4054 ( .A(n5536), .ZN(n5515) );
  AND2_X1 U4055 ( .A1(n5541), .A2(n5540), .ZN(n6621) );
  AND2_X1 U4056 ( .A1(n5541), .A2(n4554), .ZN(n5383) );
  NOR2_X1 U4057 ( .A1(n6508), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5060) );
  INV_X1 U4058 ( .A(n6144), .ZN(n6165) );
  OAI21_X1 U4059 ( .B1(n4424), .B2(n6611), .A(n4423), .ZN(n4478) );
  INV_X1 U4060 ( .A(n5841), .ZN(n5621) );
  INV_X1 U4061 ( .A(n5633), .ZN(n6624) );
  INV_X1 U4062 ( .A(n6202), .ZN(n6173) );
  AND2_X1 U4063 ( .A1(n3637), .A2(n3636), .ZN(n4408) );
  NOR2_X1 U4064 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NOR2_X1 U4065 ( .A1(n5705), .A2(n5679), .ZN(n5695) );
  OR2_X1 U4066 ( .A1(n5734), .A2(n3764), .ZN(n5724) );
  NOR2_X1 U4067 ( .A1(n5904), .A2(n3750), .ZN(n5739) );
  INV_X1 U4068 ( .A(n5650), .ZN(n5645) );
  NOR2_X1 U4069 ( .A1(n5363), .A2(n5302), .ZN(n5932) );
  INV_X1 U4070 ( .A(n6302), .ZN(n6273) );
  AND2_X1 U4071 ( .A1(n5947), .A2(n6506), .ZN(n6282) );
  AND2_X1 U4072 ( .A1(n6257), .A2(n4518), .ZN(n6297) );
  INV_X1 U4073 ( .A(n6224), .ZN(n6307) );
  NAND2_X1 U4074 ( .A1(n6506), .A2(n4383), .ZN(n4910) );
  OR2_X1 U4075 ( .A1(n4672), .A2(n4872), .ZN(n4745) );
  OAI21_X1 U4076 ( .B1(n6367), .B2(n4671), .A(n4670), .ZN(n4751) );
  INV_X1 U4077 ( .A(n4743), .ZN(n6339) );
  AND2_X1 U4078 ( .A1(n3777), .A2(n3409), .ZN(n4792) );
  AND2_X1 U4079 ( .A1(n4792), .A2(n4975), .ZN(n6349) );
  INV_X1 U4080 ( .A(n6366), .ZN(n6410) );
  NOR2_X1 U4081 ( .A1(n4977), .A2(n4976), .ZN(n6424) );
  NOR2_X2 U4082 ( .A1(n4817), .A2(n4872), .ZN(n5158) );
  INV_X1 U4083 ( .A(n5177), .ZN(n5229) );
  INV_X1 U4084 ( .A(n4947), .ZN(n6450) );
  OR3_X1 U4085 ( .A1(n4913), .A2(n4912), .A3(n5114), .ZN(n4940) );
  AND2_X1 U4086 ( .A1(n5778), .A2(n4872), .ZN(n4975) );
  INV_X1 U4087 ( .A(n5205), .ZN(n6397) );
  INV_X1 U4088 ( .A(n6448), .ZN(n6392) );
  OAI211_X1 U4089 ( .C1(n4638), .C2(n4637), .A(n6371), .B(n4636), .ZN(n4681)
         );
  INV_X1 U4090 ( .A(n6442), .ZN(n6388) );
  AND2_X1 U4091 ( .A1(n6506), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4294) );
  INV_X1 U4092 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6803) );
  AND2_X1 U4093 ( .A1(n4322), .A2(n4321), .ZN(n4323) );
  INV_X1 U4094 ( .A(n6067), .ZN(n6093) );
  NAND2_X1 U4095 ( .A1(n6080), .A2(n4298), .ZN(n6024) );
  INV_X1 U4096 ( .A(n6054), .ZN(n6094) );
  OAI211_X2 U4097 ( .C1(n4343), .C2(n4351), .A(n6168), .B(n4342), .ZN(n5541)
         );
  OR2_X1 U4098 ( .A1(n6612), .A2(n6131), .ZN(n6111) );
  NAND2_X1 U4099 ( .A1(n6131), .A2(n3265), .ZN(n6108) );
  INV_X1 U4100 ( .A(n6131), .ZN(n6141) );
  OR2_X1 U4101 ( .A1(n4422), .A2(n4421), .ZN(n6144) );
  NAND2_X1 U4102 ( .A1(n6178), .A2(n4278), .ZN(n5903) );
  NAND2_X1 U4103 ( .A1(n5903), .A2(n6207), .ZN(n6202) );
  INV_X1 U4104 ( .A(n6290), .ZN(n6304) );
  NAND2_X1 U4105 ( .A1(n3753), .A2(n3639), .ZN(n6224) );
  INV_X1 U4106 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6359) );
  AND2_X1 U4107 ( .A1(n4666), .A2(n4665), .ZN(n4749) );
  NAND2_X1 U4108 ( .A1(n4792), .A2(n4973), .ZN(n6356) );
  NAND2_X1 U4109 ( .A1(n4874), .A2(n4873), .ZN(n5100) );
  NAND2_X1 U4110 ( .A1(n4974), .A2(n4973), .ZN(n6430) );
  AOI211_X2 U4111 ( .C1(n5117), .C2(n5116), .A(n5115), .B(n5114), .ZN(n5162)
         );
  NAND2_X1 U4112 ( .A1(n4811), .A2(n4872), .ZN(n5177) );
  INV_X1 U4113 ( .A(n6454), .ZN(n5199) );
  INV_X1 U4114 ( .A(n6382), .ZN(n5214) );
  NAND2_X1 U4115 ( .A1(n4847), .A2(n4975), .ZN(n4947) );
  NAND2_X1 U4116 ( .A1(n4633), .A2(n4872), .ZN(n4783) );
  INV_X1 U4117 ( .A(n6445), .ZN(n5194) );
  INV_X1 U4118 ( .A(n4737), .ZN(n4585) );
  AND2_X1 U4119 ( .A1(n6495), .A2(n6494), .ZN(n6510) );
  INV_X1 U4120 ( .A(n6588), .ZN(n6513) );
  OR2_X1 U4121 ( .A1(n3606), .A2(STATE_REG_0__SCAN_IN), .ZN(n6520) );
  INV_X1 U4122 ( .A(n6577), .ZN(n6583) );
  OAI21_X1 U4123 ( .B1(n5577), .B2(n6024), .A(n4323), .ZN(U2799) );
  NAND2_X1 U4124 ( .A1(n4367), .A2(n4366), .ZN(U2829) );
  AND2_X2 U4125 ( .A1(n4454), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3126)
         );
  AND2_X4 U4126 ( .A1(n3126), .A2(n4603), .ZN(n3316) );
  NAND2_X1 U4127 ( .A1(n3024), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3115)
         );
  INV_X1 U4128 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3111) );
  AND2_X4 U4129 ( .A1(n3128), .A2(n4603), .ZN(n3462) );
  BUF_X4 U4130 ( .A(n3462), .Z(n4256) );
  AND2_X2 U4131 ( .A1(n3126), .A2(n3129), .ZN(n3248) );
  NAND2_X1 U4132 ( .A1(n3248), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U4133 ( .A1(n3247), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3112) );
  AND2_X2 U4135 ( .A1(n3126), .A2(n4588), .ZN(n3175) );
  NAND2_X1 U4136 ( .A1(n3175), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3119) );
  AND2_X4 U4137 ( .A1(n3127), .A2(n3128), .ZN(n3311) );
  NAND2_X1 U4138 ( .A1(n3311), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3118) );
  AND2_X2 U4139 ( .A1(n3128), .A2(n4588), .ZN(n3242) );
  NAND2_X1 U4140 ( .A1(n3242), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3117) );
  AND2_X2 U4141 ( .A1(n4588), .A2(n4446), .ZN(n3251) );
  NAND2_X1 U4142 ( .A1(n3251), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3116) );
  NOR2_X4 U4143 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U4144 ( .A1(n4121), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U4145 ( .A1(n3390), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3122) );
  AND2_X2 U4146 ( .A1(n4606), .A2(n4603), .ZN(n3250) );
  NAND2_X1 U4147 ( .A1(n3250), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3121)
         );
  NAND2_X1 U4148 ( .A1(n3238), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3120)
         );
  AND2_X2 U4149 ( .A1(n3127), .A2(n3126), .ZN(n3241) );
  NAND2_X1 U4150 ( .A1(n3241), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U4151 ( .A1(n3240), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3132)
         );
  NAND2_X1 U4152 ( .A1(n3366), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3131)
         );
  AND2_X2 U4153 ( .A1(n3129), .A2(n4606), .ZN(n3249) );
  NAND2_X1 U4154 ( .A1(n3249), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U4155 ( .A1(n3025), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3140)
         );
  NAND2_X1 U4156 ( .A1(n3242), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U4157 ( .A1(n3311), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U4158 ( .A1(n4256), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3137)
         );
  NAND2_X1 U4159 ( .A1(n3366), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3144)
         );
  NAND2_X1 U4160 ( .A1(n3249), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U4161 ( .A1(n4121), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4162 ( .A1(n3390), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U4163 ( .A1(n3175), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4164 ( .A1(n3248), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U4165 ( .A1(n3247), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4166 ( .A1(n3251), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U4167 ( .A1(n3241), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U4168 ( .A1(n3240), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3151)
         );
  NAND2_X1 U4169 ( .A1(n3238), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3150)
         );
  NAND2_X1 U4170 ( .A1(n3250), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3149)
         );
  INV_X2 U4171 ( .A(n3402), .ZN(n3412) );
  AOI22_X1 U4172 ( .A1(n3248), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4173 ( .A1(n3316), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4174 ( .A1(n3250), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3238), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4175 ( .A1(n4121), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U4176 ( .A1(n3248), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U4177 ( .A1(n3251), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U4178 ( .A1(n3238), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3168)
         );
  NAND2_X1 U4179 ( .A1(n3250), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3167)
         );
  NAND2_X1 U4180 ( .A1(n3249), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3174) );
  NAND2_X1 U4181 ( .A1(n3241), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3173) );
  NAND2_X1 U4182 ( .A1(n3390), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3172) );
  NAND2_X1 U4183 ( .A1(n3366), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3171)
         );
  NAND2_X1 U4184 ( .A1(n3175), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U4185 ( .A1(n3247), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U4186 ( .A1(n3240), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3177)
         );
  NAND2_X1 U4187 ( .A1(n4121), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4188 ( .A1(n3316), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3183)
         );
  NAND2_X1 U4189 ( .A1(n3242), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U4190 ( .A1(n3462), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3180)
         );
  NAND2_X2 U4191 ( .A1(n3790), .A2(n3273), .ZN(n3263) );
  NAND2_X1 U4192 ( .A1(n6784), .A2(n6591), .ZN(n6594) );
  INV_X1 U4193 ( .A(n6594), .ZN(n5411) );
  OAI211_X1 U4194 ( .C1(n3412), .C2(n3263), .A(STATE2_REG_0__SCAN_IN), .B(
        n5411), .ZN(n3199) );
  AOI22_X1 U4195 ( .A1(n3175), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3251), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4196 ( .A1(n3316), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4197 ( .A1(n3248), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4198 ( .A1(n3311), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4199 ( .A1(n3241), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3240), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4200 ( .A1(n3366), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4201 ( .A1(n3250), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3238), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4202 ( .A1(n4121), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3192) );
  AOI21_X1 U4203 ( .B1(n3412), .B2(n3237), .A(n3331), .ZN(n3198) );
  NOR2_X1 U4204 ( .A1(n3199), .A2(n3198), .ZN(n3236) );
  NAND2_X1 U4205 ( .A1(n3248), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4206 ( .A1(n3175), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4207 ( .A1(n3247), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4208 ( .A1(n3251), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4209 ( .A1(n3316), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3208)
         );
  NAND2_X1 U4210 ( .A1(n3242), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U4211 ( .A1(n3311), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4212 ( .A1(n3462), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3205)
         );
  NAND2_X1 U4213 ( .A1(n3366), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3212)
         );
  NAND2_X1 U4214 ( .A1(n3249), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4215 ( .A1(n4121), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4216 ( .A1(n3390), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4217 ( .A1(n3238), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4218 ( .A1(n3240), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3215)
         );
  NAND2_X1 U4219 ( .A1(n3241), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4220 ( .A1(n3250), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3213)
         );
  NAND4_X2 U4221 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3233)
         );
  INV_X1 U4222 ( .A(n3260), .ZN(n3231) );
  AOI22_X1 U4223 ( .A1(n4255), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3224) );
  AOI22_X1 U4224 ( .A1(n3248), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3223) );
  AOI22_X1 U4225 ( .A1(n3311), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4226 ( .A1(n3175), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3251), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3221) );
  NAND4_X1 U4227 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3230)
         );
  AOI22_X1 U4228 ( .A1(n3241), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3240), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4229 ( .A1(n3366), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4230 ( .A1(n3250), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3238), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4231 ( .A1(n4121), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3225) );
  NAND4_X1 U4232 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3229)
         );
  NAND2_X1 U4233 ( .A1(n4564), .A2(n3022), .ZN(n3330) );
  NOR2_X1 U4234 ( .A1(n3330), .A2(n3680), .ZN(n3232) );
  AOI21_X1 U4235 ( .B1(n3616), .B2(n3402), .A(n3232), .ZN(n3276) );
  NAND2_X1 U4236 ( .A1(n3263), .A2(n3233), .ZN(n3274) );
  NAND2_X1 U4237 ( .A1(n3274), .A2(n3331), .ZN(n3234) );
  OAI21_X1 U4238 ( .B1(n3269), .B2(n3234), .A(n4421), .ZN(n3235) );
  NAND2_X1 U4239 ( .A1(n3260), .A2(n3790), .ZN(n3258) );
  AOI22_X1 U4240 ( .A1(n3241), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3240), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4241 ( .A1(n4121), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4242 ( .A1(n3311), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4243 ( .A1(n3248), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4244 ( .A1(n3316), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4245 ( .A1(n3251), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3252) );
  NAND2_X1 U4246 ( .A1(n3255), .A2(n3609), .ZN(n3256) );
  NAND2_X1 U4247 ( .A1(n3256), .A2(n3237), .ZN(n3257) );
  NAND2_X1 U4248 ( .A1(n3258), .A2(n3257), .ZN(n3262) );
  NAND2_X1 U4249 ( .A1(n3262), .A2(n3261), .ZN(n3333) );
  AOI21_X2 U4250 ( .B1(n3333), .B2(n3614), .A(n3264), .ZN(n3277) );
  NAND2_X1 U4251 ( .A1(n3272), .A2(n3614), .ZN(n4467) );
  INV_X1 U4252 ( .A(n4467), .ZN(n5170) );
  AOI22_X1 U4253 ( .A1(n5170), .A2(n3330), .B1(n3265), .B2(n3259), .ZN(n3266)
         );
  NAND2_X1 U4254 ( .A1(n3277), .A2(n3266), .ZN(n3738) );
  NAND2_X1 U4255 ( .A1(n3268), .A2(n3267), .ZN(n3283) );
  INV_X1 U4256 ( .A(n3269), .ZN(n3270) );
  NAND2_X1 U4257 ( .A1(n3270), .A2(n3326), .ZN(n3613) );
  NAND2_X1 U4258 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6514) );
  OAI21_X1 U4259 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6514), .ZN(n3606) );
  INV_X1 U4260 ( .A(n3606), .ZN(n3271) );
  OAI211_X1 U4261 ( .C1(n3328), .C2(n3022), .A(n3274), .B(n4467), .ZN(n3275)
         );
  NOR2_X1 U4262 ( .A1(n3613), .A2(n3275), .ZN(n3278) );
  NAND3_X1 U4263 ( .A1(n3278), .A2(n3277), .A3(n3276), .ZN(n3279) );
  MUX2_X1 U4264 ( .A(n4335), .B(n3359), .S(n6632), .Z(n3280) );
  OAI21_X2 U4265 ( .B1(n3355), .B2(n6463), .A(n3281), .ZN(n3282) );
  OAI21_X1 U4266 ( .B1(n3282), .B2(n3283), .A(n3352), .ZN(n3791) );
  AOI22_X1 U4267 ( .A1(n4255), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4268 ( .A1(n4181), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4269 ( .A1(n3299), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4270 ( .A1(n4225), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3284) );
  NAND4_X1 U4271 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3293)
         );
  AOI22_X1 U4272 ( .A1(n4248), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3240), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4273 ( .A1(n4249), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3290) );
  INV_X1 U4274 ( .A(n3238), .ZN(n3294) );
  INV_X2 U4275 ( .A(n3294), .ZN(n4592) );
  AOI22_X1 U4276 ( .A1(n4157), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4277 ( .A1(n4099), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3288) );
  NAND4_X1 U4278 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  INV_X1 U4279 ( .A(n3522), .ZN(n3524) );
  AOI22_X1 U4280 ( .A1(n4181), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4255), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4281 ( .A1(n4249), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4282 ( .A1(n4157), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4283 ( .A1(n4250), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3295) );
  NAND4_X1 U4284 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3305)
         );
  AOI22_X1 U4285 ( .A1(n4248), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4286 ( .A1(n4223), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4287 ( .A1(n4099), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3301) );
  BUF_X1 U4288 ( .A(n3311), .Z(n3299) );
  AOI22_X1 U4289 ( .A1(n3299), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3300) );
  NAND4_X1 U4290 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3304)
         );
  XNOR2_X1 U4291 ( .A(n3524), .B(n3428), .ZN(n3306) );
  NAND2_X1 U4292 ( .A1(n3306), .A2(n4337), .ZN(n3424) );
  INV_X1 U4293 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4397) );
  AOI21_X1 U4294 ( .B1(n4564), .B2(n3522), .A(n6506), .ZN(n3308) );
  NAND2_X1 U4295 ( .A1(n3614), .A2(n3428), .ZN(n3307) );
  OAI211_X1 U4296 ( .C1(n3374), .C2(n4397), .A(n3308), .B(n3307), .ZN(n3423)
         );
  NAND2_X1 U4297 ( .A1(n4337), .A2(n3522), .ZN(n3310) );
  INV_X1 U4298 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4382) );
  NOR2_X1 U4299 ( .A1(n3374), .A2(n4382), .ZN(n3324) );
  AOI22_X1 U4300 ( .A1(n3299), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4301 ( .A1(n4226), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4302 ( .A1(n4223), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4303 ( .A1(n4157), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3312) );
  NAND4_X1 U4304 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3322)
         );
  AOI22_X1 U4305 ( .A1(n4181), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4255), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4306 ( .A1(n4248), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4307 ( .A1(n4225), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4308 ( .A1(n4249), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3317) );
  NAND4_X1 U4309 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  OAI22_X1 U4310 ( .A1(n3385), .A2(n3345), .B1(n3384), .B2(n3522), .ZN(n3323)
         );
  NAND2_X1 U4311 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  INV_X1 U4312 ( .A(n3328), .ZN(n3329) );
  NAND2_X1 U4313 ( .A1(n3017), .A2(n3605), .ZN(n3336) );
  NAND3_X1 U4314 ( .A1(n3636), .A2(n3614), .A3(n3640), .ZN(n3332) );
  NAND2_X1 U4315 ( .A1(n3619), .A2(n3612), .ZN(n3634) );
  INV_X1 U4316 ( .A(n4352), .ZN(n3334) );
  AND2_X1 U4317 ( .A1(n3335), .A2(n3237), .ZN(n4345) );
  NAND3_X1 U4318 ( .A1(n3336), .A2(n3634), .A3(n3732), .ZN(n3337) );
  NAND2_X1 U4319 ( .A1(n3337), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3339) );
  XNOR2_X1 U4320 ( .A(n6632), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6360)
         );
  AND2_X1 U4321 ( .A1(n4335), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3338)
         );
  AOI21_X1 U4322 ( .B1(n3359), .B2(n6360), .A(n3338), .ZN(n3340) );
  INV_X1 U4323 ( .A(n3339), .ZN(n3342) );
  INV_X1 U4324 ( .A(n3340), .ZN(n3341) );
  NAND2_X1 U4325 ( .A1(n3342), .A2(n3104), .ZN(n3343) );
  XNOR2_X2 U4326 ( .A(n3351), .B(n3344), .ZN(n4375) );
  NOR2_X1 U4327 ( .A1(n3345), .A2(n3384), .ZN(n3346) );
  INV_X1 U4328 ( .A(n3347), .ZN(n3348) );
  NOR2_X1 U4329 ( .A1(n3349), .A2(n3348), .ZN(n3350) );
  NAND2_X1 U4330 ( .A1(n3015), .A2(n3016), .ZN(n3354) );
  NAND2_X1 U4331 ( .A1(n3354), .A2(n3353), .ZN(n3377) );
  AND2_X1 U4332 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4333 ( .A1(n3356), .A2(n6474), .ZN(n4840) );
  INV_X1 U4334 ( .A(n3356), .ZN(n3357) );
  NAND2_X1 U4335 ( .A1(n3357), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4336 ( .A1(n4840), .A2(n3358), .ZN(n4384) );
  AOI22_X1 U4337 ( .A1(n3359), .A2(n4384), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4335), .ZN(n3360) );
  XNOR2_X1 U4338 ( .A(n3377), .B(n3378), .ZN(n4373) );
  AOI22_X1 U4339 ( .A1(n4255), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4340 ( .A1(n4181), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4341 ( .A1(n3299), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4342 ( .A1(n4157), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3362) );
  NAND4_X1 U4343 ( .A1(n3365), .A2(n3364), .A3(n3363), .A4(n3362), .ZN(n3372)
         );
  AOI22_X1 U4344 ( .A1(n4248), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3240), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4345 ( .A1(n4249), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4346 ( .A1(n4250), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4347 ( .A1(n4099), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3367) );
  NAND4_X1 U4348 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n3371)
         );
  NOR2_X1 U4349 ( .A1(n3400), .A2(n3384), .ZN(n3373) );
  INV_X1 U4350 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4391) );
  OAI22_X1 U4351 ( .A1(n3374), .A2(n4391), .B1(n3385), .B2(n3400), .ZN(n3375)
         );
  XNOR2_X1 U4352 ( .A(n3376), .B(n3375), .ZN(n3406) );
  NAND2_X1 U4353 ( .A1(n3405), .A2(n3406), .ZN(n3407) );
  INV_X1 U4354 ( .A(n3377), .ZN(n3379) );
  NAND3_X1 U4355 ( .A1(n6359), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4972) );
  INV_X1 U4356 ( .A(n4972), .ZN(n6357) );
  NAND2_X1 U4357 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6357), .ZN(n4978) );
  NAND2_X1 U4358 ( .A1(n6359), .A2(n4978), .ZN(n3380) );
  NOR3_X1 U4359 ( .A1(n6359), .A2(n6474), .A3(n6467), .ZN(n4635) );
  NAND2_X1 U4360 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4635), .ZN(n4580) );
  NAND2_X1 U4361 ( .A1(n3380), .A2(n4580), .ZN(n4909) );
  OAI22_X1 U4362 ( .A1(n4277), .A2(n4909), .B1(n3604), .B2(n6359), .ZN(n3381)
         );
  INV_X1 U4363 ( .A(n3381), .ZN(n3382) );
  AOI22_X1 U4364 ( .A1(n4255), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4365 ( .A1(n4181), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4366 ( .A1(n3299), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4367 ( .A1(n4157), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3386) );
  NAND4_X1 U4368 ( .A1(n3389), .A2(n3388), .A3(n3387), .A4(n3386), .ZN(n3396)
         );
  AOI22_X1 U4369 ( .A1(n4248), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4370 ( .A1(n4249), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4371 ( .A1(n4250), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4372 ( .A1(n4099), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4373 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3395)
         );
  AOI22_X1 U4374 ( .A1(n3597), .A2(n3452), .B1(n3589), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3397) );
  INV_X1 U4375 ( .A(n4370), .ZN(n4614) );
  NAND2_X1 U4376 ( .A1(n3407), .A2(n4614), .ZN(n3399) );
  INV_X1 U4377 ( .A(n3563), .ZN(n3581) );
  NAND2_X1 U4378 ( .A1(n3428), .A2(n3418), .ZN(n3411) );
  NAND2_X1 U4379 ( .A1(n3411), .A2(n3400), .ZN(n3453) );
  INV_X1 U4380 ( .A(n3452), .ZN(n3401) );
  XNOR2_X1 U4381 ( .A(n3453), .B(n3401), .ZN(n3403) );
  NAND2_X1 U4382 ( .A1(n3403), .A2(n4424), .ZN(n3404) );
  INV_X1 U4383 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6295) );
  XNOR2_X1 U4384 ( .A(n3438), .B(n6295), .ZN(n4538) );
  XNOR2_X1 U4385 ( .A(n3411), .B(n3410), .ZN(n3414) );
  INV_X1 U4386 ( .A(n3413), .ZN(n3427) );
  OAI21_X1 U4387 ( .B1(n3414), .B2(n3412), .A(n3427), .ZN(n3415) );
  NAND2_X1 U4388 ( .A1(n4369), .A2(n3563), .ZN(n3422) );
  XNOR2_X1 U4389 ( .A(n3428), .B(n3418), .ZN(n3419) );
  OAI211_X1 U4390 ( .C1(n3419), .C2(n3412), .A(n3326), .B(n3022), .ZN(n3420)
         );
  INV_X1 U4391 ( .A(n3420), .ZN(n3421) );
  NAND2_X1 U4392 ( .A1(n3422), .A2(n3421), .ZN(n4516) );
  INV_X1 U4393 ( .A(n3423), .ZN(n3425) );
  OAI21_X1 U4394 ( .B1(n3412), .B2(n3428), .A(n3427), .ZN(n3429) );
  INV_X1 U4395 ( .A(n3429), .ZN(n3430) );
  NAND2_X1 U4396 ( .A1(n4440), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3431)
         );
  INV_X1 U4397 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U4398 ( .A1(n3431), .A2(n4520), .ZN(n3432) );
  AND2_X1 U4399 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U4400 ( .A1(n4440), .A2(n6299), .ZN(n3433) );
  AND2_X1 U4401 ( .A1(n3432), .A2(n3433), .ZN(n4517) );
  NAND2_X1 U4402 ( .A1(n4516), .A2(n4517), .ZN(n3434) );
  NAND2_X2 U4403 ( .A1(n3434), .A2(n3433), .ZN(n6197) );
  NAND2_X1 U4404 ( .A1(n6197), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3437)
         );
  INV_X1 U4405 ( .A(n6197), .ZN(n3436) );
  NAND2_X1 U4406 ( .A1(n3438), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3439)
         );
  NAND2_X1 U4407 ( .A1(n4539), .A2(n3439), .ZN(n6189) );
  AOI22_X1 U4408 ( .A1(n4255), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4409 ( .A1(n4181), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4410 ( .A1(n3299), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4411 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4157), .B1(n4225), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3440) );
  NAND4_X1 U4412 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n3449)
         );
  AOI22_X1 U4413 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4248), .B1(n3240), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4414 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4218), .B1(n4249), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4415 ( .A1(n4250), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4416 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4099), .B1(n4257), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3444) );
  NAND4_X1 U4417 ( .A1(n3447), .A2(n3446), .A3(n3445), .A4(n3444), .ZN(n3448)
         );
  NAND2_X1 U4418 ( .A1(n3597), .A2(n3503), .ZN(n3451) );
  NAND2_X1 U4419 ( .A1(n3589), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3450) );
  NAND2_X1 U4420 ( .A1(n3451), .A2(n3450), .ZN(n3460) );
  NAND2_X1 U4421 ( .A1(n3821), .A2(n3563), .ZN(n3456) );
  NAND2_X1 U4422 ( .A1(n3453), .A2(n3452), .ZN(n3505) );
  XNOR2_X1 U4423 ( .A(n3505), .B(n3503), .ZN(n3454) );
  NAND2_X1 U4424 ( .A1(n3454), .A2(n4424), .ZN(n3455) );
  NAND2_X1 U4425 ( .A1(n3456), .A2(n3455), .ZN(n3457) );
  INV_X1 U4426 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6287) );
  XNOR2_X1 U4427 ( .A(n3457), .B(n6287), .ZN(n6188) );
  NAND2_X1 U4428 ( .A1(n3457), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3458)
         );
  AOI22_X1 U4429 ( .A1(n4255), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4430 ( .A1(n4181), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3465) );
  INV_X1 U4431 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U4432 ( .A1(n3299), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4433 ( .A1(n4157), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3251), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4434 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3472)
         );
  AOI22_X1 U4435 ( .A1(n4248), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4436 ( .A1(n4249), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4437 ( .A1(n4250), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4438 ( .A1(n4099), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3467) );
  NAND4_X1 U4439 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3471)
         );
  NAND2_X1 U4440 ( .A1(n3597), .A2(n3502), .ZN(n3474) );
  NAND2_X1 U4441 ( .A1(n3589), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U4442 ( .A1(n3474), .A2(n3473), .ZN(n3483) );
  XNOR2_X1 U4443 ( .A(n3485), .B(n3483), .ZN(n3822) );
  NAND2_X1 U4444 ( .A1(n3822), .A2(n3563), .ZN(n3479) );
  INV_X1 U4445 ( .A(n3503), .ZN(n3475) );
  OR2_X1 U4446 ( .A1(n3505), .A2(n3475), .ZN(n3476) );
  XNOR2_X1 U4447 ( .A(n3476), .B(n3502), .ZN(n3477) );
  NAND2_X1 U4448 ( .A1(n3477), .A2(n4424), .ZN(n3478) );
  NAND2_X1 U4449 ( .A1(n3479), .A2(n3478), .ZN(n3481) );
  INV_X1 U4450 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3480) );
  XNOR2_X1 U4451 ( .A(n3481), .B(n3480), .ZN(n4964) );
  NAND2_X1 U4452 ( .A1(n3481), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3482)
         );
  INV_X1 U4453 ( .A(n3483), .ZN(n3484) );
  AOI22_X1 U4454 ( .A1(n4255), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4455 ( .A1(n4181), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4456 ( .A1(n3299), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4457 ( .A1(n4157), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3486) );
  NAND4_X1 U4458 ( .A1(n3489), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(n3495)
         );
  AOI22_X1 U4459 ( .A1(n4248), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4460 ( .A1(n4249), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4461 ( .A1(n4250), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4462 ( .A1(n4099), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3490) );
  NAND4_X1 U4463 ( .A1(n3493), .A2(n3492), .A3(n3491), .A4(n3490), .ZN(n3494)
         );
  NAND2_X1 U4464 ( .A1(n3597), .A2(n3514), .ZN(n3497) );
  NAND2_X1 U4465 ( .A1(n3589), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U4466 ( .A1(n3497), .A2(n3496), .ZN(n3499) );
  INV_X1 U4467 ( .A(n3498), .ZN(n3501) );
  INV_X1 U4468 ( .A(n3499), .ZN(n3500) );
  NAND2_X1 U4469 ( .A1(n3501), .A2(n3500), .ZN(n3834) );
  NAND3_X1 U4470 ( .A1(n3512), .A2(n3563), .A3(n3834), .ZN(n3508) );
  NAND2_X1 U4471 ( .A1(n3503), .A2(n3502), .ZN(n3504) );
  OR2_X1 U4472 ( .A1(n3505), .A2(n3504), .ZN(n3513) );
  XNOR2_X1 U4473 ( .A(n3513), .B(n3514), .ZN(n3506) );
  NAND2_X1 U4474 ( .A1(n3506), .A2(n4424), .ZN(n3507) );
  NAND2_X1 U4475 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  INV_X1 U4476 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6266) );
  XNOR2_X1 U4477 ( .A(n3509), .B(n6266), .ZN(n6180) );
  NAND2_X1 U4478 ( .A1(n3509), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3510)
         );
  AOI22_X1 U4479 ( .A1(n3597), .A2(n3522), .B1(n3589), .B2(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3511) );
  XNOR2_X1 U4480 ( .A(n3512), .B(n3511), .ZN(n3835) );
  OR2_X1 U4481 ( .A1(n3835), .A2(n3581), .ZN(n3518) );
  INV_X1 U4482 ( .A(n3513), .ZN(n3515) );
  NAND2_X1 U4483 ( .A1(n3515), .A2(n3514), .ZN(n3525) );
  XNOR2_X1 U4484 ( .A(n3525), .B(n3522), .ZN(n3516) );
  NAND2_X1 U4485 ( .A1(n3516), .A2(n4424), .ZN(n3517) );
  NAND2_X1 U4486 ( .A1(n3518), .A2(n3517), .ZN(n3520) );
  INV_X1 U4487 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3519) );
  XNOR2_X1 U4488 ( .A(n3520), .B(n3519), .ZN(n5002) );
  NAND2_X1 U4489 ( .A1(n3520), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3521)
         );
  NAND2_X1 U4490 ( .A1(n5001), .A2(n3521), .ZN(n5236) );
  OR3_X1 U4491 ( .A1(n3525), .A2(n3524), .A3(n3412), .ZN(n3526) );
  INV_X1 U4492 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6757) );
  XNOR2_X1 U4493 ( .A(n3527), .B(n6757), .ZN(n5235) );
  NAND2_X1 U4494 ( .A1(n5236), .A2(n5235), .ZN(n5234) );
  NAND2_X1 U4495 ( .A1(n3527), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3528)
         );
  INV_X1 U4496 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6238) );
  OR2_X1 U4497 ( .A1(n5650), .A2(n6238), .ZN(n5250) );
  INV_X1 U4498 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3530) );
  NAND2_X1 U4499 ( .A1(n5650), .A2(n3530), .ZN(n5260) );
  INV_X1 U4500 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3531) );
  AND2_X1 U4501 ( .A1(n5650), .A2(n3531), .ZN(n3534) );
  OR2_X1 U4502 ( .A1(n5650), .A2(n3530), .ZN(n6169) );
  INV_X1 U4503 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5304) );
  NOR2_X1 U4504 ( .A1(n5650), .A2(n5304), .ZN(n5292) );
  XNOR2_X1 U4505 ( .A(n5650), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5353)
         );
  INV_X1 U4506 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U4507 ( .A1(n5650), .A2(n5940), .ZN(n3535) );
  INV_X1 U4508 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5360) );
  AND2_X1 U4509 ( .A1(n5650), .A2(n5360), .ZN(n3537) );
  INV_X1 U4510 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5930) );
  NOR2_X1 U4511 ( .A1(n5650), .A2(n5930), .ZN(n3539) );
  NAND2_X1 U4512 ( .A1(n5650), .A2(n5930), .ZN(n3538) );
  AND2_X1 U4513 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U4514 ( .A1(n5742), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3540) );
  INV_X1 U4515 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5908) );
  INV_X1 U4516 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5755) );
  INV_X1 U4517 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5923) );
  AND3_X1 U4518 ( .A1(n5908), .A2(n5755), .A3(n5923), .ZN(n3541) );
  NOR2_X1 U4519 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5713) );
  NOR2_X1 U4520 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5728) );
  INV_X1 U4521 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U4522 ( .A1(n5643), .A2(n3103), .ZN(n3547) );
  NAND2_X1 U4523 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3763) );
  INV_X1 U4524 ( .A(n3763), .ZN(n3544) );
  NAND2_X1 U4525 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U4526 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3765) );
  INV_X1 U4527 ( .A(n3545), .ZN(n3546) );
  NAND2_X1 U4528 ( .A1(n3547), .A2(n3546), .ZN(n5570) );
  NAND2_X1 U4529 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5591) );
  AND2_X1 U4530 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5673) );
  INV_X1 U4531 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5672) );
  INV_X1 U4532 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5694) );
  INV_X1 U4533 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3550) );
  NAND2_X1 U4534 ( .A1(n5694), .A2(n3550), .ZN(n5685) );
  NOR2_X1 U4535 ( .A1(n5592), .A2(n5685), .ZN(n5564) );
  NAND2_X1 U4536 ( .A1(n5564), .A2(n5672), .ZN(n5393) );
  NOR3_X1 U4537 ( .A1(n3549), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5393), 
        .ZN(n3551) );
  AOI21_X1 U4538 ( .B1(n5396), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n3551), 
        .ZN(n3552) );
  XNOR2_X1 U4539 ( .A(n3552), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3776)
         );
  XNOR2_X1 U4540 ( .A(n6598), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3585)
         );
  XNOR2_X1 U4541 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3562) );
  NAND2_X1 U4542 ( .A1(n3564), .A2(n3562), .ZN(n3554) );
  NAND2_X1 U4543 ( .A1(n6467), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3553) );
  NAND2_X1 U4544 ( .A1(n3554), .A2(n3553), .ZN(n3559) );
  XNOR2_X1 U4545 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3557) );
  NAND2_X1 U4546 ( .A1(n3559), .A2(n3557), .ZN(n3556) );
  NAND2_X1 U4547 ( .A1(n6474), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3555) );
  XOR2_X1 U4548 ( .A(n3585), .B(n3586), .Z(n3625) );
  INV_X1 U4549 ( .A(n3597), .ZN(n3560) );
  INV_X1 U4550 ( .A(n3557), .ZN(n3558) );
  XNOR2_X1 U4551 ( .A(n3559), .B(n3558), .ZN(n3623) );
  INV_X1 U4552 ( .A(n3623), .ZN(n3578) );
  NOR2_X1 U4553 ( .A1(n3560), .A2(n3578), .ZN(n3576) );
  INV_X1 U4554 ( .A(n3576), .ZN(n3583) );
  AOI21_X1 U4555 ( .B1(n3612), .B2(n3022), .A(n5032), .ZN(n3582) );
  XOR2_X1 U4556 ( .A(n3562), .B(n3564), .Z(n3624) );
  INV_X1 U4557 ( .A(n3624), .ZN(n3575) );
  INV_X1 U4558 ( .A(n3601), .ZN(n3574) );
  AOI21_X1 U4559 ( .B1(n3597), .B2(n4421), .A(n3325), .ZN(n3570) );
  NOR3_X1 U4560 ( .A1(n3570), .A2(n3575), .A3(n6506), .ZN(n3573) );
  INV_X1 U4561 ( .A(n3564), .ZN(n3565) );
  OAI21_X1 U4562 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6632), .A(n3565), 
        .ZN(n3568) );
  INV_X1 U4563 ( .A(n3568), .ZN(n3566) );
  NAND2_X1 U4564 ( .A1(n3597), .A2(n3566), .ZN(n3571) );
  OAI21_X1 U4565 ( .B1(n3636), .B2(n3568), .A(n3567), .ZN(n3569) );
  AOI222_X1 U4566 ( .A1(n3571), .A2(n3601), .B1(n3575), .B2(n3570), .C1(n3569), 
        .C2(n3582), .ZN(n3572) );
  AOI211_X1 U4567 ( .C1(n3575), .C2(n3574), .A(n3573), .B(n3572), .ZN(n3580)
         );
  INV_X1 U4568 ( .A(n3582), .ZN(n3577) );
  AOI211_X1 U4569 ( .C1(n3589), .C2(n3578), .A(n3577), .B(n3576), .ZN(n3579)
         );
  OAI222_X1 U4570 ( .A1(n3583), .A2(n3582), .B1(n3581), .B2(n3625), .C1(n3580), 
        .C2(n3579), .ZN(n3584) );
  OAI21_X1 U4571 ( .B1(n3589), .B2(n3625), .A(n3584), .ZN(n3591) );
  NAND2_X1 U4572 ( .A1(n3586), .A2(n3585), .ZN(n3588) );
  NAND2_X1 U4573 ( .A1(n6359), .A2(n6598), .ZN(n3587) );
  NAND2_X1 U4574 ( .A1(n3588), .A2(n3587), .ZN(n3594) );
  NOR2_X1 U4575 ( .A1(n3589), .A2(n3622), .ZN(n3590) );
  OAI22_X1 U4576 ( .A1(n3591), .A2(n3590), .B1(n3601), .B2(n3622), .ZN(n3592)
         );
  AOI21_X1 U4577 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6506), .A(n3592), 
        .ZN(n3599) );
  NAND2_X1 U4578 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4507), .ZN(n3595) );
  NAND2_X1 U4579 ( .A1(n3627), .A2(n3597), .ZN(n3598) );
  NAND2_X1 U4580 ( .A1(n3599), .A2(n3598), .ZN(n3603) );
  INV_X1 U4581 ( .A(n3627), .ZN(n3600) );
  NAND2_X1 U4582 ( .A1(n3612), .A2(n6520), .ZN(n4303) );
  AND2_X1 U4583 ( .A1(n4303), .A2(n6611), .ZN(n4464) );
  NAND2_X1 U4584 ( .A1(n3020), .A2(n4464), .ZN(n3608) );
  INV_X1 U4585 ( .A(n4345), .ZN(n3607) );
  NAND3_X1 U4586 ( .A1(n3608), .A2(n3265), .A3(n3607), .ZN(n3610) );
  NAND2_X1 U4587 ( .A1(n3610), .A2(n3609), .ZN(n3633) );
  NAND2_X1 U4588 ( .A1(n3335), .A2(n3233), .ZN(n3611) );
  NOR2_X1 U4589 ( .A1(n5786), .A2(n3612), .ZN(n3743) );
  NAND2_X1 U4590 ( .A1(n4473), .A2(n3743), .ZN(n3630) );
  AND2_X1 U4591 ( .A1(n5786), .A2(n3614), .ZN(n3615) );
  INV_X1 U4592 ( .A(n3263), .ZN(n3618) );
  AND2_X1 U4593 ( .A1(n3263), .A2(n3265), .ZN(n3617) );
  OAI22_X1 U4594 ( .A1(n3616), .A2(n3618), .B1(n4424), .B2(n3617), .ZN(n3736)
         );
  AND2_X1 U4595 ( .A1(n3637), .A2(n3736), .ZN(n3621) );
  OR2_X1 U4596 ( .A1(n3621), .A2(n3620), .ZN(n4469) );
  NAND2_X1 U4597 ( .A1(n4421), .A2(n6520), .ZN(n3628) );
  AND4_X1 U4598 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3626)
         );
  NOR2_X1 U4599 ( .A1(READY_N), .A2(n4406), .ZN(n4340) );
  NAND3_X1 U4600 ( .A1(n3628), .A2(n4340), .A3(n3259), .ZN(n3629) );
  NAND3_X1 U4601 ( .A1(n3630), .A2(n4469), .A3(n3629), .ZN(n3631) );
  NAND2_X1 U4602 ( .A1(n3631), .A2(n6503), .ZN(n3632) );
  INV_X1 U4603 ( .A(n3732), .ZN(n3635) );
  AOI22_X1 U4604 ( .A1(n3635), .A2(n3233), .B1(n3020), .B2(n4438), .ZN(n3638)
         );
  INV_X1 U4605 ( .A(n4408), .ZN(n6481) );
  NAND2_X1 U4606 ( .A1(n3637), .A2(n5032), .ZN(n4407) );
  NAND4_X1 U4607 ( .A1(n3634), .A2(n3638), .A3(n6481), .A4(n4407), .ZN(n3639)
         );
  NAND2_X1 U4608 ( .A1(n3776), .A2(n6307), .ZN(n3774) );
  INV_X1 U4609 ( .A(n3026), .ZN(n3651) );
  AOI22_X1 U4610 ( .A1(n4428), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3027), .ZN(n3730) );
  INV_X1 U4611 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U4612 ( .A1(n3641), .A2(n3034), .ZN(n3645) );
  NAND2_X1 U4613 ( .A1(n3716), .A2(EBX_REG_0__SCAN_IN), .ZN(n3644) );
  INV_X1 U4614 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U4615 ( .A1(n3026), .A2(n3642), .ZN(n3643) );
  NAND2_X1 U4616 ( .A1(n3644), .A2(n3643), .ZN(n4429) );
  XNOR2_X1 U4617 ( .A(n3645), .B(n4429), .ZN(n4439) );
  NAND2_X1 U4618 ( .A1(n4439), .A2(n4438), .ZN(n4437) );
  NAND2_X1 U4619 ( .A1(n4437), .A2(n3645), .ZN(n4530) );
  INV_X1 U4620 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6805) );
  MUX2_X1 U4621 ( .A(n3044), .B(n3725), .S(n6805), .Z(n3647) );
  OAI21_X1 U4622 ( .B1(n4438), .B2(n3435), .A(n3708), .ZN(n3646) );
  NOR2_X1 U4623 ( .A1(n3647), .A2(n3646), .ZN(n4531) );
  OR2_X1 U4624 ( .A1(n3720), .A2(EBX_REG_3__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4625 ( .A1(n3026), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3648)
         );
  OAI211_X1 U4626 ( .C1(n3027), .C2(EBX_REG_3__SCAN_IN), .A(n3716), .B(n3648), 
        .ZN(n3649) );
  AND2_X1 U4627 ( .A1(n3650), .A2(n3649), .ZN(n4513) );
  INV_X1 U4628 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U4629 ( .A1(n3725), .A2(n6787), .ZN(n3654) );
  NAND2_X1 U4630 ( .A1(n3716), .A2(n6287), .ZN(n3652) );
  OAI211_X1 U4631 ( .C1(n3027), .C2(EBX_REG_4__SCAN_IN), .A(n3652), .B(n3026), 
        .ZN(n3653) );
  INV_X1 U4632 ( .A(EBX_REG_5__SCAN_IN), .ZN(n3655) );
  MUX2_X1 U4633 ( .A(n3026), .B(n3720), .S(n3655), .Z(n3657) );
  OR2_X1 U4634 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3656)
         );
  NAND2_X1 U4635 ( .A1(n3657), .A2(n3656), .ZN(n4755) );
  MUX2_X1 U4636 ( .A(n3720), .B(n3026), .S(EBX_REG_7__SCAN_IN), .Z(n3658) );
  OAI21_X1 U4637 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4428), .A(n3658), 
        .ZN(n4951) );
  INV_X1 U4638 ( .A(EBX_REG_6__SCAN_IN), .ZN(n3659) );
  NAND2_X1 U4639 ( .A1(n3725), .A2(n3659), .ZN(n3662) );
  NAND2_X1 U4640 ( .A1(n3716), .A2(n6266), .ZN(n3660) );
  OAI211_X1 U4641 ( .C1(n3027), .C2(EBX_REG_6__SCAN_IN), .A(n3660), .B(n3026), 
        .ZN(n3661) );
  NOR2_X1 U4642 ( .A1(n4951), .A2(n4950), .ZN(n3663) );
  AND2_X2 U4643 ( .A1(n4753), .A2(n3663), .ZN(n5108) );
  OR2_X1 U4644 ( .A1(n3720), .A2(EBX_REG_9__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4645 ( .A1(n3026), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3664)
         );
  OAI211_X1 U4646 ( .C1(n3027), .C2(EBX_REG_9__SCAN_IN), .A(n3716), .B(n3664), 
        .ZN(n3665) );
  AND2_X1 U4647 ( .A1(n3666), .A2(n3665), .ZN(n5106) );
  NAND2_X1 U4648 ( .A1(n3716), .A2(n6757), .ZN(n3668) );
  INV_X1 U4649 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U4650 ( .A1(n4438), .A2(n6042), .ZN(n3667) );
  NAND3_X1 U4651 ( .A1(n3668), .A2(n3667), .A3(n3026), .ZN(n3669) );
  OAI21_X1 U4652 ( .B1(EBX_REG_8__SCAN_IN), .B2(n3717), .A(n3669), .ZN(n5107)
         );
  AND2_X1 U4653 ( .A1(n5106), .A2(n5107), .ZN(n3670) );
  NAND2_X1 U4654 ( .A1(n5108), .A2(n3670), .ZN(n5105) );
  INV_X1 U4655 ( .A(n5105), .ZN(n3675) );
  INV_X1 U4656 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6667) );
  MUX2_X1 U4657 ( .A(n3044), .B(n3725), .S(n6667), .Z(n3673) );
  NAND2_X1 U4658 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n3027), .ZN(n3671) );
  NAND2_X1 U4659 ( .A1(n3708), .A2(n3671), .ZN(n3672) );
  NOR2_X1 U4660 ( .A1(n3673), .A2(n3672), .ZN(n5245) );
  INV_X1 U4661 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5271) );
  MUX2_X1 U4662 ( .A(n3026), .B(n3720), .S(n5271), .Z(n3676) );
  OAI21_X1 U4663 ( .B1(n4428), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n3676), 
        .ZN(n5268) );
  NAND2_X1 U4664 ( .A1(n3716), .A2(n5304), .ZN(n3678) );
  INV_X1 U4665 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U4666 ( .A1(n4438), .A2(n5278), .ZN(n3677) );
  NAND3_X1 U4667 ( .A1(n3678), .A2(n3677), .A3(n3026), .ZN(n3679) );
  OAI21_X1 U4668 ( .B1(EBX_REG_12__SCAN_IN), .B2(n3717), .A(n3679), .ZN(n5275)
         );
  OR2_X1 U4669 ( .A1(n3720), .A2(EBX_REG_13__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U4670 ( .A1(n3026), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3681) );
  OAI211_X1 U4671 ( .C1(n3027), .C2(EBX_REG_13__SCAN_IN), .A(n3716), .B(n3681), 
        .ZN(n3682) );
  INV_X1 U4672 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U4673 ( .A1(n3725), .A2(n5348), .ZN(n3686) );
  NAND2_X1 U4674 ( .A1(n3716), .A2(n5360), .ZN(n3684) );
  OAI211_X1 U4675 ( .C1(n3027), .C2(EBX_REG_14__SCAN_IN), .A(n3684), .B(n3026), 
        .ZN(n3685) );
  MUX2_X1 U4676 ( .A(n3720), .B(n3026), .S(EBX_REG_15__SCAN_IN), .Z(n3688) );
  OR2_X1 U4677 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3687)
         );
  NAND2_X1 U4678 ( .A1(n3688), .A2(n3687), .ZN(n5532) );
  OR2_X1 U4679 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3690)
         );
  INV_X1 U4680 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5531) );
  MUX2_X1 U4681 ( .A(n3026), .B(n3720), .S(n5531), .Z(n3689) );
  AND2_X1 U4682 ( .A1(n3690), .A2(n3689), .ZN(n5526) );
  NAND2_X1 U4683 ( .A1(n3716), .A2(n5923), .ZN(n3692) );
  INV_X1 U4684 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U4685 ( .A1(n4438), .A2(n5389), .ZN(n3691) );
  NAND3_X1 U4686 ( .A1(n3692), .A2(n3691), .A3(n3026), .ZN(n3693) );
  OAI21_X1 U4687 ( .B1(EBX_REG_16__SCAN_IN), .B2(n3717), .A(n3693), .ZN(n5527)
         );
  NAND2_X1 U4688 ( .A1(n5526), .A2(n5527), .ZN(n3694) );
  INV_X1 U4689 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U4690 ( .A1(n3716), .A2(n5763), .ZN(n3697) );
  INV_X1 U4691 ( .A(EBX_REG_19__SCAN_IN), .ZN(n3695) );
  NAND2_X1 U4692 ( .A1(n4438), .A2(n3695), .ZN(n3696) );
  NAND3_X1 U4693 ( .A1(n3697), .A2(n3696), .A3(n3026), .ZN(n3698) );
  OAI21_X1 U4694 ( .B1(EBX_REG_19__SCAN_IN), .B2(n3717), .A(n3698), .ZN(n5514)
         );
  OR2_X1 U4695 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3700)
         );
  INV_X1 U4696 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U4697 ( .A1(n4438), .A2(n5521), .ZN(n3699) );
  OAI22_X1 U4698 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n3027), .ZN(n5505) );
  NAND2_X1 U4699 ( .A1(n5512), .A2(n5505), .ZN(n3702) );
  NAND2_X1 U4700 ( .A1(n3651), .A2(EBX_REG_20__SCAN_IN), .ZN(n3701) );
  OAI211_X1 U4701 ( .C1(n5512), .C2(n3651), .A(n3702), .B(n3701), .ZN(n3703)
         );
  OR2_X1 U4702 ( .A1(n3720), .A2(EBX_REG_21__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U4703 ( .A1(n3026), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3704) );
  OAI211_X1 U4704 ( .C1(n3027), .C2(EBX_REG_21__SCAN_IN), .A(n3716), .B(n3704), 
        .ZN(n3705) );
  NAND2_X1 U4705 ( .A1(n3706), .A2(n3705), .ZN(n5495) );
  MUX2_X1 U4706 ( .A(n3717), .B(n3716), .S(EBX_REG_22__SCAN_IN), .Z(n3710) );
  NAND2_X1 U4707 ( .A1(n3027), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3707) );
  AND2_X1 U4708 ( .A1(n3708), .A2(n3707), .ZN(n3709) );
  NAND2_X1 U4709 ( .A1(n3710), .A2(n3709), .ZN(n5488) );
  NAND2_X1 U4710 ( .A1(n5489), .A2(n5488), .ZN(n5482) );
  MUX2_X1 U4711 ( .A(n3720), .B(n3026), .S(EBX_REG_23__SCAN_IN), .Z(n3712) );
  OR2_X1 U4712 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3711)
         );
  NAND2_X1 U4713 ( .A1(n3712), .A2(n3711), .ZN(n5483) );
  OR2_X2 U4714 ( .A1(n5482), .A2(n5483), .ZN(n5485) );
  MUX2_X1 U4715 ( .A(n3725), .B(n3044), .S(EBX_REG_24__SCAN_IN), .Z(n3713) );
  NOR2_X1 U4716 ( .A1(n3713), .A2(n3108), .ZN(n5475) );
  MUX2_X1 U4717 ( .A(n3720), .B(n3026), .S(EBX_REG_25__SCAN_IN), .Z(n3715) );
  OR2_X1 U4718 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3714)
         );
  AND2_X1 U4719 ( .A1(n3715), .A2(n3714), .ZN(n5470) );
  AND2_X2 U4720 ( .A1(n5476), .A2(n5470), .ZN(n5472) );
  MUX2_X1 U4721 ( .A(n3717), .B(n3716), .S(EBX_REG_26__SCAN_IN), .Z(n3719) );
  NAND2_X1 U4722 ( .A1(n3027), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3718) );
  NAND2_X1 U4723 ( .A1(n3719), .A2(n3718), .ZN(n5462) );
  MUX2_X1 U4724 ( .A(n3720), .B(n3026), .S(EBX_REG_27__SCAN_IN), .Z(n3722) );
  OR2_X1 U4725 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3721)
         );
  NAND2_X1 U4726 ( .A1(n3722), .A2(n3721), .ZN(n5438) );
  MUX2_X1 U4727 ( .A(n3725), .B(n3044), .S(EBX_REG_28__SCAN_IN), .Z(n3724) );
  AND2_X1 U4728 ( .A1(n3027), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3723)
         );
  NOR2_X1 U4729 ( .A1(n3724), .A2(n3723), .ZN(n4299) );
  OAI22_X1 U4730 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n3027), .ZN(n5454) );
  INV_X1 U4731 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U4732 ( .A1(n3725), .A2(n5457), .ZN(n5452) );
  NOR2_X1 U4733 ( .A1(n5453), .A2(n5452), .ZN(n3726) );
  AOI21_X1 U4734 ( .B1(n4360), .B2(n3026), .A(n3726), .ZN(n5456) );
  NAND2_X1 U4735 ( .A1(n4428), .A2(EBX_REG_30__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4736 ( .A1(n3027), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3727) );
  NAND2_X1 U4737 ( .A1(n3728), .A2(n3727), .ZN(n4361) );
  OAI21_X1 U4738 ( .B1(n5456), .B2(n4361), .A(n4363), .ZN(n3729) );
  XNOR2_X1 U4739 ( .A(n3730), .B(n3729), .ZN(n3731) );
  INV_X1 U4740 ( .A(n3731), .ZN(n5447) );
  NAND2_X1 U4741 ( .A1(n3020), .A2(n4424), .ZN(n6493) );
  OAI21_X1 U4742 ( .B1(n3732), .B2(n3233), .A(n6493), .ZN(n3733) );
  NAND2_X1 U4743 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U4744 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6229) );
  NOR2_X1 U4745 ( .A1(n6240), .A2(n6229), .ZN(n3747) );
  NAND2_X1 U4746 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3745) );
  INV_X1 U4747 ( .A(n3326), .ZN(n3734) );
  AOI22_X1 U4748 ( .A1(n3269), .A2(n3651), .B1(n3734), .B2(n4428), .ZN(n3735)
         );
  NAND2_X1 U4749 ( .A1(n3736), .A2(n3735), .ZN(n3737) );
  NOR2_X1 U4750 ( .A1(n3738), .A2(n3737), .ZN(n4452) );
  INV_X1 U4751 ( .A(n5786), .ZN(n3740) );
  NOR2_X1 U4752 ( .A1(n3331), .A2(n3259), .ZN(n3739) );
  NAND2_X1 U4753 ( .A1(n3740), .A2(n3739), .ZN(n4594) );
  OAI21_X1 U4754 ( .B1(n4343), .B2(n3237), .A(n4594), .ZN(n3741) );
  INV_X1 U4755 ( .A(n3741), .ZN(n3742) );
  NAND2_X1 U4756 ( .A1(n4452), .A2(n3742), .ZN(n3746) );
  INV_X1 U4757 ( .A(n3743), .ZN(n3744) );
  NAND2_X1 U4758 ( .A1(n3753), .A2(n4466), .ZN(n6301) );
  AOI21_X1 U4759 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6298) );
  NAND2_X1 U4760 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6284) );
  NOR2_X1 U4761 ( .A1(n6298), .A2(n6284), .ZN(n6228) );
  NAND2_X1 U4762 ( .A1(n6279), .A2(n6228), .ZN(n6267) );
  NOR2_X1 U4763 ( .A1(n3745), .A2(n6267), .ZN(n6222) );
  NAND2_X1 U4764 ( .A1(n3747), .A2(n6222), .ZN(n5301) );
  NAND2_X1 U4765 ( .A1(n3753), .A2(n3746), .ZN(n3751) );
  NOR2_X1 U4766 ( .A1(n3435), .A2(n4520), .ZN(n6227) );
  INV_X1 U4767 ( .A(n6227), .ZN(n6256) );
  NOR2_X1 U4768 ( .A1(n6256), .A2(n6284), .ZN(n6269) );
  AND3_X1 U4769 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6269), .ZN(n6219) );
  NAND2_X1 U4770 ( .A1(n6219), .A2(n3747), .ZN(n5302) );
  INV_X1 U4771 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4447) );
  NOR3_X1 U4772 ( .A1(n3751), .A2(n5302), .A3(n4447), .ZN(n5300) );
  INV_X1 U4773 ( .A(n5300), .ZN(n3748) );
  NAND2_X1 U4774 ( .A1(n5301), .A2(n3748), .ZN(n5364) );
  AND2_X1 U4775 ( .A1(n3620), .A2(n4421), .ZN(n5412) );
  NAND2_X1 U4776 ( .A1(n3753), .A2(n5412), .ZN(n5363) );
  NOR2_X1 U4777 ( .A1(n3531), .A2(n5304), .ZN(n5933) );
  NAND2_X1 U4778 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5933), .ZN(n5367) );
  NOR2_X1 U4779 ( .A1(n5360), .A2(n5367), .ZN(n5917) );
  NAND3_X1 U4780 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5917), .ZN(n3758) );
  NAND2_X1 U4781 ( .A1(n3543), .A2(n5742), .ZN(n3750) );
  NAND2_X1 U4782 ( .A1(n5739), .A2(n3544), .ZN(n5721) );
  NAND2_X1 U4783 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5679) );
  NAND3_X1 U4784 ( .A1(n5695), .A2(n5673), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5398) );
  INV_X1 U4785 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U4786 ( .A1(n6664), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4787 ( .A1(n6282), .A2(REIP_REG_31__SCAN_IN), .ZN(n4284) );
  NOR2_X1 U4788 ( .A1(n3758), .A2(n5301), .ZN(n5749) );
  INV_X1 U4789 ( .A(n3750), .ZN(n3749) );
  NAND2_X1 U4790 ( .A1(n5749), .A2(n3749), .ZN(n3757) );
  NAND2_X1 U4791 ( .A1(n6257), .A2(n3750), .ZN(n3755) );
  AND2_X1 U4792 ( .A1(n6301), .A2(n3751), .ZN(n5365) );
  INV_X1 U4793 ( .A(n5365), .ZN(n3752) );
  NAND2_X1 U4794 ( .A1(n3752), .A2(n4447), .ZN(n4442) );
  INV_X1 U4795 ( .A(n3753), .ZN(n3754) );
  NAND2_X1 U4796 ( .A1(n3754), .A2(n6302), .ZN(n4441) );
  NAND2_X1 U4797 ( .A1(n4442), .A2(n4441), .ZN(n6258) );
  INV_X1 U4798 ( .A(n6258), .ZN(n4519) );
  AND2_X1 U4799 ( .A1(n6301), .A2(n4519), .ZN(n6221) );
  NAND2_X1 U4800 ( .A1(n3755), .A2(n6221), .ZN(n3756) );
  NAND2_X1 U4801 ( .A1(n3757), .A2(n3756), .ZN(n3762) );
  INV_X1 U4802 ( .A(n3758), .ZN(n3760) );
  INV_X1 U4803 ( .A(n5302), .ZN(n3759) );
  NAND2_X1 U4804 ( .A1(n3760), .A2(n3759), .ZN(n3761) );
  NAND2_X1 U4805 ( .A1(n6257), .A2(n3761), .ZN(n5752) );
  NAND2_X1 U4806 ( .A1(n3762), .A2(n5752), .ZN(n5734) );
  AND2_X1 U4807 ( .A1(n6260), .A2(n3763), .ZN(n3764) );
  NAND2_X1 U4808 ( .A1(n5363), .A2(n4447), .ZN(n4518) );
  OAI21_X1 U4809 ( .B1(n6297), .B2(n6279), .A(n3765), .ZN(n3766) );
  INV_X1 U4810 ( .A(n3766), .ZN(n3767) );
  OAI21_X1 U4811 ( .B1(n5679), .B2(n3083), .A(n6260), .ZN(n3768) );
  NAND2_X1 U4812 ( .A1(n5712), .A2(n3768), .ZN(n5671) );
  INV_X1 U4813 ( .A(n6260), .ZN(n5913) );
  AOI21_X1 U4814 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5913), .ZN(n3769) );
  OAI21_X1 U4815 ( .B1(n5671), .B2(n3769), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n3770) );
  OAI211_X1 U4816 ( .C1(n5398), .C2(n3771), .A(n4284), .B(n3770), .ZN(n3772)
         );
  AOI21_X1 U4817 ( .B1(n5447), .B2(n6290), .A(n3772), .ZN(n3773) );
  NAND2_X1 U4818 ( .A1(n3774), .A2(n3773), .ZN(U2987) );
  NAND2_X1 U4819 ( .A1(n3776), .A2(n6206), .ZN(n4288) );
  INV_X1 U4820 ( .A(n3777), .ZN(n3784) );
  NAND2_X1 U4821 ( .A1(n4345), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3817) );
  NAND2_X1 U4822 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3798) );
  INV_X1 U4823 ( .A(n3798), .ZN(n3780) );
  INV_X1 U4824 ( .A(n3810), .ZN(n3811) );
  OAI21_X1 U4825 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3780), .A(n3811), 
        .ZN(n5169) );
  AOI22_X1 U4826 ( .A1(n4242), .A2(n5169), .B1(n4272), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U4827 ( .A1(n4273), .A2(EAX_REG_3__SCAN_IN), .ZN(n3781) );
  OAI211_X1 U4828 ( .C1(n3817), .C2(n3087), .A(n3782), .B(n3781), .ZN(n3783)
         );
  AOI21_X1 U4829 ( .B1(n3784), .B2(n3778), .A(n3783), .ZN(n4511) );
  INV_X1 U4830 ( .A(n4511), .ZN(n3809) );
  NAND2_X1 U4831 ( .A1(n4369), .A2(n3778), .ZN(n3789) );
  NAND2_X1 U4832 ( .A1(n4378), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3786)
         );
  NAND2_X1 U4833 ( .A1(n3794), .A2(EAX_REG_1__SCAN_IN), .ZN(n3785) );
  OAI211_X1 U4834 ( .C1(n3817), .C2(n4454), .A(n3786), .B(n3785), .ZN(n3787)
         );
  INV_X1 U4835 ( .A(n3787), .ZN(n3788) );
  NAND2_X1 U4836 ( .A1(n3789), .A2(n3788), .ZN(n4433) );
  AOI21_X1 U4837 ( .B1(n4873), .B2(n3790), .A(n4378), .ZN(n4432) );
  INV_X1 U4838 ( .A(n3792), .ZN(n4841) );
  INV_X1 U4839 ( .A(n3778), .ZN(n3793) );
  OR2_X1 U4840 ( .A1(n3792), .A2(n3793), .ZN(n3796) );
  AOI22_X1 U4841 ( .A1(n3794), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4378), .ZN(n3795) );
  OAI211_X1 U4842 ( .C1(n3817), .C2(n6463), .A(n3796), .B(n3795), .ZN(n4431)
         );
  MUX2_X1 U4843 ( .A(n4242), .B(n4432), .S(n4431), .Z(n4434) );
  NAND2_X1 U4844 ( .A1(n3805), .A2(n4436), .ZN(n3804) );
  INV_X1 U4845 ( .A(n3817), .ZN(n3797) );
  NAND2_X1 U4846 ( .A1(n3797), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3803) );
  OAI21_X1 U4847 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3798), .ZN(n6201) );
  NAND2_X1 U4848 ( .A1(n4242), .A2(n6201), .ZN(n3800) );
  NAND2_X1 U4849 ( .A1(n4272), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3799)
         );
  NAND2_X1 U4850 ( .A1(n3800), .A2(n3799), .ZN(n3801) );
  AOI21_X1 U4851 ( .B1(n4273), .B2(EAX_REG_2__SCAN_IN), .A(n3801), .ZN(n3802)
         );
  AND2_X1 U4852 ( .A1(n3803), .A2(n3802), .ZN(n4533) );
  NAND2_X1 U4853 ( .A1(n3804), .A2(n4533), .ZN(n3807) );
  INV_X1 U4854 ( .A(n3805), .ZN(n4535) );
  INV_X1 U4855 ( .A(n4436), .ZN(n4534) );
  NAND2_X1 U4856 ( .A1(n4535), .A2(n4534), .ZN(n3806) );
  NAND2_X1 U4857 ( .A1(n3807), .A2(n3806), .ZN(n4510) );
  INV_X1 U4858 ( .A(n4510), .ZN(n3808) );
  NAND2_X1 U4859 ( .A1(n3809), .A2(n3808), .ZN(n4509) );
  INV_X1 U4860 ( .A(n3826), .ZN(n3814) );
  INV_X1 U4861 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3812) );
  NAND2_X1 U4862 ( .A1(n3812), .A2(n3811), .ZN(n3813) );
  NAND2_X1 U4863 ( .A1(n3814), .A2(n3813), .ZN(n6194) );
  NAND2_X1 U4864 ( .A1(n4378), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3816)
         );
  NAND2_X1 U4865 ( .A1(n4273), .A2(EAX_REG_4__SCAN_IN), .ZN(n3815) );
  OAI211_X1 U4866 ( .C1(n3817), .C2(n4507), .A(n3816), .B(n3815), .ZN(n3819)
         );
  MUX2_X1 U4867 ( .A(n6194), .B(n3819), .S(n3818), .Z(n3820) );
  AOI21_X1 U4868 ( .B1(n3821), .B2(n3778), .A(n3820), .ZN(n4625) );
  NAND2_X1 U4869 ( .A1(n3822), .A2(n3778), .ZN(n3825) );
  INV_X1 U4870 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5035) );
  XNOR2_X1 U4871 ( .A(n3826), .B(n5035), .ZN(n5037) );
  OAI22_X1 U4872 ( .A1(n5037), .A2(n3818), .B1(n4131), .B2(n5035), .ZN(n3823)
         );
  AOI21_X1 U4873 ( .B1(n4273), .B2(EAX_REG_5__SCAN_IN), .A(n3823), .ZN(n3824)
         );
  NAND2_X1 U4874 ( .A1(n3825), .A2(n3824), .ZN(n4711) );
  NAND2_X1 U4875 ( .A1(n4624), .A2(n4711), .ZN(n4710) );
  INV_X1 U4876 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3832) );
  AND2_X1 U4877 ( .A1(n3827), .A2(n3829), .ZN(n3828) );
  OR2_X1 U4878 ( .A1(n3828), .A2(n3852), .ZN(n6187) );
  NOR2_X1 U4879 ( .A1(n4131), .A2(n3829), .ZN(n3830) );
  AOI21_X1 U4880 ( .B1(n6187), .B2(n4242), .A(n3830), .ZN(n3831) );
  OAI21_X1 U4881 ( .B1(n3839), .B2(n3832), .A(n3831), .ZN(n3833) );
  AOI21_X1 U4882 ( .B1(n3834), .B2(n3778), .A(n3833), .ZN(n4862) );
  INV_X1 U4883 ( .A(n3835), .ZN(n3841) );
  INV_X1 U4884 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3838) );
  XNOR2_X1 U4885 ( .A(n3852), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5005) );
  INV_X1 U4886 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4956) );
  NOR2_X1 U4887 ( .A1(n4131), .A2(n4956), .ZN(n3836) );
  AOI21_X1 U4888 ( .B1(n5005), .B2(n4242), .A(n3836), .ZN(n3837) );
  OAI21_X1 U4889 ( .B1(n3839), .B2(n3838), .A(n3837), .ZN(n3840) );
  AOI21_X1 U4890 ( .B1(n3841), .B2(n3778), .A(n3840), .ZN(n4948) );
  AOI22_X1 U4891 ( .A1(n4218), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4892 ( .A1(n4157), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4893 ( .A1(n4225), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4894 ( .A1(n4226), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4895 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3851)
         );
  AOI22_X1 U4896 ( .A1(n4181), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4897 ( .A1(n4248), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4898 ( .A1(n4255), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4899 ( .A1(n4249), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4900 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3850)
         );
  OAI21_X1 U4901 ( .B1(n3851), .B2(n3850), .A(n3778), .ZN(n3856) );
  NAND2_X1 U4902 ( .A1(n4273), .A2(EAX_REG_8__SCAN_IN), .ZN(n3855) );
  XNOR2_X1 U4903 ( .A(n3857), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U4904 ( .A1(n6045), .A2(n4242), .ZN(n3854) );
  NAND2_X1 U4905 ( .A1(n4272), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3853)
         );
  NAND4_X1 U4906 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n5029)
         );
  INV_X1 U4907 ( .A(n5027), .ZN(n3873) );
  XOR2_X1 U4908 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3874), .Z(n6030) );
  INV_X1 U4909 ( .A(n6030), .ZN(n5252) );
  AOI22_X1 U4910 ( .A1(n4255), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4911 ( .A1(n4099), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4912 ( .A1(n3299), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4913 ( .A1(n4218), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4914 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3867)
         );
  AOI22_X1 U4915 ( .A1(n4157), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4916 ( .A1(n4248), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4917 ( .A1(n4181), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4918 ( .A1(n4226), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4919 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3866)
         );
  OAI21_X1 U4920 ( .B1(n3867), .B2(n3866), .A(n3778), .ZN(n3870) );
  NAND2_X1 U4921 ( .A1(n4273), .A2(EAX_REG_9__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4922 ( .A1(n4272), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3868)
         );
  NAND3_X1 U4923 ( .A1(n3870), .A2(n3869), .A3(n3868), .ZN(n3871) );
  AOI21_X1 U4924 ( .B1(n5252), .B2(n4242), .A(n3871), .ZN(n5102) );
  NAND2_X1 U4925 ( .A1(n3873), .A2(n3872), .ZN(n5101) );
  INV_X1 U4926 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3875) );
  XNOR2_X1 U4927 ( .A(n3889), .B(n3875), .ZN(n6028) );
  AOI22_X1 U4928 ( .A1(n4273), .A2(EAX_REG_10__SCAN_IN), .B1(n4272), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4929 ( .A1(n4248), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4930 ( .A1(n3311), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4931 ( .A1(n4157), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4932 ( .A1(n4218), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4933 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3885)
         );
  AOI22_X1 U4934 ( .A1(n3025), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4935 ( .A1(n4249), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4936 ( .A1(n4181), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4937 ( .A1(n4225), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4938 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884)
         );
  OAI21_X1 U4939 ( .B1(n3885), .B2(n3884), .A(n3778), .ZN(n3886) );
  OAI211_X1 U4940 ( .C1(n6028), .C2(n3818), .A(n3887), .B(n3886), .ZN(n3888)
         );
  INV_X1 U4941 ( .A(n3888), .ZN(n5243) );
  NOR2_X2 U4942 ( .A1(n5101), .A2(n5243), .ZN(n5241) );
  XOR2_X1 U4943 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3903), .Z(n6174) );
  AOI22_X1 U4944 ( .A1(n4157), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4945 ( .A1(n4248), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4946 ( .A1(n4181), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4947 ( .A1(n4225), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4948 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3899)
         );
  AOI22_X1 U4949 ( .A1(n4226), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4950 ( .A1(n4255), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4951 ( .A1(n4099), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4952 ( .A1(n3311), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4953 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3898)
         );
  OR2_X1 U4954 ( .A1(n3899), .A2(n3898), .ZN(n3900) );
  AOI22_X1 U4955 ( .A1(n3778), .A2(n3900), .B1(n4272), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3902) );
  NAND2_X1 U4956 ( .A1(n4273), .A2(EAX_REG_11__SCAN_IN), .ZN(n3901) );
  OAI211_X1 U4957 ( .C1(n6174), .C2(n3818), .A(n3902), .B(n3901), .ZN(n5257)
         );
  XNOR2_X1 U4958 ( .A(n3919), .B(n3918), .ZN(n5296) );
  AOI21_X1 U4959 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3918), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3905) );
  AND2_X1 U4960 ( .A1(n4273), .A2(EAX_REG_12__SCAN_IN), .ZN(n3904) );
  OAI22_X1 U4961 ( .A1(n5296), .A2(n3818), .B1(n3905), .B2(n3904), .ZN(n3917)
         );
  AOI22_X1 U4962 ( .A1(n4181), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4963 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4248), .B1(n4218), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4964 ( .A1(n3025), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4965 ( .A1(n4226), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4966 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3915)
         );
  AOI22_X1 U4967 ( .A1(n4223), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4968 ( .A1(n4224), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4969 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4099), .B1(n4257), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4970 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4249), .B1(n4250), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4971 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3914)
         );
  OAI21_X1 U4972 ( .B1(n3915), .B2(n3914), .A(n3778), .ZN(n3916) );
  NAND2_X1 U4973 ( .A1(n3917), .A2(n3916), .ZN(n5273) );
  XOR2_X1 U4974 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3935), .Z(n5324) );
  INV_X1 U4975 ( .A(n5324), .ZN(n5355) );
  AOI22_X1 U4976 ( .A1(n4157), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4977 ( .A1(n4255), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4978 ( .A1(n4249), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4979 ( .A1(n4225), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4980 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3929)
         );
  AOI22_X1 U4981 ( .A1(n4248), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4982 ( .A1(n4218), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4983 ( .A1(n3299), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4984 ( .A1(n4181), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3924) );
  NAND4_X1 U4985 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3928)
         );
  OAI21_X1 U4986 ( .B1(n3929), .B2(n3928), .A(n3778), .ZN(n3932) );
  NAND2_X1 U4987 ( .A1(n4273), .A2(EAX_REG_13__SCAN_IN), .ZN(n3931) );
  NAND2_X1 U4988 ( .A1(n4272), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3930)
         );
  NAND3_X1 U4989 ( .A1(n3932), .A2(n3931), .A3(n3930), .ZN(n3933) );
  AOI21_X1 U4990 ( .B1(n5355), .B2(n4242), .A(n3933), .ZN(n5314) );
  XNOR2_X1 U4991 ( .A(n3952), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5376)
         );
  AOI22_X1 U4992 ( .A1(n4181), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4993 ( .A1(n4248), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4994 ( .A1(n4218), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4995 ( .A1(n4223), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4996 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3945)
         );
  AOI22_X1 U4997 ( .A1(n4255), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4998 ( .A1(n3251), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4999 ( .A1(n4249), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U5000 ( .A1(n4226), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U5001 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3944)
         );
  OAI21_X1 U5002 ( .B1(n3945), .B2(n3944), .A(n3778), .ZN(n3948) );
  NAND2_X1 U5003 ( .A1(n4273), .A2(EAX_REG_14__SCAN_IN), .ZN(n3947) );
  NAND2_X1 U5004 ( .A1(n4272), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3946)
         );
  NAND3_X1 U5005 ( .A1(n3948), .A2(n3947), .A3(n3946), .ZN(n3949) );
  AOI21_X1 U5006 ( .B1(n5376), .B2(n4242), .A(n3949), .ZN(n5331) );
  NAND2_X1 U5007 ( .A1(n3951), .A2(n3950), .ZN(n5329) );
  AOI21_X1 U5008 ( .B1(n3953), .B2(n6666), .A(n3996), .ZN(n6000) );
  OR2_X1 U5009 ( .A1(n6000), .A2(n3818), .ZN(n3968) );
  AOI22_X1 U5010 ( .A1(n3025), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U5011 ( .A1(n4226), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U5012 ( .A1(n4249), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U5013 ( .A1(n4224), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U5014 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3963)
         );
  AOI22_X1 U5015 ( .A1(n4181), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U5016 ( .A1(n4248), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U5017 ( .A1(n4157), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U5018 ( .A1(n4250), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U5019 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3962)
         );
  OAI21_X1 U5020 ( .B1(n3963), .B2(n3962), .A(n3778), .ZN(n3966) );
  NAND2_X1 U5021 ( .A1(n4273), .A2(EAX_REG_15__SCAN_IN), .ZN(n3965) );
  NAND2_X1 U5022 ( .A1(n4272), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3964)
         );
  AND3_X1 U5023 ( .A1(n3966), .A2(n3965), .A3(n3964), .ZN(n3967) );
  INV_X1 U5024 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3969) );
  XNOR2_X1 U5025 ( .A(n3996), .B(n3969), .ZN(n5987) );
  AOI22_X1 U5026 ( .A1(n4273), .A2(EAX_REG_16__SCAN_IN), .B1(n4272), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U5027 ( .A1(n4226), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U5028 ( .A1(n3311), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U5029 ( .A1(n4099), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U5030 ( .A1(n4250), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U5031 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3979)
         );
  AOI22_X1 U5032 ( .A1(n4181), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U5033 ( .A1(n4248), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U5034 ( .A1(n4255), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U5035 ( .A1(n4157), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U5036 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3978)
         );
  OAI21_X1 U5037 ( .B1(n3979), .B2(n3978), .A(n4266), .ZN(n3980) );
  OAI211_X1 U5038 ( .C1(n5987), .C2(n3818), .A(n3981), .B(n3980), .ZN(n5386)
         );
  AOI22_X1 U5039 ( .A1(n4157), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U5040 ( .A1(n4248), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U5041 ( .A1(n4181), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U5042 ( .A1(n4226), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U5043 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3991)
         );
  AOI22_X1 U5044 ( .A1(n4255), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U5045 ( .A1(n4249), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U5046 ( .A1(n3299), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U5047 ( .A1(n4218), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3986) );
  NAND4_X1 U5048 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3990)
         );
  NOR2_X1 U5049 ( .A1(n3991), .A2(n3990), .ZN(n3995) );
  NAND2_X1 U5050 ( .A1(n4378), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3992)
         );
  NAND2_X1 U5051 ( .A1(n3818), .A2(n3992), .ZN(n3993) );
  AOI21_X1 U5052 ( .B1(n4273), .B2(EAX_REG_17__SCAN_IN), .A(n3993), .ZN(n3994)
         );
  OAI21_X1 U5053 ( .B1(n4238), .B2(n3995), .A(n3994), .ZN(n3999) );
  OAI21_X1 U5054 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3997), .A(n4029), 
        .ZN(n5978) );
  INV_X1 U5055 ( .A(n5978), .ZN(n5900) );
  NAND2_X1 U5056 ( .A1(n5900), .A2(n4242), .ZN(n3998) );
  AOI22_X1 U5057 ( .A1(n4157), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5058 ( .A1(n4218), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U5059 ( .A1(n3311), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U5060 ( .A1(n4226), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4000) );
  NAND4_X1 U5061 ( .A1(n4003), .A2(n4002), .A3(n4001), .A4(n4000), .ZN(n4009)
         );
  AOI22_X1 U5062 ( .A1(n4255), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U5063 ( .A1(n4249), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U5064 ( .A1(n4181), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U5065 ( .A1(n4248), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4004) );
  NAND4_X1 U5066 ( .A1(n4007), .A2(n4006), .A3(n4005), .A4(n4004), .ZN(n4008)
         );
  NOR2_X1 U5067 ( .A1(n4009), .A2(n4008), .ZN(n4012) );
  INV_X1 U5068 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5971) );
  OAI21_X1 U5069 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5971), .A(n3818), .ZN(
        n4010) );
  AOI21_X1 U5070 ( .B1(n4273), .B2(EAX_REG_18__SCAN_IN), .A(n4010), .ZN(n4011)
         );
  OAI21_X1 U5071 ( .B1(n4238), .B2(n4012), .A(n4011), .ZN(n4014) );
  XNOR2_X1 U5072 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4029), .ZN(n5969)
         );
  NAND2_X1 U5073 ( .A1(n4242), .A2(n5969), .ZN(n4013) );
  AOI22_X1 U5074 ( .A1(n4248), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U5075 ( .A1(n4249), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U5076 ( .A1(n4255), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U5077 ( .A1(n4181), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4015) );
  NAND4_X1 U5078 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4024)
         );
  AOI22_X1 U5079 ( .A1(n4157), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U5080 ( .A1(n3299), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5081 ( .A1(n4226), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5082 ( .A1(n4250), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4019) );
  NAND4_X1 U5083 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4023)
         );
  NOR2_X1 U5084 ( .A1(n4024), .A2(n4023), .ZN(n4028) );
  OAI21_X1 U5085 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6365), .A(n4378), 
        .ZN(n4025) );
  INV_X1 U5086 ( .A(n4025), .ZN(n4026) );
  AOI21_X1 U5087 ( .B1(n4273), .B2(EAX_REG_19__SCAN_IN), .A(n4026), .ZN(n4027)
         );
  OAI21_X1 U5088 ( .B1(n4238), .B2(n4028), .A(n4027), .ZN(n4033) );
  OAI21_X1 U5089 ( .B1(n4031), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n4065), 
        .ZN(n5878) );
  OR2_X1 U5090 ( .A1(n5878), .A2(n3818), .ZN(n4032) );
  NAND2_X1 U5091 ( .A1(n4033), .A2(n4032), .ZN(n5511) );
  AOI22_X1 U5092 ( .A1(n4181), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4157), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5093 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4249), .B1(n4099), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5094 ( .A1(n4255), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5095 ( .A1(n4218), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4035) );
  NAND4_X1 U5096 ( .A1(n4038), .A2(n4037), .A3(n4036), .A4(n4035), .ZN(n4044)
         );
  AOI22_X1 U5097 ( .A1(n3299), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5098 ( .A1(n4224), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5099 ( .A1(n4248), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5100 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4226), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U5101 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4043)
         );
  NOR2_X1 U5102 ( .A1(n4044), .A2(n4043), .ZN(n4048) );
  NOR2_X1 U5103 ( .A1(n5640), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4045) );
  OR2_X1 U5104 ( .A1(n4242), .A2(n4045), .ZN(n4046) );
  AOI21_X1 U5105 ( .B1(n4273), .B2(EAX_REG_20__SCAN_IN), .A(n4046), .ZN(n4047)
         );
  OAI21_X1 U5106 ( .B1(n4238), .B2(n4048), .A(n4047), .ZN(n4050) );
  XNOR2_X1 U5107 ( .A(n4065), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5870)
         );
  NAND2_X1 U5108 ( .A1(n5870), .A2(n4242), .ZN(n4049) );
  NAND2_X1 U5109 ( .A1(n4050), .A2(n4049), .ZN(n5501) );
  AOI22_X1 U5110 ( .A1(n4248), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5111 ( .A1(n4218), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5112 ( .A1(n4181), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5113 ( .A1(n4224), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4051) );
  NAND4_X1 U5114 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4060)
         );
  AOI22_X1 U5115 ( .A1(n4157), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5116 ( .A1(n3024), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5117 ( .A1(n4249), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5118 ( .A1(n3251), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U5119 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4059)
         );
  NOR2_X1 U5120 ( .A1(n4060), .A2(n4059), .ZN(n4064) );
  NAND2_X1 U5121 ( .A1(n4378), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4061)
         );
  NAND2_X1 U5122 ( .A1(n3818), .A2(n4061), .ZN(n4062) );
  AOI21_X1 U5123 ( .B1(n4273), .B2(EAX_REG_21__SCAN_IN), .A(n4062), .ZN(n4063)
         );
  OAI21_X1 U5124 ( .B1(n4238), .B2(n4064), .A(n4063), .ZN(n4069) );
  OR2_X1 U5125 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4067)
         );
  NAND2_X1 U5126 ( .A1(n4110), .A2(n4067), .ZN(n5860) );
  AOI22_X1 U5127 ( .A1(n3025), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5128 ( .A1(n4181), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5129 ( .A1(n3299), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5130 ( .A1(n4157), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4070) );
  NAND4_X1 U5131 ( .A1(n4073), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4079)
         );
  AOI22_X1 U5132 ( .A1(n4248), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5133 ( .A1(n4249), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5134 ( .A1(n4250), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5135 ( .A1(n4099), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4074) );
  NAND4_X1 U5136 ( .A1(n4077), .A2(n4076), .A3(n4075), .A4(n4074), .ZN(n4078)
         );
  NOR2_X1 U5137 ( .A1(n4079), .A2(n4078), .ZN(n4082) );
  AOI21_X1 U5138 ( .B1(n5626), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4080) );
  AOI21_X1 U5139 ( .B1(n4273), .B2(EAX_REG_22__SCAN_IN), .A(n4080), .ZN(n4081)
         );
  OAI21_X1 U5140 ( .B1(n4238), .B2(n4082), .A(n4081), .ZN(n4084) );
  XNOR2_X1 U5141 ( .A(n4110), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5850)
         );
  NAND2_X1 U5142 ( .A1(n5850), .A2(n4242), .ZN(n4083) );
  AOI22_X1 U5143 ( .A1(n4249), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5144 ( .A1(n3025), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5145 ( .A1(n4157), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5146 ( .A1(n4218), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4085) );
  NAND4_X1 U5147 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4094)
         );
  AOI22_X1 U5148 ( .A1(n4181), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5149 ( .A1(n3299), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5150 ( .A1(n4248), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5151 ( .A1(n4226), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4089) );
  NAND4_X1 U5152 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4093)
         );
  NOR2_X1 U5153 ( .A1(n4094), .A2(n4093), .ZN(n4115) );
  AOI22_X1 U5154 ( .A1(n4255), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5155 ( .A1(n4157), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5156 ( .A1(n3299), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5157 ( .A1(n4257), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4095) );
  NAND4_X1 U5158 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4105)
         );
  AOI22_X1 U5159 ( .A1(n4248), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5160 ( .A1(n4249), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5161 ( .A1(n4181), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5162 ( .A1(n4226), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4100) );
  NAND4_X1 U5163 ( .A1(n4103), .A2(n4102), .A3(n4101), .A4(n4100), .ZN(n4104)
         );
  NOR2_X1 U5164 ( .A1(n4105), .A2(n4104), .ZN(n4116) );
  XNOR2_X1 U5165 ( .A(n4115), .B(n4116), .ZN(n4109) );
  NOR2_X1 U5166 ( .A1(n5618), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4106) );
  OR2_X1 U5167 ( .A1(n4242), .A2(n4106), .ZN(n4107) );
  AOI21_X1 U5168 ( .B1(n4273), .B2(EAX_REG_23__SCAN_IN), .A(n4107), .ZN(n4108)
         );
  OAI21_X1 U5169 ( .B1(n4238), .B2(n4109), .A(n4108), .ZN(n4114) );
  AND2_X1 U5170 ( .A1(n4111), .A2(n5618), .ZN(n4112) );
  OR2_X1 U5171 ( .A1(n4112), .A2(n4150), .ZN(n5841) );
  NAND2_X1 U5172 ( .A1(n5621), .A2(n4242), .ZN(n4113) );
  NAND2_X1 U5173 ( .A1(n4114), .A2(n4113), .ZN(n5480) );
  NOR2_X1 U5174 ( .A1(n4116), .A2(n4115), .ZN(n4146) );
  AOI22_X1 U5175 ( .A1(n3025), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5176 ( .A1(n3248), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5177 ( .A1(n3299), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5178 ( .A1(n4157), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4117) );
  NAND4_X1 U5179 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4127)
         );
  AOI22_X1 U5180 ( .A1(n4248), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5181 ( .A1(n4249), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5182 ( .A1(n4250), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5183 ( .A1(n4121), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4122) );
  NAND4_X1 U5184 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(n4126)
         );
  INV_X1 U5185 ( .A(n4145), .ZN(n4128) );
  XNOR2_X1 U5186 ( .A(n4146), .B(n4128), .ZN(n4133) );
  INV_X1 U5187 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5829) );
  XNOR2_X1 U5188 ( .A(n4150), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5828)
         );
  NAND2_X1 U5189 ( .A1(n5828), .A2(n4242), .ZN(n4130) );
  NAND2_X1 U5190 ( .A1(n4273), .A2(EAX_REG_24__SCAN_IN), .ZN(n4129) );
  OAI211_X1 U5191 ( .C1(n5829), .C2(n4131), .A(n4130), .B(n4129), .ZN(n4132)
         );
  AOI21_X1 U5192 ( .B1(n4133), .B2(n4266), .A(n4132), .ZN(n5474) );
  AOI22_X1 U5193 ( .A1(n3248), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5194 ( .A1(n4223), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5195 ( .A1(n4157), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5196 ( .A1(n4226), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4135) );
  NAND4_X1 U5197 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4144)
         );
  AOI22_X1 U5198 ( .A1(n4249), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5199 ( .A1(n4255), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5200 ( .A1(n4248), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5201 ( .A1(n4099), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4139) );
  NAND4_X1 U5202 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4143)
         );
  NOR2_X1 U5203 ( .A1(n4144), .A2(n4143), .ZN(n4156) );
  NAND2_X1 U5204 ( .A1(n4146), .A2(n4145), .ZN(n4155) );
  XNOR2_X1 U5205 ( .A(n4156), .B(n4155), .ZN(n4149) );
  INV_X1 U5206 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5601) );
  AOI21_X1 U5207 ( .B1(n5601), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4147) );
  AOI21_X1 U5208 ( .B1(n4273), .B2(EAX_REG_25__SCAN_IN), .A(n4147), .ZN(n4148)
         );
  OAI21_X1 U5209 ( .B1(n4149), .B2(n4238), .A(n4148), .ZN(n4154) );
  OR2_X1 U5210 ( .A1(n4151), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4152)
         );
  NAND2_X1 U5211 ( .A1(n4193), .A2(n4152), .ZN(n5818) );
  NOR2_X1 U5212 ( .A1(n4156), .A2(n4155), .ZN(n4176) );
  AOI22_X1 U5213 ( .A1(n3024), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5214 ( .A1(n3248), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5215 ( .A1(n3299), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5216 ( .A1(n4157), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4158) );
  NAND4_X1 U5217 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4167)
         );
  AOI22_X1 U5218 ( .A1(n4248), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4226), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U5219 ( .A1(n4249), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5220 ( .A1(n4250), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5221 ( .A1(n4099), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4162) );
  NAND4_X1 U5222 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4166)
         );
  OR2_X1 U5223 ( .A1(n4167), .A2(n4166), .ZN(n4175) );
  INV_X1 U5224 ( .A(n4175), .ZN(n4168) );
  XNOR2_X1 U5225 ( .A(n4176), .B(n4168), .ZN(n4169) );
  NAND2_X1 U5226 ( .A1(n4169), .A2(n4266), .ZN(n4174) );
  NOR2_X1 U5227 ( .A1(n5595), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4170) );
  OR2_X1 U5228 ( .A1(n4242), .A2(n4170), .ZN(n4171) );
  AOI21_X1 U5229 ( .B1(n3794), .B2(EAX_REG_26__SCAN_IN), .A(n4171), .ZN(n4173)
         );
  XNOR2_X1 U5230 ( .A(n4193), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5808)
         );
  AOI21_X1 U5231 ( .B1(n4174), .B2(n4173), .A(n4172), .ZN(n5461) );
  NAND2_X1 U5232 ( .A1(n4176), .A2(n4175), .ZN(n4197) );
  AOI22_X1 U5233 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4248), .B1(n4218), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5234 ( .A1(n3299), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5235 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4249), .B1(n4257), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5236 ( .A1(n4226), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4177) );
  NAND4_X1 U5237 ( .A1(n4180), .A2(n4179), .A3(n4178), .A4(n4177), .ZN(n4187)
         );
  AOI22_X1 U5238 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4181), .B1(n3247), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U5239 ( .A1(n3024), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U5240 ( .A1(n3175), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U5241 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4099), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4182) );
  NAND4_X1 U5242 ( .A1(n4185), .A2(n4184), .A3(n4183), .A4(n4182), .ZN(n4186)
         );
  NOR2_X1 U5243 ( .A1(n4187), .A2(n4186), .ZN(n4198) );
  XNOR2_X1 U5244 ( .A(n4197), .B(n4198), .ZN(n4191) );
  NOR2_X1 U5245 ( .A1(n4192), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4188) );
  OR2_X1 U5246 ( .A1(n4242), .A2(n4188), .ZN(n4189) );
  AOI21_X1 U5247 ( .B1(n3794), .B2(EAX_REG_27__SCAN_IN), .A(n4189), .ZN(n4190)
         );
  OAI21_X1 U5248 ( .B1(n4191), .B2(n4238), .A(n4190), .ZN(n4196) );
  OAI21_X1 U5249 ( .B1(n4193), .B2(n5595), .A(n4192), .ZN(n4194) );
  NAND2_X1 U5250 ( .A1(n4194), .A2(n4213), .ZN(n5587) );
  NAND2_X1 U5251 ( .A1(n4196), .A2(n4195), .ZN(n5437) );
  NOR2_X1 U5252 ( .A1(n4198), .A2(n4197), .ZN(n4234) );
  AOI22_X1 U5253 ( .A1(n3316), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5254 ( .A1(n4181), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5255 ( .A1(n3311), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5256 ( .A1(n3175), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4199) );
  NAND4_X1 U5257 ( .A1(n4202), .A2(n4201), .A3(n4200), .A4(n4199), .ZN(n4208)
         );
  AOI22_X1 U5258 ( .A1(n4248), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3240), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5259 ( .A1(n4249), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5260 ( .A1(n4250), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U5261 ( .A1(n4099), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4203) );
  NAND4_X1 U5262 ( .A1(n4206), .A2(n4205), .A3(n4204), .A4(n4203), .ZN(n4207)
         );
  OR2_X1 U5263 ( .A1(n4208), .A2(n4207), .ZN(n4233) );
  XNOR2_X1 U5264 ( .A(n4234), .B(n4233), .ZN(n4212) );
  NOR2_X1 U5265 ( .A1(n5576), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4209) );
  OR2_X1 U5266 ( .A1(n4242), .A2(n4209), .ZN(n4210) );
  AOI21_X1 U5267 ( .B1(n3794), .B2(EAX_REG_28__SCAN_IN), .A(n4210), .ZN(n4211)
         );
  OAI21_X1 U5268 ( .B1(n4212), .B2(n4238), .A(n4211), .ZN(n4216) );
  AND2_X1 U5269 ( .A1(n4213), .A2(n5576), .ZN(n4214) );
  NOR2_X1 U5270 ( .A1(n4240), .A2(n4214), .ZN(n5580) );
  NAND2_X1 U5271 ( .A1(n5580), .A2(n4242), .ZN(n4215) );
  NAND2_X1 U5272 ( .A1(n4216), .A2(n4215), .ZN(n4290) );
  AOI22_X1 U5273 ( .A1(n3248), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5274 ( .A1(n4255), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5275 ( .A1(n4099), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5276 ( .A1(n4218), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4219) );
  NAND4_X1 U5277 ( .A1(n4222), .A2(n4221), .A3(n4220), .A4(n4219), .ZN(n4232)
         );
  AOI22_X1 U5278 ( .A1(n3241), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4249), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4230) );
  AOI22_X1 U5279 ( .A1(n4224), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U5280 ( .A1(n3175), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U5281 ( .A1(n4226), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4227) );
  NAND4_X1 U5282 ( .A1(n4230), .A2(n4229), .A3(n4228), .A4(n4227), .ZN(n4231)
         );
  NOR2_X1 U5283 ( .A1(n4232), .A2(n4231), .ZN(n4247) );
  NAND2_X1 U5284 ( .A1(n4234), .A2(n4233), .ZN(n4246) );
  XNOR2_X1 U5285 ( .A(n4247), .B(n4246), .ZN(n4239) );
  NAND2_X1 U5286 ( .A1(n4378), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4235)
         );
  NAND2_X1 U5287 ( .A1(n3818), .A2(n4235), .ZN(n4236) );
  AOI21_X1 U5288 ( .B1(n3794), .B2(EAX_REG_29__SCAN_IN), .A(n4236), .ZN(n4237)
         );
  OAI21_X1 U5289 ( .B1(n4239), .B2(n4238), .A(n4237), .ZN(n4245) );
  NAND2_X1 U5290 ( .A1(n4240), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4281)
         );
  OR2_X1 U5291 ( .A1(n4240), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4241)
         );
  NAND2_X1 U5292 ( .A1(n4281), .A2(n4241), .ZN(n5799) );
  INV_X1 U5293 ( .A(n5799), .ZN(n4243) );
  NAND2_X1 U5294 ( .A1(n4243), .A2(n4242), .ZN(n4244) );
  NOR2_X1 U5295 ( .A1(n4247), .A2(n4246), .ZN(n4265) );
  AOI22_X1 U5296 ( .A1(n4248), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3240), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5297 ( .A1(n4249), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4218), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5298 ( .A1(n3311), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U5299 ( .A1(n3175), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4250), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4251) );
  NAND4_X1 U5300 ( .A1(n4254), .A2(n4253), .A3(n4252), .A4(n4251), .ZN(n4263)
         );
  AOI22_X1 U5301 ( .A1(n3316), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4261) );
  AOI22_X1 U5302 ( .A1(n4181), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4256), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4260) );
  AOI22_X1 U5303 ( .A1(n4099), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4257), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4259) );
  AOI22_X1 U5304 ( .A1(n3251), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4592), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4258) );
  NAND4_X1 U5305 ( .A1(n4261), .A2(n4260), .A3(n4259), .A4(n4258), .ZN(n4262)
         );
  NOR2_X1 U5306 ( .A1(n4263), .A2(n4262), .ZN(n4264) );
  XNOR2_X1 U5307 ( .A(n4265), .B(n4264), .ZN(n4267) );
  NAND2_X1 U5308 ( .A1(n4267), .A2(n4266), .ZN(n4271) );
  INV_X1 U5309 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5424) );
  AOI21_X1 U5310 ( .B1(n5424), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4268) );
  AOI21_X1 U5311 ( .B1(n4273), .B2(EAX_REG_30__SCAN_IN), .A(n4268), .ZN(n4270)
         );
  XNOR2_X1 U5312 ( .A(n4281), .B(n5424), .ZN(n5423) );
  INV_X1 U5313 ( .A(n5423), .ZN(n4269) );
  AOI22_X1 U5314 ( .A1(n4271), .A2(n4270), .B1(n4242), .B2(n4269), .ZN(n4348)
         );
  NAND2_X1 U5315 ( .A1(n5451), .A2(n4348), .ZN(n4276) );
  AOI22_X1 U5316 ( .A1(n4273), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4272), .ZN(n4274) );
  INV_X1 U5317 ( .A(n4274), .ZN(n4275) );
  NAND2_X1 U5318 ( .A1(n4294), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6511) );
  NAND2_X1 U5319 ( .A1(n4344), .A2(n6184), .ZN(n4287) );
  NAND2_X1 U5320 ( .A1(n6316), .A2(n4277), .ZN(n6610) );
  NAND2_X1 U5321 ( .A1(n6610), .A2(n6506), .ZN(n4278) );
  NAND2_X1 U5322 ( .A1(n6506), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4280) );
  NAND2_X1 U5323 ( .A1(n6365), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U5324 ( .A1(n4280), .A2(n4279), .ZN(n6207) );
  INV_X1 U5325 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4328) );
  NAND2_X1 U5326 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4283)
         );
  OAI211_X1 U5327 ( .C1(n6202), .C2(n4305), .A(n4284), .B(n4283), .ZN(n4285)
         );
  INV_X1 U5328 ( .A(n4285), .ZN(n4286) );
  NAND3_X1 U5329 ( .A1(n4288), .A2(n4287), .A3(n4286), .ZN(U2955) );
  INV_X1 U5330 ( .A(n4406), .ZN(n4293) );
  NAND2_X1 U5331 ( .A1(n3620), .A2(n4293), .ZN(n4402) );
  INV_X1 U5332 ( .A(n6614), .ZN(n6498) );
  NOR3_X1 U5333 ( .A1(n6506), .A2(n6591), .A3(n6498), .ZN(n6496) );
  AND2_X1 U5334 ( .A1(n4294), .A2(n4242), .ZN(n4295) );
  NAND2_X1 U5335 ( .A1(n5440), .A2(n4299), .ZN(n4300) );
  NAND2_X1 U5336 ( .A1(n5453), .A2(n4300), .ZN(n5683) );
  NAND2_X1 U5337 ( .A1(n6365), .A2(n6611), .ZN(n4315) );
  NAND2_X1 U5338 ( .A1(n4315), .A2(EBX_REG_31__SCAN_IN), .ZN(n4301) );
  NOR2_X1 U5339 ( .A1(n3027), .A2(n4301), .ZN(n4302) );
  INV_X1 U5340 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6572) );
  INV_X1 U5341 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6568) );
  INV_X1 U5342 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6562) );
  INV_X1 U5343 ( .A(n4315), .ZN(n4314) );
  AND3_X1 U5344 ( .A1(n4303), .A2(n4314), .A3(n3265), .ZN(n4304) );
  INV_X1 U5345 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6551) );
  INV_X1 U5346 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6535) );
  NAND3_X1 U5347 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6060) );
  NOR2_X1 U5348 ( .A1(n6535), .A2(n6060), .ZN(n4958) );
  NAND2_X1 U5349 ( .A1(REIP_REG_5__SCAN_IN), .A2(n4958), .ZN(n4949) );
  NAND3_X1 U5350 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n6019) );
  NOR2_X1 U5351 ( .A1(n4949), .A2(n6019), .ZN(n5286) );
  NAND4_X1 U5352 ( .A1(n5286), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U5353 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5333) );
  NOR3_X1 U5354 ( .A1(n6551), .A2(n5281), .A3(n5333), .ZN(n4307) );
  NAND2_X1 U5355 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n4308) );
  INV_X1 U5356 ( .A(n5882), .ZN(n5972) );
  INV_X1 U5357 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6560) );
  NAND3_X1 U5358 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        n5862), .ZN(n5840) );
  NAND3_X1 U5359 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        n5836), .ZN(n5815) );
  NOR2_X1 U5360 ( .A1(n6572), .A2(n5815), .ZN(n5445) );
  INV_X1 U5361 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6673) );
  INV_X1 U5362 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6575) );
  NOR2_X1 U5363 ( .A1(n6673), .A2(n6575), .ZN(n4313) );
  NAND2_X1 U5364 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5854) );
  INV_X1 U5365 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U5366 ( .A1(n4307), .A2(n6080), .ZN(n5334) );
  NOR3_X1 U5367 ( .A1(n6553), .A2(n4308), .A3(n5334), .ZN(n5876) );
  NAND4_X1 U5368 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5876), .ZN(n5849) );
  NOR2_X1 U5369 ( .A1(n5854), .A2(n5849), .ZN(n4309) );
  AOI21_X1 U5370 ( .B1(REIP_REG_23__SCAN_IN), .B2(n4309), .A(n5875), .ZN(n5831) );
  NAND2_X1 U5371 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5823) );
  INV_X1 U5372 ( .A(n5823), .ZN(n4310) );
  NAND2_X1 U5373 ( .A1(REIP_REG_26__SCAN_IN), .A2(n4310), .ZN(n4311) );
  AND2_X1 U5374 ( .A1(n6082), .A2(n4311), .ZN(n4312) );
  OAI21_X1 U5375 ( .B1(n4313), .B2(n6079), .A(n5816), .ZN(n4324) );
  AOI22_X1 U5376 ( .A1(n5580), .A2(n6062), .B1(REIP_REG_28__SCAN_IN), .B2(
        n4324), .ZN(n4319) );
  INV_X1 U5377 ( .A(n6520), .ZN(n5014) );
  NAND2_X1 U5378 ( .A1(n5014), .A2(n4314), .ZN(n6492) );
  AND2_X1 U5379 ( .A1(n4424), .A2(n6492), .ZN(n4325) );
  INV_X1 U5380 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5448) );
  AND3_X1 U5381 ( .A1(n3265), .A2(n5448), .A3(n4315), .ZN(n4316) );
  OR2_X1 U5382 ( .A1(n4325), .A2(n4316), .ZN(n4317) );
  AOI22_X1 U5383 ( .A1(EBX_REG_28__SCAN_IN), .A2(n6054), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6087), .ZN(n4318) );
  NAND2_X1 U5384 ( .A1(n4319), .A2(n4318), .ZN(n4320) );
  INV_X1 U5385 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U5386 ( .A1(n4324), .A2(n6580), .ZN(n5797) );
  INV_X1 U5387 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6584) );
  AOI211_X1 U5388 ( .C1(n5797), .C2(REIP_REG_30__SCAN_IN), .A(n5875), .B(n6584), .ZN(n4330) );
  NAND3_X1 U5389 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5445), .ZN(n5798) );
  INV_X1 U5390 ( .A(n5798), .ZN(n5427) );
  NAND4_X1 U5391 ( .A1(n6584), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n5427), .ZN(n4327) );
  NAND3_X1 U5392 ( .A1(n6609), .A2(EBX_REG_31__SCAN_IN), .A3(n4325), .ZN(n4326) );
  OAI211_X1 U5393 ( .C1(n6075), .C2(n4328), .A(n4327), .B(n4326), .ZN(n4329)
         );
  AOI211_X1 U5394 ( .C1(n5447), .C2(n6067), .A(n4330), .B(n4329), .ZN(n4333)
         );
  NAND2_X1 U5395 ( .A1(n4344), .A2(n4331), .ZN(n4332) );
  NAND2_X1 U5396 ( .A1(n4333), .A2(n4332), .ZN(U2796) );
  NOR2_X1 U5397 ( .A1(n3335), .A2(n4335), .ZN(n4336) );
  NAND3_X1 U5398 ( .A1(n4337), .A2(n4336), .A3(n3237), .ZN(n4351) );
  NOR2_X1 U5399 ( .A1(n3027), .A2(READY_N), .ZN(n4338) );
  INV_X1 U5400 ( .A(n4340), .ZN(n4341) );
  OAI22_X1 U5401 ( .A1(n4473), .A2(n4407), .B1(n3634), .B2(n4341), .ZN(n4475)
         );
  NAND2_X1 U5402 ( .A1(n4475), .A2(n6503), .ZN(n4342) );
  NAND2_X1 U5403 ( .A1(n4344), .A2(n3100), .ZN(n4347) );
  AND2_X1 U5404 ( .A1(n5541), .A2(n4345), .ZN(n6622) );
  AOI22_X1 U5405 ( .A1(n6622), .A2(DATAI_31_), .B1(n6620), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n4346) );
  NAND2_X1 U5406 ( .A1(n4347), .A2(n4346), .ZN(U2860) );
  AND2_X1 U5407 ( .A1(n4466), .A2(n6503), .ZN(n4350) );
  NAND2_X1 U5408 ( .A1(n4473), .A2(n4350), .ZN(n4357) );
  INV_X1 U5409 ( .A(n4351), .ZN(n4355) );
  NOR2_X1 U5410 ( .A1(n4352), .A2(n3027), .ZN(n4354) );
  NAND2_X1 U5411 ( .A1(n4355), .A2(n4354), .ZN(n4356) );
  NAND2_X1 U5412 ( .A1(n5422), .A2(n5350), .ZN(n4367) );
  INV_X1 U5413 ( .A(n4361), .ZN(n4358) );
  AOI211_X1 U5414 ( .C1(n3651), .C2(n5453), .A(n4361), .B(n4360), .ZN(n4362)
         );
  AOI21_X1 U5415 ( .B1(n4364), .B2(n4363), .A(n4362), .ZN(n5433) );
  INV_X1 U5416 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5431) );
  INV_X1 U5417 ( .A(n4365), .ZN(n4366) );
  AND2_X1 U5418 ( .A1(n5778), .A2(n4370), .ZN(n4371) );
  NAND2_X1 U5419 ( .A1(n6367), .A2(n6365), .ZN(n6317) );
  AOI22_X1 U5420 ( .A1(n4737), .A2(n6317), .B1(n5171), .B2(n5111), .ZN(n4381)
         );
  NAND2_X1 U5421 ( .A1(n4792), .A2(n4810), .ZN(n4672) );
  NAND2_X1 U5422 ( .A1(n4672), .A2(n6367), .ZN(n4376) );
  NAND2_X1 U5423 ( .A1(n4376), .A2(n6317), .ZN(n4669) );
  NOR3_X1 U5424 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4671) );
  NAND2_X1 U5425 ( .A1(n6632), .A2(n4671), .ZN(n4735) );
  AND2_X1 U5426 ( .A1(n4384), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6361) );
  INV_X1 U5427 ( .A(n4909), .ZN(n4377) );
  INV_X1 U5428 ( .A(n4910), .ZN(n4634) );
  OAI21_X1 U5429 ( .B1(n3102), .B2(n4378), .A(n4634), .ZN(n5065) );
  AOI211_X1 U5430 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4735), .A(n6361), .B(
        n5065), .ZN(n4379) );
  INV_X1 U5431 ( .A(n4379), .ZN(n4380) );
  AOI21_X1 U5432 ( .B1(n4381), .B2(n4669), .A(n4380), .ZN(n4712) );
  NOR2_X1 U5433 ( .A1(n4712), .A2(n4382), .ZN(n4390) );
  NAND2_X1 U5434 ( .A1(n6184), .A2(DATAI_17_), .ZN(n6381) );
  NOR2_X1 U5435 ( .A1(n4745), .A2(n6381), .ZN(n4389) );
  NAND2_X1 U5436 ( .A1(n6184), .A2(DATAI_25_), .ZN(n6421) );
  INV_X1 U5437 ( .A(n6421), .ZN(n6378) );
  AND2_X1 U5438 ( .A1(n4737), .A2(n6378), .ZN(n4388) );
  NAND3_X1 U5439 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6506), .A3(n4383), .ZN(
        n4565) );
  NAND2_X1 U5440 ( .A1(n4578), .A2(n4421), .ZN(n5215) );
  NOR2_X1 U5441 ( .A1(n3023), .A2(n6316), .ZN(n6358) );
  NAND2_X1 U5442 ( .A1(n6358), .A2(n5111), .ZN(n4386) );
  NOR2_X1 U5443 ( .A1(n4384), .A2(n4378), .ZN(n6314) );
  NAND2_X1 U5444 ( .A1(n3102), .A2(n6314), .ZN(n4385) );
  INV_X1 U5445 ( .A(DATAI_1_), .ZN(n6153) );
  OAI22_X1 U5446 ( .A1(n5215), .A2(n4735), .B1(n4734), .B2(n5219), .ZN(n4387)
         );
  OR4_X1 U5447 ( .A1(n4390), .A2(n4389), .A3(n4388), .A4(n4387), .ZN(U3021) );
  NOR2_X1 U5448 ( .A1(n4712), .A2(n4391), .ZN(n4396) );
  NAND2_X1 U5449 ( .A1(n6184), .A2(DATAI_18_), .ZN(n6387) );
  NOR2_X1 U5450 ( .A1(n4745), .A2(n6387), .ZN(n4395) );
  INV_X1 U5451 ( .A(DATAI_26_), .ZN(n4392) );
  NOR2_X1 U5452 ( .A1(n6211), .A2(n4392), .ZN(n6384) );
  AND2_X1 U5453 ( .A1(n4737), .A2(n6384), .ZN(n4394) );
  NAND2_X1 U5454 ( .A1(n4578), .A2(n3259), .ZN(n5210) );
  INV_X1 U5455 ( .A(DATAI_2_), .ZN(n6155) );
  OAI22_X1 U5456 ( .A1(n5210), .A2(n4735), .B1(n4734), .B2(n5214), .ZN(n4393)
         );
  OR4_X1 U5457 ( .A1(n4396), .A2(n4395), .A3(n4394), .A4(n4393), .ZN(U3022) );
  NOR2_X1 U5458 ( .A1(n4712), .A2(n4397), .ZN(n4401) );
  NAND2_X1 U5459 ( .A1(n6184), .A2(DATAI_16_), .ZN(n6377) );
  NOR2_X1 U5460 ( .A1(n4745), .A2(n6377), .ZN(n4400) );
  NAND2_X1 U5461 ( .A1(n6184), .A2(DATAI_24_), .ZN(n6436) );
  NOR2_X1 U5462 ( .A1(n4585), .A2(n6436), .ZN(n4399) );
  NAND2_X1 U5463 ( .A1(n4578), .A2(n3265), .ZN(n5220) );
  INV_X1 U5464 ( .A(DATAI_0_), .ZN(n6151) );
  OAI22_X1 U5465 ( .A1(n5220), .A2(n4735), .B1(n4734), .B2(n5224), .ZN(n4398)
         );
  OR4_X1 U5466 ( .A1(n4401), .A2(n4400), .A3(n4399), .A4(n4398), .ZN(U3020) );
  NAND2_X1 U5467 ( .A1(n4473), .A2(n3561), .ZN(n4404) );
  NAND2_X1 U5468 ( .A1(n4402), .A2(n3018), .ZN(n4403) );
  NAND2_X1 U5469 ( .A1(n4404), .A2(n4403), .ZN(n5948) );
  OR2_X1 U5470 ( .A1(n5170), .A2(n4424), .ZN(n4419) );
  AOI21_X1 U5471 ( .B1(n4419), .B2(n6520), .A(READY_N), .ZN(n6613) );
  OR2_X1 U5472 ( .A1(n5948), .A2(n6613), .ZN(n6484) );
  AND2_X1 U5473 ( .A1(n6484), .A2(n6503), .ZN(n5954) );
  INV_X1 U5474 ( .A(MORE_REG_SCAN_IN), .ZN(n4415) );
  INV_X1 U5475 ( .A(n4466), .ZN(n4405) );
  OR2_X1 U5476 ( .A1(n4473), .A2(n4405), .ZN(n4412) );
  NAND2_X1 U5477 ( .A1(n3620), .A2(n4406), .ZN(n4411) );
  INV_X1 U5478 ( .A(n4407), .ZN(n4453) );
  OR3_X1 U5479 ( .A1(n4408), .A2(n4453), .A3(n4292), .ZN(n4409) );
  NAND2_X1 U5480 ( .A1(n4473), .A2(n4409), .ZN(n4410) );
  AND3_X1 U5481 ( .A1(n4412), .A2(n4411), .A3(n4410), .ZN(n6482) );
  INV_X1 U5482 ( .A(n6482), .ZN(n4413) );
  NAND2_X1 U5483 ( .A1(n5954), .A2(n4413), .ZN(n4414) );
  OAI21_X1 U5484 ( .B1(n5954), .B2(n4415), .A(n4414), .ZN(U3471) );
  INV_X1 U5485 ( .A(n4422), .ZN(n4423) );
  AOI211_X1 U5486 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4416), .A(n5947), .B(
        n4423), .ZN(n4417) );
  INV_X1 U5487 ( .A(n4417), .ZN(U2788) );
  INV_X1 U5488 ( .A(n6609), .ZN(n4420) );
  OAI21_X1 U5489 ( .B1(n5947), .B2(READREQUEST_REG_SCAN_IN), .A(n4420), .ZN(
        n4418) );
  OAI21_X1 U5490 ( .B1(n4420), .B2(n4419), .A(n4418), .ZN(U3474) );
  INV_X1 U5491 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U5492 ( .A1(n4478), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4425) );
  NAND2_X1 U5493 ( .A1(n4494), .A2(DATAI_9_), .ZN(n4487) );
  OAI211_X1 U5494 ( .C1(n6144), .C2(n5017), .A(n4425), .B(n4487), .ZN(U2933)
         );
  INV_X1 U5495 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U5496 ( .A1(n4478), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U5497 ( .A1(n4494), .A2(DATAI_8_), .ZN(n4492) );
  OAI211_X1 U5498 ( .C1(n5051), .C2(n6144), .A(n4426), .B(n4492), .ZN(U2932)
         );
  INV_X1 U5499 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U5500 ( .A1(n4478), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4427) );
  NAND2_X1 U5501 ( .A1(n4494), .A2(DATAI_10_), .ZN(n4484) );
  OAI211_X1 U5502 ( .C1(n5057), .C2(n6144), .A(n4427), .B(n4484), .ZN(U2934)
         );
  OR2_X1 U5503 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4430)
         );
  NAND2_X1 U5504 ( .A1(n4430), .A2(n4429), .ZN(n5417) );
  XNOR2_X1 U5505 ( .A(n4432), .B(n4431), .ZN(n6212) );
  OAI222_X1 U5506 ( .A1(n5417), .A2(n5536), .B1(n5538), .B2(n3642), .C1(n3010), 
        .C2(n6212), .ZN(U2859) );
  NOR2_X1 U5507 ( .A1(n4433), .A2(n4434), .ZN(n4435) );
  NOR2_X1 U5508 ( .A1(n4436), .A2(n4435), .ZN(n6099) );
  INV_X1 U5509 ( .A(n6099), .ZN(n4556) );
  OAI21_X1 U5510 ( .B1(n4439), .B2(n4438), .A(n4437), .ZN(n4522) );
  INV_X1 U5511 ( .A(n4522), .ZN(n6092) );
  OAI222_X1 U5512 ( .A1(n4556), .A2(n3010), .B1(n5538), .B2(n6095), .C1(n5536), 
        .C2(n6092), .ZN(U2858) );
  XNOR2_X1 U5513 ( .A(n4440), .B(n4447), .ZN(n6205) );
  AOI21_X1 U5514 ( .B1(n4441), .B2(n5363), .A(n4447), .ZN(n4444) );
  NAND2_X1 U5515 ( .A1(n6282), .A2(REIP_REG_0__SCAN_IN), .ZN(n6203) );
  OAI211_X1 U5516 ( .C1(n6304), .C2(n5417), .A(n4442), .B(n6203), .ZN(n4443)
         );
  AOI211_X1 U5517 ( .C1(n6307), .C2(n6205), .A(n4444), .B(n4443), .ZN(n4445)
         );
  INV_X1 U5518 ( .A(n4445), .ZN(U3018) );
  NOR2_X1 U5519 ( .A1(n6592), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4462)
         );
  NOR2_X1 U5520 ( .A1(n6784), .A2(n4447), .ZN(n5791) );
  INV_X1 U5521 ( .A(n5791), .ZN(n4448) );
  AOI22_X1 U5522 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6664), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4520), .ZN(n5790) );
  NOR2_X1 U5523 ( .A1(n4448), .A2(n5790), .ZN(n4461) );
  NOR2_X1 U5524 ( .A1(n3020), .A2(n4449), .ZN(n4450) );
  AND2_X1 U5525 ( .A1(n3634), .A2(n4450), .ZN(n4451) );
  NAND2_X1 U5526 ( .A1(n4452), .A2(n4451), .ZN(n5789) );
  XNOR2_X1 U5527 ( .A(n4446), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4458)
         );
  OR2_X1 U5528 ( .A1(n4466), .A2(n4453), .ZN(n4591) );
  NAND2_X1 U5529 ( .A1(n4591), .A2(n4458), .ZN(n4457) );
  NAND2_X1 U5530 ( .A1(n5412), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U5531 ( .A1(n5412), .A2(n4454), .ZN(n5785) );
  MUX2_X1 U5532 ( .A(n4455), .B(n5785), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4456) );
  OAI211_X1 U5533 ( .C1(n4458), .C2(n4594), .A(n4457), .B(n4456), .ZN(n4459)
         );
  AOI21_X1 U5534 ( .B1(n4374), .B2(n5789), .A(n4459), .ZN(n4599) );
  NOR2_X1 U5535 ( .A1(n4599), .A2(n6594), .ZN(n4460) );
  AOI211_X1 U5536 ( .C1(n4446), .C2(n4462), .A(n4461), .B(n4460), .ZN(n4477)
         );
  NAND2_X1 U5537 ( .A1(n5412), .A2(n5014), .ZN(n4463) );
  NAND2_X1 U5538 ( .A1(n4463), .A2(n3018), .ZN(n4465) );
  NAND2_X1 U5539 ( .A1(n4465), .A2(n4464), .ZN(n4472) );
  NAND2_X1 U5540 ( .A1(n4473), .A2(n4466), .ZN(n4471) );
  OR2_X1 U5541 ( .A1(n4467), .A2(n3259), .ZN(n4468) );
  AND2_X1 U5542 ( .A1(n4469), .A2(n4468), .ZN(n4470) );
  OAI211_X1 U5543 ( .C1(n4473), .C2(n4472), .A(n4471), .B(n4470), .ZN(n4474)
         );
  OR2_X1 U5544 ( .A1(n4475), .A2(n4474), .ZN(n4608) );
  INV_X1 U5545 ( .A(n4608), .ZN(n6470) );
  INV_X1 U5546 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5953) );
  NAND2_X1 U5547 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4620), .ZN(n6589) );
  OAI22_X1 U5548 ( .A1(n6470), .A2(n6501), .B1(n5953), .B2(n6589), .ZN(n4506)
         );
  AOI21_X1 U5549 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6506), .A(n4506), .ZN(
        n5795) );
  NOR2_X1 U5550 ( .A1(n4446), .A2(n6592), .ZN(n5793) );
  OAI21_X1 U5551 ( .B1(n5793), .B2(n5795), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4476) );
  OAI21_X1 U5552 ( .B1(n4477), .B2(n5795), .A(n4476), .ZN(U3459) );
  INV_X1 U5553 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4479) );
  INV_X1 U5554 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5023) );
  OAI222_X1 U5555 ( .A1(n6151), .A2(n6168), .B1(n4479), .B2(n6143), .C1(n6144), 
        .C2(n5023), .ZN(U2924) );
  INV_X1 U5556 ( .A(DATAI_15_), .ZN(n4481) );
  INV_X1 U5557 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4480) );
  INV_X1 U5558 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6113) );
  OAI222_X1 U5559 ( .A1(n4481), .A2(n6168), .B1(n4480), .B2(n6143), .C1(n6144), 
        .C2(n6113), .ZN(U2954) );
  INV_X1 U5560 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4482) );
  INV_X1 U5561 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5021) );
  OAI222_X1 U5562 ( .A1(n6153), .A2(n6168), .B1(n4482), .B2(n6143), .C1(n6144), 
        .C2(n5021), .ZN(U2925) );
  INV_X1 U5563 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n4483) );
  INV_X1 U5564 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5019) );
  OAI222_X1 U5565 ( .A1(n6155), .A2(n6168), .B1(n4483), .B2(n6143), .C1(n6144), 
        .C2(n5019), .ZN(U2926) );
  INV_X1 U5566 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U5567 ( .A1(n4498), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4485) );
  OAI211_X1 U5568 ( .C1(n6122), .C2(n6144), .A(n4485), .B(n4484), .ZN(U2949)
         );
  INV_X1 U5569 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U5570 ( .A1(n4498), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U5571 ( .A1(n4494), .A2(DATAI_13_), .ZN(n4489) );
  OAI211_X1 U5572 ( .C1(n6755), .C2(n6144), .A(n4486), .B(n4489), .ZN(U2937)
         );
  INV_X1 U5573 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U5574 ( .A1(n4498), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4488) );
  OAI211_X1 U5575 ( .C1(n6124), .C2(n6144), .A(n4488), .B(n4487), .ZN(U2948)
         );
  INV_X1 U5576 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U5577 ( .A1(n4498), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4490) );
  OAI211_X1 U5578 ( .C1(n6117), .C2(n6144), .A(n4490), .B(n4489), .ZN(U2952)
         );
  INV_X1 U5579 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U5580 ( .A1(n4498), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U5581 ( .A1(n4494), .A2(DATAI_14_), .ZN(n4496) );
  OAI211_X1 U5582 ( .C1(n5045), .C2(n6144), .A(n4491), .B(n4496), .ZN(U2938)
         );
  INV_X1 U5583 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U5584 ( .A1(n4498), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4493) );
  OAI211_X1 U5585 ( .C1(n6126), .C2(n6144), .A(n4493), .B(n4492), .ZN(U2947)
         );
  INV_X1 U5586 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U5587 ( .A1(n4498), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U5588 ( .A1(n4494), .A2(DATAI_11_), .ZN(n4499) );
  OAI211_X1 U5589 ( .C1(n6120), .C2(n6144), .A(n4495), .B(n4499), .ZN(U2950)
         );
  INV_X1 U5590 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U5591 ( .A1(n4498), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4497) );
  OAI211_X1 U5592 ( .C1(n6115), .C2(n6144), .A(n4497), .B(n4496), .ZN(U2953)
         );
  INV_X1 U5593 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U5594 ( .A1(n4498), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4500) );
  OAI211_X1 U5595 ( .C1(n5059), .C2(n6144), .A(n4500), .B(n4499), .ZN(U2935)
         );
  INV_X1 U5596 ( .A(DATAI_3_), .ZN(n4502) );
  INV_X1 U5597 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4501) );
  INV_X1 U5598 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5049) );
  OAI222_X1 U5599 ( .A1(n4502), .A2(n6168), .B1(n4501), .B2(n6143), .C1(n5049), 
        .C2(n6144), .ZN(U2927) );
  INV_X1 U5600 ( .A(n4970), .ZN(n4867) );
  NOR2_X1 U5601 ( .A1(n4503), .A2(n4867), .ZN(n4504) );
  XNOR2_X1 U5602 ( .A(n4504), .B(n4507), .ZN(n6064) );
  INV_X1 U5603 ( .A(n3634), .ZN(n4505) );
  NAND2_X1 U5604 ( .A1(n6064), .A2(n4505), .ZN(n4607) );
  NAND2_X1 U5605 ( .A1(n5411), .A2(n4506), .ZN(n4508) );
  INV_X1 U5606 ( .A(n5795), .ZN(n6596) );
  OAI22_X1 U5607 ( .A1(n4607), .A2(n4508), .B1(n4507), .B2(n6596), .ZN(U3455)
         );
  NAND2_X1 U5608 ( .A1(n4510), .A2(n4511), .ZN(n4512) );
  NAND2_X1 U5609 ( .A1(n4509), .A2(n4512), .ZN(n5176) );
  OR2_X1 U5610 ( .A1(n3041), .A2(n4513), .ZN(n4514) );
  AND2_X1 U5611 ( .A1(n4514), .A2(n4629), .ZN(n6289) );
  INV_X1 U5612 ( .A(n5538), .ZN(n4864) );
  AOI22_X1 U5613 ( .A1(n5515), .A2(n6289), .B1(n4864), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4515) );
  OAI21_X1 U5614 ( .B1(n5176), .B2(n3010), .A(n4515), .ZN(U2856) );
  XNOR2_X1 U5615 ( .A(n4517), .B(n4516), .ZN(n4529) );
  NAND3_X1 U5616 ( .A1(n6260), .A2(n4518), .A3(n4520), .ZN(n4524) );
  INV_X1 U5617 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6599) );
  OAI22_X1 U5618 ( .A1(n6302), .A2(n6599), .B1(n4520), .B2(n4519), .ZN(n4521)
         );
  AOI21_X1 U5619 ( .B1(n6290), .B2(n4522), .A(n4521), .ZN(n4523) );
  OAI211_X1 U5620 ( .C1(n4529), .C2(n6224), .A(n4524), .B(n4523), .ZN(U3017)
         );
  INV_X1 U5621 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4525) );
  OAI22_X1 U5622 ( .A1(n5903), .A2(n4525), .B1(n6302), .B2(n6599), .ZN(n4527)
         );
  NOR2_X1 U5623 ( .A1(n6202), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4526)
         );
  AOI211_X1 U5624 ( .C1(n6099), .C2(n6184), .A(n4527), .B(n4526), .ZN(n4528)
         );
  OAI21_X1 U5625 ( .B1(n4529), .B2(n6178), .A(n4528), .ZN(U2985) );
  AOI21_X1 U5626 ( .B1(n4531), .B2(n4530), .A(n3041), .ZN(n4532) );
  INV_X1 U5627 ( .A(n4532), .ZN(n6303) );
  NAND3_X1 U5628 ( .A1(n4535), .A2(n4534), .A3(n4533), .ZN(n4536) );
  AND2_X1 U5629 ( .A1(n4510), .A2(n4536), .ZN(n6198) );
  INV_X1 U5630 ( .A(n6198), .ZN(n4555) );
  OAI222_X1 U5631 ( .A1(n6303), .A2(n5536), .B1(n5538), .B2(n6805), .C1(n4555), 
        .C2(n3010), .ZN(U2857) );
  AND2_X1 U5632 ( .A1(n6273), .A2(REIP_REG_3__SCAN_IN), .ZN(n6288) );
  NOR2_X1 U5633 ( .A1(n6202), .A2(n5169), .ZN(n4537) );
  AOI211_X1 U5634 ( .C1(n6208), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6288), 
        .B(n4537), .ZN(n4543) );
  OAI21_X1 U5635 ( .B1(n4538), .B2(n4540), .A(n4539), .ZN(n4541) );
  INV_X1 U5636 ( .A(n4541), .ZN(n6291) );
  NAND2_X1 U5637 ( .A1(n6291), .A2(n6206), .ZN(n4542) );
  OAI211_X1 U5638 ( .C1(n6211), .C2(n5176), .A(n4543), .B(n4542), .ZN(U2983)
         );
  NAND2_X1 U5639 ( .A1(n6184), .A2(DATAI_19_), .ZN(n6391) );
  NAND2_X1 U5640 ( .A1(n6184), .A2(DATAI_27_), .ZN(n6442) );
  NAND3_X1 U5641 ( .A1(n4368), .A2(n4973), .A3(n4370), .ZN(n4677) );
  NAND2_X1 U5642 ( .A1(n4578), .A2(n3331), .ZN(n5227) );
  NAND2_X1 U5643 ( .A1(n4374), .A2(n4375), .ZN(n6363) );
  INV_X1 U5644 ( .A(n6363), .ZN(n4640) );
  INV_X1 U5645 ( .A(n4580), .ZN(n4544) );
  AOI21_X1 U5646 ( .B1(n4812), .B2(n4640), .A(n4544), .ZN(n4548) );
  INV_X1 U5647 ( .A(n4548), .ZN(n4545) );
  AOI22_X1 U5648 ( .A1(n4545), .A2(n6367), .B1(n4635), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4579) );
  OAI22_X1 U5649 ( .A1(n5227), .A2(n4580), .B1(n4579), .B2(n5232), .ZN(n4546)
         );
  AOI21_X1 U5650 ( .B1(n6388), .B2(n4660), .A(n4546), .ZN(n4552) );
  OAI21_X1 U5651 ( .B1(n4547), .B2(n6211), .A(n6317), .ZN(n4549) );
  NAND2_X1 U5652 ( .A1(n4549), .A2(n4548), .ZN(n4550) );
  OAI211_X1 U5653 ( .C1(n4635), .C2(n6367), .A(n4550), .B(n4983), .ZN(n4582)
         );
  NAND2_X1 U5654 ( .A1(n4582), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4551)
         );
  OAI211_X1 U5655 ( .C1(n4585), .C2(n6391), .A(n4552), .B(n4551), .ZN(U3143)
         );
  NAND2_X1 U5656 ( .A1(n3263), .A2(n3335), .ZN(n4553) );
  INV_X1 U5657 ( .A(n4553), .ZN(n4554) );
  INV_X1 U5658 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6142) );
  OAI222_X1 U5659 ( .A1(n5886), .A2(n6212), .B1(n5290), .B2(n6151), .C1(n5541), 
        .C2(n6142), .ZN(U2891) );
  INV_X1 U5660 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6136) );
  OAI222_X1 U5661 ( .A1(n4555), .A2(n5886), .B1(n5290), .B2(n6155), .C1(n5541), 
        .C2(n6136), .ZN(U2889) );
  INV_X1 U5662 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6138) );
  OAI222_X1 U5663 ( .A1(n4556), .A2(n5886), .B1(n5290), .B2(n6153), .C1(n5541), 
        .C2(n6138), .ZN(U2890) );
  INV_X1 U5664 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6134) );
  OAI222_X1 U5665 ( .A1(n5176), .A2(n5886), .B1(n5290), .B2(n4502), .C1(n5541), 
        .C2(n6134), .ZN(U2888) );
  NAND2_X1 U5666 ( .A1(n6184), .A2(DATAI_21_), .ZN(n6401) );
  INV_X1 U5667 ( .A(DATAI_29_), .ZN(n4557) );
  NOR2_X1 U5668 ( .A1(n6211), .A2(n4557), .ZN(n6398) );
  NAND2_X1 U5669 ( .A1(n4578), .A2(n3022), .ZN(n5205) );
  INV_X1 U5670 ( .A(DATAI_5_), .ZN(n6160) );
  OAI22_X1 U5671 ( .A1(n5205), .A2(n4580), .B1(n4579), .B2(n5209), .ZN(n4558)
         );
  AOI21_X1 U5672 ( .B1(n6398), .B2(n4660), .A(n4558), .ZN(n4560) );
  NAND2_X1 U5673 ( .A1(n4582), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4559)
         );
  OAI211_X1 U5674 ( .C1(n4585), .C2(n6401), .A(n4560), .B(n4559), .ZN(U3145)
         );
  OAI22_X1 U5675 ( .A1(n5210), .A2(n4580), .B1(n4579), .B2(n5214), .ZN(n4561)
         );
  AOI21_X1 U5676 ( .B1(n6384), .B2(n4660), .A(n4561), .ZN(n4563) );
  NAND2_X1 U5677 ( .A1(n4582), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4562)
         );
  OAI211_X1 U5678 ( .C1(n4585), .C2(n6387), .A(n4563), .B(n4562), .ZN(U3142)
         );
  INV_X1 U5679 ( .A(DATAI_4_), .ZN(n6158) );
  NAND2_X1 U5680 ( .A1(n6184), .A2(DATAI_20_), .ZN(n6395) );
  INV_X1 U5681 ( .A(n6395), .ZN(n6444) );
  NOR2_X2 U5682 ( .A1(n4565), .A2(n4564), .ZN(n6443) );
  INV_X1 U5683 ( .A(n6443), .ZN(n5190) );
  NAND2_X1 U5684 ( .A1(n6184), .A2(DATAI_28_), .ZN(n6448) );
  OAI22_X1 U5685 ( .A1(n5190), .A2(n4580), .B1(n6448), .B2(n4677), .ZN(n4566)
         );
  AOI21_X1 U5686 ( .B1(n6444), .B2(n4737), .A(n4566), .ZN(n4568) );
  NAND2_X1 U5687 ( .A1(n4582), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4567)
         );
  OAI211_X1 U5688 ( .C1(n4579), .C2(n5194), .A(n4568), .B(n4567), .ZN(U3144)
         );
  OAI22_X1 U5689 ( .A1(n5215), .A2(n4580), .B1(n4579), .B2(n5219), .ZN(n4569)
         );
  AOI21_X1 U5690 ( .B1(n6378), .B2(n4660), .A(n4569), .ZN(n4571) );
  NAND2_X1 U5691 ( .A1(n4582), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4570)
         );
  OAI211_X1 U5692 ( .C1(n4585), .C2(n6381), .A(n4571), .B(n4570), .ZN(U3141)
         );
  INV_X1 U5693 ( .A(n6436), .ZN(n6374) );
  OAI22_X1 U5694 ( .A1(n5220), .A2(n4580), .B1(n4579), .B2(n5224), .ZN(n4572)
         );
  AOI21_X1 U5695 ( .B1(n6374), .B2(n4660), .A(n4572), .ZN(n4574) );
  NAND2_X1 U5696 ( .A1(n4582), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4573)
         );
  OAI211_X1 U5697 ( .C1(n4585), .C2(n6377), .A(n4574), .B(n4573), .ZN(U3140)
         );
  NAND2_X1 U5698 ( .A1(n6184), .A2(DATAI_22_), .ZN(n6405) );
  NAND2_X1 U5699 ( .A1(n6184), .A2(DATAI_30_), .ZN(n6459) );
  INV_X1 U5700 ( .A(n6459), .ZN(n6402) );
  NAND2_X1 U5701 ( .A1(n4578), .A2(n3237), .ZN(n5195) );
  INV_X1 U5702 ( .A(DATAI_6_), .ZN(n6162) );
  OAI22_X1 U5703 ( .A1(n5195), .A2(n4580), .B1(n4579), .B2(n5199), .ZN(n4575)
         );
  AOI21_X1 U5704 ( .B1(n6402), .B2(n4660), .A(n4575), .ZN(n4577) );
  NAND2_X1 U5705 ( .A1(n4582), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4576)
         );
  OAI211_X1 U5706 ( .C1(n4585), .C2(n6405), .A(n4577), .B(n4576), .ZN(U3146)
         );
  NAND2_X1 U5707 ( .A1(n6184), .A2(DATAI_23_), .ZN(n6415) );
  NAND2_X1 U5708 ( .A1(n6184), .A2(DATAI_31_), .ZN(n6355) );
  INV_X1 U5709 ( .A(n6355), .ZN(n6411) );
  NAND2_X1 U5710 ( .A1(n4578), .A2(n3335), .ZN(n5200) );
  INV_X1 U5711 ( .A(DATAI_7_), .ZN(n6164) );
  OAI22_X1 U5712 ( .A1(n5200), .A2(n4580), .B1(n4579), .B2(n5204), .ZN(n4581)
         );
  AOI21_X1 U5713 ( .B1(n6411), .B2(n4660), .A(n4581), .ZN(n4584) );
  NAND2_X1 U5714 ( .A1(n4582), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4583)
         );
  OAI211_X1 U5715 ( .C1(n4585), .C2(n6415), .A(n4584), .B(n4583), .ZN(U3147)
         );
  NAND2_X1 U5716 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4587) );
  INV_X1 U5717 ( .A(n4587), .ZN(n4586) );
  MUX2_X1 U5718 ( .A(n4587), .B(n4586), .S(n6598), .Z(n4597) );
  INV_X1 U5719 ( .A(n5412), .ZN(n6462) );
  MUX2_X1 U5720 ( .A(n4588), .B(n6598), .S(n4446), .Z(n4589) );
  NOR2_X1 U5721 ( .A1(n4589), .A2(n4603), .ZN(n4590) );
  NAND2_X1 U5722 ( .A1(n4591), .A2(n4590), .ZN(n4596) );
  INV_X1 U5723 ( .A(n4588), .ZN(n4593) );
  OAI211_X1 U5724 ( .C1(n6598), .C2(n4446), .A(n3294), .B(n4593), .ZN(n6593)
         );
  OR2_X1 U5725 ( .A1(n4594), .A2(n6593), .ZN(n4595) );
  OAI211_X1 U5726 ( .C1(n4597), .C2(n6462), .A(n4596), .B(n4595), .ZN(n4598)
         );
  AOI21_X1 U5727 ( .B1(n3023), .B2(n5789), .A(n4598), .ZN(n6595) );
  MUX2_X1 U5728 ( .A(n3087), .B(n6595), .S(n4608), .Z(n6477) );
  INV_X1 U5729 ( .A(n6477), .ZN(n4602) );
  NAND2_X1 U5730 ( .A1(n4608), .A2(n4599), .ZN(n4600) );
  OAI21_X1 U5731 ( .B1(n4608), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4600), 
        .ZN(n6472) );
  INV_X1 U5732 ( .A(n6472), .ZN(n4601) );
  NAND3_X1 U5733 ( .A1(n4602), .A2(n4601), .A3(n6784), .ZN(n4605) );
  AND2_X1 U5734 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5953), .ZN(n4610) );
  NAND2_X1 U5735 ( .A1(n4603), .A2(n4610), .ZN(n4604) );
  NOR2_X1 U5736 ( .A1(n6488), .A2(n4606), .ZN(n4621) );
  OAI21_X1 U5737 ( .B1(n4608), .B2(n4507), .A(n4607), .ZN(n4609) );
  NAND2_X1 U5738 ( .A1(n4609), .A2(n6784), .ZN(n4612) );
  NAND2_X1 U5739 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4610), .ZN(n4611) );
  NAND2_X1 U5740 ( .A1(n4612), .A2(n4611), .ZN(n6486) );
  NOR3_X1 U5741 ( .A1(n4621), .A2(n6486), .A3(FLUSH_REG_SCAN_IN), .ZN(n4613)
         );
  NOR2_X1 U5742 ( .A1(n5778), .A2(n4614), .ZN(n4615) );
  NAND2_X1 U5743 ( .A1(n4368), .A2(n4615), .ZN(n4763) );
  NAND2_X1 U5744 ( .A1(n4633), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4756) );
  INV_X1 U5745 ( .A(n4756), .ZN(n4616) );
  NOR2_X1 U5746 ( .A1(n4616), .A2(n4847), .ZN(n4784) );
  NAND2_X1 U5747 ( .A1(n4974), .A2(n5781), .ZN(n4969) );
  AOI21_X1 U5748 ( .B1(n4784), .B2(n4969), .A(n6316), .ZN(n4618) );
  AND2_X1 U5749 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6591), .ZN(n5782) );
  OAI22_X1 U5750 ( .A1(n3777), .A2(n6317), .B1(n5171), .B2(n5782), .ZN(n4617)
         );
  OAI21_X1 U5751 ( .B1(n4618), .B2(n4617), .A(n6312), .ZN(n4619) );
  OAI21_X1 U5752 ( .B1(n6312), .B2(n6359), .A(n4619), .ZN(U3462) );
  INV_X1 U5753 ( .A(n4620), .ZN(n6508) );
  NOR3_X1 U5754 ( .A1(n4621), .A2(n6486), .A3(n6508), .ZN(n6497) );
  OAI22_X1 U5755 ( .A1(n4873), .A2(n6316), .B1(n3792), .B2(n5782), .ZN(n4622)
         );
  OAI21_X1 U5756 ( .B1(n6497), .B2(n4622), .A(n6312), .ZN(n4623) );
  OAI21_X1 U5757 ( .B1(n6312), .B2(n6632), .A(n4623), .ZN(U3465) );
  AND2_X1 U5758 ( .A1(n4509), .A2(n4625), .ZN(n4626) );
  NOR2_X1 U5759 ( .A1(n4624), .A2(n4626), .ZN(n6191) );
  INV_X1 U5760 ( .A(n6191), .ZN(n4632) );
  AOI22_X1 U5761 ( .A1(n5383), .A2(DATAI_4_), .B1(n6620), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4627) );
  OAI21_X1 U5762 ( .B1(n4632), .B2(n5886), .A(n4627), .ZN(U2887) );
  NAND2_X1 U5763 ( .A1(n4629), .A2(n4628), .ZN(n4630) );
  AND2_X1 U5764 ( .A1(n4754), .A2(n4630), .ZN(n6281) );
  AOI22_X1 U5765 ( .A1(n5515), .A2(n6281), .B1(n4864), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4631) );
  OAI21_X1 U5766 ( .B1(n4632), .B2(n3010), .A(n4631), .ZN(U2855) );
  AOI21_X1 U5767 ( .B1(n4783), .B2(n4677), .A(n6365), .ZN(n4638) );
  NAND2_X1 U5768 ( .A1(n6367), .A2(n6363), .ZN(n4637) );
  OAI21_X1 U5769 ( .B1(n6360), .B2(n4378), .A(n4634), .ZN(n5183) );
  NOR2_X1 U5770 ( .A1(n6314), .A2(n5183), .ZN(n6371) );
  NAND2_X1 U5771 ( .A1(n6632), .A2(n4635), .ZN(n4678) );
  AOI21_X1 U5772 ( .B1(n4678), .B2(STATE2_REG_3__SCAN_IN), .A(n6359), .ZN(
        n4636) );
  NAND2_X1 U5773 ( .A1(n4681), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4643)
         );
  INV_X1 U5774 ( .A(n6415), .ZN(n6348) );
  NAND2_X1 U5775 ( .A1(n3023), .A2(n6367), .ZN(n5120) );
  INV_X1 U5776 ( .A(n5120), .ZN(n4916) );
  INV_X1 U5777 ( .A(n6361), .ZN(n5113) );
  NOR2_X1 U5778 ( .A1(n5113), .A2(n6359), .ZN(n4639) );
  AOI22_X1 U5779 ( .A1(n4916), .A2(n4640), .B1(n6360), .B2(n4639), .ZN(n4684)
         );
  OAI22_X1 U5780 ( .A1(n5200), .A2(n4678), .B1(n4684), .B2(n5204), .ZN(n4641)
         );
  AOI21_X1 U5781 ( .B1(n6348), .B2(n4660), .A(n4641), .ZN(n4642) );
  OAI211_X1 U5782 ( .C1(n4783), .C2(n6355), .A(n4643), .B(n4642), .ZN(U3139)
         );
  NAND2_X1 U5783 ( .A1(n4681), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4646)
         );
  INV_X1 U5784 ( .A(n6405), .ZN(n6449) );
  OAI22_X1 U5785 ( .A1(n5195), .A2(n4678), .B1(n4684), .B2(n5199), .ZN(n4644)
         );
  AOI21_X1 U5786 ( .B1(n6449), .B2(n4660), .A(n4644), .ZN(n4645) );
  OAI211_X1 U5787 ( .C1(n4783), .C2(n6459), .A(n4646), .B(n4645), .ZN(U3138)
         );
  NAND2_X1 U5788 ( .A1(n4681), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4649)
         );
  INV_X1 U5789 ( .A(n6381), .ZN(n6416) );
  OAI22_X1 U5790 ( .A1(n5215), .A2(n4678), .B1(n4684), .B2(n5219), .ZN(n4647)
         );
  AOI21_X1 U5791 ( .B1(n6416), .B2(n4660), .A(n4647), .ZN(n4648) );
  OAI211_X1 U5792 ( .C1(n4783), .C2(n6421), .A(n4649), .B(n4648), .ZN(U3133)
         );
  NAND2_X1 U5793 ( .A1(n4681), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4652)
         );
  INV_X1 U5794 ( .A(n6377), .ZN(n6431) );
  OAI22_X1 U5795 ( .A1(n5220), .A2(n4678), .B1(n4684), .B2(n5224), .ZN(n4650)
         );
  AOI21_X1 U5796 ( .B1(n6431), .B2(n4660), .A(n4650), .ZN(n4651) );
  OAI211_X1 U5797 ( .C1(n4783), .C2(n6436), .A(n4652), .B(n4651), .ZN(U3132)
         );
  NAND2_X1 U5798 ( .A1(n4681), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4655)
         );
  INV_X1 U5799 ( .A(n6391), .ZN(n6437) );
  OAI22_X1 U5800 ( .A1(n5227), .A2(n4678), .B1(n4684), .B2(n5232), .ZN(n4653)
         );
  AOI21_X1 U5801 ( .B1(n6437), .B2(n4660), .A(n4653), .ZN(n4654) );
  OAI211_X1 U5802 ( .C1(n4783), .C2(n6442), .A(n4655), .B(n4654), .ZN(U3135)
         );
  INV_X1 U5803 ( .A(n6398), .ZN(n5156) );
  NAND2_X1 U5804 ( .A1(n4681), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4658)
         );
  INV_X1 U5805 ( .A(n6401), .ZN(n5159) );
  OAI22_X1 U5806 ( .A1(n5205), .A2(n4678), .B1(n4684), .B2(n5209), .ZN(n4656)
         );
  AOI21_X1 U5807 ( .B1(n5159), .B2(n4660), .A(n4656), .ZN(n4657) );
  OAI211_X1 U5808 ( .C1(n4783), .C2(n5156), .A(n4658), .B(n4657), .ZN(U3137)
         );
  INV_X1 U5809 ( .A(n6384), .ZN(n5138) );
  NAND2_X1 U5810 ( .A1(n4681), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4662)
         );
  INV_X1 U5811 ( .A(n6387), .ZN(n5140) );
  OAI22_X1 U5812 ( .A1(n5210), .A2(n4678), .B1(n4684), .B2(n5214), .ZN(n4659)
         );
  AOI21_X1 U5813 ( .B1(n5140), .B2(n4660), .A(n4659), .ZN(n4661) );
  OAI211_X1 U5814 ( .C1(n4783), .C2(n5138), .A(n4662), .B(n4661), .ZN(U3134)
         );
  NAND3_X1 U5815 ( .A1(n5171), .A2(n5111), .A3(n4841), .ZN(n4664) );
  INV_X1 U5816 ( .A(n4671), .ZN(n4663) );
  NOR2_X1 U5817 ( .A1(n6632), .A2(n4663), .ZN(n4744) );
  INV_X1 U5818 ( .A(n4744), .ZN(n4705) );
  NAND2_X1 U5819 ( .A1(n4664), .A2(n4705), .ZN(n4667) );
  NAND2_X1 U5820 ( .A1(n4669), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U5821 ( .A1(n4671), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4665) );
  INV_X1 U5822 ( .A(n4667), .ZN(n4668) );
  AOI21_X1 U5823 ( .B1(n4669), .B2(n4668), .A(n4843), .ZN(n4670) );
  NAND2_X1 U5824 ( .A1(n4751), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4676) );
  OR2_X1 U5825 ( .A1(n4672), .A2(n4873), .ZN(n4743) );
  OAI22_X1 U5826 ( .A1(n4743), .A2(n6401), .B1(n5205), .B2(n4705), .ZN(n4674)
         );
  NOR2_X1 U5827 ( .A1(n4745), .A2(n5156), .ZN(n4673) );
  NOR2_X1 U5828 ( .A1(n4674), .A2(n4673), .ZN(n4675) );
  OAI211_X1 U5829 ( .C1(n4749), .C2(n5209), .A(n4676), .B(n4675), .ZN(U3033)
         );
  INV_X1 U5830 ( .A(n4783), .ZN(n4680) );
  OAI22_X1 U5831 ( .A1(n5190), .A2(n4678), .B1(n6395), .B2(n4677), .ZN(n4679)
         );
  AOI21_X1 U5832 ( .B1(n6392), .B2(n4680), .A(n4679), .ZN(n4683) );
  NAND2_X1 U5833 ( .A1(n4681), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4682)
         );
  OAI211_X1 U5834 ( .C1(n4684), .C2(n5194), .A(n4683), .B(n4682), .ZN(U3136)
         );
  NAND2_X1 U5835 ( .A1(n4751), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4688) );
  OAI22_X1 U5836 ( .A1(n4743), .A2(n6381), .B1(n5215), .B2(n4705), .ZN(n4686)
         );
  NOR2_X1 U5837 ( .A1(n4745), .A2(n6421), .ZN(n4685) );
  NOR2_X1 U5838 ( .A1(n4686), .A2(n4685), .ZN(n4687) );
  OAI211_X1 U5839 ( .C1(n4749), .C2(n5219), .A(n4688), .B(n4687), .ZN(U3029)
         );
  NAND2_X1 U5840 ( .A1(n4751), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4692) );
  OAI22_X1 U5841 ( .A1(n4743), .A2(n6377), .B1(n5220), .B2(n4705), .ZN(n4690)
         );
  NOR2_X1 U5842 ( .A1(n4745), .A2(n6436), .ZN(n4689) );
  NOR2_X1 U5843 ( .A1(n4690), .A2(n4689), .ZN(n4691) );
  OAI211_X1 U5844 ( .C1(n4749), .C2(n5224), .A(n4692), .B(n4691), .ZN(U3028)
         );
  NAND2_X1 U5845 ( .A1(n4751), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4696) );
  OAI22_X1 U5846 ( .A1(n4743), .A2(n6415), .B1(n5200), .B2(n4705), .ZN(n4694)
         );
  NOR2_X1 U5847 ( .A1(n4745), .A2(n6355), .ZN(n4693) );
  NOR2_X1 U5848 ( .A1(n4694), .A2(n4693), .ZN(n4695) );
  OAI211_X1 U5849 ( .C1(n4749), .C2(n5204), .A(n4696), .B(n4695), .ZN(U3035)
         );
  NAND2_X1 U5850 ( .A1(n4751), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4700) );
  OAI22_X1 U5851 ( .A1(n4743), .A2(n6391), .B1(n5227), .B2(n4705), .ZN(n4698)
         );
  NOR2_X1 U5852 ( .A1(n4745), .A2(n6442), .ZN(n4697) );
  NOR2_X1 U5853 ( .A1(n4698), .A2(n4697), .ZN(n4699) );
  OAI211_X1 U5854 ( .C1(n4749), .C2(n5232), .A(n4700), .B(n4699), .ZN(U3031)
         );
  NAND2_X1 U5855 ( .A1(n4751), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4704) );
  OAI22_X1 U5856 ( .A1(n4743), .A2(n6387), .B1(n5210), .B2(n4705), .ZN(n4702)
         );
  NOR2_X1 U5857 ( .A1(n4745), .A2(n5138), .ZN(n4701) );
  NOR2_X1 U5858 ( .A1(n4702), .A2(n4701), .ZN(n4703) );
  OAI211_X1 U5859 ( .C1(n4749), .C2(n5214), .A(n4704), .B(n4703), .ZN(U3030)
         );
  NAND2_X1 U5860 ( .A1(n4751), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4709) );
  OAI22_X1 U5861 ( .A1(n4743), .A2(n6405), .B1(n5195), .B2(n4705), .ZN(n4707)
         );
  NOR2_X1 U5862 ( .A1(n4745), .A2(n6459), .ZN(n4706) );
  NOR2_X1 U5863 ( .A1(n4707), .A2(n4706), .ZN(n4708) );
  OAI211_X1 U5864 ( .C1(n4749), .C2(n5199), .A(n4709), .B(n4708), .ZN(U3034)
         );
  OAI21_X1 U5865 ( .B1(n4624), .B2(n4711), .A(n4710), .ZN(n5043) );
  INV_X1 U5866 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6130) );
  OAI222_X1 U5867 ( .A1(n5043), .A2(n5886), .B1(n5290), .B2(n6160), .C1(n5541), 
        .C2(n6130), .ZN(U2886) );
  INV_X1 U5868 ( .A(n4712), .ZN(n4741) );
  OAI22_X1 U5869 ( .A1(n5227), .A2(n4735), .B1(n4734), .B2(n5232), .ZN(n4713)
         );
  INV_X1 U5870 ( .A(n4713), .ZN(n4715) );
  NAND2_X1 U5871 ( .A1(n4737), .A2(n6388), .ZN(n4714) );
  OAI211_X1 U5872 ( .C1(n4745), .C2(n6391), .A(n4715), .B(n4714), .ZN(n4716)
         );
  AOI21_X1 U5873 ( .B1(n4741), .B2(INSTQUEUE_REG_0__3__SCAN_IN), .A(n4716), 
        .ZN(n4717) );
  INV_X1 U5874 ( .A(n4717), .ZN(U3023) );
  OAI22_X1 U5875 ( .A1(n5205), .A2(n4735), .B1(n4734), .B2(n5209), .ZN(n4718)
         );
  INV_X1 U5876 ( .A(n4718), .ZN(n4720) );
  NAND2_X1 U5877 ( .A1(n4737), .A2(n6398), .ZN(n4719) );
  OAI211_X1 U5878 ( .C1(n4745), .C2(n6401), .A(n4720), .B(n4719), .ZN(n4721)
         );
  AOI21_X1 U5879 ( .B1(n4741), .B2(INSTQUEUE_REG_0__5__SCAN_IN), .A(n4721), 
        .ZN(n4722) );
  INV_X1 U5880 ( .A(n4722), .ZN(U3025) );
  INV_X1 U5881 ( .A(n4734), .ZN(n4723) );
  NAND2_X1 U5882 ( .A1(n6445), .A2(n4723), .ZN(n4726) );
  INV_X1 U5883 ( .A(n4735), .ZN(n4724) );
  AOI22_X1 U5884 ( .A1(n6443), .A2(n4724), .B1(n6392), .B2(n4737), .ZN(n4725)
         );
  OAI211_X1 U5885 ( .C1(n4745), .C2(n6395), .A(n4726), .B(n4725), .ZN(n4727)
         );
  AOI21_X1 U5886 ( .B1(n4741), .B2(INSTQUEUE_REG_0__4__SCAN_IN), .A(n4727), 
        .ZN(n4728) );
  INV_X1 U5887 ( .A(n4728), .ZN(U3024) );
  OAI22_X1 U5888 ( .A1(n5200), .A2(n4735), .B1(n4734), .B2(n5204), .ZN(n4729)
         );
  INV_X1 U5889 ( .A(n4729), .ZN(n4731) );
  NAND2_X1 U5890 ( .A1(n4737), .A2(n6411), .ZN(n4730) );
  OAI211_X1 U5891 ( .C1(n4745), .C2(n6415), .A(n4731), .B(n4730), .ZN(n4732)
         );
  AOI21_X1 U5892 ( .B1(n4741), .B2(INSTQUEUE_REG_0__7__SCAN_IN), .A(n4732), 
        .ZN(n4733) );
  INV_X1 U5893 ( .A(n4733), .ZN(U3027) );
  OAI22_X1 U5894 ( .A1(n5195), .A2(n4735), .B1(n4734), .B2(n5199), .ZN(n4736)
         );
  INV_X1 U5895 ( .A(n4736), .ZN(n4739) );
  NAND2_X1 U5896 ( .A1(n4737), .A2(n6402), .ZN(n4738) );
  OAI211_X1 U5897 ( .C1(n4745), .C2(n6405), .A(n4739), .B(n4738), .ZN(n4740)
         );
  AOI21_X1 U5898 ( .B1(n4741), .B2(INSTQUEUE_REG_0__6__SCAN_IN), .A(n4740), 
        .ZN(n4742) );
  INV_X1 U5899 ( .A(n4742), .ZN(U3026) );
  AOI22_X1 U5900 ( .A1(n6339), .A2(n6444), .B1(n6443), .B2(n4744), .ZN(n4748)
         );
  INV_X1 U5901 ( .A(n4745), .ZN(n4746) );
  NAND2_X1 U5902 ( .A1(n4746), .A2(n6392), .ZN(n4747) );
  OAI211_X1 U5903 ( .C1(n5194), .C2(n4749), .A(n4748), .B(n4747), .ZN(n4750)
         );
  AOI21_X1 U5904 ( .B1(n4751), .B2(INSTQUEUE_REG_1__4__SCAN_IN), .A(n4750), 
        .ZN(n4752) );
  INV_X1 U5905 ( .A(n4752), .ZN(U3032) );
  AOI21_X1 U5906 ( .B1(n4755), .B2(n4754), .A(n4753), .ZN(n6271) );
  INV_X1 U5907 ( .A(n6271), .ZN(n5039) );
  OAI222_X1 U5908 ( .A1(n5039), .A2(n5536), .B1(n5538), .B2(n3655), .C1(n3010), 
        .C2(n5043), .ZN(U2854) );
  NAND2_X1 U5909 ( .A1(n6467), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4760) );
  INV_X1 U5910 ( .A(n4760), .ZN(n4868) );
  NAND2_X1 U5911 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4868), .ZN(n4908) );
  NOR2_X1 U5912 ( .A1(n6632), .A2(n4908), .ZN(n4780) );
  AOI21_X1 U5913 ( .B1(n4812), .B2(n5068), .A(n4780), .ZN(n4762) );
  INV_X1 U5914 ( .A(n4762), .ZN(n4758) );
  NAND2_X1 U5915 ( .A1(n6367), .A2(n4756), .ZN(n4761) );
  AOI21_X1 U5916 ( .B1(n6316), .B2(n4908), .A(n4843), .ZN(n4757) );
  OAI21_X1 U5917 ( .B1(n4758), .B2(n4761), .A(n4757), .ZN(n4779) );
  NAND2_X1 U5918 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4759) );
  OAI22_X1 U5919 ( .A1(n4762), .A2(n4761), .B1(n4760), .B2(n4759), .ZN(n4778)
         );
  AOI22_X1 U5920 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4779), .B1(n6439), 
        .B2(n4778), .ZN(n4765) );
  NOR2_X2 U5921 ( .A1(n4763), .A2(n4872), .ZN(n4944) );
  AOI22_X1 U5922 ( .A1(n6438), .A2(n4780), .B1(n6388), .B2(n4944), .ZN(n4764)
         );
  OAI211_X1 U5923 ( .C1(n6391), .C2(n4783), .A(n4765), .B(n4764), .ZN(U3127)
         );
  AOI22_X1 U5924 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4779), .B1(n6382), 
        .B2(n4778), .ZN(n4767) );
  AOI22_X1 U5925 ( .A1(n6383), .A2(n4780), .B1(n6384), .B2(n4944), .ZN(n4766)
         );
  OAI211_X1 U5926 ( .C1(n6387), .C2(n4783), .A(n4767), .B(n4766), .ZN(U3126)
         );
  AOI22_X1 U5927 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4779), .B1(n6418), 
        .B2(n4778), .ZN(n4769) );
  AOI22_X1 U5928 ( .A1(n6417), .A2(n4780), .B1(n6378), .B2(n4944), .ZN(n4768)
         );
  OAI211_X1 U5929 ( .C1(n6381), .C2(n4783), .A(n4769), .B(n4768), .ZN(U3125)
         );
  AOI22_X1 U5930 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4779), .B1(n6433), 
        .B2(n4778), .ZN(n4771) );
  AOI22_X1 U5931 ( .A1(n6432), .A2(n4780), .B1(n6374), .B2(n4944), .ZN(n4770)
         );
  OAI211_X1 U5932 ( .C1(n6377), .C2(n4783), .A(n4771), .B(n4770), .ZN(U3124)
         );
  AOI22_X1 U5933 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4779), .B1(n6454), 
        .B2(n4778), .ZN(n4773) );
  AOI22_X1 U5934 ( .A1(n6452), .A2(n4780), .B1(n6402), .B2(n4944), .ZN(n4772)
         );
  OAI211_X1 U5935 ( .C1(n6405), .C2(n4783), .A(n4773), .B(n4772), .ZN(U3130)
         );
  AOI22_X1 U5936 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4779), .B1(n6396), 
        .B2(n4778), .ZN(n4775) );
  AOI22_X1 U5937 ( .A1(n6397), .A2(n4780), .B1(n6398), .B2(n4944), .ZN(n4774)
         );
  OAI211_X1 U5938 ( .C1(n6401), .C2(n4783), .A(n4775), .B(n4774), .ZN(U3129)
         );
  AOI22_X1 U5939 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4779), .B1(n6407), 
        .B2(n4778), .ZN(n4777) );
  AOI22_X1 U5940 ( .A1(n6409), .A2(n4780), .B1(n6411), .B2(n4944), .ZN(n4776)
         );
  OAI211_X1 U5941 ( .C1(n6415), .C2(n4783), .A(n4777), .B(n4776), .ZN(U3131)
         );
  AOI22_X1 U5942 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4779), .B1(n6445), 
        .B2(n4778), .ZN(n4782) );
  AOI22_X1 U5943 ( .A1(n6443), .A2(n4780), .B1(n6392), .B2(n4944), .ZN(n4781)
         );
  OAI211_X1 U5944 ( .C1(n6395), .C2(n4783), .A(n4782), .B(n4781), .ZN(U3128)
         );
  NAND3_X1 U5945 ( .A1(n4784), .A2(n5781), .A3(n3409), .ZN(n4785) );
  NAND2_X1 U5946 ( .A1(n4785), .A2(n6367), .ZN(n4791) );
  NOR2_X1 U5947 ( .A1(n4374), .A2(n6090), .ZN(n4839) );
  NAND2_X1 U5948 ( .A1(n5171), .A2(n4839), .ZN(n6319) );
  OR2_X1 U5949 ( .A1(n6319), .A2(n3792), .ZN(n4787) );
  INV_X1 U5950 ( .A(n4840), .ZN(n4786) );
  NAND2_X1 U5951 ( .A1(n4786), .A2(n6359), .ZN(n6343) );
  NAND3_X1 U5952 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6359), .A3(n6474), .ZN(n6313) );
  OAI22_X1 U5953 ( .A1(n4791), .A2(n4788), .B1(n6313), .B2(n4378), .ZN(n6351)
         );
  INV_X1 U5954 ( .A(n6351), .ZN(n4809) );
  INV_X1 U5955 ( .A(n4788), .ZN(n4790) );
  AOI21_X1 U5956 ( .B1(n6316), .B2(n6313), .A(n4843), .ZN(n4789) );
  OAI21_X1 U5957 ( .B1(n4791), .B2(n4790), .A(n4789), .ZN(n6352) );
  NOR2_X1 U5958 ( .A1(n6356), .A2(n6459), .ZN(n4794) );
  INV_X1 U5959 ( .A(n6349), .ZN(n4805) );
  OAI22_X1 U5960 ( .A1(n4805), .A2(n6405), .B1(n5195), .B2(n6343), .ZN(n4793)
         );
  AOI211_X1 U5961 ( .C1(n6352), .C2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n4794), 
        .B(n4793), .ZN(n4795) );
  OAI21_X1 U5962 ( .B1(n4809), .B2(n5199), .A(n4795), .ZN(U3050) );
  NOR2_X1 U5963 ( .A1(n6356), .A2(n5156), .ZN(n4797) );
  OAI22_X1 U5964 ( .A1(n4805), .A2(n6401), .B1(n5205), .B2(n6343), .ZN(n4796)
         );
  AOI211_X1 U5965 ( .C1(n6352), .C2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4797), 
        .B(n4796), .ZN(n4798) );
  OAI21_X1 U5966 ( .B1(n4809), .B2(n5209), .A(n4798), .ZN(U3049) );
  NOR2_X1 U5967 ( .A1(n6356), .A2(n6436), .ZN(n4800) );
  OAI22_X1 U5968 ( .A1(n4805), .A2(n6377), .B1(n5220), .B2(n6343), .ZN(n4799)
         );
  AOI211_X1 U5969 ( .C1(n6352), .C2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4800), 
        .B(n4799), .ZN(n4801) );
  OAI21_X1 U5970 ( .B1(n4809), .B2(n5224), .A(n4801), .ZN(U3044) );
  NOR2_X1 U5971 ( .A1(n6356), .A2(n5138), .ZN(n4803) );
  OAI22_X1 U5972 ( .A1(n4805), .A2(n6387), .B1(n5210), .B2(n6343), .ZN(n4802)
         );
  AOI211_X1 U5973 ( .C1(n6352), .C2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n4803), 
        .B(n4802), .ZN(n4804) );
  OAI21_X1 U5974 ( .B1(n4809), .B2(n5214), .A(n4804), .ZN(U3046) );
  NOR2_X1 U5975 ( .A1(n6356), .A2(n6421), .ZN(n4807) );
  OAI22_X1 U5976 ( .A1(n4805), .A2(n6381), .B1(n5215), .B2(n6343), .ZN(n4806)
         );
  AOI211_X1 U5977 ( .C1(n6352), .C2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4807), 
        .B(n4806), .ZN(n4808) );
  OAI21_X1 U5978 ( .B1(n4809), .B2(n5219), .A(n4808), .ZN(U3045) );
  INV_X1 U5979 ( .A(n4817), .ZN(n4811) );
  OAI21_X1 U5980 ( .B1(n4817), .B2(n6365), .A(n6367), .ZN(n4816) );
  NAND3_X1 U5981 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6474), .A3(n6467), .ZN(n5112) );
  NOR2_X1 U5982 ( .A1(n6632), .A2(n5112), .ZN(n4834) );
  AOI21_X1 U5983 ( .B1(n4812), .B2(n5111), .A(n4834), .ZN(n4815) );
  INV_X1 U5984 ( .A(n4815), .ZN(n4814) );
  AOI21_X1 U5985 ( .B1(n6316), .B2(n5112), .A(n4843), .ZN(n4813) );
  OAI21_X1 U5986 ( .B1(n4816), .B2(n4814), .A(n4813), .ZN(n4833) );
  OAI22_X1 U5987 ( .A1(n4816), .A2(n4815), .B1(n4378), .B2(n5112), .ZN(n4832)
         );
  AOI22_X1 U5988 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4833), .B1(n6407), 
        .B2(n4832), .ZN(n4819) );
  AOI22_X1 U5989 ( .A1(n5158), .A2(n6411), .B1(n6409), .B2(n4834), .ZN(n4818)
         );
  OAI211_X1 U5990 ( .C1(n6415), .C2(n5177), .A(n4819), .B(n4818), .ZN(U3099)
         );
  AOI22_X1 U5991 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4833), .B1(n6454), 
        .B2(n4832), .ZN(n4821) );
  AOI22_X1 U5992 ( .A1(n5158), .A2(n6402), .B1(n6452), .B2(n4834), .ZN(n4820)
         );
  OAI211_X1 U5993 ( .C1(n6405), .C2(n5177), .A(n4821), .B(n4820), .ZN(U3098)
         );
  AOI22_X1 U5994 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4833), .B1(n6396), 
        .B2(n4832), .ZN(n4823) );
  AOI22_X1 U5995 ( .A1(n5158), .A2(n6398), .B1(n6397), .B2(n4834), .ZN(n4822)
         );
  OAI211_X1 U5996 ( .C1(n6401), .C2(n5177), .A(n4823), .B(n4822), .ZN(U3097)
         );
  AOI22_X1 U5997 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4833), .B1(n6445), 
        .B2(n4832), .ZN(n4825) );
  AOI22_X1 U5998 ( .A1(n5158), .A2(n6392), .B1(n6443), .B2(n4834), .ZN(n4824)
         );
  OAI211_X1 U5999 ( .C1(n6395), .C2(n5177), .A(n4825), .B(n4824), .ZN(U3096)
         );
  AOI22_X1 U6000 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4833), .B1(n6439), 
        .B2(n4832), .ZN(n4827) );
  AOI22_X1 U6001 ( .A1(n5158), .A2(n6388), .B1(n6438), .B2(n4834), .ZN(n4826)
         );
  OAI211_X1 U6002 ( .C1(n6391), .C2(n5177), .A(n4827), .B(n4826), .ZN(U3095)
         );
  AOI22_X1 U6003 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4833), .B1(n6382), 
        .B2(n4832), .ZN(n4829) );
  AOI22_X1 U6004 ( .A1(n5158), .A2(n6384), .B1(n6383), .B2(n4834), .ZN(n4828)
         );
  OAI211_X1 U6005 ( .C1(n6387), .C2(n5177), .A(n4829), .B(n4828), .ZN(U3094)
         );
  AOI22_X1 U6006 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4833), .B1(n6418), 
        .B2(n4832), .ZN(n4831) );
  AOI22_X1 U6007 ( .A1(n5158), .A2(n6378), .B1(n6417), .B2(n4834), .ZN(n4830)
         );
  OAI211_X1 U6008 ( .C1(n6381), .C2(n5177), .A(n4831), .B(n4830), .ZN(U3093)
         );
  AOI22_X1 U6009 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4833), .B1(n6433), 
        .B2(n4832), .ZN(n4836) );
  AOI22_X1 U6010 ( .A1(n5158), .A2(n6374), .B1(n6432), .B2(n4834), .ZN(n4835)
         );
  OAI211_X1 U6011 ( .C1(n6377), .C2(n5177), .A(n4836), .B(n4835), .ZN(U3092)
         );
  INV_X1 U6012 ( .A(n4847), .ZN(n4838) );
  INV_X1 U6013 ( .A(n5781), .ZN(n4837) );
  OAI21_X1 U6014 ( .B1(n4838), .B2(n4837), .A(n6367), .ZN(n4846) );
  NOR2_X1 U6015 ( .A1(n4840), .A2(n6359), .ZN(n6451) );
  AOI21_X1 U6016 ( .B1(n5187), .B2(n4841), .A(n6451), .ZN(n4842) );
  NAND3_X1 U6017 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6474), .ZN(n5184) );
  OAI22_X1 U6018 ( .A1(n4846), .A2(n4842), .B1(n5184), .B2(n4378), .ZN(n6453)
         );
  INV_X1 U6019 ( .A(n6453), .ZN(n4860) );
  INV_X1 U6020 ( .A(n4842), .ZN(n4845) );
  AOI21_X1 U6021 ( .B1(n6316), .B2(n5184), .A(n4843), .ZN(n4844) );
  OAI21_X1 U6022 ( .B1(n4846), .B2(n4845), .A(n4844), .ZN(n6455) );
  AOI22_X1 U6023 ( .A1(n6397), .A2(n6451), .B1(n6450), .B2(n5159), .ZN(n4848)
         );
  OAI21_X1 U6024 ( .B1(n5156), .B2(n6458), .A(n4848), .ZN(n4849) );
  AOI21_X1 U6025 ( .B1(n6455), .B2(INSTQUEUE_REG_11__5__SCAN_IN), .A(n4849), 
        .ZN(n4850) );
  OAI21_X1 U6026 ( .B1(n4860), .B2(n5209), .A(n4850), .ZN(U3113) );
  AOI22_X1 U6027 ( .A1(n6383), .A2(n6451), .B1(n6450), .B2(n5140), .ZN(n4851)
         );
  OAI21_X1 U6028 ( .B1(n5138), .B2(n6458), .A(n4851), .ZN(n4852) );
  AOI21_X1 U6029 ( .B1(n6455), .B2(INSTQUEUE_REG_11__2__SCAN_IN), .A(n4852), 
        .ZN(n4853) );
  OAI21_X1 U6030 ( .B1(n4860), .B2(n5214), .A(n4853), .ZN(U3110) );
  AOI22_X1 U6031 ( .A1(n6417), .A2(n6451), .B1(n6450), .B2(n6416), .ZN(n4854)
         );
  OAI21_X1 U6032 ( .B1(n6421), .B2(n6458), .A(n4854), .ZN(n4855) );
  AOI21_X1 U6033 ( .B1(n6455), .B2(INSTQUEUE_REG_11__1__SCAN_IN), .A(n4855), 
        .ZN(n4856) );
  OAI21_X1 U6034 ( .B1(n4860), .B2(n5219), .A(n4856), .ZN(U3109) );
  AOI22_X1 U6035 ( .A1(n6409), .A2(n6451), .B1(n6450), .B2(n6348), .ZN(n4857)
         );
  OAI21_X1 U6036 ( .B1(n6355), .B2(n6458), .A(n4857), .ZN(n4858) );
  AOI21_X1 U6037 ( .B1(n6455), .B2(INSTQUEUE_REG_11__7__SCAN_IN), .A(n4858), 
        .ZN(n4859) );
  OAI21_X1 U6038 ( .B1(n4860), .B2(n5204), .A(n4859), .ZN(U3115) );
  NAND2_X1 U6039 ( .A1(n4710), .A2(n4862), .ZN(n4863) );
  AND2_X1 U6040 ( .A1(n4861), .A2(n4863), .ZN(n6183) );
  INV_X1 U6041 ( .A(n6183), .ZN(n4882) );
  XNOR2_X1 U6042 ( .A(n4753), .B(n4950), .ZN(n6261) );
  AOI22_X1 U6043 ( .A1(n5515), .A2(n6261), .B1(n4864), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4865) );
  OAI21_X1 U6044 ( .B1(n4882), .B2(n3010), .A(n4865), .ZN(U2853) );
  NOR2_X1 U6045 ( .A1(n5778), .A2(n6365), .ZN(n4866) );
  AOI21_X1 U6046 ( .B1(n4974), .B2(n4866), .A(n6316), .ZN(n4877) );
  NAND2_X1 U6047 ( .A1(n5068), .A2(n4867), .ZN(n5063) );
  OR2_X1 U6048 ( .A1(n5063), .A2(n3792), .ZN(n4870) );
  NAND2_X1 U6049 ( .A1(n4868), .A2(n6359), .ZN(n5062) );
  NOR2_X1 U6050 ( .A1(n6632), .A2(n5062), .ZN(n4902) );
  INV_X1 U6051 ( .A(n4902), .ZN(n4869) );
  NAND2_X1 U6052 ( .A1(n4870), .A2(n4869), .ZN(n4875) );
  INV_X1 U6053 ( .A(n5062), .ZN(n4871) );
  AOI22_X1 U6054 ( .A1(n4877), .A2(n4875), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4871), .ZN(n4906) );
  NAND2_X1 U6055 ( .A1(n4874), .A2(n4872), .ZN(n6366) );
  INV_X1 U6056 ( .A(n4875), .ZN(n4876) );
  AOI22_X1 U6057 ( .A1(n4877), .A2(n4876), .B1(n5062), .B2(n6316), .ZN(n4878)
         );
  NAND2_X1 U6058 ( .A1(n4983), .A2(n4878), .ZN(n4901) );
  AOI22_X1 U6059 ( .A1(n6417), .A2(n4902), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n4901), .ZN(n4879) );
  OAI21_X1 U6060 ( .B1(n5100), .B2(n6421), .A(n4879), .ZN(n4880) );
  AOI21_X1 U6061 ( .B1(n6416), .B2(n6410), .A(n4880), .ZN(n4881) );
  OAI21_X1 U6062 ( .B1(n4906), .B2(n5219), .A(n4881), .ZN(U3061) );
  OAI222_X1 U6063 ( .A1(n4882), .A2(n5886), .B1(n5290), .B2(n6162), .C1(n5541), 
        .C2(n3832), .ZN(U2885) );
  AOI22_X1 U6064 ( .A1(n6443), .A2(n4902), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n4901), .ZN(n4883) );
  OAI21_X1 U6065 ( .B1(n5100), .B2(n6448), .A(n4883), .ZN(n4884) );
  AOI21_X1 U6066 ( .B1(n6444), .B2(n6410), .A(n4884), .ZN(n4885) );
  OAI21_X1 U6067 ( .B1(n4906), .B2(n5194), .A(n4885), .ZN(U3064) );
  AOI22_X1 U6068 ( .A1(n6397), .A2(n4902), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n4901), .ZN(n4886) );
  OAI21_X1 U6069 ( .B1(n5100), .B2(n5156), .A(n4886), .ZN(n4887) );
  AOI21_X1 U6070 ( .B1(n5159), .B2(n6410), .A(n4887), .ZN(n4888) );
  OAI21_X1 U6071 ( .B1(n4906), .B2(n5209), .A(n4888), .ZN(U3065) );
  AOI22_X1 U6072 ( .A1(n6383), .A2(n4902), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n4901), .ZN(n4889) );
  OAI21_X1 U6073 ( .B1(n5100), .B2(n5138), .A(n4889), .ZN(n4890) );
  AOI21_X1 U6074 ( .B1(n5140), .B2(n6410), .A(n4890), .ZN(n4891) );
  OAI21_X1 U6075 ( .B1(n4906), .B2(n5214), .A(n4891), .ZN(U3062) );
  AOI22_X1 U6076 ( .A1(n6452), .A2(n4902), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n4901), .ZN(n4892) );
  OAI21_X1 U6077 ( .B1(n5100), .B2(n6459), .A(n4892), .ZN(n4893) );
  AOI21_X1 U6078 ( .B1(n6449), .B2(n6410), .A(n4893), .ZN(n4894) );
  OAI21_X1 U6079 ( .B1(n4906), .B2(n5199), .A(n4894), .ZN(U3066) );
  AOI22_X1 U6080 ( .A1(n6409), .A2(n4902), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n4901), .ZN(n4895) );
  OAI21_X1 U6081 ( .B1(n5100), .B2(n6355), .A(n4895), .ZN(n4896) );
  AOI21_X1 U6082 ( .B1(n6348), .B2(n6410), .A(n4896), .ZN(n4897) );
  OAI21_X1 U6083 ( .B1(n4906), .B2(n5204), .A(n4897), .ZN(U3067) );
  AOI22_X1 U6084 ( .A1(n6438), .A2(n4902), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n4901), .ZN(n4898) );
  OAI21_X1 U6085 ( .B1(n5100), .B2(n6442), .A(n4898), .ZN(n4899) );
  AOI21_X1 U6086 ( .B1(n6437), .B2(n6410), .A(n4899), .ZN(n4900) );
  OAI21_X1 U6087 ( .B1(n4906), .B2(n5232), .A(n4900), .ZN(U3063) );
  AOI22_X1 U6088 ( .A1(n6432), .A2(n4902), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n4901), .ZN(n4903) );
  OAI21_X1 U6089 ( .B1(n5100), .B2(n6436), .A(n4903), .ZN(n4904) );
  AOI21_X1 U6090 ( .B1(n6431), .B2(n6410), .A(n4904), .ZN(n4905) );
  OAI21_X1 U6091 ( .B1(n4906), .B2(n5224), .A(n4905), .ZN(U3060) );
  INV_X1 U6092 ( .A(n4944), .ZN(n4929) );
  AOI21_X1 U6093 ( .B1(n4947), .B2(n4929), .A(n6365), .ZN(n4907) );
  AOI211_X1 U6094 ( .C1(n5068), .C2(n4970), .A(n6316), .B(n4907), .ZN(n4913)
         );
  NOR2_X1 U6095 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4908), .ZN(n4914)
         );
  INV_X1 U6096 ( .A(n6314), .ZN(n5180) );
  OAI21_X1 U6097 ( .B1(n6591), .B2(n4914), .A(n5180), .ZN(n4912) );
  OR2_X1 U6098 ( .A1(n6360), .A2(n4909), .ZN(n5118) );
  AOI21_X1 U6099 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5118), .A(n4910), .ZN(
        n4911) );
  INV_X1 U6100 ( .A(n4911), .ZN(n5114) );
  NAND2_X1 U6101 ( .A1(n4940), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4919)
         );
  INV_X1 U6102 ( .A(n4914), .ZN(n4942) );
  INV_X1 U6103 ( .A(n5118), .ZN(n4915) );
  AOI22_X1 U6104 ( .A1(n4916), .A2(n5068), .B1(n6361), .B2(n4915), .ZN(n4941)
         );
  OAI22_X1 U6105 ( .A1(n5195), .A2(n4942), .B1(n4941), .B2(n5199), .ZN(n4917)
         );
  AOI21_X1 U6106 ( .B1(n6449), .B2(n4944), .A(n4917), .ZN(n4918) );
  OAI211_X1 U6107 ( .C1(n4947), .C2(n6459), .A(n4919), .B(n4918), .ZN(U3122)
         );
  NAND2_X1 U6108 ( .A1(n4940), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4922)
         );
  OAI22_X1 U6109 ( .A1(n5205), .A2(n4942), .B1(n4941), .B2(n5209), .ZN(n4920)
         );
  AOI21_X1 U6110 ( .B1(n5159), .B2(n4944), .A(n4920), .ZN(n4921) );
  OAI211_X1 U6111 ( .C1(n4947), .C2(n5156), .A(n4922), .B(n4921), .ZN(U3121)
         );
  NAND2_X1 U6112 ( .A1(n4940), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4925)
         );
  OAI22_X1 U6113 ( .A1(n5210), .A2(n4942), .B1(n4941), .B2(n5214), .ZN(n4923)
         );
  AOI21_X1 U6114 ( .B1(n5140), .B2(n4944), .A(n4923), .ZN(n4924) );
  OAI211_X1 U6115 ( .C1(n4947), .C2(n5138), .A(n4925), .B(n4924), .ZN(U3118)
         );
  NAND2_X1 U6116 ( .A1(n4940), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4928)
         );
  OAI22_X1 U6117 ( .A1(n5215), .A2(n4942), .B1(n4941), .B2(n5219), .ZN(n4926)
         );
  AOI21_X1 U6118 ( .B1(n6416), .B2(n4944), .A(n4926), .ZN(n4927) );
  OAI211_X1 U6119 ( .C1(n4947), .C2(n6421), .A(n4928), .B(n4927), .ZN(U3117)
         );
  NAND2_X1 U6120 ( .A1(n4940), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4933)
         );
  INV_X1 U6121 ( .A(n4941), .ZN(n4931) );
  OAI22_X1 U6122 ( .A1(n5190), .A2(n4942), .B1(n6395), .B2(n4929), .ZN(n4930)
         );
  AOI21_X1 U6123 ( .B1(n6445), .B2(n4931), .A(n4930), .ZN(n4932) );
  OAI211_X1 U6124 ( .C1(n4947), .C2(n6448), .A(n4933), .B(n4932), .ZN(U3120)
         );
  NAND2_X1 U6125 ( .A1(n4940), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4936)
         );
  OAI22_X1 U6126 ( .A1(n5220), .A2(n4942), .B1(n4941), .B2(n5224), .ZN(n4934)
         );
  AOI21_X1 U6127 ( .B1(n6431), .B2(n4944), .A(n4934), .ZN(n4935) );
  OAI211_X1 U6128 ( .C1(n4947), .C2(n6436), .A(n4936), .B(n4935), .ZN(U3116)
         );
  NAND2_X1 U6129 ( .A1(n4940), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4939)
         );
  OAI22_X1 U6130 ( .A1(n5227), .A2(n4942), .B1(n4941), .B2(n5232), .ZN(n4937)
         );
  AOI21_X1 U6131 ( .B1(n6437), .B2(n4944), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6132 ( .C1(n4947), .C2(n6442), .A(n4939), .B(n4938), .ZN(U3119)
         );
  NAND2_X1 U6133 ( .A1(n4940), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4946)
         );
  OAI22_X1 U6134 ( .A1(n5200), .A2(n4942), .B1(n4941), .B2(n5204), .ZN(n4943)
         );
  AOI21_X1 U6135 ( .B1(n6348), .B2(n4944), .A(n4943), .ZN(n4945) );
  OAI211_X1 U6136 ( .C1(n4947), .C2(n6355), .A(n4946), .B(n4945), .ZN(U3123)
         );
  XOR2_X1 U6137 ( .A(n4861), .B(n4948), .Z(n5007) );
  INV_X1 U6138 ( .A(n5007), .ZN(n5010) );
  INV_X1 U6139 ( .A(n6080), .ZN(n6086) );
  AND2_X1 U6140 ( .A1(n6082), .A2(n6018), .ZN(n6052) );
  INV_X1 U6141 ( .A(n4950), .ZN(n4953) );
  INV_X1 U6142 ( .A(n4951), .ZN(n4952) );
  AOI21_X1 U6143 ( .B1(n4753), .B2(n4953), .A(n4952), .ZN(n4954) );
  OR2_X1 U6144 ( .A1(n5108), .A2(n4954), .ZN(n5011) );
  INV_X1 U6145 ( .A(n5011), .ZN(n6249) );
  AOI22_X1 U6146 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6054), .B1(n6067), .B2(n6249), 
        .ZN(n4955) );
  OAI211_X1 U6147 ( .C1(n6075), .C2(n4956), .A(n4955), .B(n6302), .ZN(n4957)
         );
  AOI21_X1 U6148 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6052), .A(n4957), .ZN(n4962)
         );
  NAND2_X1 U6149 ( .A1(n5163), .A2(n4958), .ZN(n5034) );
  INV_X1 U6150 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6537) );
  NOR2_X1 U6151 ( .A1(n5034), .A2(n6537), .ZN(n6055) );
  INV_X1 U6152 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6541) );
  INV_X1 U6153 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6539) );
  NOR2_X1 U6154 ( .A1(n6541), .A2(n6539), .ZN(n6040) );
  AOI21_X1 U6155 ( .B1(n6541), .B2(n6539), .A(n6040), .ZN(n4960) );
  INV_X1 U6156 ( .A(n5005), .ZN(n4959) );
  AOI22_X1 U6157 ( .A1(n6055), .A2(n4960), .B1(n4959), .B2(n6062), .ZN(n4961)
         );
  OAI211_X1 U6158 ( .C1(n5010), .C2(n6024), .A(n4962), .B(n4961), .ZN(U2820)
         );
  OAI222_X1 U6159 ( .A1(n5886), .A2(n5010), .B1(n5290), .B2(n6164), .C1(n5541), 
        .C2(n3838), .ZN(U2884) );
  OAI21_X1 U6160 ( .B1(n4965), .B2(n4964), .A(n4963), .ZN(n6270) );
  OAI22_X1 U6161 ( .A1(n5903), .A2(n5035), .B1(n6302), .B2(n6537), .ZN(n4967)
         );
  NOR2_X1 U6162 ( .A1(n5043), .A2(n6211), .ZN(n4966) );
  AOI211_X1 U6163 ( .C1(n6173), .C2(n5037), .A(n4967), .B(n4966), .ZN(n4968)
         );
  OAI21_X1 U6164 ( .B1(n6178), .B2(n6270), .A(n4968), .ZN(U2981) );
  NAND2_X1 U6165 ( .A1(n4969), .A2(n6367), .ZN(n4979) );
  OR2_X1 U6166 ( .A1(n6363), .A2(n4970), .ZN(n6368) );
  OR2_X1 U6167 ( .A1(n6368), .A2(n3792), .ZN(n4971) );
  AND2_X1 U6168 ( .A1(n4971), .A2(n4978), .ZN(n4981) );
  OAI22_X1 U6169 ( .A1(n4979), .A2(n4981), .B1(n4972), .B2(n4378), .ZN(n6426)
         );
  INV_X1 U6170 ( .A(n6426), .ZN(n5000) );
  INV_X1 U6171 ( .A(n6430), .ZN(n4998) );
  INV_X1 U6172 ( .A(n4975), .ZN(n4976) );
  INV_X1 U6173 ( .A(n4978), .ZN(n6425) );
  INV_X1 U6174 ( .A(n4979), .ZN(n4980) );
  NAND2_X1 U6175 ( .A1(n4981), .A2(n4980), .ZN(n4982) );
  OAI211_X1 U6176 ( .C1(n6367), .C2(n6357), .A(n4983), .B(n4982), .ZN(n6427)
         );
  AOI22_X1 U6177 ( .A1(n6452), .A2(n6425), .B1(INSTQUEUE_REG_7__6__SCAN_IN), 
        .B2(n6427), .ZN(n4984) );
  OAI21_X1 U6178 ( .B1(n6405), .B2(n5155), .A(n4984), .ZN(n4985) );
  AOI21_X1 U6179 ( .B1(n6402), .B2(n4998), .A(n4985), .ZN(n4986) );
  OAI21_X1 U6180 ( .B1(n5000), .B2(n5199), .A(n4986), .ZN(U3082) );
  AOI22_X1 U6181 ( .A1(n6383), .A2(n6425), .B1(INSTQUEUE_REG_7__2__SCAN_IN), 
        .B2(n6427), .ZN(n4987) );
  OAI21_X1 U6182 ( .B1(n6387), .B2(n5155), .A(n4987), .ZN(n4988) );
  AOI21_X1 U6183 ( .B1(n6384), .B2(n4998), .A(n4988), .ZN(n4989) );
  OAI21_X1 U6184 ( .B1(n5000), .B2(n5214), .A(n4989), .ZN(U3078) );
  AOI22_X1 U6185 ( .A1(n6432), .A2(n6425), .B1(INSTQUEUE_REG_7__0__SCAN_IN), 
        .B2(n6427), .ZN(n4990) );
  OAI21_X1 U6186 ( .B1(n6377), .B2(n5155), .A(n4990), .ZN(n4991) );
  AOI21_X1 U6187 ( .B1(n6374), .B2(n4998), .A(n4991), .ZN(n4992) );
  OAI21_X1 U6188 ( .B1(n5000), .B2(n5224), .A(n4992), .ZN(U3076) );
  AOI22_X1 U6189 ( .A1(n6409), .A2(n6425), .B1(INSTQUEUE_REG_7__7__SCAN_IN), 
        .B2(n6427), .ZN(n4993) );
  OAI21_X1 U6190 ( .B1(n6415), .B2(n5155), .A(n4993), .ZN(n4994) );
  AOI21_X1 U6191 ( .B1(n6411), .B2(n4998), .A(n4994), .ZN(n4995) );
  OAI21_X1 U6192 ( .B1(n5000), .B2(n5204), .A(n4995), .ZN(U3083) );
  AOI22_X1 U6193 ( .A1(n6397), .A2(n6425), .B1(INSTQUEUE_REG_7__5__SCAN_IN), 
        .B2(n6427), .ZN(n4996) );
  OAI21_X1 U6194 ( .B1(n6401), .B2(n5155), .A(n4996), .ZN(n4997) );
  AOI21_X1 U6195 ( .B1(n6398), .B2(n4998), .A(n4997), .ZN(n4999) );
  OAI21_X1 U6196 ( .B1(n5000), .B2(n5209), .A(n4999), .ZN(U3081) );
  OAI21_X1 U6197 ( .B1(n5003), .B2(n5002), .A(n3019), .ZN(n6250) );
  NAND2_X1 U6198 ( .A1(n6273), .A2(REIP_REG_7__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U6199 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5004)
         );
  OAI211_X1 U6200 ( .C1(n6202), .C2(n5005), .A(n6247), .B(n5004), .ZN(n5006)
         );
  AOI21_X1 U6201 ( .B1(n5007), .B2(n6184), .A(n5006), .ZN(n5008) );
  OAI21_X1 U6202 ( .B1(n6250), .B2(n6178), .A(n5008), .ZN(U2979) );
  INV_X1 U6203 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5009) );
  OAI222_X1 U6204 ( .A1(n5011), .A2(n5536), .B1(n3010), .B2(n5010), .C1(n5009), 
        .C2(n5538), .ZN(U2852) );
  NAND2_X1 U6205 ( .A1(n5012), .A2(n5412), .ZN(n5013) );
  AOI22_X1 U6206 ( .A1(n6612), .A2(UWORD_REG_9__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5016) );
  OAI21_X1 U6207 ( .B1(n5017), .B2(n6108), .A(n5016), .ZN(U2898) );
  AOI22_X1 U6208 ( .A1(n6612), .A2(UWORD_REG_2__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5018) );
  OAI21_X1 U6209 ( .B1(n5019), .B2(n6108), .A(n5018), .ZN(U2905) );
  AOI22_X1 U6210 ( .A1(n6612), .A2(UWORD_REG_1__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5020) );
  OAI21_X1 U6211 ( .B1(n5021), .B2(n6108), .A(n5020), .ZN(U2906) );
  AOI22_X1 U6212 ( .A1(n6612), .A2(UWORD_REG_0__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5022) );
  OAI21_X1 U6213 ( .B1(n5023), .B2(n6108), .A(n5022), .ZN(U2907) );
  INV_X1 U6214 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5025) );
  AOI22_X1 U6215 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n5060), .B1(n6139), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5024) );
  OAI21_X1 U6216 ( .B1(n5025), .B2(n6108), .A(n5024), .ZN(U2902) );
  OAI21_X1 U6217 ( .B1(n5026), .B2(n5029), .A(n5028), .ZN(n6044) );
  AOI22_X1 U6218 ( .A1(n5383), .A2(DATAI_8_), .B1(n6620), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5030) );
  OAI21_X1 U6219 ( .B1(n6044), .B2(n5886), .A(n5030), .ZN(U2883) );
  XOR2_X1 U6220 ( .A(n5107), .B(n5108), .Z(n6242) );
  AOI22_X1 U6221 ( .A1(n5515), .A2(n6242), .B1(n4864), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5031) );
  OAI21_X1 U6222 ( .B1(n6044), .B2(n3010), .A(n5031), .ZN(U2851) );
  NAND2_X1 U6223 ( .A1(n6609), .A2(n5032), .ZN(n5033) );
  NAND2_X1 U6224 ( .A1(n6537), .A2(n5034), .ZN(n5041) );
  OAI22_X1 U6225 ( .A1(n3655), .A2(n6094), .B1(n5035), .B2(n6075), .ZN(n5036)
         );
  AOI211_X1 U6226 ( .C1(n6062), .C2(n5037), .A(n5036), .B(n6282), .ZN(n5038)
         );
  OAI21_X1 U6227 ( .B1(n6093), .B2(n5039), .A(n5038), .ZN(n5040) );
  AOI21_X1 U6228 ( .B1(n6052), .B2(n5041), .A(n5040), .ZN(n5042) );
  OAI21_X1 U6229 ( .B1(n5415), .B2(n5043), .A(n5042), .ZN(U2822) );
  AOI22_X1 U6230 ( .A1(n5060), .A2(UWORD_REG_14__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5044) );
  OAI21_X1 U6231 ( .B1(n5045), .B2(n6108), .A(n5044), .ZN(U2893) );
  INV_X1 U6232 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5047) );
  AOI22_X1 U6233 ( .A1(n5060), .A2(UWORD_REG_12__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5046) );
  OAI21_X1 U6234 ( .B1(n5047), .B2(n6108), .A(n5046), .ZN(U2895) );
  AOI22_X1 U6235 ( .A1(n5060), .A2(UWORD_REG_3__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5048) );
  OAI21_X1 U6236 ( .B1(n5049), .B2(n6108), .A(n5048), .ZN(U2904) );
  AOI22_X1 U6237 ( .A1(n5060), .A2(UWORD_REG_8__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5050) );
  OAI21_X1 U6238 ( .B1(n5051), .B2(n6108), .A(n5050), .ZN(U2899) );
  INV_X1 U6239 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U6240 ( .A1(n5060), .A2(UWORD_REG_6__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5052) );
  OAI21_X1 U6241 ( .B1(n5053), .B2(n6108), .A(n5052), .ZN(U2901) );
  INV_X1 U6242 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5055) );
  AOI22_X1 U6243 ( .A1(n5060), .A2(UWORD_REG_7__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5054) );
  OAI21_X1 U6244 ( .B1(n5055), .B2(n6108), .A(n5054), .ZN(U2900) );
  AOI22_X1 U6245 ( .A1(n5060), .A2(UWORD_REG_10__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5056) );
  OAI21_X1 U6246 ( .B1(n5057), .B2(n6108), .A(n5056), .ZN(U2897) );
  AOI22_X1 U6247 ( .A1(n5060), .A2(UWORD_REG_11__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5058) );
  OAI21_X1 U6248 ( .B1(n5059), .B2(n6108), .A(n5058), .ZN(U2896) );
  AOI22_X1 U6249 ( .A1(n5060), .A2(UWORD_REG_13__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5061) );
  OAI21_X1 U6250 ( .B1(n6755), .B2(n6108), .A(n5061), .ZN(U2894) );
  NOR2_X1 U6251 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5062), .ZN(n5075)
         );
  INV_X1 U6252 ( .A(n5100), .ZN(n5070) );
  OAI21_X1 U6253 ( .B1(n5070), .B2(n6349), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5064) );
  AND2_X1 U6254 ( .A1(n5064), .A2(n5063), .ZN(n5066) );
  AOI211_X1 U6255 ( .C1(n6367), .C2(n5066), .A(n6314), .B(n5065), .ZN(n5067)
         );
  INV_X1 U6256 ( .A(n5094), .ZN(n5074) );
  INV_X1 U6257 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5073) );
  AOI22_X1 U6258 ( .A1(n6358), .A2(n5068), .B1(n6361), .B2(n3102), .ZN(n5095)
         );
  INV_X1 U6259 ( .A(n5095), .ZN(n5069) );
  AOI22_X1 U6260 ( .A1(n6445), .A2(n5069), .B1(n5075), .B2(n6443), .ZN(n5072)
         );
  AOI22_X1 U6261 ( .A1(n5070), .A2(n6444), .B1(n6349), .B2(n6392), .ZN(n5071)
         );
  OAI211_X1 U6262 ( .C1(n5074), .C2(n5073), .A(n5072), .B(n5071), .ZN(U3056)
         );
  NAND2_X1 U6263 ( .A1(n5094), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5078) );
  INV_X1 U6264 ( .A(n5075), .ZN(n5096) );
  OAI22_X1 U6265 ( .A1(n5227), .A2(n5096), .B1(n5095), .B2(n5232), .ZN(n5076)
         );
  AOI21_X1 U6266 ( .B1(n6349), .B2(n6388), .A(n5076), .ZN(n5077) );
  OAI211_X1 U6267 ( .C1(n5100), .C2(n6391), .A(n5078), .B(n5077), .ZN(U3055)
         );
  NAND2_X1 U6268 ( .A1(n5094), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5081) );
  OAI22_X1 U6269 ( .A1(n5200), .A2(n5096), .B1(n5095), .B2(n5204), .ZN(n5079)
         );
  AOI21_X1 U6270 ( .B1(n6349), .B2(n6411), .A(n5079), .ZN(n5080) );
  OAI211_X1 U6271 ( .C1(n5100), .C2(n6415), .A(n5081), .B(n5080), .ZN(U3059)
         );
  NAND2_X1 U6272 ( .A1(n5094), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5084) );
  OAI22_X1 U6273 ( .A1(n5195), .A2(n5096), .B1(n5095), .B2(n5199), .ZN(n5082)
         );
  AOI21_X1 U6274 ( .B1(n6349), .B2(n6402), .A(n5082), .ZN(n5083) );
  OAI211_X1 U6275 ( .C1(n5100), .C2(n6405), .A(n5084), .B(n5083), .ZN(U3058)
         );
  NAND2_X1 U6276 ( .A1(n5094), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5087) );
  OAI22_X1 U6277 ( .A1(n5220), .A2(n5096), .B1(n5095), .B2(n5224), .ZN(n5085)
         );
  AOI21_X1 U6278 ( .B1(n6349), .B2(n6374), .A(n5085), .ZN(n5086) );
  OAI211_X1 U6279 ( .C1(n6377), .C2(n5100), .A(n5087), .B(n5086), .ZN(U3052)
         );
  NAND2_X1 U6280 ( .A1(n5094), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5090) );
  OAI22_X1 U6281 ( .A1(n5210), .A2(n5096), .B1(n5095), .B2(n5214), .ZN(n5088)
         );
  AOI21_X1 U6282 ( .B1(n6349), .B2(n6384), .A(n5088), .ZN(n5089) );
  OAI211_X1 U6283 ( .C1(n5100), .C2(n6387), .A(n5090), .B(n5089), .ZN(U3054)
         );
  NAND2_X1 U6284 ( .A1(n5094), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5093) );
  OAI22_X1 U6285 ( .A1(n5215), .A2(n5096), .B1(n5095), .B2(n5219), .ZN(n5091)
         );
  AOI21_X1 U6286 ( .B1(n6349), .B2(n6378), .A(n5091), .ZN(n5092) );
  OAI211_X1 U6287 ( .C1(n5100), .C2(n6381), .A(n5093), .B(n5092), .ZN(U3053)
         );
  NAND2_X1 U6288 ( .A1(n5094), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5099) );
  OAI22_X1 U6289 ( .A1(n5205), .A2(n5096), .B1(n5095), .B2(n5209), .ZN(n5097)
         );
  AOI21_X1 U6290 ( .B1(n6349), .B2(n6398), .A(n5097), .ZN(n5098) );
  OAI211_X1 U6291 ( .C1(n5100), .C2(n6401), .A(n5099), .B(n5098), .ZN(U3057)
         );
  NAND2_X1 U6292 ( .A1(n5028), .A2(n5102), .ZN(n5103) );
  NAND2_X1 U6293 ( .A1(n5101), .A2(n5103), .ZN(n6031) );
  AOI22_X1 U6294 ( .A1(n5383), .A2(DATAI_9_), .B1(n6620), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5104) );
  OAI21_X1 U6295 ( .B1(n6031), .B2(n5886), .A(n5104), .ZN(U2882) );
  AOI21_X1 U6296 ( .B1(n5108), .B2(n5107), .A(n5106), .ZN(n5109) );
  NOR2_X1 U6297 ( .A1(n3675), .A2(n5109), .ZN(n6233) );
  AOI22_X1 U6298 ( .A1(n5515), .A2(n6233), .B1(n4864), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5110) );
  OAI21_X1 U6299 ( .B1(n6031), .B2(n3010), .A(n5110), .ZN(U2850) );
  OAI21_X1 U6300 ( .B1(n5158), .B2(n6424), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5117) );
  AOI21_X1 U6301 ( .B1(n5111), .B2(n3023), .A(n6316), .ZN(n5116) );
  NOR2_X1 U6302 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5112), .ZN(n5153)
         );
  OAI21_X1 U6303 ( .B1(n6591), .B2(n5153), .A(n5113), .ZN(n5115) );
  INV_X1 U6304 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5124) );
  OAI22_X1 U6305 ( .A1(n5120), .A2(n5119), .B1(n5180), .B2(n5118), .ZN(n5152)
         );
  AOI22_X1 U6306 ( .A1(n6409), .A2(n5153), .B1(n6407), .B2(n5152), .ZN(n5121)
         );
  OAI21_X1 U6307 ( .B1(n6355), .B2(n5155), .A(n5121), .ZN(n5122) );
  AOI21_X1 U6308 ( .B1(n6348), .B2(n5158), .A(n5122), .ZN(n5123) );
  OAI21_X1 U6309 ( .B1(n5162), .B2(n5124), .A(n5123), .ZN(U3091) );
  INV_X1 U6310 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U6311 ( .A1(n6438), .A2(n5153), .B1(n6439), .B2(n5152), .ZN(n5125)
         );
  OAI21_X1 U6312 ( .B1(n6442), .B2(n5155), .A(n5125), .ZN(n5126) );
  AOI21_X1 U6313 ( .B1(n6437), .B2(n5158), .A(n5126), .ZN(n5127) );
  OAI21_X1 U6314 ( .B1(n5162), .B2(n5128), .A(n5127), .ZN(U3087) );
  INV_X1 U6315 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5132) );
  AOI22_X1 U6316 ( .A1(n6417), .A2(n5153), .B1(n6418), .B2(n5152), .ZN(n5129)
         );
  OAI21_X1 U6317 ( .B1(n6421), .B2(n5155), .A(n5129), .ZN(n5130) );
  AOI21_X1 U6318 ( .B1(n6416), .B2(n5158), .A(n5130), .ZN(n5131) );
  OAI21_X1 U6319 ( .B1(n5162), .B2(n5132), .A(n5131), .ZN(U3085) );
  INV_X1 U6320 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5136) );
  AOI22_X1 U6321 ( .A1(n6452), .A2(n5153), .B1(n6454), .B2(n5152), .ZN(n5133)
         );
  OAI21_X1 U6322 ( .B1(n6459), .B2(n5155), .A(n5133), .ZN(n5134) );
  AOI21_X1 U6323 ( .B1(n6449), .B2(n5158), .A(n5134), .ZN(n5135) );
  OAI21_X1 U6324 ( .B1(n5162), .B2(n5136), .A(n5135), .ZN(U3090) );
  INV_X1 U6325 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5142) );
  AOI22_X1 U6326 ( .A1(n6383), .A2(n5153), .B1(n6382), .B2(n5152), .ZN(n5137)
         );
  OAI21_X1 U6327 ( .B1(n5138), .B2(n5155), .A(n5137), .ZN(n5139) );
  AOI21_X1 U6328 ( .B1(n5140), .B2(n5158), .A(n5139), .ZN(n5141) );
  OAI21_X1 U6329 ( .B1(n5162), .B2(n5142), .A(n5141), .ZN(U3086) );
  INV_X1 U6330 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5146) );
  AOI22_X1 U6331 ( .A1(n6432), .A2(n5153), .B1(n6433), .B2(n5152), .ZN(n5143)
         );
  OAI21_X1 U6332 ( .B1(n6436), .B2(n5155), .A(n5143), .ZN(n5144) );
  AOI21_X1 U6333 ( .B1(n6431), .B2(n5158), .A(n5144), .ZN(n5145) );
  OAI21_X1 U6334 ( .B1(n5162), .B2(n5146), .A(n5145), .ZN(U3084) );
  INV_X1 U6335 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5151) );
  INV_X1 U6336 ( .A(n5152), .ZN(n5148) );
  AOI22_X1 U6337 ( .A1(n6443), .A2(n5153), .B1(n6392), .B2(n6424), .ZN(n5147)
         );
  OAI21_X1 U6338 ( .B1(n5194), .B2(n5148), .A(n5147), .ZN(n5149) );
  AOI21_X1 U6339 ( .B1(n6444), .B2(n5158), .A(n5149), .ZN(n5150) );
  OAI21_X1 U6340 ( .B1(n5162), .B2(n5151), .A(n5150), .ZN(U3088) );
  INV_X1 U6341 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5161) );
  AOI22_X1 U6342 ( .A1(n6397), .A2(n5153), .B1(n6396), .B2(n5152), .ZN(n5154)
         );
  OAI21_X1 U6343 ( .B1(n5156), .B2(n5155), .A(n5154), .ZN(n5157) );
  AOI21_X1 U6344 ( .B1(n5159), .B2(n5158), .A(n5157), .ZN(n5160) );
  OAI21_X1 U6345 ( .B1(n5162), .B2(n5161), .A(n5160), .ZN(U3089) );
  NAND2_X1 U6346 ( .A1(n5163), .A2(n6060), .ZN(n5165) );
  NAND2_X1 U6347 ( .A1(n5165), .A2(n6080), .ZN(n6066) );
  NAND2_X1 U6348 ( .A1(n6067), .A2(n6289), .ZN(n5168) );
  NAND2_X1 U6349 ( .A1(n5163), .A2(n6599), .ZN(n6088) );
  NAND2_X1 U6350 ( .A1(n6088), .A2(REIP_REG_2__SCAN_IN), .ZN(n5164) );
  NOR2_X1 U6351 ( .A1(n5165), .A2(n5164), .ZN(n5166) );
  AOI21_X1 U6352 ( .B1(n6087), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5166), 
        .ZN(n5167) );
  OAI211_X1 U6353 ( .C1(n6101), .C2(n5169), .A(n5168), .B(n5167), .ZN(n5174)
         );
  INV_X1 U6354 ( .A(EBX_REG_3__SCAN_IN), .ZN(n5172) );
  AND2_X1 U6355 ( .A1(n6609), .A2(n5170), .ZN(n6065) );
  INV_X1 U6356 ( .A(n6065), .ZN(n6091) );
  OAI22_X1 U6357 ( .A1(n5172), .A2(n6094), .B1(n6091), .B2(n5171), .ZN(n5173)
         );
  AOI211_X1 U6358 ( .C1(n6066), .C2(REIP_REG_3__SCAN_IN), .A(n5174), .B(n5173), 
        .ZN(n5175) );
  OAI21_X1 U6359 ( .B1(n5415), .B2(n5176), .A(n5175), .ZN(U2824) );
  INV_X1 U6360 ( .A(n6458), .ZN(n5178) );
  OAI21_X1 U6361 ( .B1(n5229), .B2(n5178), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5179) );
  NAND2_X1 U6362 ( .A1(n5179), .A2(n6367), .ZN(n5188) );
  INV_X1 U6363 ( .A(n5188), .ZN(n5182) );
  NOR2_X1 U6364 ( .A1(n5180), .A2(n6359), .ZN(n5181) );
  NOR2_X1 U6365 ( .A1(n6361), .A2(n5183), .ZN(n6321) );
  NOR2_X1 U6366 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5184), .ZN(n5189)
         );
  OAI22_X1 U6367 ( .A1(n4378), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n6591), .B2(n5189), .ZN(n5185) );
  INV_X1 U6368 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6369 ( .A1(n5225), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5193)
         );
  INV_X1 U6370 ( .A(n5189), .ZN(n5226) );
  OAI22_X1 U6371 ( .A1(n5190), .A2(n5226), .B1(n6395), .B2(n6458), .ZN(n5191)
         );
  AOI21_X1 U6372 ( .B1(n6392), .B2(n5229), .A(n5191), .ZN(n5192) );
  OAI211_X1 U6373 ( .C1(n5233), .C2(n5194), .A(n5193), .B(n5192), .ZN(U3104)
         );
  NAND2_X1 U6374 ( .A1(n5225), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5198)
         );
  OAI22_X1 U6375 ( .A1(n5195), .A2(n5226), .B1(n6458), .B2(n6405), .ZN(n5196)
         );
  AOI21_X1 U6376 ( .B1(n6402), .B2(n5229), .A(n5196), .ZN(n5197) );
  OAI211_X1 U6377 ( .C1(n5233), .C2(n5199), .A(n5198), .B(n5197), .ZN(U3106)
         );
  NAND2_X1 U6378 ( .A1(n5225), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5203)
         );
  OAI22_X1 U6379 ( .A1(n5200), .A2(n5226), .B1(n6458), .B2(n6415), .ZN(n5201)
         );
  AOI21_X1 U6380 ( .B1(n6411), .B2(n5229), .A(n5201), .ZN(n5202) );
  OAI211_X1 U6381 ( .C1(n5233), .C2(n5204), .A(n5203), .B(n5202), .ZN(U3107)
         );
  NAND2_X1 U6382 ( .A1(n5225), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5208)
         );
  OAI22_X1 U6383 ( .A1(n5205), .A2(n5226), .B1(n6458), .B2(n6401), .ZN(n5206)
         );
  AOI21_X1 U6384 ( .B1(n6398), .B2(n5229), .A(n5206), .ZN(n5207) );
  OAI211_X1 U6385 ( .C1(n5233), .C2(n5209), .A(n5208), .B(n5207), .ZN(U3105)
         );
  NAND2_X1 U6386 ( .A1(n5225), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5213)
         );
  OAI22_X1 U6387 ( .A1(n5210), .A2(n5226), .B1(n6458), .B2(n6387), .ZN(n5211)
         );
  AOI21_X1 U6388 ( .B1(n6384), .B2(n5229), .A(n5211), .ZN(n5212) );
  OAI211_X1 U6389 ( .C1(n5233), .C2(n5214), .A(n5213), .B(n5212), .ZN(U3102)
         );
  NAND2_X1 U6390 ( .A1(n5225), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5218)
         );
  OAI22_X1 U6391 ( .A1(n5215), .A2(n5226), .B1(n6458), .B2(n6381), .ZN(n5216)
         );
  AOI21_X1 U6392 ( .B1(n6378), .B2(n5229), .A(n5216), .ZN(n5217) );
  OAI211_X1 U6393 ( .C1(n5233), .C2(n5219), .A(n5218), .B(n5217), .ZN(U3101)
         );
  NAND2_X1 U6394 ( .A1(n5225), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5223)
         );
  OAI22_X1 U6395 ( .A1(n5220), .A2(n5226), .B1(n6458), .B2(n6377), .ZN(n5221)
         );
  AOI21_X1 U6396 ( .B1(n6374), .B2(n5229), .A(n5221), .ZN(n5222) );
  OAI211_X1 U6397 ( .C1(n5233), .C2(n5224), .A(n5223), .B(n5222), .ZN(U3100)
         );
  NAND2_X1 U6398 ( .A1(n5225), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5231)
         );
  OAI22_X1 U6399 ( .A1(n5227), .A2(n5226), .B1(n6458), .B2(n6391), .ZN(n5228)
         );
  AOI21_X1 U6400 ( .B1(n6388), .B2(n5229), .A(n5228), .ZN(n5230) );
  OAI211_X1 U6401 ( .C1(n5233), .C2(n5232), .A(n5231), .B(n5230), .ZN(U3103)
         );
  OAI21_X1 U6402 ( .B1(n5236), .B2(n5235), .A(n5234), .ZN(n5237) );
  INV_X1 U6403 ( .A(n5237), .ZN(n6243) );
  NAND2_X1 U6404 ( .A1(n6243), .A2(n6206), .ZN(n5240) );
  AND2_X1 U6405 ( .A1(n6273), .A2(REIP_REG_8__SCAN_IN), .ZN(n6241) );
  NOR2_X1 U6406 ( .A1(n6202), .A2(n6045), .ZN(n5238) );
  AOI211_X1 U6407 ( .C1(n6208), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6241), 
        .B(n5238), .ZN(n5239) );
  OAI211_X1 U6408 ( .C1(n6211), .C2(n6044), .A(n5240), .B(n5239), .ZN(U2978)
         );
  AOI21_X1 U6409 ( .B1(n5243), .B2(n5101), .A(n5242), .ZN(n5266) );
  INV_X1 U6410 ( .A(n5266), .ZN(n6025) );
  AOI22_X1 U6411 ( .A1(n5383), .A2(DATAI_10_), .B1(n6620), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5244) );
  OAI21_X1 U6412 ( .B1(n6025), .B2(n5886), .A(n5244), .ZN(U2881) );
  NAND2_X1 U6413 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  NAND2_X1 U6414 ( .A1(n5269), .A2(n5247), .ZN(n6225) );
  OAI222_X1 U6415 ( .A1(n6025), .A2(n3010), .B1(n5538), .B2(n6667), .C1(n6225), 
        .C2(n5536), .ZN(U2849) );
  NAND2_X1 U6416 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  XNOR2_X1 U6417 ( .A(n5248), .B(n5251), .ZN(n6235) );
  NAND2_X1 U6418 ( .A1(n6235), .A2(n6206), .ZN(n5255) );
  AND2_X1 U6419 ( .A1(n6273), .A2(REIP_REG_9__SCAN_IN), .ZN(n6232) );
  NOR2_X1 U6420 ( .A1(n6202), .A2(n5252), .ZN(n5253) );
  AOI211_X1 U6421 ( .C1(n6208), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6232), 
        .B(n5253), .ZN(n5254) );
  OAI211_X1 U6422 ( .C1(n6211), .C2(n6031), .A(n5255), .B(n5254), .ZN(U2977)
         );
  NOR2_X1 U6423 ( .A1(n5242), .A2(n5257), .ZN(n5258) );
  OR2_X1 U6424 ( .A1(n5256), .A2(n5258), .ZN(n6012) );
  AOI22_X1 U6425 ( .A1(n5383), .A2(DATAI_11_), .B1(n6620), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5259) );
  OAI21_X1 U6426 ( .B1(n6012), .B2(n5886), .A(n5259), .ZN(U2880) );
  NAND2_X1 U6427 ( .A1(n6169), .A2(n5260), .ZN(n5262) );
  XOR2_X1 U6428 ( .A(n5262), .B(n5261), .Z(n6223) );
  INV_X1 U6429 ( .A(n6028), .ZN(n5264) );
  AOI22_X1 U6430 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6273), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5263) );
  OAI21_X1 U6431 ( .B1(n5264), .B2(n6202), .A(n5263), .ZN(n5265) );
  AOI21_X1 U6432 ( .B1(n5266), .B2(n6184), .A(n5265), .ZN(n5267) );
  OAI21_X1 U6433 ( .B1(n6223), .B2(n6178), .A(n5267), .ZN(U2976) );
  AND2_X1 U6434 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  OR2_X1 U6435 ( .A1(n5270), .A2(n5276), .ZN(n6011) );
  OAI222_X1 U6436 ( .A1(n6012), .A2(n3010), .B1(n5538), .B2(n5271), .C1(n5536), 
        .C2(n6011), .ZN(U2848) );
  OR2_X1 U6437 ( .A1(n5256), .A2(n5273), .ZN(n5274) );
  AND2_X1 U6438 ( .A1(n5272), .A2(n5274), .ZN(n5298) );
  NOR2_X1 U6439 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  OR2_X1 U6440 ( .A1(n5317), .A2(n5277), .ZN(n5306) );
  OAI22_X1 U6441 ( .A1(n5306), .A2(n5536), .B1(n5278), .B2(n5538), .ZN(n5279)
         );
  AOI21_X1 U6442 ( .B1(n5298), .B2(n5350), .A(n5279), .ZN(n5280) );
  INV_X1 U6443 ( .A(n5280), .ZN(U2847) );
  INV_X1 U6444 ( .A(n5298), .ZN(n5291) );
  INV_X1 U6445 ( .A(n5281), .ZN(n5282) );
  AOI21_X1 U6446 ( .B1(n6080), .B2(n5282), .A(n5875), .ZN(n6013) );
  NOR2_X1 U6447 ( .A1(n6101), .A2(n5296), .ZN(n5285) );
  AOI22_X1 U6448 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6054), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6087), .ZN(n5283) );
  OAI211_X1 U6449 ( .C1(n5306), .C2(n6093), .A(n5283), .B(n6302), .ZN(n5284)
         );
  AOI211_X1 U6450 ( .C1(n6013), .C2(REIP_REG_12__SCAN_IN), .A(n5285), .B(n5284), .ZN(n5289) );
  INV_X1 U6451 ( .A(n5286), .ZN(n5287) );
  NOR2_X1 U6452 ( .A1(n6079), .A2(n5287), .ZN(n6021) );
  NAND4_X1 U6453 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n6021), .ZN(n5332) );
  NOR2_X1 U6454 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5332), .ZN(n5325) );
  INV_X1 U6455 ( .A(n5325), .ZN(n5288) );
  OAI211_X1 U6456 ( .C1(n5291), .C2(n6024), .A(n5289), .B(n5288), .ZN(U2815)
         );
  INV_X1 U6457 ( .A(DATAI_12_), .ZN(n6167) );
  INV_X1 U6458 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6802) );
  OAI222_X1 U6459 ( .A1(n5291), .A2(n5886), .B1(n5290), .B2(n6167), .C1(n5541), 
        .C2(n6802), .ZN(U2879) );
  NOR2_X1 U6460 ( .A1(n5292), .A2(n3042), .ZN(n5293) );
  XNOR2_X1 U6461 ( .A(n5294), .B(n5293), .ZN(n5311) );
  NAND2_X1 U6462 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5295)
         );
  NAND2_X1 U6463 ( .A1(n6273), .A2(REIP_REG_12__SCAN_IN), .ZN(n5305) );
  OAI211_X1 U6464 ( .C1(n6202), .C2(n5296), .A(n5295), .B(n5305), .ZN(n5297)
         );
  AOI21_X1 U6465 ( .B1(n5298), .B2(n6184), .A(n5297), .ZN(n5299) );
  OAI21_X1 U6466 ( .B1(n5311), .B2(n6178), .A(n5299), .ZN(U2974) );
  NOR3_X1 U6467 ( .A1(n6279), .A2(n5932), .A3(n5300), .ZN(n5303) );
  INV_X1 U6468 ( .A(n6221), .ZN(n5750) );
  AOI22_X1 U6469 ( .A1(n6257), .A2(n5302), .B1(n5750), .B2(n5301), .ZN(n5912)
         );
  OAI21_X1 U6470 ( .B1(n5933), .B2(n5303), .A(n5912), .ZN(n5309) );
  OAI21_X1 U6471 ( .B1(n5916), .B2(n3531), .A(n5304), .ZN(n5308) );
  OAI21_X1 U6472 ( .B1(n6304), .B2(n5306), .A(n5305), .ZN(n5307) );
  AOI21_X1 U6473 ( .B1(n5309), .B2(n5308), .A(n5307), .ZN(n5310) );
  OAI21_X1 U6474 ( .B1(n5311), .B2(n6224), .A(n5310), .ZN(U3006) );
  AOI21_X1 U6475 ( .B1(n5314), .B2(n5272), .A(n3951), .ZN(n5357) );
  INV_X1 U6476 ( .A(n5357), .ZN(n5328) );
  AOI22_X1 U6477 ( .A1(n5383), .A2(DATAI_13_), .B1(n6620), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5315) );
  OAI21_X1 U6478 ( .B1(n5328), .B2(n5886), .A(n5315), .ZN(U2878) );
  OAI21_X1 U6479 ( .B1(n5317), .B2(n5316), .A(n5336), .ZN(n5318) );
  INV_X1 U6480 ( .A(n5318), .ZN(n5936) );
  AOI22_X1 U6481 ( .A1(n5936), .A2(n5515), .B1(n4864), .B2(EBX_REG_13__SCAN_IN), .ZN(n5319) );
  OAI21_X1 U6482 ( .B1(n5328), .B2(n3010), .A(n5319), .ZN(U2846) );
  INV_X1 U6483 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6549) );
  NOR3_X1 U6484 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6549), .A3(n5332), .ZN(n5323) );
  INV_X1 U6485 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5321) );
  AOI22_X1 U6486 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6087), .B1(n6067), 
        .B2(n5936), .ZN(n5320) );
  OAI211_X1 U6487 ( .C1(n6094), .C2(n5321), .A(n5320), .B(n6302), .ZN(n5322)
         );
  AOI211_X1 U6488 ( .C1(n6062), .C2(n5324), .A(n5323), .B(n5322), .ZN(n5327)
         );
  OAI21_X1 U6489 ( .B1(n5325), .B2(n6013), .A(REIP_REG_13__SCAN_IN), .ZN(n5326) );
  OAI211_X1 U6490 ( .C1(n5328), .C2(n6024), .A(n5327), .B(n5326), .ZN(U2814)
         );
  INV_X1 U6491 ( .A(n5329), .ZN(n5330) );
  AOI21_X1 U6492 ( .B1(n5331), .B2(n5313), .A(n5330), .ZN(n5378) );
  INV_X1 U6493 ( .A(n5378), .ZN(n5347) );
  NOR3_X1 U6494 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5333), .A3(n5332), .ZN(n5344) );
  NAND2_X1 U6495 ( .A1(n6082), .A2(n5334), .ZN(n6009) );
  NOR2_X1 U6496 ( .A1(n6551), .A2(n6009), .ZN(n5343) );
  INV_X1 U6497 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5341) );
  INV_X1 U6498 ( .A(n5376), .ZN(n5339) );
  NAND2_X1 U6499 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  NAND2_X1 U6500 ( .A1(n5533), .A2(n5337), .ZN(n5362) );
  OAI22_X1 U6501 ( .A1(n5348), .A2(n6094), .B1(n6093), .B2(n5362), .ZN(n5338)
         );
  AOI211_X1 U6502 ( .C1(n6062), .C2(n5339), .A(n5338), .B(n6273), .ZN(n5340)
         );
  OAI21_X1 U6503 ( .B1(n5341), .B2(n6075), .A(n5340), .ZN(n5342) );
  NOR3_X1 U6504 ( .A1(n5344), .A2(n5343), .A3(n5342), .ZN(n5345) );
  OAI21_X1 U6505 ( .B1(n5347), .B2(n6024), .A(n5345), .ZN(U2813) );
  AOI22_X1 U6506 ( .A1(n5383), .A2(DATAI_14_), .B1(n6620), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5346) );
  OAI21_X1 U6507 ( .B1(n5347), .B2(n5886), .A(n5346), .ZN(U2877) );
  OAI22_X1 U6508 ( .A1(n5362), .A2(n5536), .B1(n5348), .B2(n5538), .ZN(n5349)
         );
  AOI21_X1 U6509 ( .B1(n5378), .B2(n5350), .A(n5349), .ZN(n5351) );
  INV_X1 U6510 ( .A(n5351), .ZN(U2845) );
  XOR2_X1 U6511 ( .A(n5352), .B(n5353), .Z(n5937) );
  NAND2_X1 U6512 ( .A1(n6273), .A2(REIP_REG_13__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U6513 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5354)
         );
  OAI211_X1 U6514 ( .C1(n6202), .C2(n5355), .A(n5934), .B(n5354), .ZN(n5356)
         );
  AOI21_X1 U6515 ( .B1(n5357), .B2(n6184), .A(n5356), .ZN(n5358) );
  OAI21_X1 U6516 ( .B1(n5937), .B2(n6178), .A(n5358), .ZN(U2973) );
  XNOR2_X1 U6517 ( .A(n5650), .B(n5360), .ZN(n5361) );
  XNOR2_X1 U6518 ( .A(n5359), .B(n5361), .ZN(n5380) );
  INV_X1 U6519 ( .A(n5362), .ZN(n5372) );
  AND2_X1 U6520 ( .A1(n6273), .A2(REIP_REG_14__SCAN_IN), .ZN(n5374) );
  NOR2_X1 U6521 ( .A1(n5916), .A2(n5367), .ZN(n5370) );
  INV_X1 U6522 ( .A(n5363), .ZN(n5368) );
  INV_X1 U6523 ( .A(n5912), .ZN(n6215) );
  NAND3_X1 U6524 ( .A1(n5933), .A2(n5940), .A3(n5364), .ZN(n5939) );
  OAI21_X1 U6525 ( .B1(n5365), .B2(n5933), .A(n5939), .ZN(n5366) );
  AOI211_X1 U6526 ( .C1(n5368), .C2(n5367), .A(n6215), .B(n5366), .ZN(n5938)
         );
  INV_X1 U6527 ( .A(n5938), .ZN(n5369) );
  MUX2_X1 U6528 ( .A(n5370), .B(n5369), .S(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .Z(n5371) );
  AOI211_X1 U6529 ( .C1(n6290), .C2(n5372), .A(n5374), .B(n5371), .ZN(n5373)
         );
  OAI21_X1 U6530 ( .B1(n5380), .B2(n6224), .A(n5373), .ZN(U3004) );
  AOI21_X1 U6531 ( .B1(n6208), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5374), 
        .ZN(n5375) );
  OAI21_X1 U6532 ( .B1(n5376), .B2(n6202), .A(n5375), .ZN(n5377) );
  AOI21_X1 U6533 ( .B1(n5378), .B2(n6184), .A(n5377), .ZN(n5379) );
  OAI21_X1 U6534 ( .B1(n5380), .B2(n6178), .A(n5379), .ZN(U2972) );
  NOR2_X1 U6535 ( .A1(n5381), .A2(n3110), .ZN(n6007) );
  INV_X1 U6536 ( .A(n6007), .ZN(n5539) );
  AOI22_X1 U6537 ( .A1(n5383), .A2(DATAI_15_), .B1(n6620), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U6538 ( .B1(n5539), .B2(n5886), .A(n5384), .ZN(U2876) );
  NOR2_X1 U6539 ( .A1(n5381), .A2(n5386), .ZN(n5387) );
  OR2_X1 U6540 ( .A1(n5385), .A2(n5387), .ZN(n5995) );
  INV_X1 U6541 ( .A(n5527), .ZN(n5388) );
  XNOR2_X1 U6542 ( .A(n5535), .B(n5388), .ZN(n5991) );
  OAI22_X1 U6543 ( .A1(n5991), .A2(n5536), .B1(n5389), .B2(n5538), .ZN(n5390)
         );
  INV_X1 U6544 ( .A(n5390), .ZN(n5391) );
  OAI21_X1 U6545 ( .B1(n5995), .B2(n3010), .A(n5391), .ZN(U2843) );
  INV_X1 U6546 ( .A(n5393), .ZN(n5394) );
  XOR2_X1 U6547 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5397), .Z(n5408) );
  INV_X1 U6548 ( .A(n5398), .ZN(n5403) );
  INV_X1 U6549 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6550 ( .A1(n6282), .A2(REIP_REG_30__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6551 ( .A1(n5712), .A2(n5913), .ZN(n5399) );
  OAI211_X1 U6552 ( .C1(n5671), .C2(n5672), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5399), .ZN(n5400) );
  NAND2_X1 U6553 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5404)
         );
  OAI211_X1 U6554 ( .C1(n6202), .C2(n5423), .A(n5405), .B(n5404), .ZN(n5406)
         );
  AOI21_X1 U6555 ( .B1(n5422), .B2(n6184), .A(n5406), .ZN(n5407) );
  OAI21_X1 U6556 ( .B1(n5408), .B2(n6178), .A(n5407), .ZN(U2956) );
  INV_X1 U6557 ( .A(n5789), .ZN(n5409) );
  OAI22_X1 U6558 ( .A1(n3792), .A2(n5409), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5786), .ZN(n6460) );
  OAI22_X1 U6559 ( .A1(n6784), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6592), .ZN(n5410) );
  AOI21_X1 U6560 ( .B1(n6460), .B2(n5411), .A(n5410), .ZN(n5414) );
  AOI21_X1 U6561 ( .B1(n5412), .B2(n5411), .A(n5795), .ZN(n5413) );
  OAI22_X1 U6562 ( .A1(n5414), .A2(n5795), .B1(n5413), .B2(n6463), .ZN(U3461)
         );
  INV_X1 U6563 ( .A(n6212), .ZN(n5416) );
  AOI22_X1 U6564 ( .A1(n6098), .A2(n5416), .B1(REIP_REG_0__SCAN_IN), .B2(n6082), .ZN(n5421) );
  NAND2_X1 U6565 ( .A1(n6075), .A2(n6101), .ZN(n5419) );
  OAI22_X1 U6566 ( .A1(n3642), .A2(n6094), .B1(n6093), .B2(n5417), .ZN(n5418)
         );
  AOI21_X1 U6567 ( .B1(n5419), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5418), 
        .ZN(n5420) );
  OAI211_X1 U6568 ( .C1(n3792), .C2(n6091), .A(n5421), .B(n5420), .ZN(U2827)
         );
  INV_X1 U6569 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5428) );
  NOR3_X1 U6570 ( .A1(n5875), .A2(n5797), .A3(n5428), .ZN(n5426) );
  OAI22_X1 U6571 ( .A1(n5424), .A2(n6075), .B1(n5423), .B2(n6101), .ZN(n5425)
         );
  NOR2_X1 U6572 ( .A1(n5426), .A2(n5425), .ZN(n5430) );
  NAND3_X1 U6573 ( .A1(REIP_REG_29__SCAN_IN), .A2(n5428), .A3(n5427), .ZN(
        n5429) );
  OAI211_X1 U6574 ( .C1(n6094), .C2(n5431), .A(n5430), .B(n5429), .ZN(n5432)
         );
  AOI21_X1 U6575 ( .B1(n5433), .B2(n6067), .A(n5432), .ZN(n5434) );
  OAI21_X1 U6576 ( .B1(n5544), .B2(n6024), .A(n5434), .ZN(U2797) );
  AOI21_X1 U6577 ( .B1(n5437), .B2(n5435), .A(n4289), .ZN(n5589) );
  INV_X1 U6578 ( .A(n5589), .ZN(n5551) );
  OAI22_X1 U6579 ( .A1(n5816), .A2(n6575), .B1(n4192), .B2(n6075), .ZN(n5444)
         );
  NAND2_X1 U6580 ( .A1(n5464), .A2(n5438), .ZN(n5439) );
  NAND2_X1 U6581 ( .A1(n5440), .A2(n5439), .ZN(n5692) );
  NOR2_X1 U6582 ( .A1(n5587), .A2(n6101), .ZN(n5441) );
  AOI21_X1 U6583 ( .B1(n6054), .B2(EBX_REG_27__SCAN_IN), .A(n5441), .ZN(n5442)
         );
  OAI21_X1 U6584 ( .B1(n5692), .B2(n6093), .A(n5442), .ZN(n5443) );
  AOI211_X1 U6585 ( .C1(n5445), .C2(n6575), .A(n5444), .B(n5443), .ZN(n5446)
         );
  OAI21_X1 U6586 ( .B1(n5551), .B2(n6024), .A(n5446), .ZN(U2800) );
  OAI22_X1 U6587 ( .A1(n3731), .A2(n5536), .B1(n5448), .B2(n5538), .ZN(U2828)
         );
  NOR2_X1 U6588 ( .A1(n3101), .A2(n5449), .ZN(n5450) );
  OAI211_X1 U6589 ( .C1(n3651), .C2(n5454), .A(n5453), .B(n5452), .ZN(n5455)
         );
  NAND2_X1 U6590 ( .A1(n5456), .A2(n5455), .ZN(n5803) );
  OAI222_X1 U6591 ( .A1(n3010), .A2(n5804), .B1(n5538), .B2(n5457), .C1(n5803), 
        .C2(n5536), .ZN(U2830) );
  INV_X1 U6592 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5458) );
  OAI222_X1 U6593 ( .A1(n3010), .A2(n5577), .B1(n5538), .B2(n5458), .C1(n5683), 
        .C2(n5536), .ZN(U2831) );
  INV_X1 U6594 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5459) );
  OAI222_X1 U6595 ( .A1(n5459), .A2(n5538), .B1(n5536), .B2(n5692), .C1(n5551), 
        .C2(n3010), .ZN(U2832) );
  INV_X1 U6596 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5465) );
  OR2_X1 U6597 ( .A1(n5472), .A2(n5462), .ZN(n5463) );
  NAND2_X1 U6598 ( .A1(n5464), .A2(n5463), .ZN(n5810) );
  OAI222_X1 U6599 ( .A1(n3010), .A2(n5811), .B1(n5538), .B2(n5465), .C1(n5810), 
        .C2(n5536), .ZN(U2833) );
  NOR2_X1 U6601 ( .A1(n5467), .A2(n5468), .ZN(n5469) );
  OR2_X1 U6602 ( .A1(n5460), .A2(n5469), .ZN(n5821) );
  INV_X1 U6603 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5473) );
  NOR2_X1 U6604 ( .A1(n5476), .A2(n5470), .ZN(n5471) );
  OR2_X1 U6605 ( .A1(n5472), .A2(n5471), .ZN(n5820) );
  OAI222_X1 U6606 ( .A1(n3010), .A2(n5821), .B1(n5538), .B2(n5473), .C1(n5820), 
        .C2(n5536), .ZN(U2834) );
  AOI21_X1 U6607 ( .B1(n5474), .B2(n3029), .A(n5467), .ZN(n5613) );
  INV_X1 U6608 ( .A(n5613), .ZN(n5834) );
  INV_X1 U6609 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5478) );
  AND2_X1 U6610 ( .A1(n5485), .A2(n5475), .ZN(n5477) );
  OR2_X1 U6611 ( .A1(n5477), .A2(n5476), .ZN(n5838) );
  OAI222_X1 U6612 ( .A1(n3010), .A2(n5834), .B1(n5538), .B2(n5478), .C1(n5838), 
        .C2(n5536), .ZN(U2835) );
  NAND2_X1 U6613 ( .A1(n5479), .A2(n5480), .ZN(n5481) );
  NAND2_X1 U6614 ( .A1(n3029), .A2(n5481), .ZN(n5845) );
  INV_X1 U6615 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6616 ( .A1(n5482), .A2(n5483), .ZN(n5484) );
  NAND2_X1 U6617 ( .A1(n5485), .A2(n5484), .ZN(n5844) );
  OAI222_X1 U6618 ( .A1(n3010), .A2(n5845), .B1(n5538), .B2(n5486), .C1(n5844), 
        .C2(n5536), .ZN(U2836) );
  OAI21_X1 U6619 ( .B1(n3030), .B2(n5487), .A(n5479), .ZN(n5851) );
  INV_X1 U6620 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5491) );
  OR2_X1 U6621 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  NAND2_X1 U6622 ( .A1(n5482), .A2(n5490), .ZN(n5852) );
  OAI222_X1 U6623 ( .A1(n3010), .A2(n5851), .B1(n5538), .B2(n5491), .C1(n5852), 
        .C2(n5536), .ZN(U2837) );
  NOR2_X1 U6624 ( .A1(n5492), .A2(n5493), .ZN(n5494) );
  OR2_X1 U6625 ( .A1(n3030), .A2(n5494), .ZN(n5633) );
  XNOR2_X1 U6626 ( .A(n5496), .B(n5495), .ZN(n5865) );
  INV_X1 U6627 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5497) );
  OAI22_X1 U6628 ( .A1(n5865), .A2(n5536), .B1(n5497), .B2(n5538), .ZN(n5498)
         );
  INV_X1 U6629 ( .A(n5498), .ZN(n5499) );
  OAI21_X1 U6630 ( .B1(n5633), .B2(n3010), .A(n5499), .ZN(U2838) );
  AND2_X1 U6631 ( .A1(n5500), .A2(n5501), .ZN(n5502) );
  NOR2_X1 U6632 ( .A1(n5492), .A2(n5502), .ZN(n5890) );
  INV_X1 U6633 ( .A(n5890), .ZN(n5508) );
  INV_X1 U6634 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5507) );
  INV_X1 U6635 ( .A(n5512), .ZN(n5504) );
  MUX2_X1 U6636 ( .A(n5504), .B(n3026), .S(n5503), .Z(n5506) );
  XNOR2_X1 U6637 ( .A(n5506), .B(n5505), .ZN(n5866) );
  OAI222_X1 U6638 ( .A1(n3010), .A2(n5508), .B1(n5538), .B2(n5507), .C1(n5866), 
        .C2(n5536), .ZN(U2839) );
  INV_X1 U6639 ( .A(n5500), .ZN(n5510) );
  AOI21_X1 U6640 ( .B1(n5511), .B2(n5509), .A(n5510), .ZN(n5893) );
  INV_X1 U6641 ( .A(n5893), .ZN(n5517) );
  MUX2_X1 U6642 ( .A(n5512), .B(n5521), .S(n3651), .Z(n5513) );
  NAND2_X1 U6643 ( .A1(n5529), .A2(n5513), .ZN(n5520) );
  XNOR2_X1 U6644 ( .A(n5520), .B(n3057), .ZN(n5761) );
  INV_X1 U6645 ( .A(n5761), .ZN(n5880) );
  AOI22_X1 U6646 ( .A1(n5880), .A2(n5515), .B1(n4864), .B2(EBX_REG_19__SCAN_IN), .ZN(n5516) );
  OAI21_X1 U6647 ( .B1(n5517), .B2(n3010), .A(n5516), .ZN(U2840) );
  OAI21_X1 U6648 ( .B1(n3031), .B2(n5518), .A(n5509), .ZN(n5973) );
  OR2_X1 U6649 ( .A1(n5529), .A2(n5513), .ZN(n5519) );
  NAND2_X1 U6650 ( .A1(n5520), .A2(n5519), .ZN(n5977) );
  OAI22_X1 U6651 ( .A1(n5977), .A2(n5536), .B1(n5521), .B2(n5538), .ZN(n5522)
         );
  INV_X1 U6652 ( .A(n5522), .ZN(n5523) );
  OAI21_X1 U6653 ( .B1(n5973), .B2(n3010), .A(n5523), .ZN(U2841) );
  NOR2_X1 U6654 ( .A1(n5385), .A2(n5524), .ZN(n5525) );
  OR2_X1 U6655 ( .A1(n3031), .A2(n5525), .ZN(n5899) );
  INV_X1 U6656 ( .A(n5535), .ZN(n5528) );
  AOI21_X1 U6657 ( .B1(n5528), .B2(n5527), .A(n5526), .ZN(n5530) );
  OR2_X1 U6658 ( .A1(n5530), .A2(n5529), .ZN(n5985) );
  OAI222_X1 U6659 ( .A1(n3010), .A2(n5899), .B1(n5538), .B2(n5531), .C1(n5536), 
        .C2(n5985), .ZN(U2842) );
  INV_X1 U6660 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U6661 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U6662 ( .A1(n5535), .A2(n5534), .ZN(n5998) );
  OAI222_X1 U6663 ( .A1(n5539), .A2(n3010), .B1(n5538), .B2(n5537), .C1(n5998), 
        .C2(n5536), .ZN(U2844) );
  AOI22_X1 U6664 ( .A1(n6622), .A2(DATAI_30_), .B1(n6620), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5543) );
  AND2_X1 U6665 ( .A1(n3325), .A2(n3335), .ZN(n5540) );
  NAND2_X1 U6666 ( .A1(n6621), .A2(DATAI_14_), .ZN(n5542) );
  OAI211_X1 U6667 ( .C1(n5544), .C2(n5886), .A(n5543), .B(n5542), .ZN(U2861)
         );
  AOI22_X1 U6668 ( .A1(n6621), .A2(DATAI_13_), .B1(n6620), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U6669 ( .A1(n6622), .A2(DATAI_29_), .ZN(n5545) );
  OAI211_X1 U6670 ( .C1(n5804), .C2(n5886), .A(n5546), .B(n5545), .ZN(U2862)
         );
  AOI22_X1 U6671 ( .A1(n6621), .A2(DATAI_12_), .B1(n6620), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6672 ( .A1(n6622), .A2(DATAI_28_), .ZN(n5547) );
  OAI211_X1 U6673 ( .C1(n5577), .C2(n5886), .A(n5548), .B(n5547), .ZN(U2863)
         );
  AOI22_X1 U6674 ( .A1(n6622), .A2(DATAI_27_), .B1(n6620), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U6675 ( .A1(n6621), .A2(DATAI_11_), .ZN(n5549) );
  OAI211_X1 U6676 ( .C1(n5551), .C2(n5886), .A(n5550), .B(n5549), .ZN(U2864)
         );
  AOI22_X1 U6677 ( .A1(n6621), .A2(DATAI_10_), .B1(n6620), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U6678 ( .A1(n6622), .A2(DATAI_26_), .ZN(n5552) );
  OAI211_X1 U6679 ( .C1(n5811), .C2(n5886), .A(n5553), .B(n5552), .ZN(U2865)
         );
  AOI22_X1 U6680 ( .A1(n6621), .A2(DATAI_9_), .B1(n6620), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U6681 ( .A1(n6622), .A2(DATAI_25_), .ZN(n5554) );
  OAI211_X1 U6682 ( .C1(n5821), .C2(n5886), .A(n5555), .B(n5554), .ZN(U2866)
         );
  AOI22_X1 U6683 ( .A1(n6621), .A2(DATAI_8_), .B1(n6620), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U6684 ( .A1(n6622), .A2(DATAI_24_), .ZN(n5556) );
  OAI211_X1 U6685 ( .C1(n5834), .C2(n5886), .A(n5557), .B(n5556), .ZN(U2867)
         );
  AOI22_X1 U6686 ( .A1(n6621), .A2(DATAI_7_), .B1(n6620), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U6687 ( .A1(n6622), .A2(DATAI_23_), .ZN(n5558) );
  OAI211_X1 U6688 ( .C1(n5845), .C2(n5886), .A(n5559), .B(n5558), .ZN(U2868)
         );
  AOI22_X1 U6689 ( .A1(n6622), .A2(DATAI_18_), .B1(n6620), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6690 ( .A1(n6621), .A2(DATAI_2_), .ZN(n5560) );
  OAI211_X1 U6691 ( .C1(n5973), .C2(n5886), .A(n5561), .B(n5560), .ZN(U2873)
         );
  INV_X1 U6692 ( .A(n5562), .ZN(n5563) );
  AOI21_X1 U6693 ( .B1(n5564), .B2(n5392), .A(n5563), .ZN(n5565) );
  XNOR2_X1 U6694 ( .A(n5565), .B(n5672), .ZN(n5678) );
  INV_X1 U6695 ( .A(n5804), .ZN(n5568) );
  NAND2_X1 U6696 ( .A1(n6282), .A2(REIP_REG_29__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U6697 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5566)
         );
  OAI211_X1 U6698 ( .C1(n6202), .C2(n5799), .A(n5669), .B(n5566), .ZN(n5567)
         );
  AOI21_X1 U6699 ( .B1(n5568), .B2(n6184), .A(n5567), .ZN(n5569) );
  OAI21_X1 U6700 ( .B1(n5678), .B2(n6178), .A(n5569), .ZN(U2957) );
  INV_X1 U6701 ( .A(n5392), .ZN(n5594) );
  NAND3_X1 U6702 ( .A1(n5594), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5650), .ZN(n5574) );
  INV_X1 U6703 ( .A(n5592), .ZN(n5572) );
  INV_X1 U6704 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5571) );
  NAND3_X1 U6705 ( .A1(n5570), .A2(n5572), .A3(n5571), .ZN(n5582) );
  INV_X1 U6706 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5573) );
  AOI22_X1 U6707 ( .A1(n5574), .A2(n5582), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5573), .ZN(n5575) );
  XNOR2_X1 U6708 ( .A(n5575), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5688)
         );
  NAND2_X1 U6709 ( .A1(n6282), .A2(REIP_REG_28__SCAN_IN), .ZN(n5682) );
  OAI21_X1 U6710 ( .B1(n5903), .B2(n5576), .A(n5682), .ZN(n5579) );
  NOR2_X1 U6711 ( .A1(n5577), .A2(n6211), .ZN(n5578) );
  OAI21_X1 U6712 ( .B1(n6178), .B2(n5688), .A(n5581), .ZN(U2958) );
  INV_X1 U6713 ( .A(n5582), .ZN(n5583) );
  NOR2_X1 U6714 ( .A1(n5584), .A2(n5583), .ZN(n5585) );
  XNOR2_X1 U6715 ( .A(n5585), .B(n5694), .ZN(n5697) );
  NAND2_X1 U6716 ( .A1(n6282), .A2(REIP_REG_27__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U6717 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5586)
         );
  OAI211_X1 U6718 ( .C1(n6202), .C2(n5587), .A(n5691), .B(n5586), .ZN(n5588)
         );
  AOI21_X1 U6719 ( .B1(n5589), .B2(n6184), .A(n5588), .ZN(n5590) );
  OAI21_X1 U6720 ( .B1(n5697), .B2(n6178), .A(n5590), .ZN(U2959) );
  NAND2_X1 U6721 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  XNOR2_X1 U6722 ( .A(n5594), .B(n5593), .ZN(n5703) );
  NAND2_X1 U6723 ( .A1(n6282), .A2(REIP_REG_26__SCAN_IN), .ZN(n5698) );
  OAI21_X1 U6724 ( .B1(n5903), .B2(n5595), .A(n5698), .ZN(n5597) );
  NOR2_X1 U6725 ( .A1(n5811), .A2(n6211), .ZN(n5596) );
  AOI211_X1 U6726 ( .C1(n6173), .C2(n5808), .A(n5597), .B(n5596), .ZN(n5598)
         );
  OAI21_X1 U6727 ( .B1(n5703), .B2(n6178), .A(n5598), .ZN(U2960) );
  OAI21_X1 U6728 ( .B1(n5570), .B2(n5599), .A(n3549), .ZN(n5600) );
  INV_X1 U6729 ( .A(n5600), .ZN(n5710) );
  INV_X1 U6730 ( .A(n5821), .ZN(n5604) );
  NOR2_X1 U6731 ( .A1(n6202), .A2(n5818), .ZN(n5603) );
  NAND2_X1 U6732 ( .A1(n6282), .A2(REIP_REG_25__SCAN_IN), .ZN(n5704) );
  OAI21_X1 U6733 ( .B1(n5903), .B2(n5601), .A(n5704), .ZN(n5602) );
  AOI211_X1 U6734 ( .C1(n5604), .C2(n6184), .A(n5603), .B(n5602), .ZN(n5605)
         );
  OAI21_X1 U6735 ( .B1(n5710), .B2(n6178), .A(n5605), .ZN(U2961) );
  AOI21_X1 U6736 ( .B1(n3033), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5645), 
        .ZN(n5606) );
  OR2_X2 U6737 ( .A1(n5606), .A2(n5643), .ZN(n5638) );
  XNOR2_X1 U6738 ( .A(n5650), .B(n5607), .ZN(n5637) );
  OAI22_X1 U6739 ( .A1(n5638), .A2(n5637), .B1(n5650), .B2(n5607), .ZN(n5631)
         );
  INV_X1 U6740 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5738) );
  XNOR2_X1 U6741 ( .A(n5650), .B(n5738), .ZN(n5632) );
  INV_X1 U6742 ( .A(n5608), .ZN(n5630) );
  NOR2_X1 U6743 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5623)
         );
  NAND2_X1 U6744 ( .A1(n5630), .A2(n5623), .ZN(n5615) );
  OAI21_X1 U6745 ( .B1(n5645), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5608), 
        .ZN(n5625) );
  NAND3_X1 U6746 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5609) );
  XNOR2_X1 U6747 ( .A(n5610), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5719)
         );
  NAND2_X1 U6748 ( .A1(n6273), .A2(REIP_REG_24__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6749 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5611)
         );
  OAI211_X1 U6750 ( .C1(n6202), .C2(n5828), .A(n5711), .B(n5611), .ZN(n5612)
         );
  AOI21_X1 U6751 ( .B1(n5613), .B2(n6184), .A(n5612), .ZN(n5614) );
  OAI21_X1 U6752 ( .B1(n5719), .B2(n6178), .A(n5614), .ZN(U2962) );
  NAND3_X1 U6753 ( .A1(n5650), .A2(n3544), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5616) );
  OAI21_X1 U6754 ( .B1(n5638), .B2(n5616), .A(n5615), .ZN(n5617) );
  XNOR2_X1 U6755 ( .A(n5617), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5726)
         );
  NAND2_X1 U6756 ( .A1(n6282), .A2(REIP_REG_23__SCAN_IN), .ZN(n5720) );
  OAI21_X1 U6757 ( .B1(n5903), .B2(n5618), .A(n5720), .ZN(n5620) );
  NOR2_X1 U6758 ( .A1(n5845), .A2(n6211), .ZN(n5619) );
  AOI211_X1 U6759 ( .C1(n6173), .C2(n5621), .A(n5620), .B(n5619), .ZN(n5622)
         );
  OAI21_X1 U6760 ( .B1(n5726), .B2(n6178), .A(n5622), .ZN(U2963) );
  AOI21_X1 U6761 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5650), .A(n5623), 
        .ZN(n5624) );
  XNOR2_X1 U6762 ( .A(n5625), .B(n5624), .ZN(n5733) );
  NAND2_X1 U6763 ( .A1(n6282), .A2(REIP_REG_22__SCAN_IN), .ZN(n5727) );
  OAI21_X1 U6764 ( .B1(n5903), .B2(n5626), .A(n5727), .ZN(n5628) );
  NOR2_X1 U6765 ( .A1(n5851), .A2(n6211), .ZN(n5627) );
  AOI211_X1 U6766 ( .C1(n6173), .C2(n5850), .A(n5628), .B(n5627), .ZN(n5629)
         );
  OAI21_X1 U6767 ( .B1(n5733), .B2(n6178), .A(n5629), .ZN(U2964) );
  AOI21_X1 U6768 ( .B1(n5632), .B2(n5631), .A(n5630), .ZN(n5741) );
  NAND2_X1 U6769 ( .A1(n6282), .A2(REIP_REG_21__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U6770 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5634)
         );
  OAI211_X1 U6771 ( .C1(n6202), .C2(n5860), .A(n5735), .B(n5634), .ZN(n5635)
         );
  AOI21_X1 U6772 ( .B1(n6624), .B2(n6184), .A(n5635), .ZN(n5636) );
  OAI21_X1 U6773 ( .B1(n5741), .B2(n6178), .A(n5636), .ZN(U2965) );
  XNOR2_X1 U6774 ( .A(n5638), .B(n5637), .ZN(n5759) );
  NAND2_X1 U6775 ( .A1(n6173), .A2(n5870), .ZN(n5639) );
  NAND2_X1 U6776 ( .A1(n6282), .A2(REIP_REG_20__SCAN_IN), .ZN(n5746) );
  OAI211_X1 U6777 ( .C1(n5903), .C2(n5640), .A(n5639), .B(n5746), .ZN(n5641)
         );
  AOI21_X1 U6778 ( .B1(n5890), .B2(n6184), .A(n5641), .ZN(n5642) );
  OAI21_X1 U6779 ( .B1(n5759), .B2(n6178), .A(n5642), .ZN(U2966) );
  AOI21_X1 U6780 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5644), .A(n5643), 
        .ZN(n5646) );
  XNOR2_X1 U6781 ( .A(n5646), .B(n5645), .ZN(n5768) );
  NAND2_X1 U6782 ( .A1(n6282), .A2(REIP_REG_19__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U6783 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5647)
         );
  OAI211_X1 U6784 ( .C1(n6202), .C2(n5878), .A(n5760), .B(n5647), .ZN(n5648)
         );
  AOI21_X1 U6785 ( .B1(n5893), .B2(n6184), .A(n5648), .ZN(n5649) );
  OAI21_X1 U6786 ( .B1(n5768), .B2(n6178), .A(n5649), .ZN(U2967) );
  NAND2_X1 U6787 ( .A1(n6282), .A2(REIP_REG_18__SCAN_IN), .ZN(n5774) );
  AND2_X1 U6788 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5897)
         );
  NAND2_X1 U6789 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5897), .ZN(n5653) );
  NOR2_X1 U6790 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5896)
         );
  NAND3_X1 U6791 ( .A1(n5896), .A2(n5908), .A3(n5651), .ZN(n5652) );
  OAI21_X1 U6792 ( .B1(n5653), .B2(n5651), .A(n5652), .ZN(n5654) );
  XOR2_X1 U6793 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5654), .Z(n5776) );
  NAND2_X1 U6794 ( .A1(n6206), .A2(n5776), .ZN(n5655) );
  OAI211_X1 U6795 ( .C1(n5903), .C2(n5971), .A(n5774), .B(n5655), .ZN(n5656)
         );
  AOI21_X1 U6796 ( .B1(n6173), .B2(n5969), .A(n5656), .ZN(n5657) );
  OAI21_X1 U6797 ( .B1(n5973), .B2(n6211), .A(n5657), .ZN(U2968) );
  NOR2_X1 U6798 ( .A1(n5896), .A2(n5897), .ZN(n5658) );
  XNOR2_X1 U6799 ( .A(n5651), .B(n5658), .ZN(n5915) );
  INV_X1 U6800 ( .A(n5995), .ZN(n6105) );
  INV_X1 U6801 ( .A(n5987), .ZN(n5660) );
  AOI22_X1 U6802 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6273), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5659) );
  OAI21_X1 U6803 ( .B1(n5660), .B2(n6202), .A(n5659), .ZN(n5661) );
  AOI21_X1 U6804 ( .B1(n6105), .B2(n6184), .A(n5661), .ZN(n5662) );
  OAI21_X1 U6805 ( .B1(n5915), .B2(n6178), .A(n5662), .ZN(U2970) );
  XNOR2_X1 U6806 ( .A(n5650), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5664)
         );
  XNOR2_X1 U6807 ( .A(n5663), .B(n5664), .ZN(n5924) );
  INV_X1 U6808 ( .A(n6000), .ZN(n5666) );
  AOI22_X1 U6809 ( .A1(n6208), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6282), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5665) );
  OAI21_X1 U6810 ( .B1(n5666), .B2(n6202), .A(n5665), .ZN(n5667) );
  AOI21_X1 U6811 ( .B1(n6007), .B2(n6184), .A(n5667), .ZN(n5668) );
  OAI21_X1 U6812 ( .B1(n5924), .B2(n6178), .A(n5668), .ZN(U2971) );
  INV_X1 U6813 ( .A(n5669), .ZN(n5670) );
  AOI21_X1 U6814 ( .B1(n5671), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5670), 
        .ZN(n5675) );
  NAND3_X1 U6815 ( .A1(n5695), .A2(n5673), .A3(n5672), .ZN(n5674) );
  OAI211_X1 U6816 ( .C1(n5803), .C2(n6304), .A(n5675), .B(n5674), .ZN(n5676)
         );
  INV_X1 U6817 ( .A(n5676), .ZN(n5677) );
  OAI21_X1 U6818 ( .B1(n5678), .B2(n6224), .A(n5677), .ZN(U2989) );
  NAND2_X1 U6819 ( .A1(n6260), .A2(n5679), .ZN(n5680) );
  NAND2_X1 U6820 ( .A1(n5712), .A2(n5680), .ZN(n5689) );
  NAND2_X1 U6821 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5681) );
  OAI211_X1 U6822 ( .C1(n5683), .C2(n6304), .A(n5682), .B(n5681), .ZN(n5684)
         );
  INV_X1 U6823 ( .A(n5684), .ZN(n5687) );
  NAND3_X1 U6824 ( .A1(n5695), .A2(n5685), .A3(n3083), .ZN(n5686) );
  OAI211_X1 U6825 ( .C1(n5688), .C2(n6224), .A(n5687), .B(n5686), .ZN(U2990)
         );
  NAND2_X1 U6826 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5690) );
  OAI211_X1 U6827 ( .C1(n5692), .C2(n6304), .A(n5691), .B(n5690), .ZN(n5693)
         );
  AOI21_X1 U6828 ( .B1(n5695), .B2(n5694), .A(n5693), .ZN(n5696) );
  OAI21_X1 U6829 ( .B1(n5697), .B2(n6224), .A(n5696), .ZN(U2991) );
  INV_X1 U6830 ( .A(n5712), .ZN(n5708) );
  OAI21_X1 U6831 ( .B1(n5810), .B2(n6304), .A(n5698), .ZN(n5701) );
  XNOR2_X1 U6832 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5699) );
  NOR2_X1 U6833 ( .A1(n5705), .A2(n5699), .ZN(n5700) );
  AOI211_X1 U6834 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5708), .A(n5701), .B(n5700), .ZN(n5702) );
  OAI21_X1 U6835 ( .B1(n5703), .B2(n6224), .A(n5702), .ZN(U2992) );
  OAI21_X1 U6836 ( .B1(n5820), .B2(n6304), .A(n5704), .ZN(n5707) );
  NOR2_X1 U6837 ( .A1(n5705), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5706)
         );
  AOI211_X1 U6838 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5708), .A(n5707), .B(n5706), .ZN(n5709) );
  OAI21_X1 U6839 ( .B1(n5710), .B2(n6224), .A(n5709), .ZN(U2993) );
  INV_X1 U6840 ( .A(n5838), .ZN(n5717) );
  INV_X1 U6841 ( .A(n5711), .ZN(n5716) );
  INV_X1 U6842 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5714) );
  AOI211_X1 U6843 ( .C1(n5714), .C2(n5721), .A(n5713), .B(n5712), .ZN(n5715)
         );
  AOI211_X1 U6844 ( .C1(n6290), .C2(n5717), .A(n5716), .B(n5715), .ZN(n5718)
         );
  OAI21_X1 U6845 ( .B1(n5719), .B2(n6224), .A(n5718), .ZN(U2994) );
  OAI21_X1 U6846 ( .B1(n5844), .B2(n6304), .A(n5720), .ZN(n5723) );
  NOR2_X1 U6847 ( .A1(n5721), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5722)
         );
  AOI211_X1 U6848 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5724), .A(n5723), .B(n5722), .ZN(n5725) );
  OAI21_X1 U6849 ( .B1(n5726), .B2(n6224), .A(n5725), .ZN(U2995) );
  OAI21_X1 U6850 ( .B1(n5852), .B2(n6304), .A(n5727), .ZN(n5731) );
  INV_X1 U6851 ( .A(n5739), .ZN(n5729) );
  NOR3_X1 U6852 ( .A1(n5729), .A2(n5728), .A3(n3544), .ZN(n5730) );
  AOI211_X1 U6853 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5734), .A(n5731), .B(n5730), .ZN(n5732) );
  OAI21_X1 U6854 ( .B1(n5733), .B2(n6224), .A(n5732), .ZN(U2996) );
  NAND2_X1 U6855 ( .A1(n5734), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5736) );
  OAI211_X1 U6856 ( .C1(n6304), .C2(n5865), .A(n5736), .B(n5735), .ZN(n5737)
         );
  AOI21_X1 U6857 ( .B1(n5739), .B2(n5738), .A(n5737), .ZN(n5740) );
  OAI21_X1 U6858 ( .B1(n5741), .B2(n6224), .A(n5740), .ZN(U2997) );
  INV_X1 U6859 ( .A(n5742), .ZN(n5743) );
  NOR2_X1 U6860 ( .A1(n5904), .A2(n5743), .ZN(n5764) );
  OAI21_X1 U6861 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5744), .ZN(n5745) );
  INV_X1 U6862 ( .A(n5745), .ZN(n5748) );
  OAI21_X1 U6863 ( .B1(n5866), .B2(n6304), .A(n5746), .ZN(n5747) );
  AOI21_X1 U6864 ( .B1(n5764), .B2(n5748), .A(n5747), .ZN(n5758) );
  NAND2_X1 U6865 ( .A1(n5749), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U6866 ( .A1(n5751), .A2(n5750), .ZN(n5753) );
  NAND2_X1 U6867 ( .A1(n5753), .A2(n5752), .ZN(n5907) );
  AND2_X1 U6868 ( .A1(n6297), .A2(n5908), .ZN(n5754) );
  NOR2_X1 U6869 ( .A1(n5907), .A2(n5754), .ZN(n5769) );
  NAND2_X1 U6870 ( .A1(n6260), .A2(n5755), .ZN(n5756) );
  NAND2_X1 U6871 ( .A1(n5769), .A2(n5756), .ZN(n5765) );
  NAND2_X1 U6872 ( .A1(n5765), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5757) );
  OAI211_X1 U6873 ( .C1(n5759), .C2(n6224), .A(n5758), .B(n5757), .ZN(U2998)
         );
  OAI21_X1 U6874 ( .B1(n5761), .B2(n6304), .A(n5760), .ZN(n5762) );
  AOI21_X1 U6875 ( .B1(n5764), .B2(n5763), .A(n5762), .ZN(n5767) );
  NAND2_X1 U6876 ( .A1(n5765), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5766) );
  OAI211_X1 U6877 ( .C1(n5768), .C2(n6224), .A(n5767), .B(n5766), .ZN(U2999)
         );
  NOR2_X1 U6878 ( .A1(n5908), .A2(n5904), .ZN(n5771) );
  INV_X1 U6879 ( .A(n5769), .ZN(n5770) );
  MUX2_X1 U6880 ( .A(n5771), .B(n5770), .S(INSTADDRPOINTER_REG_18__SCAN_IN), 
        .Z(n5772) );
  INV_X1 U6881 ( .A(n5772), .ZN(n5773) );
  NAND2_X1 U6882 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  AOI21_X1 U6883 ( .B1(n6307), .B2(n5776), .A(n5775), .ZN(n5777) );
  OAI21_X1 U6884 ( .B1(n5977), .B2(n6304), .A(n5777), .ZN(U3000) );
  OAI21_X1 U6885 ( .B1(n5778), .B2(STATEBS16_REG_SCAN_IN), .A(n6367), .ZN(
        n5779) );
  OAI22_X1 U6886 ( .A1(n5779), .A2(n5781), .B1(n6090), .B2(n5782), .ZN(n5780)
         );
  MUX2_X1 U6887 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5780), .S(n6312), 
        .Z(U3464) );
  XNOR2_X1 U6888 ( .A(n4368), .B(n5781), .ZN(n5783) );
  INV_X1 U6889 ( .A(n4374), .ZN(n6076) );
  OAI22_X1 U6890 ( .A1(n5783), .A2(n6316), .B1(n6076), .B2(n5782), .ZN(n5784)
         );
  MUX2_X1 U6891 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5784), .S(n6312), 
        .Z(U3463) );
  INV_X1 U6892 ( .A(n5785), .ZN(n5788) );
  NOR3_X1 U6893 ( .A1(n5786), .A2(n4446), .A3(n4606), .ZN(n5787) );
  INV_X1 U6894 ( .A(n4606), .ZN(n5792) );
  AOI22_X1 U6895 ( .A1(n5793), .A2(n5792), .B1(n5791), .B2(n5790), .ZN(n5794)
         );
  OAI21_X1 U6896 ( .B1(n6464), .B2(n6594), .A(n5794), .ZN(n5796) );
  MUX2_X1 U6897 ( .A(n5796), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n5795), 
        .Z(U3460) );
  AND2_X1 U6898 ( .A1(n6139), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6899 ( .B1(n6580), .B2(n5798), .A(n5797), .ZN(n5802) );
  INV_X1 U6900 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5800) );
  OAI22_X1 U6901 ( .A1(n5800), .A2(n6075), .B1(n5799), .B2(n6101), .ZN(n5801)
         );
  AOI211_X1 U6902 ( .C1(n6054), .C2(EBX_REG_29__SCAN_IN), .A(n5802), .B(n5801), 
        .ZN(n5807) );
  OAI22_X1 U6903 ( .A1(n5804), .A2(n6024), .B1(n5803), .B2(n6093), .ZN(n5805)
         );
  INV_X1 U6904 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U6905 ( .A1(n5807), .A2(n5806), .ZN(U2798) );
  AOI22_X1 U6906 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6087), .B1(n5808), 
        .B2(n6062), .ZN(n5809) );
  INV_X1 U6907 ( .A(n5809), .ZN(n5813) );
  OAI22_X1 U6908 ( .A1(n5811), .A2(n6024), .B1(n5810), .B2(n6093), .ZN(n5812)
         );
  AOI211_X1 U6909 ( .C1(EBX_REG_26__SCAN_IN), .C2(n6054), .A(n5813), .B(n5812), 
        .ZN(n5814) );
  OAI221_X1 U6910 ( .B1(n5816), .B2(n6572), .C1(n5816), .C2(n5815), .A(n5814), 
        .ZN(U2801) );
  AOI22_X1 U6911 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6054), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6087), .ZN(n5827) );
  INV_X1 U6912 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5817) );
  INV_X1 U6913 ( .A(n5831), .ZN(n5839) );
  OAI22_X1 U6914 ( .A1(n5818), .A2(n6101), .B1(n5817), .B2(n5839), .ZN(n5819)
         );
  INV_X1 U6915 ( .A(n5819), .ZN(n5826) );
  OAI22_X1 U6916 ( .A1(n5821), .A2(n6024), .B1(n5820), .B2(n6093), .ZN(n5822)
         );
  INV_X1 U6917 ( .A(n5822), .ZN(n5825) );
  OAI211_X1 U6918 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5836), .B(n5823), .ZN(n5824) );
  NAND4_X1 U6919 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(U2802)
         );
  INV_X1 U6920 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6570) );
  OAI22_X1 U6921 ( .A1(n5829), .A2(n6075), .B1(n6101), .B2(n5828), .ZN(n5830)
         );
  AOI21_X1 U6922 ( .B1(EBX_REG_24__SCAN_IN), .B2(n6054), .A(n5830), .ZN(n5833)
         );
  NAND2_X1 U6923 ( .A1(n5831), .A2(REIP_REG_24__SCAN_IN), .ZN(n5832) );
  OAI211_X1 U6924 ( .C1(n5834), .C2(n6024), .A(n5833), .B(n5832), .ZN(n5835)
         );
  AOI21_X1 U6925 ( .B1(n5836), .B2(n6570), .A(n5835), .ZN(n5837) );
  OAI21_X1 U6926 ( .B1(n5838), .B2(n6093), .A(n5837), .ZN(U2803) );
  AOI21_X1 U6927 ( .B1(n6568), .B2(n5840), .A(n5839), .ZN(n5843) );
  OAI22_X1 U6928 ( .A1(n5618), .A2(n6075), .B1(n5841), .B2(n6101), .ZN(n5842)
         );
  AOI211_X1 U6929 ( .C1(n6054), .C2(EBX_REG_23__SCAN_IN), .A(n5843), .B(n5842), 
        .ZN(n5848) );
  OAI22_X1 U6930 ( .A1(n5845), .A2(n6024), .B1(n5844), .B2(n6093), .ZN(n5846)
         );
  INV_X1 U6931 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U6932 ( .A1(n5848), .A2(n5847), .ZN(U2804) );
  AOI22_X1 U6933 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6054), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6087), .ZN(n5858) );
  AND2_X1 U6934 ( .A1(n6082), .A2(n5849), .ZN(n5868) );
  AOI22_X1 U6935 ( .A1(n5850), .A2(n6062), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5868), .ZN(n5857) );
  INV_X1 U6936 ( .A(n5851), .ZN(n5887) );
  INV_X1 U6937 ( .A(n5852), .ZN(n5853) );
  AOI22_X1 U6938 ( .A1(n5887), .A2(n4331), .B1(n5853), .B2(n6067), .ZN(n5856)
         );
  OAI211_X1 U6939 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5862), .B(n5854), .ZN(n5855) );
  NAND4_X1 U6940 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(U2805)
         );
  INV_X1 U6941 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6564) );
  AOI22_X1 U6942 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6054), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6087), .ZN(n5859) );
  OAI21_X1 U6943 ( .B1(n5860), .B2(n6101), .A(n5859), .ZN(n5861) );
  AOI221_X1 U6944 ( .B1(n5868), .B2(REIP_REG_21__SCAN_IN), .C1(n5862), .C2(
        n6564), .A(n5861), .ZN(n5864) );
  NAND2_X1 U6945 ( .A1(n6624), .A2(n4331), .ZN(n5863) );
  OAI211_X1 U6946 ( .C1(n6093), .C2(n5865), .A(n5864), .B(n5863), .ZN(U2806)
         );
  AOI22_X1 U6947 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6054), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6087), .ZN(n5874) );
  INV_X1 U6948 ( .A(n5866), .ZN(n5867) );
  AOI22_X1 U6949 ( .A1(n5890), .A2(n4331), .B1(n5867), .B2(n6067), .ZN(n5873)
         );
  OAI21_X1 U6950 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5869), .A(n5868), .ZN(n5872) );
  NAND2_X1 U6951 ( .A1(n5870), .A2(n6062), .ZN(n5871) );
  NAND4_X1 U6952 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(U2807)
         );
  NOR2_X1 U6953 ( .A1(n5876), .A2(n5875), .ZN(n5982) );
  AOI22_X1 U6954 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6054), .B1(
        REIP_REG_19__SCAN_IN), .B2(n5982), .ZN(n5877) );
  OAI21_X1 U6955 ( .B1(n5878), .B2(n6101), .A(n5877), .ZN(n5879) );
  AOI211_X1 U6956 ( .C1(n6087), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6273), 
        .B(n5879), .ZN(n5885) );
  AOI22_X1 U6957 ( .A1(n5893), .A2(n4331), .B1(n6067), .B2(n5880), .ZN(n5884)
         );
  NAND2_X1 U6958 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5881) );
  OAI211_X1 U6959 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5882), .B(n5881), .ZN(n5883) );
  NAND3_X1 U6960 ( .A1(n5885), .A2(n5884), .A3(n5883), .ZN(U2808) );
  AOI22_X1 U6961 ( .A1(n5887), .A2(n6623), .B1(n6622), .B2(DATAI_22_), .ZN(
        n5889) );
  AOI22_X1 U6962 ( .A1(n6621), .A2(DATAI_6_), .B1(n6620), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U6963 ( .A1(n5889), .A2(n5888), .ZN(U2869) );
  AOI22_X1 U6964 ( .A1(n5890), .A2(n6623), .B1(n6622), .B2(DATAI_20_), .ZN(
        n5892) );
  AOI22_X1 U6965 ( .A1(n6621), .A2(DATAI_4_), .B1(n6620), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U6966 ( .A1(n5892), .A2(n5891), .ZN(U2871) );
  AOI22_X1 U6967 ( .A1(n5893), .A2(n6623), .B1(n6622), .B2(DATAI_19_), .ZN(
        n5895) );
  AOI22_X1 U6968 ( .A1(n6621), .A2(DATAI_3_), .B1(n6620), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6969 ( .A1(n5895), .A2(n5894), .ZN(U2872) );
  INV_X1 U6970 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5979) );
  MUX2_X1 U6971 ( .A(n5897), .B(n5896), .S(n5651), .Z(n5898) );
  XNOR2_X1 U6972 ( .A(n5898), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5911)
         );
  INV_X1 U6973 ( .A(n5911), .ZN(n5901) );
  AOI222_X1 U6974 ( .A1(n5901), .A2(n6206), .B1(n6184), .B2(n6102), .C1(n5900), 
        .C2(n6173), .ZN(n5902) );
  NAND2_X1 U6975 ( .A1(n6282), .A2(REIP_REG_17__SCAN_IN), .ZN(n5905) );
  OAI211_X1 U6976 ( .C1(n5979), .C2(n5903), .A(n5902), .B(n5905), .ZN(U2969)
         );
  INV_X1 U6977 ( .A(n5904), .ZN(n5909) );
  OAI21_X1 U6978 ( .B1(n5985), .B2(n6304), .A(n5905), .ZN(n5906) );
  AOI221_X1 U6979 ( .B1(n5909), .B2(n5908), .C1(n5907), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5906), .ZN(n5910) );
  OAI21_X1 U6980 ( .B1(n5911), .B2(n6224), .A(n5910), .ZN(U3001) );
  OAI21_X1 U6981 ( .B1(n5913), .B2(n5917), .A(n5912), .ZN(n5914) );
  INV_X1 U6982 ( .A(n5914), .ZN(n5931) );
  INV_X1 U6983 ( .A(n5915), .ZN(n5921) );
  INV_X1 U6984 ( .A(n5916), .ZN(n6214) );
  NAND2_X1 U6985 ( .A1(n5917), .A2(n6214), .ZN(n5925) );
  AOI221_X1 U6986 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5930), .C2(n5923), .A(n5925), 
        .ZN(n5918) );
  AOI21_X1 U6987 ( .B1(n6273), .B2(REIP_REG_16__SCAN_IN), .A(n5918), .ZN(n5919) );
  OAI21_X1 U6988 ( .B1(n5991), .B2(n6304), .A(n5919), .ZN(n5920) );
  AOI21_X1 U6989 ( .B1(n5921), .B2(n6307), .A(n5920), .ZN(n5922) );
  OAI21_X1 U6990 ( .B1(n5931), .B2(n5923), .A(n5922), .ZN(U3002) );
  INV_X1 U6991 ( .A(n5924), .ZN(n5928) );
  NOR2_X1 U6992 ( .A1(n5925), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5927)
         );
  OAI22_X1 U6993 ( .A1(n6304), .A2(n5998), .B1(n6553), .B2(n6302), .ZN(n5926)
         );
  AOI211_X1 U6994 ( .C1(n5928), .C2(n6307), .A(n5927), .B(n5926), .ZN(n5929)
         );
  OAI21_X1 U6995 ( .B1(n5931), .B2(n5930), .A(n5929), .ZN(U3003) );
  INV_X1 U6996 ( .A(n5932), .ZN(n5946) );
  NAND2_X1 U6997 ( .A1(n5933), .A2(n5940), .ZN(n5945) );
  INV_X1 U6998 ( .A(n5934), .ZN(n5935) );
  AOI21_X1 U6999 ( .B1(n5936), .B2(n6290), .A(n5935), .ZN(n5944) );
  INV_X1 U7000 ( .A(n5937), .ZN(n5942) );
  AOI21_X1 U7001 ( .B1(n5940), .B2(n5939), .A(n5938), .ZN(n5941) );
  AOI21_X1 U7002 ( .B1(n5942), .B2(n6307), .A(n5941), .ZN(n5943) );
  OAI211_X1 U7003 ( .C1(n5946), .C2(n5945), .A(n5944), .B(n5943), .ZN(U3005)
         );
  AND2_X1 U7004 ( .A1(n6803), .A2(STATE_REG_1__SCAN_IN), .ZN(n6559) );
  INV_X1 U7005 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6641) );
  INV_X1 U7006 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6521) );
  AOI221_X1 U7007 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n6521), .C2(STATE_REG_0__SCAN_IN), .A(n6559), .ZN(n6588) );
  OAI21_X1 U7008 ( .B1(n6559), .B2(n6641), .A(n6513), .ZN(U2789) );
  INV_X1 U7009 ( .A(n5947), .ZN(n5950) );
  OAI21_X1 U7010 ( .B1(n5948), .B2(n6501), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5949) );
  OAI21_X1 U7011 ( .B1(n5950), .B2(n6506), .A(n5949), .ZN(U2790) );
  INV_X2 U7012 ( .A(n6559), .ZN(n6619) );
  NOR2_X1 U7013 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5952) );
  OAI21_X1 U7014 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5952), .A(n6619), .ZN(n5951)
         );
  OAI21_X1 U7015 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6619), .A(n5951), .ZN(
        U2791) );
  OAI21_X1 U7016 ( .B1(BS16_N), .B2(n5952), .A(n6588), .ZN(n6586) );
  OAI21_X1 U7017 ( .B1(n6588), .B2(n6365), .A(n6586), .ZN(U2792) );
  OAI21_X1 U7018 ( .B1(n5954), .B2(n5953), .A(n6178), .ZN(U2793) );
  NOR4_X1 U7019 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5958) );
  NOR4_X1 U7020 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5957) );
  NOR4_X1 U7021 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5956) );
  NOR4_X1 U7022 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n5955) );
  NAND4_X1 U7023 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n5964)
         );
  NOR4_X1 U7024 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n5962) );
  AOI211_X1 U7025 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_28__SCAN_IN), .B(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n5961) );
  NOR4_X1 U7026 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n5960) );
  NOR4_X1 U7027 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n5959) );
  NAND4_X1 U7028 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n5963)
         );
  NOR2_X1 U7029 ( .A1(n5964), .A2(n5963), .ZN(n6603) );
  INV_X1 U7030 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6670) );
  NOR3_X1 U7031 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5966) );
  OAI21_X1 U7032 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5966), .A(n6603), .ZN(n5965)
         );
  OAI21_X1 U7033 ( .B1(n6603), .B2(n6670), .A(n5965), .ZN(U2794) );
  INV_X1 U7034 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6587) );
  AOI21_X1 U7035 ( .B1(n6599), .B2(n6587), .A(n5966), .ZN(n5968) );
  INV_X1 U7036 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5967) );
  INV_X1 U7037 ( .A(n6603), .ZN(n6606) );
  AOI22_X1 U7038 ( .A1(n6603), .A2(n5968), .B1(n5967), .B2(n6606), .ZN(U2795)
         );
  AOI22_X1 U7039 ( .A1(n5969), .A2(n6062), .B1(REIP_REG_18__SCAN_IN), .B2(
        n5982), .ZN(n5970) );
  OAI211_X1 U7040 ( .C1(n6075), .C2(n5971), .A(n5970), .B(n6302), .ZN(n5975)
         );
  OAI22_X1 U7041 ( .A1(n5973), .A2(n6024), .B1(REIP_REG_18__SCAN_IN), .B2(
        n5972), .ZN(n5974) );
  AOI211_X1 U7042 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6054), .A(n5975), .B(n5974), 
        .ZN(n5976) );
  OAI21_X1 U7043 ( .B1(n6093), .B2(n5977), .A(n5976), .ZN(U2809) );
  OAI22_X1 U7044 ( .A1(n5979), .A2(n6075), .B1(n5978), .B2(n6101), .ZN(n5980)
         );
  AOI211_X1 U7045 ( .C1(n6054), .C2(EBX_REG_17__SCAN_IN), .A(n6273), .B(n5980), 
        .ZN(n5984) );
  INV_X1 U7046 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6556) );
  INV_X1 U7047 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6558) );
  OAI21_X1 U7048 ( .B1(n5989), .B2(n6556), .A(n6558), .ZN(n5981) );
  AOI22_X1 U7049 ( .A1(n6102), .A2(n4331), .B1(n5982), .B2(n5981), .ZN(n5983)
         );
  OAI211_X1 U7050 ( .C1(n5985), .C2(n6093), .A(n5984), .B(n5983), .ZN(U2810)
         );
  NAND2_X1 U7051 ( .A1(n5986), .A2(n6553), .ZN(n6002) );
  AOI22_X1 U7052 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n6087), .B1(n5987), 
        .B2(n6062), .ZN(n5988) );
  OAI211_X1 U7053 ( .C1(REIP_REG_16__SCAN_IN), .C2(n5989), .A(n6302), .B(n5988), .ZN(n5990) );
  AOI21_X1 U7054 ( .B1(n6054), .B2(EBX_REG_16__SCAN_IN), .A(n5990), .ZN(n5994)
         );
  INV_X1 U7055 ( .A(n5991), .ZN(n5992) );
  NAND2_X1 U7056 ( .A1(n6067), .A2(n5992), .ZN(n5993) );
  OAI211_X1 U7057 ( .C1(n5995), .C2(n6024), .A(n5994), .B(n5993), .ZN(n5996)
         );
  INV_X1 U7058 ( .A(n5996), .ZN(n5997) );
  OAI221_X1 U7059 ( .B1(n6556), .B2(n6009), .C1(n6556), .C2(n6002), .A(n5997), 
        .ZN(U2811) );
  INV_X1 U7060 ( .A(n5998), .ZN(n5999) );
  NAND2_X1 U7061 ( .A1(n6067), .A2(n5999), .ZN(n6005) );
  AOI22_X1 U7062 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6054), .B1(n6000), .B2(n6062), .ZN(n6001) );
  NAND3_X1 U7063 ( .A1(n6302), .A2(n6002), .A3(n6001), .ZN(n6003) );
  AOI21_X1 U7064 ( .B1(n6087), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6003), 
        .ZN(n6004) );
  NAND2_X1 U7065 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  AOI21_X1 U7066 ( .B1(n6007), .B2(n4331), .A(n6006), .ZN(n6008) );
  OAI21_X1 U7067 ( .B1(n6553), .B2(n6009), .A(n6008), .ZN(U2812) );
  NAND2_X1 U7068 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6020) );
  INV_X1 U7069 ( .A(n6021), .ZN(n6033) );
  NOR3_X1 U7070 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6020), .A3(n6033), .ZN(n6010) );
  AOI211_X1 U7071 ( .C1(n6087), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6273), 
        .B(n6010), .ZN(n6017) );
  INV_X1 U7072 ( .A(n6011), .ZN(n6213) );
  AOI22_X1 U7073 ( .A1(n6174), .A2(n6062), .B1(n6067), .B2(n6213), .ZN(n6016)
         );
  INV_X1 U7074 ( .A(n6012), .ZN(n6175) );
  AOI22_X1 U7075 ( .A1(n6175), .A2(n4331), .B1(n6013), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7076 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6054), .ZN(n6014) );
  NAND4_X1 U7077 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(U2816)
         );
  INV_X1 U7078 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6546) );
  OAI21_X1 U7079 ( .B1(n6019), .B2(n6018), .A(n6082), .ZN(n6050) );
  OAI22_X1 U7080 ( .A1(n6667), .A2(n6094), .B1(n6093), .B2(n6225), .ZN(n6027)
         );
  AOI21_X1 U7081 ( .B1(n6087), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6282), 
        .ZN(n6023) );
  OAI211_X1 U7082 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n6021), .B(n6020), .ZN(n6022) );
  OAI211_X1 U7083 ( .C1(n6025), .C2(n6024), .A(n6023), .B(n6022), .ZN(n6026)
         );
  AOI211_X1 U7084 ( .C1(n6028), .C2(n6062), .A(n6027), .B(n6026), .ZN(n6029)
         );
  OAI21_X1 U7085 ( .B1(n6546), .B2(n6050), .A(n6029), .ZN(U2817) );
  INV_X1 U7086 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6039) );
  AOI22_X1 U7087 ( .A1(n6030), .A2(n6062), .B1(n6067), .B2(n6233), .ZN(n6038)
         );
  INV_X1 U7088 ( .A(n6031), .ZN(n6036) );
  AOI21_X1 U7089 ( .B1(n6087), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6282), 
        .ZN(n6032) );
  OAI21_X1 U7090 ( .B1(n6033), .B2(REIP_REG_9__SCAN_IN), .A(n6032), .ZN(n6035)
         );
  INV_X1 U7091 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6544) );
  NOR2_X1 U7092 ( .A1(n6050), .A2(n6544), .ZN(n6034) );
  AOI211_X1 U7093 ( .C1(n6036), .C2(n4331), .A(n6035), .B(n6034), .ZN(n6037)
         );
  OAI211_X1 U7094 ( .C1(n6039), .C2(n6094), .A(n6038), .B(n6037), .ZN(U2818)
         );
  AOI21_X1 U7095 ( .B1(n6040), .B2(n6055), .A(REIP_REG_8__SCAN_IN), .ZN(n6051)
         );
  INV_X1 U7096 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6041) );
  OAI22_X1 U7097 ( .A1(n6042), .A2(n6094), .B1(n6041), .B2(n6075), .ZN(n6043)
         );
  AOI211_X1 U7098 ( .C1(n6067), .C2(n6242), .A(n6273), .B(n6043), .ZN(n6049)
         );
  INV_X1 U7099 ( .A(n6044), .ZN(n6047) );
  INV_X1 U7100 ( .A(n6045), .ZN(n6046) );
  AOI22_X1 U7101 ( .A1(n6047), .A2(n4331), .B1(n6046), .B2(n6062), .ZN(n6048)
         );
  OAI211_X1 U7102 ( .C1(n6051), .C2(n6050), .A(n6049), .B(n6048), .ZN(U2819)
         );
  INV_X1 U7103 ( .A(n6187), .ZN(n6053) );
  AOI22_X1 U7104 ( .A1(n6053), .A2(n6062), .B1(REIP_REG_6__SCAN_IN), .B2(n6052), .ZN(n6059) );
  AOI22_X1 U7105 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6054), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6087), .ZN(n6058) );
  AOI21_X1 U7106 ( .B1(n6067), .B2(n6261), .A(n6273), .ZN(n6057) );
  AOI22_X1 U7107 ( .A1(n6183), .A2(n4331), .B1(n6055), .B2(n6539), .ZN(n6056)
         );
  NAND4_X1 U7108 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(U2821)
         );
  NOR3_X1 U7109 ( .A1(n6079), .A2(n6060), .A3(REIP_REG_4__SCAN_IN), .ZN(n6061)
         );
  AOI211_X1 U7110 ( .C1(n6087), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6273), 
        .B(n6061), .ZN(n6073) );
  NAND2_X1 U7111 ( .A1(n6191), .A2(n6098), .ZN(n6071) );
  INV_X1 U7112 ( .A(n6194), .ZN(n6063) );
  AOI22_X1 U7113 ( .A1(n6065), .A2(n6064), .B1(n6063), .B2(n6062), .ZN(n6070)
         );
  NAND2_X1 U7114 ( .A1(n6066), .A2(REIP_REG_4__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7115 ( .A1(n6067), .A2(n6281), .ZN(n6068) );
  AND4_X1 U7116 ( .A1(n6071), .A2(n6070), .A3(n6069), .A4(n6068), .ZN(n6072)
         );
  OAI211_X1 U7117 ( .C1(n6787), .C2(n6094), .A(n6073), .B(n6072), .ZN(U2823)
         );
  INV_X1 U7118 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6074) );
  OAI22_X1 U7119 ( .A1(n6091), .A2(n6076), .B1(n6075), .B2(n6074), .ZN(n6078)
         );
  OAI22_X1 U7120 ( .A1(n6805), .A2(n6094), .B1(n6093), .B2(n6303), .ZN(n6077)
         );
  AOI211_X1 U7121 ( .C1(n6198), .C2(n6098), .A(n6078), .B(n6077), .ZN(n6085)
         );
  NOR2_X1 U7122 ( .A1(n6079), .A2(n6599), .ZN(n6083) );
  NAND3_X1 U7123 ( .A1(n6080), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6081) );
  OAI211_X1 U7124 ( .C1(n6083), .C2(REIP_REG_2__SCAN_IN), .A(n6082), .B(n6081), 
        .ZN(n6084) );
  OAI211_X1 U7125 ( .C1(n6101), .C2(n6201), .A(n6085), .B(n6084), .ZN(U2825)
         );
  AOI22_X1 U7126 ( .A1(n6087), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6086), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6089) );
  OAI211_X1 U7127 ( .C1(n6091), .C2(n6090), .A(n6089), .B(n6088), .ZN(n6097)
         );
  OAI22_X1 U7128 ( .A1(n6095), .A2(n6094), .B1(n6093), .B2(n6092), .ZN(n6096)
         );
  AOI211_X1 U7129 ( .C1(n6099), .C2(n6098), .A(n6097), .B(n6096), .ZN(n6100)
         );
  OAI21_X1 U7130 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6101), .A(n6100), 
        .ZN(U2826) );
  AOI22_X1 U7131 ( .A1(n6102), .A2(n6623), .B1(n6622), .B2(DATAI_17_), .ZN(
        n6104) );
  AOI22_X1 U7132 ( .A1(n6621), .A2(DATAI_1_), .B1(n6620), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7133 ( .A1(n6104), .A2(n6103), .ZN(U2874) );
  AOI22_X1 U7134 ( .A1(n6105), .A2(n6623), .B1(n6622), .B2(DATAI_16_), .ZN(
        n6107) );
  AOI22_X1 U7135 ( .A1(n6621), .A2(DATAI_0_), .B1(n6620), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7136 ( .A1(n6107), .A2(n6106), .ZN(U2875) );
  INV_X1 U7137 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6669) );
  INV_X1 U7138 ( .A(n6108), .ZN(n6109) );
  AOI22_X1 U7139 ( .A1(n6109), .A2(EAX_REG_20__SCAN_IN), .B1(n6612), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7140 ( .B1(n6669), .B2(n6111), .A(n6110), .ZN(U2903) );
  AOI22_X1 U7141 ( .A1(n6612), .A2(LWORD_REG_15__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7142 ( .B1(n6113), .B2(n6141), .A(n6112), .ZN(U2908) );
  AOI22_X1 U7143 ( .A1(n6612), .A2(LWORD_REG_14__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6114) );
  OAI21_X1 U7144 ( .B1(n6115), .B2(n6141), .A(n6114), .ZN(U2909) );
  AOI22_X1 U7145 ( .A1(n6612), .A2(LWORD_REG_13__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U7146 ( .B1(n6117), .B2(n6141), .A(n6116), .ZN(U2910) );
  AOI22_X1 U7147 ( .A1(n6612), .A2(LWORD_REG_12__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6118) );
  OAI21_X1 U7148 ( .B1(n6802), .B2(n6141), .A(n6118), .ZN(U2911) );
  AOI22_X1 U7149 ( .A1(n6612), .A2(LWORD_REG_11__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6119) );
  OAI21_X1 U7150 ( .B1(n6120), .B2(n6141), .A(n6119), .ZN(U2912) );
  AOI22_X1 U7151 ( .A1(n6612), .A2(LWORD_REG_10__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6121) );
  OAI21_X1 U7152 ( .B1(n6122), .B2(n6141), .A(n6121), .ZN(U2913) );
  AOI22_X1 U7153 ( .A1(n6612), .A2(LWORD_REG_9__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7154 ( .B1(n6124), .B2(n6141), .A(n6123), .ZN(U2914) );
  AOI22_X1 U7155 ( .A1(DATAO_REG_8__SCAN_IN), .A2(n6139), .B1(n6612), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U7156 ( .B1(n6126), .B2(n6141), .A(n6125), .ZN(U2915) );
  AOI22_X1 U7157 ( .A1(n6612), .A2(LWORD_REG_7__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6127) );
  OAI21_X1 U7158 ( .B1(n3838), .B2(n6141), .A(n6127), .ZN(U2916) );
  AOI22_X1 U7159 ( .A1(n6612), .A2(LWORD_REG_6__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6128) );
  OAI21_X1 U7160 ( .B1(n3832), .B2(n6141), .A(n6128), .ZN(U2917) );
  AOI22_X1 U7161 ( .A1(n6612), .A2(LWORD_REG_5__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6129) );
  OAI21_X1 U7162 ( .B1(n6130), .B2(n6141), .A(n6129), .ZN(U2918) );
  AOI222_X1 U7163 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6612), .B1(n6131), .B2(
        EAX_REG_4__SCAN_IN), .C1(n6139), .C2(DATAO_REG_4__SCAN_IN), .ZN(n6132)
         );
  INV_X1 U7164 ( .A(n6132), .ZN(U2919) );
  AOI22_X1 U7165 ( .A1(DATAO_REG_3__SCAN_IN), .A2(n6139), .B1(n6612), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n6133) );
  OAI21_X1 U7166 ( .B1(n6134), .B2(n6141), .A(n6133), .ZN(U2920) );
  AOI22_X1 U7167 ( .A1(n6612), .A2(LWORD_REG_2__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6135) );
  OAI21_X1 U7168 ( .B1(n6136), .B2(n6141), .A(n6135), .ZN(U2921) );
  AOI22_X1 U7169 ( .A1(n6612), .A2(LWORD_REG_1__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6137) );
  OAI21_X1 U7170 ( .B1(n6138), .B2(n6141), .A(n6137), .ZN(U2922) );
  AOI22_X1 U7171 ( .A1(n6612), .A2(LWORD_REG_0__SCAN_IN), .B1(n6139), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7172 ( .B1(n6142), .B2(n6141), .A(n6140), .ZN(U2923) );
  AOI22_X1 U7173 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n4478), .B1(n6165), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6145) );
  OAI21_X1 U7174 ( .B1(n6168), .B2(n6158), .A(n6145), .ZN(U2928) );
  AOI22_X1 U7175 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n4478), .B1(n6165), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6146) );
  OAI21_X1 U7176 ( .B1(n6168), .B2(n6160), .A(n6146), .ZN(U2929) );
  AOI22_X1 U7177 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n4478), .B1(n6165), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6147) );
  OAI21_X1 U7178 ( .B1(n6168), .B2(n6162), .A(n6147), .ZN(U2930) );
  AOI22_X1 U7179 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4478), .B1(n6165), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6148) );
  OAI21_X1 U7180 ( .B1(n6168), .B2(n6164), .A(n6148), .ZN(U2931) );
  AOI22_X1 U7181 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n4478), .B1(n6165), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6149) );
  OAI21_X1 U7182 ( .B1(n6168), .B2(n6167), .A(n6149), .ZN(U2936) );
  AOI22_X1 U7183 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n4478), .B1(n6165), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n6150) );
  OAI21_X1 U7184 ( .B1(n6168), .B2(n6151), .A(n6150), .ZN(U2939) );
  AOI22_X1 U7185 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n4478), .B1(n6165), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n6152) );
  OAI21_X1 U7186 ( .B1(n6168), .B2(n6153), .A(n6152), .ZN(U2940) );
  AOI22_X1 U7187 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n4498), .B1(n6165), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n6154) );
  OAI21_X1 U7188 ( .B1(n6168), .B2(n6155), .A(n6154), .ZN(U2941) );
  AOI22_X1 U7189 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n4498), .B1(n6165), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n6156) );
  OAI21_X1 U7190 ( .B1(n6168), .B2(n4502), .A(n6156), .ZN(U2942) );
  AOI22_X1 U7191 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n4498), .B1(n6165), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n6157) );
  OAI21_X1 U7192 ( .B1(n6168), .B2(n6158), .A(n6157), .ZN(U2943) );
  AOI22_X1 U7193 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4498), .B1(n6165), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n6159) );
  OAI21_X1 U7194 ( .B1(n6168), .B2(n6160), .A(n6159), .ZN(U2944) );
  AOI22_X1 U7195 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n4498), .B1(n6165), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6161) );
  OAI21_X1 U7196 ( .B1(n6168), .B2(n6162), .A(n6161), .ZN(U2945) );
  AOI22_X1 U7197 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4498), .B1(n6165), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6163) );
  OAI21_X1 U7198 ( .B1(n6168), .B2(n6164), .A(n6163), .ZN(U2946) );
  AOI22_X1 U7199 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n4498), .B1(n6165), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6166) );
  OAI21_X1 U7200 ( .B1(n6168), .B2(n6167), .A(n6166), .ZN(U2951) );
  NAND2_X1 U7201 ( .A1(n6170), .A2(n6169), .ZN(n6172) );
  XNOR2_X1 U7202 ( .A(n5650), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6171)
         );
  XNOR2_X1 U7203 ( .A(n6172), .B(n6171), .ZN(n6218) );
  AOI22_X1 U7204 ( .A1(n6273), .A2(REIP_REG_11__SCAN_IN), .B1(n6208), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6177) );
  AOI22_X1 U7205 ( .A1(n6175), .A2(n6184), .B1(n6174), .B2(n6173), .ZN(n6176)
         );
  OAI211_X1 U7206 ( .C1(n6218), .C2(n6178), .A(n6177), .B(n6176), .ZN(U2975)
         );
  AOI22_X1 U7207 ( .A1(n6273), .A2(REIP_REG_6__SCAN_IN), .B1(n6208), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6186) );
  OAI21_X1 U7208 ( .B1(n6181), .B2(n6180), .A(n6179), .ZN(n6182) );
  INV_X1 U7209 ( .A(n6182), .ZN(n6263) );
  AOI22_X1 U7210 ( .A1(n6263), .A2(n6206), .B1(n6184), .B2(n6183), .ZN(n6185)
         );
  OAI211_X1 U7211 ( .C1(n6202), .C2(n6187), .A(n6186), .B(n6185), .ZN(U2980)
         );
  AOI22_X1 U7212 ( .A1(n6273), .A2(REIP_REG_4__SCAN_IN), .B1(n6208), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6193) );
  INV_X1 U7213 ( .A(n6190), .ZN(n6280) );
  AOI22_X1 U7214 ( .A1(n6280), .A2(n6206), .B1(n6191), .B2(n6184), .ZN(n6192)
         );
  OAI211_X1 U7215 ( .C1(n6202), .C2(n6194), .A(n6193), .B(n6192), .ZN(U2982)
         );
  AOI22_X1 U7216 ( .A1(n6273), .A2(REIP_REG_2__SCAN_IN), .B1(n6208), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6200) );
  XOR2_X1 U7217 ( .A(n3021), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6196) );
  XNOR2_X1 U7218 ( .A(n6197), .B(n6196), .ZN(n6308) );
  AOI22_X1 U7219 ( .A1(n6308), .A2(n6206), .B1(n6184), .B2(n6198), .ZN(n6199)
         );
  OAI211_X1 U7220 ( .C1(n6202), .C2(n6201), .A(n6200), .B(n6199), .ZN(U2984)
         );
  INV_X1 U7221 ( .A(n6203), .ZN(n6204) );
  AOI21_X1 U7222 ( .B1(n6206), .B2(n6205), .A(n6204), .ZN(n6210) );
  OAI21_X1 U7223 ( .B1(n6208), .B2(n6207), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6209) );
  OAI211_X1 U7224 ( .C1(n6212), .C2(n6211), .A(n6210), .B(n6209), .ZN(U2986)
         );
  AOI22_X1 U7225 ( .A1(n6290), .A2(n6213), .B1(n6282), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6217) );
  AOI22_X1 U7226 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6215), .B1(n6214), .B2(n3531), .ZN(n6216) );
  OAI211_X1 U7227 ( .C1(n6218), .C2(n6224), .A(n6217), .B(n6216), .ZN(U3007)
         );
  INV_X1 U7228 ( .A(n6257), .ZN(n6220) );
  OAI22_X1 U7229 ( .A1(n6222), .A2(n6221), .B1(n6220), .B2(n6219), .ZN(n6251)
         );
  AOI21_X1 U7230 ( .B1(n6260), .B2(n6240), .A(n6251), .ZN(n6239) );
  OAI222_X1 U7231 ( .A1(n6225), .A2(n6304), .B1(n6302), .B2(n6546), .C1(n6224), 
        .C2(n6223), .ZN(n6226) );
  INV_X1 U7232 ( .A(n6226), .ZN(n6231) );
  AOI21_X1 U7233 ( .B1(n6227), .B2(n6297), .A(n6279), .ZN(n6283) );
  NAND2_X1 U7234 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6228), .ZN(n6259)
         );
  NOR2_X1 U7235 ( .A1(n6283), .A2(n6259), .ZN(n6262) );
  NAND2_X1 U7236 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6262), .ZN(n6255)
         );
  NOR2_X1 U7237 ( .A1(n6240), .A2(n6255), .ZN(n6234) );
  OAI211_X1 U7238 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6234), .B(n6229), .ZN(n6230) );
  OAI211_X1 U7239 ( .C1(n6239), .C2(n3530), .A(n6231), .B(n6230), .ZN(U3008)
         );
  AOI21_X1 U7240 ( .B1(n6290), .B2(n6233), .A(n6232), .ZN(n6237) );
  AOI22_X1 U7241 ( .A1(n6235), .A2(n6307), .B1(n6234), .B2(n6238), .ZN(n6236)
         );
  OAI211_X1 U7242 ( .C1(n6239), .C2(n6238), .A(n6237), .B(n6236), .ZN(U3009)
         );
  OAI21_X1 U7243 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6240), .ZN(n6246) );
  AOI21_X1 U7244 ( .B1(n6290), .B2(n6242), .A(n6241), .ZN(n6245) );
  AOI22_X1 U7245 ( .A1(n6243), .A2(n6307), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6251), .ZN(n6244) );
  OAI211_X1 U7246 ( .C1(n6255), .C2(n6246), .A(n6245), .B(n6244), .ZN(U3010)
         );
  INV_X1 U7247 ( .A(n6247), .ZN(n6248) );
  AOI21_X1 U7248 ( .B1(n6290), .B2(n6249), .A(n6248), .ZN(n6254) );
  INV_X1 U7249 ( .A(n6250), .ZN(n6252) );
  AOI22_X1 U7250 ( .A1(n6252), .A2(n6307), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6251), .ZN(n6253) );
  OAI211_X1 U7251 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6255), .A(n6254), 
        .B(n6253), .ZN(U3011) );
  AOI22_X1 U7252 ( .A1(n6301), .A2(n6258), .B1(n6257), .B2(n6256), .ZN(n6310)
         );
  INV_X1 U7253 ( .A(n6310), .ZN(n6278) );
  AOI21_X1 U7254 ( .B1(n6260), .B2(n6259), .A(n6278), .ZN(n6277) );
  AOI22_X1 U7255 ( .A1(n6290), .A2(n6261), .B1(n6282), .B2(REIP_REG_6__SCAN_IN), .ZN(n6265) );
  AOI22_X1 U7256 ( .A1(n6263), .A2(n6307), .B1(n6262), .B2(n6266), .ZN(n6264)
         );
  OAI211_X1 U7257 ( .C1(n6277), .C2(n6266), .A(n6265), .B(n6264), .ZN(U3012)
         );
  INV_X1 U7258 ( .A(n6267), .ZN(n6268) );
  AOI211_X1 U7259 ( .C1(n6269), .C2(n6297), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .B(n6268), .ZN(n6276) );
  INV_X1 U7260 ( .A(n6270), .ZN(n6272) );
  AOI22_X1 U7261 ( .A1(n6272), .A2(n6307), .B1(n6290), .B2(n6271), .ZN(n6275)
         );
  NAND2_X1 U7262 ( .A1(n6273), .A2(REIP_REG_5__SCAN_IN), .ZN(n6274) );
  OAI211_X1 U7263 ( .C1(n6277), .C2(n6276), .A(n6275), .B(n6274), .ZN(U3013)
         );
  AOI21_X1 U7264 ( .B1(n6279), .B2(n6298), .A(n6278), .ZN(n6296) );
  AOI222_X1 U7265 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6282), .B1(n6290), .B2(
        n6281), .C1(n6307), .C2(n6280), .ZN(n6286) );
  NOR2_X1 U7266 ( .A1(n6298), .A2(n6283), .ZN(n6292) );
  OAI211_X1 U7267 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6292), .B(n6284), .ZN(n6285) );
  OAI211_X1 U7268 ( .C1(n6296), .C2(n6287), .A(n6286), .B(n6285), .ZN(U3014)
         );
  AOI21_X1 U7269 ( .B1(n6290), .B2(n6289), .A(n6288), .ZN(n6294) );
  AOI22_X1 U7270 ( .A1(n6292), .A2(n6295), .B1(n6291), .B2(n6307), .ZN(n6293)
         );
  OAI211_X1 U7271 ( .C1(n6296), .C2(n6295), .A(n6294), .B(n6293), .ZN(U3015)
         );
  NAND2_X1 U7272 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6297), .ZN(n6311)
         );
  AOI21_X1 U7273 ( .B1(n6299), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6298), 
        .ZN(n6300) );
  NOR2_X1 U7274 ( .A1(n6301), .A2(n6300), .ZN(n6306) );
  INV_X1 U7275 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6532) );
  OAI22_X1 U7276 ( .A1(n6304), .A2(n6303), .B1(n6532), .B2(n6302), .ZN(n6305)
         );
  AOI211_X1 U7277 ( .C1(n6308), .C2(n6307), .A(n6306), .B(n6305), .ZN(n6309)
         );
  OAI221_X1 U7278 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6311), .C1(n3435), .C2(n6310), .A(n6309), .ZN(U3016) );
  NOR2_X1 U7279 ( .A1(n6479), .A2(n6312), .ZN(U3019) );
  NOR2_X1 U7280 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6313), .ZN(n6338)
         );
  NAND3_X1 U7281 ( .A1(n6314), .A2(n6360), .A3(n6359), .ZN(n6315) );
  OAI21_X1 U7282 ( .B1(n6319), .B2(n6316), .A(n6315), .ZN(n6337) );
  AOI22_X1 U7283 ( .A1(n6432), .A2(n6338), .B1(n6433), .B2(n6337), .ZN(n6324)
         );
  INV_X1 U7284 ( .A(n6356), .ZN(n6318) );
  OAI21_X1 U7285 ( .B1(n6339), .B2(n6318), .A(n6317), .ZN(n6320) );
  AOI21_X1 U7286 ( .B1(n6320), .B2(n6319), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6322) );
  AOI22_X1 U7287 ( .A1(n6340), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6374), 
        .B2(n6339), .ZN(n6323) );
  OAI211_X1 U7288 ( .C1(n6377), .C2(n6356), .A(n6324), .B(n6323), .ZN(U3036)
         );
  AOI22_X1 U7289 ( .A1(n6417), .A2(n6338), .B1(n6418), .B2(n6337), .ZN(n6326)
         );
  AOI22_X1 U7290 ( .A1(n6340), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6378), 
        .B2(n6339), .ZN(n6325) );
  OAI211_X1 U7291 ( .C1(n6356), .C2(n6381), .A(n6326), .B(n6325), .ZN(U3037)
         );
  AOI22_X1 U7292 ( .A1(n6383), .A2(n6338), .B1(n6382), .B2(n6337), .ZN(n6328)
         );
  AOI22_X1 U7293 ( .A1(n6340), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6384), 
        .B2(n6339), .ZN(n6327) );
  OAI211_X1 U7294 ( .C1(n6356), .C2(n6387), .A(n6328), .B(n6327), .ZN(U3038)
         );
  AOI22_X1 U7295 ( .A1(n6438), .A2(n6338), .B1(n6439), .B2(n6337), .ZN(n6330)
         );
  AOI22_X1 U7296 ( .A1(n6340), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6388), 
        .B2(n6339), .ZN(n6329) );
  OAI211_X1 U7297 ( .C1(n6356), .C2(n6391), .A(n6330), .B(n6329), .ZN(U3039)
         );
  AOI22_X1 U7298 ( .A1(n6445), .A2(n6337), .B1(n6443), .B2(n6338), .ZN(n6332)
         );
  AOI22_X1 U7299 ( .A1(n6340), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6392), 
        .B2(n6339), .ZN(n6331) );
  OAI211_X1 U7300 ( .C1(n6356), .C2(n6395), .A(n6332), .B(n6331), .ZN(U3040)
         );
  AOI22_X1 U7301 ( .A1(n6397), .A2(n6338), .B1(n6396), .B2(n6337), .ZN(n6334)
         );
  AOI22_X1 U7302 ( .A1(n6340), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6398), 
        .B2(n6339), .ZN(n6333) );
  OAI211_X1 U7303 ( .C1(n6356), .C2(n6401), .A(n6334), .B(n6333), .ZN(U3041)
         );
  AOI22_X1 U7304 ( .A1(n6452), .A2(n6338), .B1(n6454), .B2(n6337), .ZN(n6336)
         );
  AOI22_X1 U7305 ( .A1(n6340), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6402), 
        .B2(n6339), .ZN(n6335) );
  OAI211_X1 U7306 ( .C1(n6356), .C2(n6405), .A(n6336), .B(n6335), .ZN(U3042)
         );
  AOI22_X1 U7307 ( .A1(n6409), .A2(n6338), .B1(n6407), .B2(n6337), .ZN(n6342)
         );
  AOI22_X1 U7308 ( .A1(n6340), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6411), 
        .B2(n6339), .ZN(n6341) );
  OAI211_X1 U7309 ( .C1(n6356), .C2(n6415), .A(n6342), .B(n6341), .ZN(U3043)
         );
  INV_X1 U7310 ( .A(n6343), .ZN(n6350) );
  AOI22_X1 U7311 ( .A1(n6438), .A2(n6350), .B1(n6349), .B2(n6437), .ZN(n6345)
         );
  AOI22_X1 U7312 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6352), .B1(n6439), 
        .B2(n6351), .ZN(n6344) );
  OAI211_X1 U7313 ( .C1(n6356), .C2(n6442), .A(n6345), .B(n6344), .ZN(U3047)
         );
  AOI22_X1 U7314 ( .A1(n6443), .A2(n6350), .B1(n6349), .B2(n6444), .ZN(n6347)
         );
  AOI22_X1 U7315 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6352), .B1(n6445), 
        .B2(n6351), .ZN(n6346) );
  OAI211_X1 U7316 ( .C1(n6356), .C2(n6448), .A(n6347), .B(n6346), .ZN(U3048)
         );
  AOI22_X1 U7317 ( .A1(n6409), .A2(n6350), .B1(n6349), .B2(n6348), .ZN(n6354)
         );
  AOI22_X1 U7318 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6352), .B1(n6407), 
        .B2(n6351), .ZN(n6353) );
  OAI211_X1 U7319 ( .C1(n6356), .C2(n6355), .A(n6354), .B(n6353), .ZN(U3051)
         );
  NAND2_X1 U7320 ( .A1(n6632), .A2(n6357), .ZN(n6369) );
  INV_X1 U7321 ( .A(n6369), .ZN(n6408) );
  INV_X1 U7322 ( .A(n6358), .ZN(n6364) );
  NAND3_X1 U7323 ( .A1(n6361), .A2(n6360), .A3(n6359), .ZN(n6362) );
  OAI21_X1 U7324 ( .B1(n6364), .B2(n6363), .A(n6362), .ZN(n6406) );
  AOI22_X1 U7325 ( .A1(n6432), .A2(n6408), .B1(n6433), .B2(n6406), .ZN(n6376)
         );
  AOI21_X1 U7326 ( .B1(n6366), .B2(n6430), .A(n6365), .ZN(n6373) );
  NAND2_X1 U7327 ( .A1(n6368), .A2(n6367), .ZN(n6372) );
  AOI21_X1 U7328 ( .B1(n6369), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6370) );
  OAI211_X1 U7329 ( .C1(n6373), .C2(n6372), .A(n6371), .B(n6370), .ZN(n6412)
         );
  AOI22_X1 U7330 ( .A1(n6412), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6374), 
        .B2(n6410), .ZN(n6375) );
  OAI211_X1 U7331 ( .C1(n6377), .C2(n6430), .A(n6376), .B(n6375), .ZN(U3068)
         );
  AOI22_X1 U7332 ( .A1(n6417), .A2(n6408), .B1(n6418), .B2(n6406), .ZN(n6380)
         );
  AOI22_X1 U7333 ( .A1(n6412), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6378), 
        .B2(n6410), .ZN(n6379) );
  OAI211_X1 U7334 ( .C1(n6381), .C2(n6430), .A(n6380), .B(n6379), .ZN(U3069)
         );
  AOI22_X1 U7335 ( .A1(n6383), .A2(n6408), .B1(n6382), .B2(n6406), .ZN(n6386)
         );
  AOI22_X1 U7336 ( .A1(n6412), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6384), 
        .B2(n6410), .ZN(n6385) );
  OAI211_X1 U7337 ( .C1(n6387), .C2(n6430), .A(n6386), .B(n6385), .ZN(U3070)
         );
  AOI22_X1 U7338 ( .A1(n6438), .A2(n6408), .B1(n6439), .B2(n6406), .ZN(n6390)
         );
  AOI22_X1 U7339 ( .A1(n6412), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6388), 
        .B2(n6410), .ZN(n6389) );
  OAI211_X1 U7340 ( .C1(n6391), .C2(n6430), .A(n6390), .B(n6389), .ZN(U3071)
         );
  AOI22_X1 U7341 ( .A1(n6445), .A2(n6406), .B1(n6443), .B2(n6408), .ZN(n6394)
         );
  AOI22_X1 U7342 ( .A1(n6412), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6392), 
        .B2(n6410), .ZN(n6393) );
  OAI211_X1 U7343 ( .C1(n6395), .C2(n6430), .A(n6394), .B(n6393), .ZN(U3072)
         );
  AOI22_X1 U7344 ( .A1(n6397), .A2(n6408), .B1(n6396), .B2(n6406), .ZN(n6400)
         );
  AOI22_X1 U7345 ( .A1(n6412), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6398), 
        .B2(n6410), .ZN(n6399) );
  OAI211_X1 U7346 ( .C1(n6401), .C2(n6430), .A(n6400), .B(n6399), .ZN(U3073)
         );
  AOI22_X1 U7347 ( .A1(n6452), .A2(n6408), .B1(n6454), .B2(n6406), .ZN(n6404)
         );
  AOI22_X1 U7348 ( .A1(n6412), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6402), 
        .B2(n6410), .ZN(n6403) );
  OAI211_X1 U7349 ( .C1(n6405), .C2(n6430), .A(n6404), .B(n6403), .ZN(U3074)
         );
  AOI22_X1 U7350 ( .A1(n6409), .A2(n6408), .B1(n6407), .B2(n6406), .ZN(n6414)
         );
  AOI22_X1 U7351 ( .A1(n6412), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6411), 
        .B2(n6410), .ZN(n6413) );
  OAI211_X1 U7352 ( .C1(n6415), .C2(n6430), .A(n6414), .B(n6413), .ZN(U3075)
         );
  AOI22_X1 U7353 ( .A1(n6417), .A2(n6425), .B1(n6416), .B2(n6424), .ZN(n6420)
         );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6427), .B1(n6418), 
        .B2(n6426), .ZN(n6419) );
  OAI211_X1 U7355 ( .C1(n6421), .C2(n6430), .A(n6420), .B(n6419), .ZN(U3077)
         );
  AOI22_X1 U7356 ( .A1(n6438), .A2(n6425), .B1(n6437), .B2(n6424), .ZN(n6423)
         );
  AOI22_X1 U7357 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6427), .B1(n6439), 
        .B2(n6426), .ZN(n6422) );
  OAI211_X1 U7358 ( .C1(n6442), .C2(n6430), .A(n6423), .B(n6422), .ZN(U3079)
         );
  AOI22_X1 U7359 ( .A1(n6443), .A2(n6425), .B1(n6444), .B2(n6424), .ZN(n6429)
         );
  AOI22_X1 U7360 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6427), .B1(n6445), 
        .B2(n6426), .ZN(n6428) );
  OAI211_X1 U7361 ( .C1(n6448), .C2(n6430), .A(n6429), .B(n6428), .ZN(U3080)
         );
  AOI22_X1 U7362 ( .A1(n6432), .A2(n6451), .B1(n6450), .B2(n6431), .ZN(n6435)
         );
  AOI22_X1 U7363 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6455), .B1(n6433), 
        .B2(n6453), .ZN(n6434) );
  OAI211_X1 U7364 ( .C1(n6436), .C2(n6458), .A(n6435), .B(n6434), .ZN(U3108)
         );
  AOI22_X1 U7365 ( .A1(n6438), .A2(n6451), .B1(n6450), .B2(n6437), .ZN(n6441)
         );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6455), .B1(n6439), 
        .B2(n6453), .ZN(n6440) );
  OAI211_X1 U7367 ( .C1(n6442), .C2(n6458), .A(n6441), .B(n6440), .ZN(U3111)
         );
  AOI22_X1 U7368 ( .A1(n6450), .A2(n6444), .B1(n6443), .B2(n6451), .ZN(n6447)
         );
  AOI22_X1 U7369 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6455), .B1(n6445), 
        .B2(n6453), .ZN(n6446) );
  OAI211_X1 U7370 ( .C1(n6448), .C2(n6458), .A(n6447), .B(n6446), .ZN(U3112)
         );
  AOI22_X1 U7371 ( .A1(n6452), .A2(n6451), .B1(n6450), .B2(n6449), .ZN(n6457)
         );
  AOI22_X1 U7372 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6455), .B1(n6454), 
        .B2(n6453), .ZN(n6456) );
  OAI211_X1 U7373 ( .C1(n6459), .C2(n6458), .A(n6457), .B(n6456), .ZN(U3114)
         );
  INV_X1 U7374 ( .A(n6460), .ZN(n6461) );
  OAI211_X1 U7375 ( .C1(n6463), .C2(n6462), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n6461), .ZN(n6466) );
  INV_X1 U7376 ( .A(n6464), .ZN(n6465) );
  OAI21_X1 U7377 ( .B1(n6467), .B2(n6466), .A(n6465), .ZN(n6469) );
  NAND2_X1 U7378 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  OAI21_X1 U7379 ( .B1(n6470), .B2(n6469), .A(n6468), .ZN(n6475) );
  NAND2_X1 U7380 ( .A1(n6474), .A2(n6475), .ZN(n6471) );
  NAND2_X1 U7381 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  OAI21_X1 U7382 ( .B1(n6475), .B2(n6474), .A(n6473), .ZN(n6476) );
  OAI21_X1 U7383 ( .B1(n6477), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6476), 
        .ZN(n6480) );
  NAND2_X1 U7384 ( .A1(n6477), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6478) );
  NAND3_X1 U7385 ( .A1(n6480), .A2(n6479), .A3(n6478), .ZN(n6489) );
  NOR2_X1 U7386 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6483) );
  OAI211_X1 U7387 ( .C1(n6484), .C2(n6483), .A(n6482), .B(n6481), .ZN(n6485)
         );
  NOR2_X1 U7388 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  NAND2_X1 U7389 ( .A1(n6502), .A2(n6503), .ZN(n6491) );
  NAND2_X1 U7390 ( .A1(n6612), .A2(READY_N), .ZN(n6490) );
  NAND2_X1 U7391 ( .A1(n6491), .A2(n6490), .ZN(n6495) );
  OR2_X1 U7392 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  OAI21_X1 U7393 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6611), .A(n6590), .ZN(
        n6505) );
  AOI221_X1 U7394 ( .B1(n6497), .B2(STATE2_REG_0__SCAN_IN), .C1(n6505), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6496), .ZN(n6500) );
  OAI211_X1 U7395 ( .C1(n6498), .C2(n6592), .A(n6506), .B(n6590), .ZN(n6499)
         );
  OAI211_X1 U7396 ( .C1(n6502), .C2(n6501), .A(n6500), .B(n6499), .ZN(U3148)
         );
  NOR2_X1 U7397 ( .A1(n6506), .A2(n6594), .ZN(n6504) );
  AOI21_X1 U7398 ( .B1(n6504), .B2(n6611), .A(n6503), .ZN(n6509) );
  OAI221_X1 U7399 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n4242), .C1(n6506), .C2(
        n6505), .A(STATE2_REG_1__SCAN_IN), .ZN(n6507) );
  OAI221_X1 U7400 ( .B1(n6510), .B2(n6509), .C1(n6590), .C2(n6508), .A(n6507), 
        .ZN(U3149) );
  OAI221_X1 U7401 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6611), .A(n6589), .ZN(n6512) );
  OAI21_X1 U7402 ( .B1(n6614), .B2(n6512), .A(n6511), .ZN(U3150) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6513), .ZN(U3151) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6513), .ZN(U3152) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6513), .ZN(U3153) );
  INV_X1 U7406 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6797) );
  NOR2_X1 U7407 ( .A1(n6588), .A2(n6797), .ZN(U3154) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6513), .ZN(U3155) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6513), .ZN(U3156) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6513), .ZN(U3157) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6513), .ZN(U3158) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6513), .ZN(U3159) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6513), .ZN(U3160) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6513), .ZN(U3161) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6513), .ZN(U3162) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6513), .ZN(U3163) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6513), .ZN(U3164) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6513), .ZN(U3165) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6513), .ZN(U3166) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6513), .ZN(U3167) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6513), .ZN(U3168) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6513), .ZN(U3169) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6513), .ZN(U3170) );
  AND2_X1 U7424 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6513), .ZN(U3171) );
  AND2_X1 U7425 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6513), .ZN(U3172) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6513), .ZN(U3173) );
  AND2_X1 U7427 ( .A1(n6513), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  AND2_X1 U7428 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6513), .ZN(U3175) );
  AND2_X1 U7429 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6513), .ZN(U3176) );
  AND2_X1 U7430 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6513), .ZN(U3177) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6513), .ZN(U3178) );
  AND2_X1 U7432 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6513), .ZN(U3179) );
  AND2_X1 U7433 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6513), .ZN(U3180) );
  INV_X1 U7434 ( .A(n6514), .ZN(n6523) );
  AOI22_X1 U7435 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6527) );
  AND2_X1 U7436 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6518) );
  INV_X1 U7437 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6516) );
  INV_X1 U7438 ( .A(NA_N), .ZN(n6524) );
  AOI211_X1 U7439 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6524), .A(
        STATE_REG_0__SCAN_IN), .B(n6523), .ZN(n6529) );
  AOI221_X1 U7440 ( .B1(n6518), .B2(n6619), .C1(n6516), .C2(n6619), .A(n6529), 
        .ZN(n6515) );
  OAI21_X1 U7441 ( .B1(n6523), .B2(n6527), .A(n6515), .ZN(U3181) );
  NOR2_X1 U7442 ( .A1(n6803), .A2(n6516), .ZN(n6525) );
  NAND2_X1 U7443 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6517) );
  OAI21_X1 U7444 ( .B1(n6525), .B2(n6518), .A(n6517), .ZN(n6519) );
  OAI211_X1 U7445 ( .C1(n6521), .C2(n6611), .A(n6520), .B(n6519), .ZN(U3182)
         );
  AOI221_X1 U7446 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6611), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6522) );
  AOI221_X1 U7447 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6522), .C2(HOLD), .A(n6803), .ZN(n6528) );
  AOI21_X1 U7448 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n6526) );
  OAI22_X1 U7449 ( .A1(n6529), .A2(n6528), .B1(n6527), .B2(n6526), .ZN(U3183)
         );
  NAND2_X1 U7450 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6559), .ZN(n6579) );
  NOR2_X2 U7451 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6619), .ZN(n6577) );
  AOI22_X1 U7452 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6619), .ZN(n6530) );
  OAI21_X1 U7453 ( .B1(n6599), .B2(n6579), .A(n6530), .ZN(U3184) );
  AOI22_X1 U7454 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6619), .ZN(n6531) );
  OAI21_X1 U7455 ( .B1(n6532), .B2(n6579), .A(n6531), .ZN(U3185) );
  INV_X1 U7456 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6533) );
  INV_X1 U7457 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6806) );
  OAI222_X1 U7458 ( .A1(n6579), .A2(n6533), .B1(n6806), .B2(n6559), .C1(n6535), 
        .C2(n6583), .ZN(U3186) );
  AOI22_X1 U7459 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6619), .ZN(n6534) );
  OAI21_X1 U7460 ( .B1(n6535), .B2(n6579), .A(n6534), .ZN(U3187) );
  AOI22_X1 U7461 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6619), .ZN(n6536) );
  OAI21_X1 U7462 ( .B1(n6537), .B2(n6579), .A(n6536), .ZN(U3188) );
  AOI22_X1 U7463 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6619), .ZN(n6538) );
  OAI21_X1 U7464 ( .B1(n6539), .B2(n6579), .A(n6538), .ZN(U3189) );
  AOI22_X1 U7465 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6619), .ZN(n6540) );
  OAI21_X1 U7466 ( .B1(n6541), .B2(n6579), .A(n6540), .ZN(U3190) );
  INV_X1 U7467 ( .A(n6579), .ZN(n6581) );
  AOI22_X1 U7468 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6619), .ZN(n6542) );
  OAI21_X1 U7469 ( .B1(n6544), .B2(n6583), .A(n6542), .ZN(U3191) );
  AOI22_X1 U7470 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6619), .ZN(n6543) );
  OAI21_X1 U7471 ( .B1(n6544), .B2(n6579), .A(n6543), .ZN(U3192) );
  AOI22_X1 U7472 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6619), .ZN(n6545) );
  OAI21_X1 U7473 ( .B1(n6546), .B2(n6579), .A(n6545), .ZN(U3193) );
  AOI22_X1 U7474 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6619), .ZN(n6547) );
  OAI21_X1 U7475 ( .B1(n6549), .B2(n6583), .A(n6547), .ZN(U3194) );
  AOI22_X1 U7476 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6619), .ZN(n6548) );
  OAI21_X1 U7477 ( .B1(n6549), .B2(n6579), .A(n6548), .ZN(U3195) );
  AOI22_X1 U7478 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6619), .ZN(n6550) );
  OAI21_X1 U7479 ( .B1(n6551), .B2(n6583), .A(n6550), .ZN(U3196) );
  AOI22_X1 U7480 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6619), .ZN(n6552) );
  OAI21_X1 U7481 ( .B1(n6553), .B2(n6583), .A(n6552), .ZN(U3197) );
  AOI22_X1 U7482 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6619), .ZN(n6554) );
  OAI21_X1 U7483 ( .B1(n6556), .B2(n6583), .A(n6554), .ZN(U3198) );
  AOI22_X1 U7484 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6619), .ZN(n6555) );
  OAI21_X1 U7485 ( .B1(n6556), .B2(n6579), .A(n6555), .ZN(U3199) );
  AOI22_X1 U7486 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6619), .ZN(n6557) );
  OAI21_X1 U7487 ( .B1(n6558), .B2(n6579), .A(n6557), .ZN(U3200) );
  INV_X1 U7488 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6779) );
  OAI222_X1 U7489 ( .A1(n6579), .A2(n6560), .B1(n6779), .B2(n6559), .C1(n6562), 
        .C2(n6583), .ZN(U3201) );
  AOI22_X1 U7490 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6619), .ZN(n6561) );
  OAI21_X1 U7491 ( .B1(n6562), .B2(n6579), .A(n6561), .ZN(U3202) );
  AOI22_X1 U7492 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6619), .ZN(n6563) );
  OAI21_X1 U7493 ( .B1(n6564), .B2(n6583), .A(n6563), .ZN(U3203) );
  INV_X1 U7494 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6628) );
  AOI22_X1 U7495 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6619), .ZN(n6565) );
  OAI21_X1 U7496 ( .B1(n6628), .B2(n6583), .A(n6565), .ZN(U3204) );
  AOI22_X1 U7497 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6619), .ZN(n6566) );
  OAI21_X1 U7498 ( .B1(n6628), .B2(n6579), .A(n6566), .ZN(U3205) );
  AOI22_X1 U7499 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6619), .ZN(n6567) );
  OAI21_X1 U7500 ( .B1(n6568), .B2(n6579), .A(n6567), .ZN(U3206) );
  AOI22_X1 U7501 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6619), .ZN(n6569) );
  OAI21_X1 U7502 ( .B1(n6570), .B2(n6579), .A(n6569), .ZN(U3207) );
  AOI22_X1 U7503 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6619), .ZN(n6571) );
  OAI21_X1 U7504 ( .B1(n6572), .B2(n6583), .A(n6571), .ZN(U3208) );
  AOI22_X1 U7505 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6619), .ZN(n6573) );
  OAI21_X1 U7506 ( .B1(n6575), .B2(n6583), .A(n6573), .ZN(U3209) );
  AOI22_X1 U7507 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6619), .ZN(n6574) );
  OAI21_X1 U7508 ( .B1(n6575), .B2(n6579), .A(n6574), .ZN(U3210) );
  AOI22_X1 U7509 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6619), .ZN(n6576) );
  OAI21_X1 U7510 ( .B1(n6580), .B2(n6583), .A(n6576), .ZN(U3211) );
  AOI22_X1 U7511 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6619), .ZN(n6578) );
  OAI21_X1 U7512 ( .B1(n6580), .B2(n6579), .A(n6578), .ZN(U3212) );
  AOI22_X1 U7513 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6581), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6619), .ZN(n6582) );
  OAI21_X1 U7514 ( .B1(n6584), .B2(n6583), .A(n6582), .ZN(U3213) );
  MUX2_X1 U7515 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6619), .Z(U3445) );
  MUX2_X1 U7516 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6619), .Z(U3446) );
  MUX2_X1 U7517 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6619), .Z(U3447) );
  MUX2_X1 U7518 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6619), .Z(U3448) );
  OAI21_X1 U7519 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6588), .A(n6586), .ZN(
        n6585) );
  INV_X1 U7520 ( .A(n6585), .ZN(U3451) );
  OAI21_X1 U7521 ( .B1(n6588), .B2(n6587), .A(n6586), .ZN(U3452) );
  OAI221_X1 U7522 ( .B1(n6591), .B2(STATE2_REG_0__SCAN_IN), .C1(n6591), .C2(
        n6590), .A(n6589), .ZN(U3453) );
  OAI22_X1 U7523 ( .A1(n6595), .A2(n6594), .B1(n6593), .B2(n6592), .ZN(n6597)
         );
  MUX2_X1 U7524 ( .A(n6598), .B(n6597), .S(n6596), .Z(U3456) );
  AOI21_X1 U7525 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6600) );
  AOI22_X1 U7526 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6600), .B2(n6599), .ZN(n6602) );
  INV_X1 U7527 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U7528 ( .A1(n6603), .A2(n6602), .B1(n6601), .B2(n6606), .ZN(U3468)
         );
  INV_X1 U7529 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6607) );
  INV_X1 U7530 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6605) );
  NOR2_X1 U7531 ( .A1(n6606), .A2(REIP_REG_1__SCAN_IN), .ZN(n6604) );
  AOI22_X1 U7532 ( .A1(n6607), .A2(n6606), .B1(n6605), .B2(n6604), .ZN(U3469)
         );
  NAND2_X1 U7533 ( .A1(n6619), .A2(W_R_N_REG_SCAN_IN), .ZN(n6608) );
  OAI21_X1 U7534 ( .B1(n6619), .B2(READREQUEST_REG_SCAN_IN), .A(n6608), .ZN(
        U3470) );
  AOI211_X1 U7535 ( .C1(n6612), .C2(n6611), .A(n6610), .B(n6609), .ZN(n6618)
         );
  OAI211_X1 U7536 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3412), .A(n6613), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6615) );
  AOI21_X1 U7537 ( .B1(n6615), .B2(STATE2_REG_0__SCAN_IN), .A(n6614), .ZN(
        n6617) );
  NAND2_X1 U7538 ( .A1(n6618), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6616) );
  OAI21_X1 U7539 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(U3472) );
  MUX2_X1 U7540 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6619), .Z(U3473) );
  AOI22_X1 U7541 ( .A1(n6621), .A2(DATAI_5_), .B1(n6620), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6626) );
  AOI22_X1 U7542 ( .A1(n6624), .A2(n6623), .B1(n6622), .B2(DATAI_21_), .ZN(
        n6625) );
  NAND2_X1 U7543 ( .A1(n6626), .A2(n6625), .ZN(n6819) );
  INV_X1 U7544 ( .A(DATAI_25_), .ZN(n6629) );
  AOI22_X1 U7545 ( .A1(n6629), .A2(keyinput65), .B1(n6628), .B2(keyinput76), 
        .ZN(n6627) );
  OAI221_X1 U7546 ( .B1(n6629), .B2(keyinput65), .C1(n6628), .C2(keyinput76), 
        .A(n6627), .ZN(n6638) );
  INV_X1 U7547 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U7548 ( .A1(n6787), .A2(keyinput98), .B1(n6788), .B2(keyinput87), 
        .ZN(n6630) );
  OAI221_X1 U7549 ( .B1(n6787), .B2(keyinput98), .C1(n6788), .C2(keyinput87), 
        .A(n6630), .ZN(n6637) );
  INV_X1 U7550 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6795) );
  AOI22_X1 U7551 ( .A1(n6795), .A2(keyinput91), .B1(keyinput97), .B2(n6632), 
        .ZN(n6631) );
  OAI221_X1 U7552 ( .B1(n6795), .B2(keyinput91), .C1(n6632), .C2(keyinput97), 
        .A(n6631), .ZN(n6636) );
  INV_X1 U7553 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6634) );
  AOI22_X1 U7554 ( .A1(n6634), .A2(keyinput99), .B1(keyinput78), .B2(n3435), 
        .ZN(n6633) );
  OAI221_X1 U7555 ( .B1(n6634), .B2(keyinput99), .C1(n3435), .C2(keyinput78), 
        .A(n6633), .ZN(n6635) );
  NOR4_X1 U7556 ( .A1(n6638), .A2(n6637), .A3(n6636), .A4(n6635), .ZN(n6681)
         );
  INV_X1 U7557 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6640) );
  AOI22_X1 U7558 ( .A1(n6640), .A2(keyinput74), .B1(keyinput84), .B2(n6757), 
        .ZN(n6639) );
  OAI221_X1 U7559 ( .B1(n6640), .B2(keyinput74), .C1(n6757), .C2(keyinput84), 
        .A(n6639), .ZN(n6644) );
  XNOR2_X1 U7560 ( .A(n6641), .B(keyinput107), .ZN(n6643) );
  XOR2_X1 U7561 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .B(keyinput80), .Z(n6642)
         );
  OR3_X1 U7562 ( .A1(n6644), .A2(n6643), .A3(n6642), .ZN(n6651) );
  INV_X1 U7563 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6646) );
  INV_X1 U7564 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6758) );
  AOI22_X1 U7565 ( .A1(n6646), .A2(keyinput95), .B1(n6758), .B2(keyinput67), 
        .ZN(n6645) );
  OAI221_X1 U7566 ( .B1(n6646), .B2(keyinput95), .C1(n6758), .C2(keyinput67), 
        .A(n6645), .ZN(n6650) );
  INV_X1 U7567 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U7568 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(keyinput75), .B1(
        n6648), .B2(keyinput69), .ZN(n6647) );
  OAI221_X1 U7569 ( .B1(INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput75), .C1(
        n6648), .C2(keyinput69), .A(n6647), .ZN(n6649) );
  NOR3_X1 U7570 ( .A1(n6651), .A2(n6650), .A3(n6649), .ZN(n6680) );
  INV_X1 U7571 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6653) );
  AOI22_X1 U7572 ( .A1(n6653), .A2(keyinput88), .B1(keyinput122), .B2(n6779), 
        .ZN(n6652) );
  OAI221_X1 U7573 ( .B1(n6653), .B2(keyinput88), .C1(n6779), .C2(keyinput122), 
        .A(n6652), .ZN(n6662) );
  INV_X1 U7574 ( .A(DATAI_24_), .ZN(n6769) );
  INV_X1 U7575 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U7576 ( .A1(n6769), .A2(keyinput126), .B1(n6655), .B2(keyinput109), 
        .ZN(n6654) );
  OAI221_X1 U7577 ( .B1(n6769), .B2(keyinput126), .C1(n6655), .C2(keyinput109), 
        .A(n6654), .ZN(n6661) );
  XOR2_X1 U7578 ( .A(n6803), .B(keyinput72), .Z(n6659) );
  XNOR2_X1 U7579 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput108), .ZN(n6658) );
  XNOR2_X1 U7580 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(keyinput117), .ZN(
        n6657) );
  XNOR2_X1 U7581 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .B(keyinput92), .ZN(n6656) );
  NAND4_X1 U7582 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n6660)
         );
  NOR3_X1 U7583 ( .A1(n6662), .A2(n6661), .A3(n6660), .ZN(n6679) );
  AOI22_X1 U7584 ( .A1(n5128), .A2(keyinput123), .B1(keyinput66), .B2(n6664), 
        .ZN(n6663) );
  OAI221_X1 U7585 ( .B1(n5128), .B2(keyinput123), .C1(n6664), .C2(keyinput66), 
        .A(n6663), .ZN(n6677) );
  AOI22_X1 U7586 ( .A1(n6667), .A2(keyinput82), .B1(keyinput77), .B2(n6666), 
        .ZN(n6665) );
  OAI221_X1 U7587 ( .B1(n6667), .B2(keyinput82), .C1(n6666), .C2(keyinput77), 
        .A(n6665), .ZN(n6676) );
  AOI22_X1 U7588 ( .A1(n6670), .A2(keyinput70), .B1(keyinput100), .B2(n6669), 
        .ZN(n6668) );
  OAI221_X1 U7589 ( .B1(n6670), .B2(keyinput70), .C1(n6669), .C2(keyinput100), 
        .A(n6668), .ZN(n6675) );
  INV_X1 U7590 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6672) );
  AOI22_X1 U7591 ( .A1(n6673), .A2(keyinput125), .B1(n6672), .B2(keyinput115), 
        .ZN(n6671) );
  OAI221_X1 U7592 ( .B1(n6673), .B2(keyinput125), .C1(n6672), .C2(keyinput115), 
        .A(n6671), .ZN(n6674) );
  NOR4_X1 U7593 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6678)
         );
  NAND4_X1 U7594 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6817)
         );
  AOI22_X1 U7595 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput89), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput93), .ZN(n6682) );
  OAI221_X1 U7596 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput89), .C1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput93), .A(n6682), .ZN(n6689)
         );
  AOI22_X1 U7597 ( .A1(EAX_REG_29__SCAN_IN), .A2(keyinput114), .B1(
        INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput121), .ZN(n6683) );
  OAI221_X1 U7598 ( .B1(EAX_REG_29__SCAN_IN), .B2(keyinput114), .C1(
        INSTQUEUE_REG_13__0__SCAN_IN), .C2(keyinput121), .A(n6683), .ZN(n6688)
         );
  AOI22_X1 U7599 ( .A1(DATAI_6_), .A2(keyinput83), .B1(BS16_N), .B2(keyinput79), .ZN(n6684) );
  OAI221_X1 U7600 ( .B1(DATAI_6_), .B2(keyinput83), .C1(BS16_N), .C2(
        keyinput79), .A(n6684), .ZN(n6687) );
  AOI22_X1 U7601 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput127), .B1(
        INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput85), .ZN(n6685) );
  OAI221_X1 U7602 ( .B1(INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput127), .C1(
        INSTQUEUE_REG_13__5__SCAN_IN), .C2(keyinput85), .A(n6685), .ZN(n6686)
         );
  NOR4_X1 U7603 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n6717)
         );
  AOI22_X1 U7604 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput90), .B1(
        INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput113), .ZN(n6690) );
  OAI221_X1 U7605 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput90), 
        .C1(INSTQUEUE_REG_8__1__SCAN_IN), .C2(keyinput113), .A(n6690), .ZN(
        n6697) );
  AOI22_X1 U7606 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput104), .B1(
        STATE2_REG_1__SCAN_IN), .B2(keyinput73), .ZN(n6691) );
  OAI221_X1 U7607 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput104), .C1(
        STATE2_REG_1__SCAN_IN), .C2(keyinput73), .A(n6691), .ZN(n6696) );
  AOI22_X1 U7608 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(keyinput86), .B1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput112), .ZN(n6692) );
  OAI221_X1 U7609 ( .B1(DATAWIDTH_REG_28__SCAN_IN), .B2(keyinput86), .C1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput112), .A(n6692), .ZN(
        n6695) );
  AOI22_X1 U7610 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(keyinput124), 
        .B1(INSTQUEUE_REG_7__4__SCAN_IN), .B2(keyinput81), .ZN(n6693) );
  OAI221_X1 U7611 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(keyinput124), 
        .C1(INSTQUEUE_REG_7__4__SCAN_IN), .C2(keyinput81), .A(n6693), .ZN(
        n6694) );
  NOR4_X1 U7612 ( .A1(n6697), .A2(n6696), .A3(n6695), .A4(n6694), .ZN(n6716)
         );
  AOI22_X1 U7613 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput106), .B1(
        DATAO_REG_3__SCAN_IN), .B2(keyinput101), .ZN(n6698) );
  OAI221_X1 U7614 ( .B1(DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput106), .C1(
        DATAO_REG_3__SCAN_IN), .C2(keyinput101), .A(n6698), .ZN(n6705) );
  AOI22_X1 U7615 ( .A1(EAX_REG_12__SCAN_IN), .A2(keyinput116), .B1(
        EBX_REG_30__SCAN_IN), .B2(keyinput64), .ZN(n6699) );
  OAI221_X1 U7616 ( .B1(EAX_REG_12__SCAN_IN), .B2(keyinput116), .C1(
        EBX_REG_30__SCAN_IN), .C2(keyinput64), .A(n6699), .ZN(n6704) );
  AOI22_X1 U7617 ( .A1(DATAO_REG_8__SCAN_IN), .A2(keyinput96), .B1(
        INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput105), .ZN(n6700) );
  OAI221_X1 U7618 ( .B1(DATAO_REG_8__SCAN_IN), .B2(keyinput96), .C1(
        INSTQUEUE_REG_5__0__SCAN_IN), .C2(keyinput105), .A(n6700), .ZN(n6703)
         );
  AOI22_X1 U7619 ( .A1(UWORD_REG_5__SCAN_IN), .A2(keyinput103), .B1(
        EBX_REG_2__SCAN_IN), .B2(keyinput68), .ZN(n6701) );
  OAI221_X1 U7620 ( .B1(UWORD_REG_5__SCAN_IN), .B2(keyinput103), .C1(
        EBX_REG_2__SCAN_IN), .C2(keyinput68), .A(n6701), .ZN(n6702) );
  NOR4_X1 U7621 ( .A1(n6705), .A2(n6704), .A3(n6703), .A4(n6702), .ZN(n6715)
         );
  AOI22_X1 U7622 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput71), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput102), .ZN(n6706) );
  OAI221_X1 U7623 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput71), .C1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput102), .A(n6706), .ZN(
        n6713) );
  AOI22_X1 U7624 ( .A1(ADDRESS_REG_2__SCAN_IN), .A2(keyinput94), .B1(
        EAX_REG_17__SCAN_IN), .B2(keyinput110), .ZN(n6707) );
  OAI221_X1 U7625 ( .B1(ADDRESS_REG_2__SCAN_IN), .B2(keyinput94), .C1(
        EAX_REG_17__SCAN_IN), .C2(keyinput110), .A(n6707), .ZN(n6712) );
  AOI22_X1 U7626 ( .A1(EBX_REG_1__SCAN_IN), .A2(keyinput111), .B1(
        INSTADDRPOINTER_REG_26__SCAN_IN), .B2(keyinput119), .ZN(n6708) );
  OAI221_X1 U7627 ( .B1(EBX_REG_1__SCAN_IN), .B2(keyinput111), .C1(
        INSTADDRPOINTER_REG_26__SCAN_IN), .C2(keyinput119), .A(n6708), .ZN(
        n6711) );
  AOI22_X1 U7628 ( .A1(DATAO_REG_4__SCAN_IN), .A2(keyinput118), .B1(
        EBX_REG_5__SCAN_IN), .B2(keyinput120), .ZN(n6709) );
  OAI221_X1 U7629 ( .B1(DATAO_REG_4__SCAN_IN), .B2(keyinput118), .C1(
        EBX_REG_5__SCAN_IN), .C2(keyinput120), .A(n6709), .ZN(n6710) );
  NOR4_X1 U7630 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6714)
         );
  NAND4_X1 U7631 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6816)
         );
  OAI22_X1 U7632 ( .A1(EBX_REG_30__SCAN_IN), .A2(keyinput0), .B1(
        INSTADDRPOINTER_REG_16__SCAN_IN), .B2(keyinput60), .ZN(n6718) );
  AOI221_X1 U7633 ( .B1(EBX_REG_30__SCAN_IN), .B2(keyinput0), .C1(keyinput60), 
        .C2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6718), .ZN(n6725) );
  OAI22_X1 U7634 ( .A1(EBX_REG_1__SCAN_IN), .A2(keyinput47), .B1(keyinput42), 
        .B2(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6719) );
  AOI221_X1 U7635 ( .B1(EBX_REG_1__SCAN_IN), .B2(keyinput47), .C1(
        DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput42), .A(n6719), .ZN(n6724) );
  OAI22_X1 U7636 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(keyinput38), .B1(
        keyinput40), .B2(REIP_REG_20__SCAN_IN), .ZN(n6720) );
  AOI221_X1 U7637 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput38), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput40), .A(n6720), .ZN(n6723) );
  OAI22_X1 U7638 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(keyinput11), .B1(
        INSTADDRPOINTER_REG_26__SCAN_IN), .B2(keyinput55), .ZN(n6721) );
  AOI221_X1 U7639 ( .B1(INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput11), .C1(
        keyinput55), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6721), .ZN(
        n6722) );
  NAND4_X1 U7640 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n6753)
         );
  OAI22_X1 U7641 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(keyinput10), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput2), .ZN(n6726) );
  AOI221_X1 U7642 ( .B1(INSTQUEUE_REG_2__7__SCAN_IN), .B2(keyinput10), .C1(
        keyinput2), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n6726), .ZN(n6733) );
  OAI22_X1 U7643 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(keyinput49), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput32), .ZN(n6727) );
  AOI221_X1 U7644 ( .B1(INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput49), .C1(
        keyinput32), .C2(DATAO_REG_8__SCAN_IN), .A(n6727), .ZN(n6732) );
  OAI22_X1 U7645 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(keyinput41), .B1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput26), .ZN(n6728) );
  AOI221_X1 U7646 ( .B1(INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput41), .C1(
        keyinput26), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n6728), .ZN(
        n6731) );
  OAI22_X1 U7647 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(keyinput31), .B1(
        REIP_REG_16__SCAN_IN), .B2(keyinput7), .ZN(n6729) );
  AOI221_X1 U7648 ( .B1(INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput31), .C1(
        keyinput7), .C2(REIP_REG_16__SCAN_IN), .A(n6729), .ZN(n6730) );
  NAND4_X1 U7649 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n6752)
         );
  OAI22_X1 U7650 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(keyinput35), .B1(
        keyinput12), .B2(REIP_REG_22__SCAN_IN), .ZN(n6734) );
  AOI221_X1 U7651 ( .B1(INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput35), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput12), .A(n6734), .ZN(n6741) );
  OAI22_X1 U7652 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(keyinput45), .B1(
        keyinput43), .B2(ADS_N_REG_SCAN_IN), .ZN(n6735) );
  AOI221_X1 U7653 ( .B1(INSTQUEUE_REG_15__2__SCAN_IN), .B2(keyinput45), .C1(
        ADS_N_REG_SCAN_IN), .C2(keyinput43), .A(n6735), .ZN(n6740) );
  OAI22_X1 U7654 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(keyinput24), .B1(
        keyinput48), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6736) );
  AOI221_X1 U7655 ( .B1(INSTQUEUE_REG_6__2__SCAN_IN), .B2(keyinput24), .C1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput48), .A(n6736), .ZN(
        n6739) );
  OAI22_X1 U7656 ( .A1(DATAI_6_), .A2(keyinput19), .B1(UWORD_REG_5__SCAN_IN), 
        .B2(keyinput39), .ZN(n6737) );
  AOI221_X1 U7657 ( .B1(DATAI_6_), .B2(keyinput19), .C1(keyinput39), .C2(
        UWORD_REG_5__SCAN_IN), .A(n6737), .ZN(n6738) );
  NAND4_X1 U7658 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n6751)
         );
  OAI22_X1 U7659 ( .A1(EBX_REG_5__SCAN_IN), .A2(keyinput56), .B1(keyinput6), 
        .B2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6742) );
  AOI221_X1 U7660 ( .B1(EBX_REG_5__SCAN_IN), .B2(keyinput56), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput6), .A(n6742), .ZN(n6749) );
  OAI22_X1 U7661 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(keyinput5), .B1(
        EBX_REG_10__SCAN_IN), .B2(keyinput18), .ZN(n6743) );
  AOI221_X1 U7662 ( .B1(INSTQUEUE_REG_12__5__SCAN_IN), .B2(keyinput5), .C1(
        keyinput18), .C2(EBX_REG_10__SCAN_IN), .A(n6743), .ZN(n6748) );
  OAI22_X1 U7663 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput53), .B1(
        keyinput13), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6744) );
  AOI221_X1 U7664 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput53), .C1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput13), .A(n6744), .ZN(n6747) );
  OAI22_X1 U7665 ( .A1(EAX_REG_17__SCAN_IN), .A2(keyinput46), .B1(keyinput1), 
        .B2(DATAI_25_), .ZN(n6745) );
  AOI221_X1 U7666 ( .B1(EAX_REG_17__SCAN_IN), .B2(keyinput46), .C1(DATAI_25_), 
        .C2(keyinput1), .A(n6745), .ZN(n6746) );
  NAND4_X1 U7667 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(n6750)
         );
  NOR4_X1 U7668 ( .A1(n6753), .A2(n6752), .A3(n6751), .A4(n6750), .ZN(n6815)
         );
  AOI22_X1 U7669 ( .A1(n3435), .A2(keyinput14), .B1(keyinput50), .B2(n6755), 
        .ZN(n6754) );
  OAI221_X1 U7670 ( .B1(n3435), .B2(keyinput14), .C1(n6755), .C2(keyinput50), 
        .A(n6754), .ZN(n6765) );
  AOI22_X1 U7671 ( .A1(n6758), .A2(keyinput3), .B1(keyinput20), .B2(n6757), 
        .ZN(n6756) );
  OAI221_X1 U7672 ( .B1(n6758), .B2(keyinput3), .C1(n6757), .C2(keyinput20), 
        .A(n6756), .ZN(n6764) );
  XNOR2_X1 U7673 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput61), .ZN(n6762) );
  XNOR2_X1 U7674 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .B(keyinput17), .ZN(n6761)
         );
  XNOR2_X1 U7675 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .B(keyinput16), .ZN(n6760) );
  XNOR2_X1 U7676 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput25), .ZN(n6759) );
  NAND4_X1 U7677 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6763)
         );
  NOR3_X1 U7678 ( .A1(n6765), .A2(n6764), .A3(n6763), .ZN(n6813) );
  AOI22_X1 U7679 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(keyinput29), .B1(
        INSTQUEUE_REG_3__4__SCAN_IN), .B2(keyinput51), .ZN(n6766) );
  OAI221_X1 U7680 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput29), .C1(
        INSTQUEUE_REG_3__4__SCAN_IN), .C2(keyinput51), .A(n6766), .ZN(n6776)
         );
  AOI22_X1 U7681 ( .A1(DATAO_REG_3__SCAN_IN), .A2(keyinput37), .B1(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(keyinput33), .ZN(n6767) );
  OAI221_X1 U7682 ( .B1(DATAO_REG_3__SCAN_IN), .B2(keyinput37), .C1(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(keyinput33), .A(n6767), .ZN(
        n6775) );
  AOI22_X1 U7683 ( .A1(n6770), .A2(keyinput63), .B1(keyinput62), .B2(n6769), 
        .ZN(n6768) );
  OAI221_X1 U7684 ( .B1(n6770), .B2(keyinput63), .C1(n6769), .C2(keyinput62), 
        .A(n6768), .ZN(n6774) );
  INV_X1 U7685 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U7686 ( .A1(DATAO_REG_20__SCAN_IN), .A2(keyinput36), .B1(n6772), 
        .B2(keyinput21), .ZN(n6771) );
  OAI221_X1 U7687 ( .B1(DATAO_REG_20__SCAN_IN), .B2(keyinput36), .C1(n6772), 
        .C2(keyinput21), .A(n6771), .ZN(n6773) );
  NOR4_X1 U7688 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6812)
         );
  INV_X1 U7689 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6778) );
  AOI22_X1 U7690 ( .A1(n6778), .A2(keyinput57), .B1(keyinput59), .B2(n5128), 
        .ZN(n6777) );
  OAI221_X1 U7691 ( .B1(n6778), .B2(keyinput57), .C1(n5128), .C2(keyinput59), 
        .A(n6777), .ZN(n6781) );
  XNOR2_X1 U7692 ( .A(n6779), .B(keyinput58), .ZN(n6780) );
  NOR2_X1 U7693 ( .A1(n6781), .A2(n6780), .ZN(n6793) );
  INV_X1 U7694 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6783) );
  AOI22_X1 U7695 ( .A1(n6784), .A2(keyinput9), .B1(keyinput54), .B2(n6783), 
        .ZN(n6782) );
  OAI221_X1 U7696 ( .B1(n6784), .B2(keyinput9), .C1(n6783), .C2(keyinput54), 
        .A(n6782), .ZN(n6785) );
  INV_X1 U7697 ( .A(n6785), .ZN(n6792) );
  AOI22_X1 U7698 ( .A1(n6788), .A2(keyinput23), .B1(keyinput34), .B2(n6787), 
        .ZN(n6786) );
  OAI221_X1 U7699 ( .B1(n6788), .B2(keyinput23), .C1(n6787), .C2(keyinput34), 
        .A(n6786), .ZN(n6789) );
  INV_X1 U7700 ( .A(n6789), .ZN(n6791) );
  XNOR2_X1 U7701 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .B(keyinput28), .ZN(n6790) );
  AND4_X1 U7702 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6811)
         );
  INV_X1 U7703 ( .A(BS16_N), .ZN(n6796) );
  AOI22_X1 U7704 ( .A1(n6796), .A2(keyinput15), .B1(n6795), .B2(keyinput27), 
        .ZN(n6794) );
  OAI221_X1 U7705 ( .B1(n6796), .B2(keyinput15), .C1(n6795), .C2(keyinput27), 
        .A(n6794), .ZN(n6800) );
  XOR2_X1 U7706 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput44), .Z(n6799)
         );
  XNOR2_X1 U7707 ( .A(n6797), .B(keyinput22), .ZN(n6798) );
  OR3_X1 U7708 ( .A1(n6800), .A2(n6799), .A3(n6798), .ZN(n6809) );
  AOI22_X1 U7709 ( .A1(n6803), .A2(keyinput8), .B1(keyinput52), .B2(n6802), 
        .ZN(n6801) );
  OAI221_X1 U7710 ( .B1(n6803), .B2(keyinput8), .C1(n6802), .C2(keyinput52), 
        .A(n6801), .ZN(n6808) );
  AOI22_X1 U7711 ( .A1(n6806), .A2(keyinput30), .B1(n6805), .B2(keyinput4), 
        .ZN(n6804) );
  OAI221_X1 U7712 ( .B1(n6806), .B2(keyinput30), .C1(n6805), .C2(keyinput4), 
        .A(n6804), .ZN(n6807) );
  NOR3_X1 U7713 ( .A1(n6809), .A2(n6808), .A3(n6807), .ZN(n6810) );
  AND4_X1 U7714 ( .A1(n6813), .A2(n6812), .A3(n6811), .A4(n6810), .ZN(n6814)
         );
  OAI211_X1 U7715 ( .C1(n6817), .C2(n6816), .A(n6815), .B(n6814), .ZN(n6818)
         );
  XNOR2_X1 U7716 ( .A(n6819), .B(n6818), .ZN(U2870) );
  NAND4_X2 U34700 ( .A1(n3153), .A2(n3156), .A3(n3154), .A4(n3155), .ZN(n3272)
         );
  CLKBUF_X1 U34680 ( .A(n3316), .Z(n3024) );
  INV_X2 U3480 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4454) );
  AND4_X1 U3490 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n3136)
         );
  CLKBUF_X1 U3605 ( .A(n5466), .Z(n5467) );
  CLKBUF_X1 U4134 ( .A(n4372), .Z(n3023) );
  CLKBUF_X1 U6600 ( .A(n3791), .Z(n3792) );
endmodule

