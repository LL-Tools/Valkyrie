

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5022, n5023, n5024, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135;

  AOI222_X1 U5087 ( .A1(n9810), .A2(n10993), .B1(n10992), .B2(n10990), .C1(
        n10998), .C2(n7335), .ZN(n10951) );
  INV_X4 U5088 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OR2_X1 U5089 ( .A1(n6243), .A2(n6242), .ZN(n9257) );
  NAND2_X2 U5090 ( .A1(n8400), .A2(n8399), .ZN(n10067) );
  INV_X1 U5091 ( .A(n6226), .ZN(n6311) );
  AND2_X1 U5092 ( .A1(n6701), .A2(n6700), .ZN(n6830) );
  INV_X2 U5093 ( .A(n7237), .ZN(n9039) );
  INV_X2 U5094 ( .A(n8826), .ZN(n8848) );
  XNOR2_X1 U5095 ( .A(n5959), .B(n5958), .ZN(n7290) );
  NAND4_X2 U5096 ( .A1(n6599), .A2(n6598), .A3(n6597), .A4(n6596), .ZN(n7085)
         );
  INV_X1 U5097 ( .A(n6681), .ZN(n8320) );
  NOR2_X1 U5098 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5771) );
  NOR2_X1 U5099 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n6497) );
  AOI222_X1 U5100 ( .A1(n10998), .A2(n7190), .B1(n10863), .B2(n10990), .C1(
        n9812), .C2(n10993), .ZN(n10823) );
  AOI222_X1 U5101 ( .A1(n10998), .A2(n9921), .B1(n9920), .B2(n10990), .C1(
        n9954), .C2(n10993), .ZN(n10080) );
  AOI222_X1 U5102 ( .A1(n10998), .A2(n9894), .B1(n9893), .B2(n10990), .C1(
        n9920), .C2(n10993), .ZN(n10070) );
  NAND2_X2 U5103 ( .A1(n7113), .A2(n7112), .ZN(n10998) );
  AND2_X2 U5104 ( .A1(n8744), .A2(n9816), .ZN(n10990) );
  NAND2_X1 U5105 ( .A1(n7263), .A2(n7264), .ZN(n8889) );
  INV_X2 U5106 ( .A(n8447), .ZN(n8546) );
  INV_X1 U5107 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10552) );
  AND2_X1 U5108 ( .A1(n6379), .A2(n6378), .ZN(n6445) );
  INV_X1 U5109 ( .A(n5922), .ZN(n8834) );
  INV_X1 U5110 ( .A(n7255), .ZN(n10852) );
  OAI21_X1 U5112 ( .B1(n7956), .B2(n5032), .A(n5624), .ZN(n8141) );
  NAND2_X1 U5113 ( .A1(n8805), .A2(n8795), .ZN(n7153) );
  INV_X2 U5114 ( .A(n6680), .ZN(n5752) );
  INV_X2 U5115 ( .A(n11019), .ZN(n11014) );
  XNOR2_X1 U5116 ( .A(n5882), .B(n5881), .ZN(n7063) );
  NAND2_X1 U5117 ( .A1(n6473), .A2(n6472), .ZN(n5022) );
  OR2_X1 U5118 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5023) );
  NAND2_X1 U5119 ( .A1(n6636), .A2(n7593), .ZN(n7101) );
  INV_X1 U5120 ( .A(n9188), .ZN(n5345) );
  XNOR2_X2 U5121 ( .A(n6406), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6636) );
  INV_X2 U5122 ( .A(n6472), .ZN(n10145) );
  XNOR2_X2 U5123 ( .A(n7197), .B(n7085), .ZN(n7186) );
  OAI211_X2 U5124 ( .C1(n7291), .C2(n6658), .A(n6928), .B(n6927), .ZN(n7275)
         );
  NAND2_X2 U5125 ( .A1(n5970), .A2(n5969), .ZN(n7768) );
  INV_X1 U5126 ( .A(n7275), .ZN(n10894) );
  XNOR2_X2 U5127 ( .A(n6390), .B(n6389), .ZN(n8023) );
  NAND2_X2 U5128 ( .A1(n7065), .A2(n7064), .ZN(n10935) );
  XNOR2_X2 U5129 ( .A(n6285), .B(n6284), .ZN(n8412) );
  AND2_X2 U5130 ( .A1(n7593), .A2(n9926), .ZN(n6877) );
  AND2_X1 U5131 ( .A1(n5049), .A2(n5186), .ZN(n5882) );
  NOR4_X2 U5132 ( .A1(n8796), .A2(n8774), .A3(n8772), .A4(n8773), .ZN(n8776)
         );
  OAI222_X1 U5133 ( .A1(n6750), .A2(n9691), .B1(n9684), .B2(n7063), .C1(n6461), 
        .C2(n9687), .ZN(P2_U3352) );
  OAI222_X1 U5134 ( .A1(n10144), .A2(n10543), .B1(n10147), .B2(n7063), .C1(
        P1_U3084), .C2(n6460), .ZN(P1_U3347) );
  OR2_X1 U5135 ( .A1(n7063), .A2(n8447), .ZN(n7065) );
  NAND2_X2 U5136 ( .A1(n7294), .A2(n7293), .ZN(n10967) );
  XNOR2_X2 U5137 ( .A(n5809), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10778) );
  NAND2_X1 U5138 ( .A1(n9905), .A2(n8711), .ZN(n9891) );
  AOI21_X1 U5139 ( .B1(n9919), .B2(n5380), .A(n5379), .ZN(n5378) );
  NAND2_X1 U5140 ( .A1(n7107), .A2(n8577), .ZN(n10859) );
  NAND2_X2 U5141 ( .A1(n5806), .A2(n9034), .ZN(n6226) );
  INV_X4 U5142 ( .A(n9157), .ZN(n9152) );
  INV_X1 U5143 ( .A(n9811), .ZN(n7104) );
  NAND2_X1 U5144 ( .A1(n5639), .A2(n6837), .ZN(n5603) );
  NAND3_X2 U5145 ( .A1(n6689), .A2(n7153), .A3(n6688), .ZN(n7103) );
  INV_X2 U5146 ( .A(n9128), .ZN(n6825) );
  AND2_X4 U5147 ( .A1(n9172), .A2(n10145), .ZN(n6834) );
  INV_X1 U5148 ( .A(n8880), .ZN(n9034) );
  NAND2_X1 U5149 ( .A1(n5649), .A2(n5829), .ZN(n5651) );
  AND2_X1 U5150 ( .A1(n5598), .A2(n5767), .ZN(n5597) );
  AND2_X1 U5151 ( .A1(n5769), .A2(n5599), .ZN(n5598) );
  AOI211_X1 U5152 ( .C1(n11009), .C2(n10058), .A(n8507), .B(n8506), .ZN(n8508)
         );
  AND2_X1 U5153 ( .A1(n10059), .A2(n5268), .ZN(n5267) );
  OAI21_X1 U5154 ( .B1(n8810), .B2(n8809), .A(n8808), .ZN(n5105) );
  AND2_X1 U5155 ( .A1(n8502), .A2(n5269), .ZN(n10060) );
  AOI21_X1 U5156 ( .B1(n8505), .B2(n11062), .A(n5270), .ZN(n5269) );
  OAI21_X1 U5157 ( .B1(n5491), .B2(n9047), .A(n9046), .ZN(n5489) );
  AND2_X1 U5158 ( .A1(n8495), .A2(n8494), .ZN(n8505) );
  OAI21_X1 U5159 ( .B1(n8845), .B2(n8855), .A(n8844), .ZN(n8846) );
  NAND2_X1 U5160 ( .A1(n9891), .A2(n9892), .ZN(n9890) );
  NAND2_X1 U5161 ( .A1(n5609), .A2(n5608), .ZN(n9931) );
  OAI21_X1 U5162 ( .B1(n5109), .B2(n9915), .A(n5378), .ZN(n9906) );
  NAND2_X1 U5163 ( .A1(n5109), .A2(n8624), .ZN(n9918) );
  AOI21_X1 U5164 ( .B1(n9939), .B2(n5378), .A(n5376), .ZN(n5375) );
  INV_X1 U5165 ( .A(n8789), .ZN(n8726) );
  AOI21_X1 U5166 ( .B1(n9094), .B2(n9093), .A(n9092), .ZN(n9099) );
  NAND2_X1 U5167 ( .A1(n9951), .A2(n8619), .ZN(n9940) );
  AOI21_X1 U5168 ( .B1(n5345), .B2(n5402), .A(n5066), .ZN(n5401) );
  INV_X1 U5169 ( .A(n9015), .ZN(n5402) );
  NAND2_X1 U5170 ( .A1(n5377), .A2(n9907), .ZN(n5376) );
  NAND2_X1 U5171 ( .A1(n8548), .A2(n8547), .ZN(n10049) );
  NAND2_X1 U5172 ( .A1(n5378), .A2(n9915), .ZN(n5377) );
  NAND2_X1 U5173 ( .A1(n8423), .A2(n8422), .ZN(n10057) );
  NAND2_X1 U5174 ( .A1(n5789), .A2(n5788), .ZN(n9595) );
  AND2_X1 U5175 ( .A1(n8769), .A2(n5602), .ZN(n5601) );
  AND2_X1 U5176 ( .A1(n10067), .A2(n9740), .ZN(n8610) );
  XNOR2_X1 U5177 ( .A(n5763), .B(n8439), .ZN(n8420) );
  NAND2_X1 U5178 ( .A1(n8387), .A2(n8386), .ZN(n10072) );
  NAND2_X1 U5179 ( .A1(n5568), .A2(n7733), .ZN(n8015) );
  AND2_X1 U5180 ( .A1(n7732), .A2(n5051), .ZN(n5568) );
  NAND2_X1 U5181 ( .A1(n8350), .A2(n8349), .ZN(n10087) );
  NAND2_X1 U5182 ( .A1(n8336), .A2(n8335), .ZN(n10093) );
  NAND2_X1 U5183 ( .A1(n6155), .A2(n6154), .ZN(n9642) );
  NAND2_X1 U5184 ( .A1(n8249), .A2(n8248), .ZN(n10112) );
  NAND2_X1 U5185 ( .A1(n6136), .A2(n6135), .ZN(n9645) );
  NAND2_X1 U5186 ( .A1(n6119), .A2(n6118), .ZN(n9653) );
  OAI21_X1 U5187 ( .B1(n6058), .B2(n5702), .A(n5701), .ZN(n6077) );
  AND2_X1 U5188 ( .A1(n7146), .A2(n7095), .ZN(n7097) );
  AND2_X1 U5189 ( .A1(n8932), .A2(n8928), .ZN(n8864) );
  NAND2_X1 U5190 ( .A1(n7637), .A2(n7636), .ZN(n11054) );
  AND2_X1 U5191 ( .A1(n8588), .A2(n8591), .ZN(n8751) );
  OAI21_X1 U5192 ( .B1(n6025), .B2(n6024), .A(n5693), .ZN(n6040) );
  NAND2_X1 U5193 ( .A1(n10859), .A2(n7108), .ZN(n7109) );
  NAND2_X1 U5194 ( .A1(n7203), .A2(n7202), .ZN(n7289) );
  NAND2_X2 U5195 ( .A1(n7229), .A2(n7237), .ZN(n5834) );
  AND3_X1 U5196 ( .A1(n5906), .A2(n5905), .A3(n5904), .ZN(n7473) );
  XNOR2_X1 U5197 ( .A(n5933), .B(n5932), .ZN(n7200) );
  NAND2_X1 U5198 ( .A1(n7188), .A2(n7105), .ZN(n8581) );
  NAND2_X1 U5199 ( .A1(n5133), .A2(n5668), .ZN(n5933) );
  NAND2_X1 U5200 ( .A1(n7186), .A2(n7189), .ZN(n7188) );
  AND3_X1 U5201 ( .A1(n5876), .A2(n5875), .A3(n5874), .ZN(n10904) );
  NAND4_X2 U5202 ( .A1(n6709), .A2(n6708), .A3(n6707), .A4(n6706), .ZN(n10863)
         );
  NAND4_X1 U5203 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6938), .ZN(n9811)
         );
  NAND4_X1 U5204 ( .A1(n6901), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n10862)
         );
  NAND4_X1 U5205 ( .A1(n7222), .A2(n7221), .A3(n7220), .A4(n7219), .ZN(n10992)
         );
  CLKBUF_X3 U5206 ( .A(n6825), .Z(n9143) );
  AND2_X2 U5207 ( .A1(n6642), .A2(n6637), .ZN(n9159) );
  NAND2_X1 U5208 ( .A1(n5801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U5209 ( .A1(n6834), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6597) );
  INV_X1 U5210 ( .A(n7381), .ZN(n9054) );
  OR2_X1 U5211 ( .A1(n7101), .A2(n6638), .ZN(n9128) );
  AND4_X1 U5212 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n8486)
         );
  AND2_X1 U5213 ( .A1(n6473), .A2(n10145), .ZN(n6833) );
  OAI211_X1 U5214 ( .C1(n8447), .C2(n6824), .A(n6823), .B(n5045), .ZN(n7183)
         );
  AND4_X1 U5215 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), .ZN(n7381)
         );
  NAND2_X1 U5216 ( .A1(n6683), .A2(n5237), .ZN(n7197) );
  NAND2_X1 U5217 ( .A1(n6393), .A2(n6431), .ZN(n6879) );
  INV_X2 U5218 ( .A(n6600), .ZN(n5024) );
  NAND2_X4 U5219 ( .A1(n6355), .A2(n9690), .ZN(n6743) );
  AND2_X1 U5220 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  AND2_X1 U5221 ( .A1(n7780), .A2(n8843), .ZN(n8880) );
  MUX2_X1 U5222 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6469), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n6471) );
  NAND2_X1 U5223 ( .A1(n6470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U5224 ( .A1(n5787), .A2(n5786), .ZN(n9690) );
  NAND2_X1 U5225 ( .A1(n6468), .A2(n6414), .ZN(n9816) );
  NAND2_X1 U5226 ( .A1(n5817), .A2(n9680), .ZN(n9686) );
  NAND2_X1 U5227 ( .A1(n6419), .A2(n6418), .ZN(n10675) );
  XNOR2_X1 U5228 ( .A(n6606), .B(n10353), .ZN(n7593) );
  MUX2_X1 U5229 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5815), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5817) );
  XNOR2_X1 U5230 ( .A(n5651), .B(n10436), .ZN(n5808) );
  MUX2_X1 U5231 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5785), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5787) );
  NAND2_X2 U5232 ( .A1(n6680), .A2(P2_U3152), .ZN(n9684) );
  XNOR2_X1 U5233 ( .A(n6607), .B(n10568), .ZN(n9926) );
  AND2_X1 U5234 ( .A1(n5597), .A2(n5159), .ZN(n5158) );
  INV_X1 U5235 ( .A(n5902), .ZN(n5768) );
  INV_X1 U5236 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6570) );
  INV_X1 U5237 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10565) );
  INV_X1 U5238 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10568) );
  INV_X1 U5239 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10353) );
  INV_X1 U5240 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9849) );
  NOR2_X1 U5241 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6375) );
  INV_X1 U5242 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10190) );
  NOR2_X1 U5243 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6378) );
  NOR2_X1 U5244 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6379) );
  INV_X1 U5245 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10572) );
  INV_X1 U5246 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5797) );
  INV_X1 U5247 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6078) );
  AOI21_X1 U5248 ( .B1(n9727), .B2(n9724), .A(n9723), .ZN(n9768) );
  INV_X4 U5250 ( .A(n5022), .ZN(n5026) );
  INV_X1 U5251 ( .A(n7237), .ZN(n5027) );
  INV_X4 U5252 ( .A(n5947), .ZN(n5921) );
  NAND2_X1 U5253 ( .A1(n5819), .A2(n9686), .ZN(n5947) );
  OAI211_X2 U5254 ( .C1(n8826), .C2(n7063), .A(n5886), .B(n5885), .ZN(n8916)
         );
  OR2_X4 U5255 ( .A1(n6315), .A2(n9034), .ZN(n7237) );
  NAND2_X4 U5256 ( .A1(n5336), .A2(n5818), .ZN(n6365) );
  NAND2_X1 U5257 ( .A1(n5806), .A2(n9034), .ZN(n5028) );
  OAI21_X2 U5258 ( .B1(n5588), .B2(n5587), .A(n5591), .ZN(n9205) );
  NAND2_X2 U5259 ( .A1(n8307), .A2(n10922), .ZN(n6315) );
  INV_X1 U5260 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5767) );
  INV_X1 U5261 ( .A(SI_13_), .ZN(n5694) );
  XNOR2_X1 U5262 ( .A(n9595), .B(n9213), .ZN(n9188) );
  NAND2_X1 U5263 ( .A1(n5209), .A2(n8659), .ZN(n8666) );
  OAI21_X1 U5264 ( .B1(n8655), .B2(n8654), .A(n5072), .ZN(n5209) );
  AND2_X1 U5265 ( .A1(n9002), .A2(n5166), .ZN(n5165) );
  INV_X1 U5266 ( .A(SI_16_), .ZN(n10217) );
  AOI21_X1 U5267 ( .B1(n5583), .B2(n5586), .A(n5037), .ZN(n5581) );
  OR2_X1 U5268 ( .A1(n6206), .A2(n10490), .ZN(n6232) );
  OAI21_X1 U5269 ( .B1(n8851), .B2(n9029), .A(n9024), .ZN(n8883) );
  OR2_X1 U5270 ( .A1(n9600), .A2(n9443), .ZN(n9015) );
  OR2_X1 U5271 ( .A1(n9653), .A2(n9573), .ZN(n9173) );
  OR2_X1 U5272 ( .A1(n7820), .A2(n7788), .ZN(n8933) );
  NAND2_X1 U5273 ( .A1(n11024), .A2(n9328), .ZN(n8928) );
  NAND2_X1 U5274 ( .A1(n7229), .A2(n10836), .ZN(n8890) );
  AND2_X1 U5275 ( .A1(n5317), .A2(n5776), .ZN(n5427) );
  INV_X1 U5276 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5769) );
  INV_X1 U5277 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U5278 ( .A1(n6326), .A2(n6325), .ZN(n6328) );
  NAND2_X1 U5279 ( .A1(n8800), .A2(n9926), .ZN(n5196) );
  NOR2_X1 U5280 ( .A1(n5397), .A2(n6383), .ZN(n6384) );
  INV_X1 U5281 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6381) );
  INV_X1 U5282 ( .A(n7958), .ZN(n5626) );
  INV_X1 U5283 ( .A(n5616), .ZN(n5615) );
  OAI21_X1 U5284 ( .B1(n8753), .B2(n5617), .A(n7533), .ZN(n5616) );
  NAND2_X1 U5285 ( .A1(n5484), .A2(n8533), .ZN(n8535) );
  AND2_X1 U5286 ( .A1(n6282), .A2(n5756), .ZN(n6281) );
  NAND2_X1 U5287 ( .A1(n5743), .A2(n5742), .ZN(n6223) );
  NAND2_X1 U5288 ( .A1(n5706), .A2(n5705), .ZN(n6097) );
  AND2_X1 U5289 ( .A1(n5698), .A2(n5697), .ZN(n6039) );
  AND2_X1 U5290 ( .A1(n6310), .A2(n6309), .ZN(n9213) );
  INV_X1 U5291 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5790) );
  INV_X1 U5292 ( .A(n5108), .ZN(n5968) );
  NAND2_X1 U5293 ( .A1(n9426), .A2(n9015), .ZN(n9411) );
  INV_X1 U5294 ( .A(n5360), .ZN(n5359) );
  AOI21_X1 U5295 ( .B1(n5361), .B2(n9182), .A(n9183), .ZN(n5360) );
  INV_X1 U5296 ( .A(n5365), .ZN(n5364) );
  OAI21_X1 U5297 ( .B1(n9182), .B2(n8988), .A(n9181), .ZN(n5365) );
  AND2_X1 U5298 ( .A1(n8870), .A2(n8273), .ZN(n5352) );
  NAND2_X1 U5299 ( .A1(n5948), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5994) );
  AOI21_X1 U5300 ( .B1(n5403), .B2(n5408), .A(n5034), .ZN(n5406) );
  INV_X1 U5301 ( .A(n5411), .ZN(n5403) );
  NAND2_X1 U5302 ( .A1(n5435), .A2(n5434), .ZN(n5433) );
  INV_X1 U5303 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5434) );
  INV_X1 U5304 ( .A(n5436), .ZN(n5435) );
  NAND2_X1 U5305 ( .A1(n5798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U5306 ( .A1(n8402), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U5307 ( .A1(n8525), .A2(n6636), .ZN(n6647) );
  INV_X1 U5308 ( .A(n8734), .ZN(n8739) );
  AOI21_X1 U5309 ( .B1(n8733), .B2(n8740), .A(n8788), .ZN(n8734) );
  MUX2_X1 U5310 ( .A(n8730), .B(n8729), .S(n8741), .Z(n8733) );
  INV_X1 U5311 ( .A(n7593), .ZN(n8801) );
  AND2_X1 U5312 ( .A1(n10048), .A2(n9800), .ZN(n8796) );
  INV_X1 U5313 ( .A(n5219), .ZN(n5217) );
  NOR2_X1 U5314 ( .A1(n9899), .A2(n10067), .ZN(n9875) );
  NOR2_X1 U5315 ( .A1(n5040), .A2(n7995), .ZN(n7992) );
  NAND2_X1 U5316 ( .A1(n6681), .A2(n5752), .ZN(n8447) );
  XNOR2_X1 U5317 ( .A(n6405), .B(n6404), .ZN(n6595) );
  INV_X1 U5318 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U5319 ( .A1(n6403), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U5320 ( .A1(n5571), .A2(n5570), .ZN(n6403) );
  NAND2_X1 U5321 ( .A1(n6653), .A2(n10879), .ZN(n9773) );
  NAND2_X1 U5322 ( .A1(n5452), .A2(n5451), .ZN(n5450) );
  AND2_X1 U5323 ( .A1(n10421), .A2(n10420), .ZN(n5451) );
  NAND2_X1 U5324 ( .A1(n10419), .A2(n10418), .ZN(n5452) );
  INV_X1 U5325 ( .A(keyinput_151), .ZN(n5448) );
  OAI21_X1 U5326 ( .B1(n10232), .B2(n10231), .A(n10230), .ZN(n10236) );
  XNOR2_X1 U5327 ( .A(n10229), .B(SI_9_), .ZN(n10230) );
  NAND2_X1 U5328 ( .A1(n5292), .A2(n5291), .ZN(n5290) );
  AOI22_X1 U5329 ( .A1(n10436), .A2(n10242), .B1(keyinput_31), .B2(SI_1_), 
        .ZN(n5291) );
  NAND2_X1 U5330 ( .A1(n5294), .A2(n5293), .ZN(n5292) );
  XNOR2_X1 U5331 ( .A(P2_U3152), .B(keyinput_34), .ZN(n5288) );
  INV_X1 U5332 ( .A(n10243), .ZN(n5289) );
  OAI21_X1 U5333 ( .B1(n5445), .B2(n10456), .A(n5443), .ZN(n10462) );
  INV_X1 U5334 ( .A(n5444), .ZN(n5443) );
  AOI21_X1 U5335 ( .B1(n10451), .B2(n10450), .A(n5446), .ZN(n5445) );
  AND2_X1 U5336 ( .A1(n5303), .A2(n5302), .ZN(n5301) );
  NAND2_X1 U5337 ( .A1(n10273), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U5338 ( .A1(n10483), .A2(keyinput_52), .ZN(n5303) );
  NAND2_X1 U5339 ( .A1(n5306), .A2(n5305), .ZN(n5304) );
  NAND2_X1 U5340 ( .A1(keyinput_51), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5305)
         );
  NAND2_X1 U5341 ( .A1(n10480), .A2(n10272), .ZN(n5306) );
  AOI21_X1 U5342 ( .B1(n10488), .B2(keyinput_183), .A(n10487), .ZN(n5466) );
  OAI21_X1 U5343 ( .B1(n5472), .B2(n5469), .A(n5468), .ZN(n5467) );
  NAND2_X1 U5344 ( .A1(n5173), .A2(n9028), .ZN(n5172) );
  OAI21_X1 U5345 ( .B1(n7264), .B2(n5174), .A(n8894), .ZN(n5173) );
  NAND2_X1 U5346 ( .A1(n8893), .A2(n7263), .ZN(n5174) );
  NAND2_X1 U5347 ( .A1(n8895), .A2(n9010), .ZN(n5175) );
  NAND2_X1 U5348 ( .A1(n10500), .A2(keyinput_192), .ZN(n5482) );
  INV_X1 U5349 ( .A(n8650), .ZN(n5212) );
  NAND2_X1 U5350 ( .A1(n5285), .A2(n10293), .ZN(n5284) );
  OAI21_X1 U5351 ( .B1(n10289), .B2(n10288), .A(n5286), .ZN(n5285) );
  AOI21_X1 U5352 ( .B1(n5479), .B2(n5476), .A(n5473), .ZN(n10507) );
  AND3_X1 U5353 ( .A1(n8971), .A2(n5149), .A3(n9561), .ZN(n5155) );
  NAND2_X1 U5354 ( .A1(n8967), .A2(n5150), .ZN(n5149) );
  OAI21_X1 U5355 ( .B1(n5071), .B2(n5188), .A(n8764), .ZN(n8669) );
  NAND2_X1 U5356 ( .A1(n8662), .A2(n8735), .ZN(n5188) );
  OR2_X1 U5357 ( .A1(n5275), .A2(n5274), .ZN(n5273) );
  INV_X1 U5358 ( .A(n10312), .ZN(n5274) );
  AOI21_X1 U5359 ( .B1(n10306), .B2(n5277), .A(n5276), .ZN(n5275) );
  NAND2_X1 U5360 ( .A1(n5462), .A2(n5460), .ZN(n5459) );
  NOR2_X1 U5361 ( .A1(n10524), .A2(n5461), .ZN(n5460) );
  OAI21_X1 U5362 ( .B1(n5465), .B2(n5464), .A(n5463), .ZN(n5462) );
  XNOR2_X1 U5363 ( .A(n10525), .B(keyinput_212), .ZN(n5461) );
  NAND2_X1 U5364 ( .A1(n8637), .A2(n8638), .ZN(n8644) );
  AND2_X1 U5365 ( .A1(n5164), .A2(n9453), .ZN(n5163) );
  OR2_X1 U5366 ( .A1(n5167), .A2(n9005), .ZN(n5164) );
  INV_X1 U5367 ( .A(n9001), .ZN(n5167) );
  NAND2_X1 U5368 ( .A1(n5165), .A2(n9503), .ZN(n5162) );
  INV_X1 U5369 ( .A(n8645), .ZN(n8565) );
  INV_X1 U5370 ( .A(SI_25_), .ZN(n10395) );
  NAND2_X1 U5371 ( .A1(n5208), .A2(n8741), .ZN(n5207) );
  AND2_X1 U5372 ( .A1(n8716), .A2(n9892), .ZN(n5198) );
  NAND2_X1 U5373 ( .A1(n8719), .A2(n9868), .ZN(n5202) );
  INV_X1 U5374 ( .A(n5256), .ZN(n5252) );
  INV_X1 U5375 ( .A(n8563), .ZN(n5251) );
  INV_X1 U5376 ( .A(n8583), .ZN(n5395) );
  AND2_X1 U5377 ( .A1(n5514), .A2(n5715), .ZN(n5506) );
  INV_X1 U5378 ( .A(SI_14_), .ZN(n10222) );
  NAND2_X1 U5379 ( .A1(n5681), .A2(n10228), .ZN(n5684) );
  INV_X1 U5380 ( .A(SI_9_), .ZN(n10425) );
  INV_X1 U5381 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5486) );
  INV_X1 U5382 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U5383 ( .A1(n5296), .A2(n5295), .ZN(n10351) );
  OAI21_X1 U5384 ( .B1(n10579), .B2(n10580), .A(n5454), .ZN(n5453) );
  AND2_X1 U5385 ( .A1(n10582), .A2(n5455), .ZN(n5454) );
  AOI21_X1 U5386 ( .B1(n10578), .B2(n10577), .A(n10576), .ZN(n10579) );
  OAI21_X1 U5387 ( .B1(n9021), .B2(n9188), .A(n5170), .ZN(n5169) );
  NOR2_X1 U5388 ( .A1(n9193), .A2(n5171), .ZN(n5170) );
  NAND2_X1 U5389 ( .A1(n9019), .A2(n9020), .ZN(n5171) );
  NOR2_X2 U5390 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5791) );
  OR2_X1 U5391 ( .A1(n9607), .A2(n9250), .ZN(n9011) );
  INV_X1 U5392 ( .A(n8997), .ZN(n5431) );
  OR2_X1 U5393 ( .A1(n9615), .A2(n9261), .ZN(n8997) );
  NOR2_X1 U5394 ( .A1(n9630), .A2(n9635), .ZN(n5330) );
  OR2_X1 U5395 ( .A1(n9510), .A2(n9517), .ZN(n5358) );
  INV_X1 U5396 ( .A(n5418), .ZN(n5417) );
  OAI21_X1 U5397 ( .B1(n9561), .B2(n5419), .A(n9543), .ZN(n5418) );
  INV_X1 U5398 ( .A(n8816), .ZN(n5419) );
  OR2_X1 U5399 ( .A1(n9642), .A2(n9273), .ZN(n8977) );
  NOR2_X1 U5400 ( .A1(n7557), .A2(n5409), .ZN(n5408) );
  INV_X1 U5401 ( .A(n8910), .ZN(n5409) );
  NAND2_X1 U5402 ( .A1(n6320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U5403 ( .A1(n5537), .A2(n5540), .ZN(n7443) );
  AND2_X1 U5404 ( .A1(n5541), .A2(n7437), .ZN(n5540) );
  INV_X1 U5405 ( .A(n9172), .ZN(n6473) );
  NOR2_X1 U5406 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n5023), .ZN(n5632) );
  INV_X1 U5407 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U5408 ( .A1(n8778), .A2(n5241), .ZN(n8497) );
  NAND2_X1 U5409 ( .A1(n9890), .A2(n5055), .ZN(n5241) );
  INV_X1 U5410 ( .A(n8610), .ZN(n9867) );
  NAND2_X1 U5411 ( .A1(n9940), .A2(n9941), .ZN(n9939) );
  INV_X1 U5412 ( .A(n5611), .ZN(n5610) );
  OAI21_X1 U5413 ( .B1(n8346), .B2(n5612), .A(n8358), .ZN(n5611) );
  INV_X1 U5414 ( .A(n8347), .ZN(n5612) );
  OR2_X1 U5415 ( .A1(n10087), .A2(n9711), .ZN(n8620) );
  OR2_X1 U5416 ( .A1(n9998), .A2(n9985), .ZN(n8695) );
  INV_X1 U5417 ( .A(n8680), .ZN(n5249) );
  AND2_X1 U5418 ( .A1(n8679), .A2(n5247), .ZN(n5246) );
  NAND2_X1 U5419 ( .A1(n5248), .A2(n8680), .ZN(n5247) );
  INV_X1 U5420 ( .A(n8681), .ZN(n5248) );
  NOR2_X1 U5421 ( .A1(n10119), .A2(n8191), .ZN(n5235) );
  NOR2_X1 U5422 ( .A1(n10112), .A2(n5234), .ZN(n5233) );
  INV_X1 U5423 ( .A(n5235), .ZN(n5234) );
  OR2_X1 U5424 ( .A1(n10119), .A2(n10029), .ZN(n8681) );
  NOR2_X1 U5425 ( .A1(n7738), .A2(n5226), .ZN(n5225) );
  OR2_X1 U5426 ( .A1(n7614), .A2(n10987), .ZN(n5226) );
  NAND2_X1 U5427 ( .A1(n10987), .A2(n7499), .ZN(n8645) );
  OR2_X1 U5428 ( .A1(n5603), .A2(n7089), .ZN(n5605) );
  NAND2_X1 U5429 ( .A1(n8499), .A2(n8725), .ZN(n8462) );
  INV_X1 U5430 ( .A(n8773), .ZN(n8461) );
  NAND2_X1 U5431 ( .A1(n5030), .A2(n5631), .ZN(n5629) );
  NAND2_X1 U5432 ( .A1(n5074), .A2(n5030), .ZN(n5628) );
  NAND2_X1 U5433 ( .A1(n8531), .A2(n8530), .ZN(n5484) );
  OR2_X1 U5434 ( .A1(n5761), .A2(n5760), .ZN(n8438) );
  AOI21_X1 U5435 ( .B1(n5519), .B2(n5521), .A(n5518), .ZN(n5517) );
  INV_X1 U5436 ( .A(n5735), .ZN(n5518) );
  AND2_X1 U5437 ( .A1(n5742), .A2(n5741), .ZN(n6217) );
  NAND2_X1 U5438 ( .A1(n6153), .A2(n5722), .ZN(n6169) );
  AND2_X1 U5439 ( .A1(n5727), .A2(n5726), .ZN(n6168) );
  INV_X1 U5440 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10571) );
  OR2_X1 U5441 ( .A1(n6151), .A2(n6150), .ZN(n6153) );
  NOR2_X1 U5442 ( .A1(n5714), .A2(n5515), .ZN(n5514) );
  INV_X1 U5443 ( .A(n5710), .ZN(n5515) );
  INV_X1 U5444 ( .A(n5511), .ZN(n5510) );
  OAI21_X1 U5445 ( .B1(n5714), .B2(n5512), .A(n5713), .ZN(n5511) );
  NAND2_X1 U5446 ( .A1(n6096), .A2(n5710), .ZN(n5512) );
  INV_X1 U5447 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6374) );
  XNOR2_X1 U5448 ( .A(n5700), .B(n10222), .ZN(n6057) );
  NAND2_X1 U5449 ( .A1(n5699), .A2(n5698), .ZN(n6058) );
  OR3_X1 U5450 ( .A1(n6677), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_11__SCAN_IN), .ZN(n6873) );
  OAI21_X1 U5451 ( .B1(n5933), .B2(n5260), .A(n5258), .ZN(n5967) );
  INV_X1 U5452 ( .A(n5261), .ZN(n5260) );
  AOI21_X1 U5453 ( .B1(n5261), .B2(n5259), .A(n5494), .ZN(n5258) );
  INV_X1 U5454 ( .A(n5932), .ZN(n5259) );
  NOR2_X1 U5455 ( .A1(n6499), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6571) );
  AOI21_X1 U5456 ( .B1(n5183), .B2(n5186), .A(n5048), .ZN(n5263) );
  NOR2_X1 U5457 ( .A1(n5185), .A2(n5184), .ZN(n5183) );
  INV_X1 U5458 ( .A(n5668), .ZN(n5182) );
  INV_X1 U5459 ( .A(n5049), .ZN(n5185) );
  NAND2_X1 U5460 ( .A1(n6422), .A2(n5065), .ZN(n5649) );
  OR2_X1 U5461 ( .A1(n6268), .A2(n10284), .ZN(n6302) );
  XNOR2_X1 U5462 ( .A(n6243), .B(n6221), .ZN(n9221) );
  INV_X1 U5463 ( .A(n6232), .ZN(n6227) );
  AOI21_X1 U5464 ( .B1(n6036), .B2(n5578), .A(n5036), .ZN(n5577) );
  NOR2_X1 U5465 ( .A1(n5594), .A2(n5590), .ZN(n5589) );
  INV_X1 U5466 ( .A(n6247), .ZN(n5590) );
  INV_X1 U5467 ( .A(n6265), .ZN(n5594) );
  NAND2_X1 U5468 ( .A1(n5593), .A2(n6265), .ZN(n5592) );
  INV_X1 U5469 ( .A(n9249), .ZN(n5593) );
  AND2_X1 U5470 ( .A1(n6280), .A2(n6279), .ZN(n9305) );
  AND4_X1 U5471 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n8511)
         );
  AND4_X1 U5472 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n7788)
         );
  NAND2_X1 U5473 ( .A1(n5921), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5821) );
  NOR2_X1 U5474 ( .A1(n10773), .A2(n6715), .ZN(n10791) );
  AOI21_X1 U5475 ( .B1(n7402), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7401), .ZN(
        n9335) );
  AOI21_X1 U5476 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7423), .A(n7422), .ZN(
        n7425) );
  NOR2_X1 U5477 ( .A1(n5968), .A2(n5031), .ZN(n6041) );
  INV_X1 U5478 ( .A(n5636), .ZN(n5132) );
  NOR2_X1 U5479 ( .A1(n9611), .A2(n9477), .ZN(n9186) );
  NAND2_X1 U5480 ( .A1(n9438), .A2(n9437), .ZN(n9436) );
  NOR2_X1 U5481 ( .A1(n9485), .A2(n9615), .ZN(n9455) );
  NAND2_X1 U5482 ( .A1(n8821), .A2(n5043), .ZN(n9489) );
  INV_X1 U5483 ( .A(n9490), .ZN(n5362) );
  NAND2_X1 U5484 ( .A1(n9509), .A2(n9503), .ZN(n5363) );
  AND2_X1 U5485 ( .A1(n8996), .A2(n9474), .ZN(n9490) );
  INV_X1 U5486 ( .A(n5358), .ZN(n9509) );
  NOR2_X1 U5487 ( .A1(n9551), .A2(n9635), .ZN(n9527) );
  AOI21_X1 U5488 ( .B1(n9560), .B2(n9571), .A(n9176), .ZN(n9540) );
  NOR2_X1 U5489 ( .A1(n9645), .A2(n9175), .ZN(n9176) );
  AND2_X1 U5490 ( .A1(n9173), .A2(n8274), .ZN(n8870) );
  NOR2_X1 U5491 ( .A1(n8203), .A2(n11101), .ZN(n8204) );
  OR2_X1 U5492 ( .A1(n5642), .A2(n9067), .ZN(n8203) );
  NOR2_X1 U5493 ( .A1(n7769), .A2(n5333), .ZN(n7816) );
  INV_X1 U5494 ( .A(n5335), .ZN(n5333) );
  NOR2_X1 U5495 ( .A1(n7746), .A2(n8864), .ZN(n7747) );
  AND2_X1 U5496 ( .A1(n5052), .A2(n8924), .ZN(n5426) );
  NOR2_X1 U5497 ( .A1(n7467), .A2(n5412), .ZN(n5411) );
  INV_X1 U5498 ( .A(n7465), .ZN(n5412) );
  OAI211_X1 U5499 ( .C1(n7229), .C2(n10831), .A(n10832), .B(n5337), .ZN(n7354)
         );
  OAI21_X1 U5500 ( .B1(n7265), .B2(n10836), .A(n7254), .ZN(n5337) );
  INV_X1 U5501 ( .A(n7229), .ZN(n7265) );
  NAND2_X1 U5502 ( .A1(n5522), .A2(n8849), .ZN(n8851) );
  NAND2_X1 U5503 ( .A1(n9678), .A2(n8848), .ZN(n5522) );
  INV_X1 U5504 ( .A(n9191), .ZN(n9589) );
  OAI21_X1 U5505 ( .B1(n9426), .B2(n9188), .A(n5401), .ZN(n9194) );
  NAND2_X1 U5506 ( .A1(n6205), .A2(n6204), .ZN(n9625) );
  OAI211_X1 U5507 ( .C1(n7200), .C2(n8826), .A(n5939), .B(n5938), .ZN(n10959)
         );
  INV_X1 U5508 ( .A(n7473), .ZN(n10925) );
  AND2_X1 U5509 ( .A1(n6332), .A2(n6331), .ZN(n10183) );
  AND2_X1 U5510 ( .A1(n6721), .A2(n10760), .ZN(n10185) );
  NOR2_X1 U5511 ( .A1(n5373), .A2(n5436), .ZN(n5372) );
  NAND4_X1 U5512 ( .A1(n5317), .A2(n5768), .A3(n5158), .A4(n5776), .ZN(n5784)
         );
  INV_X1 U5513 ( .A(n5373), .ZN(n5159) );
  XNOR2_X1 U5514 ( .A(n6319), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9045) );
  INV_X1 U5515 ( .A(n5565), .ZN(n5564) );
  OAI21_X1 U5516 ( .B1(n9789), .B2(n5566), .A(n9693), .ZN(n5565) );
  INV_X1 U5517 ( .A(n9163), .ZN(n5563) );
  XNOR2_X1 U5518 ( .A(n6696), .B(n6695), .ZN(n5524) );
  OR2_X1 U5519 ( .A1(n9776), .A2(n9779), .ZN(n5553) );
  AND2_X1 U5520 ( .A1(n9777), .A2(n5079), .ZN(n5547) );
  NAND2_X1 U5521 ( .A1(n9746), .A2(n5535), .ZN(n5534) );
  INV_X1 U5522 ( .A(n9707), .ZN(n5535) );
  OAI21_X1 U5523 ( .B1(n9768), .B2(n9766), .A(n9764), .ZN(n9124) );
  OR2_X1 U5524 ( .A1(n5531), .A2(n5528), .ZN(n5527) );
  INV_X1 U5525 ( .A(n5534), .ZN(n5531) );
  NOR2_X1 U5526 ( .A1(n5536), .A2(n5529), .ZN(n5528) );
  INV_X1 U5527 ( .A(n8229), .ZN(n5545) );
  NOR2_X1 U5528 ( .A1(n9124), .A2(n9123), .ZN(n9706) );
  NAND2_X1 U5529 ( .A1(n9124), .A2(n9123), .ZN(n9704) );
  NAND2_X1 U5530 ( .A1(n9706), .A2(n9704), .ZN(n5533) );
  NAND2_X1 U5531 ( .A1(n9102), .A2(n9103), .ZN(n5555) );
  NOR2_X1 U5532 ( .A1(n9099), .A2(n9098), .ZN(n9776) );
  NAND2_X1 U5533 ( .A1(n9099), .A2(n9098), .ZN(n9777) );
  AND2_X1 U5534 ( .A1(n8168), .A2(n8167), .ZN(n8174) );
  OR2_X1 U5535 ( .A1(n10734), .A2(n10733), .ZN(n5120) );
  NAND2_X1 U5536 ( .A1(n10683), .A2(n6542), .ZN(n6586) );
  NAND2_X1 U5537 ( .A1(n6848), .A2(n5087), .ZN(n6853) );
  NAND2_X1 U5538 ( .A1(n6853), .A2(n6852), .ZN(n7003) );
  NOR2_X1 U5539 ( .A1(n10722), .A2(n10723), .ZN(n10721) );
  NAND2_X1 U5540 ( .A1(n8540), .A2(n8539), .ZN(n9852) );
  NAND2_X1 U5541 ( .A1(n9875), .A2(n5218), .ZN(n9859) );
  NOR2_X1 U5542 ( .A1(n10053), .A2(n5219), .ZN(n5218) );
  NAND2_X1 U5543 ( .A1(n8727), .A2(n8726), .ZN(n8773) );
  AND2_X1 U5544 ( .A1(n8469), .A2(n8429), .ZN(n9164) );
  NAND2_X1 U5545 ( .A1(n5240), .A2(n8771), .ZN(n8499) );
  INV_X1 U5546 ( .A(n8497), .ZN(n5240) );
  AND2_X1 U5547 ( .A1(n8778), .A2(n8720), .ZN(n9868) );
  CLKBUF_X1 U5548 ( .A(n9913), .Z(n9914) );
  AND2_X1 U5550 ( .A1(n8620), .A2(n8619), .ZN(n9953) );
  NAND2_X1 U5551 ( .A1(n9960), .A2(n8346), .ZN(n9959) );
  NOR2_X1 U5552 ( .A1(n9993), .A2(n10097), .ZN(n9977) );
  INV_X1 U5553 ( .A(n5625), .ZN(n5624) );
  OAI21_X1 U5554 ( .B1(n5029), .B2(n5032), .A(n5063), .ZN(n5625) );
  AND2_X1 U5555 ( .A1(n8661), .A2(n8670), .ZN(n8764) );
  NAND2_X1 U5556 ( .A1(n7880), .A2(n7879), .ZN(n7995) );
  NAND2_X1 U5557 ( .A1(n7956), .A2(n5029), .ZN(n7983) );
  AOI21_X1 U5558 ( .B1(n5615), .B2(n5617), .A(n5056), .ZN(n5614) );
  NAND2_X1 U5559 ( .A1(n7097), .A2(n7096), .ZN(n7287) );
  NAND2_X1 U5560 ( .A1(n7271), .A2(n7277), .ZN(n5618) );
  AND2_X1 U5561 ( .A1(n8589), .A2(n7110), .ZN(n8750) );
  INV_X1 U5562 ( .A(n11111), .ZN(n10968) );
  INV_X1 U5563 ( .A(n11109), .ZN(n11053) );
  AND2_X1 U5564 ( .A1(n6429), .A2(n6431), .ZN(n10150) );
  MUX2_X1 U5565 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6413), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n6414) );
  XNOR2_X1 U5566 ( .A(n6040), .B(n6039), .ZN(n7877) );
  XNOR2_X1 U5567 ( .A(n5967), .B(n5640), .ZN(n7495) );
  NAND2_X1 U5568 ( .A1(n8491), .A2(n5920), .ZN(n7366) );
  AND2_X1 U5569 ( .A1(n5944), .A2(n5920), .ZN(n5595) );
  AND4_X1 U5570 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(n7749)
         );
  OR2_X1 U5571 ( .A1(n5947), .A2(n5971), .ZN(n5974) );
  AND2_X1 U5572 ( .A1(n6004), .A2(n5981), .ZN(n5596) );
  AND2_X1 U5573 ( .A1(n9595), .A2(n5574), .ZN(n5573) );
  NAND2_X1 U5574 ( .A1(n9319), .A2(n9306), .ZN(n5574) );
  NAND2_X1 U5575 ( .A1(n5934), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5811) );
  AND4_X1 U5576 ( .A1(n6179), .A2(n6178), .A3(n6177), .A4(n6176), .ZN(n9549)
         );
  AND4_X1 U5577 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n8073)
         );
  NAND2_X1 U5578 ( .A1(n6029), .A2(n6028), .ZN(n11065) );
  NAND2_X1 U5579 ( .A1(n6100), .A2(n6099), .ZN(n9658) );
  INV_X1 U5580 ( .A(n7011), .ZN(n5832) );
  OR2_X1 U5581 ( .A1(n6359), .A2(n6358), .ZN(n7014) );
  AOI22_X1 U5582 ( .A1(n9037), .A2(n9038), .B1(n9040), .B2(n9039), .ZN(n5491)
         );
  NAND2_X1 U5583 ( .A1(n5047), .A2(n8879), .ZN(n5177) );
  NAND2_X1 U5584 ( .A1(n8879), .A2(n8843), .ZN(n5421) );
  INV_X1 U5585 ( .A(n9213), .ZN(n9430) );
  INV_X1 U5586 ( .A(n7749), .ZN(n9328) );
  AND2_X1 U5587 ( .A1(n9415), .A2(n9414), .ZN(n9598) );
  NAND2_X1 U5588 ( .A1(n9411), .A2(n5345), .ZN(n9410) );
  NAND2_X1 U5589 ( .A1(n7469), .A2(n8903), .ZN(n7480) );
  NAND2_X1 U5590 ( .A1(n9193), .A2(n5343), .ZN(n5342) );
  OR2_X1 U5591 ( .A1(n9193), .A2(n5638), .ZN(n5341) );
  NAND2_X1 U5592 ( .A1(n5347), .A2(n5345), .ZN(n5343) );
  OR2_X1 U5593 ( .A1(n9405), .A2(n5346), .ZN(n5135) );
  NAND2_X1 U5594 ( .A1(n9193), .A2(n5347), .ZN(n5346) );
  NAND2_X1 U5595 ( .A1(n9405), .A2(n5344), .ZN(n5134) );
  NOR2_X1 U5596 ( .A1(n9193), .A2(n5345), .ZN(n5344) );
  NAND2_X1 U5597 ( .A1(n6651), .A2(n6648), .ZN(n9785) );
  NAND2_X1 U5598 ( .A1(n5194), .A2(n8743), .ZN(n8807) );
  MUX2_X1 U5599 ( .A(n8803), .B(n8802), .S(n8801), .Z(n8810) );
  AND2_X1 U5600 ( .A1(n5193), .A2(n5192), .ZN(n8802) );
  CLKBUF_X1 U5601 ( .A(n6415), .Z(n6419) );
  XNOR2_X1 U5602 ( .A(n6441), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6682) );
  OR2_X1 U5603 ( .A1(n9851), .A2(n10702), .ZN(n5112) );
  AOI21_X1 U5604 ( .B1(n10744), .B2(n9850), .A(n5111), .ZN(n5110) );
  OR2_X1 U5605 ( .A1(n10146), .A2(n8447), .ZN(n8449) );
  INV_X1 U5606 ( .A(n5222), .ZN(n8503) );
  INV_X1 U5607 ( .A(n9926), .ZN(n9850) );
  OR2_X1 U5608 ( .A1(n11057), .A2(n6652), .ZN(n10879) );
  AND2_X1 U5609 ( .A1(n11019), .A2(n7119), .ZN(n11009) );
  NAND2_X1 U5610 ( .A1(n6412), .A2(n5627), .ZN(n6470) );
  NOR2_X1 U5611 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5627) );
  BUF_X1 U5612 ( .A(n6595), .Z(n8805) );
  INV_X1 U5613 ( .A(SI_31_), .ZN(n5279) );
  AOI221_X1 U5614 ( .B1(SI_27_), .B2(keyinput_133), .C1(keyinput_131), .C2(
        SI_29_), .A(n10397), .ZN(n10404) );
  AND2_X1 U5615 ( .A1(n5280), .A2(n5278), .ZN(n10205) );
  XNOR2_X1 U5616 ( .A(n5281), .B(keyinput_0), .ZN(n5280) );
  XNOR2_X1 U5617 ( .A(n5279), .B(keyinput_1), .ZN(n5278) );
  INV_X1 U5618 ( .A(P2_WR_REG_SCAN_IN), .ZN(n5281) );
  AOI21_X1 U5619 ( .B1(n5449), .B2(n5447), .A(n10424), .ZN(n10433) );
  XNOR2_X1 U5620 ( .A(n10425), .B(n5448), .ZN(n5447) );
  NAND2_X1 U5621 ( .A1(n5450), .A2(n10422), .ZN(n5449) );
  NAND2_X1 U5622 ( .A1(n10240), .A2(n10241), .ZN(n5294) );
  NOR2_X1 U5623 ( .A1(n10238), .A2(n10239), .ZN(n5293) );
  NAND2_X1 U5624 ( .A1(n10443), .A2(n10442), .ZN(n10447) );
  OAI22_X1 U5625 ( .A1(n10452), .A2(keyinput_166), .B1(n10453), .B2(
        P2_REG3_REG_23__SCAN_IN), .ZN(n5446) );
  OAI22_X1 U5626 ( .A1(n10458), .A2(n10457), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        keyinput_168), .ZN(n5444) );
  AOI21_X1 U5627 ( .B1(n5290), .B2(n5289), .A(n5288), .ZN(n10245) );
  NAND2_X1 U5628 ( .A1(n10465), .A2(n10464), .ZN(n10468) );
  AOI211_X1 U5629 ( .C1(n10478), .C2(n10479), .A(n10477), .B(n10476), .ZN(
        n5472) );
  NAND2_X1 U5630 ( .A1(n5471), .A2(n5470), .ZN(n5469) );
  NAND2_X1 U5631 ( .A1(n10481), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U5632 ( .A1(n10480), .A2(keyinput_179), .ZN(n5471) );
  AOI22_X1 U5633 ( .A1(n10483), .A2(n10482), .B1(keyinput_180), .B2(
        P2_REG3_REG_4__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U5634 ( .A1(n5300), .A2(n10277), .ZN(n10281) );
  OAI21_X1 U5635 ( .B1(n10271), .B2(n5304), .A(n5301), .ZN(n5300) );
  NAND2_X1 U5636 ( .A1(n5175), .A2(n5172), .ZN(n8902) );
  INV_X1 U5637 ( .A(n5287), .ZN(n5286) );
  OAI22_X1 U5638 ( .A1(n10500), .A2(keyinput_64), .B1(n10290), .B2(
        P2_B_REG_SCAN_IN), .ZN(n5287) );
  NAND2_X1 U5639 ( .A1(n5483), .A2(n5480), .ZN(n5479) );
  AND2_X1 U5640 ( .A1(n5482), .A2(n5481), .ZN(n5480) );
  NAND2_X1 U5641 ( .A1(n10501), .A2(P2_B_REG_SCAN_IN), .ZN(n5481) );
  AND2_X1 U5642 ( .A1(n5478), .A2(n5477), .ZN(n5476) );
  NAND2_X1 U5643 ( .A1(n10503), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U5644 ( .A1(n10502), .A2(keyinput_193), .ZN(n5478) );
  NAND2_X1 U5645 ( .A1(n5475), .A2(n5474), .ZN(n5473) );
  NAND2_X1 U5646 ( .A1(keyinput_194), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U5647 ( .A1(n10505), .A2(n10504), .ZN(n5475) );
  NAND2_X1 U5648 ( .A1(n5145), .A2(n5058), .ZN(n5144) );
  INV_X1 U5649 ( .A(n8928), .ZN(n5147) );
  INV_X1 U5650 ( .A(n8926), .ZN(n5148) );
  INV_X1 U5651 ( .A(n5283), .ZN(n5282) );
  OAI22_X1 U5652 ( .A1(n10505), .A2(n10294), .B1(P2_DATAO_REG_30__SCAN_IN), 
        .B2(keyinput_66), .ZN(n5283) );
  NAND2_X1 U5653 ( .A1(n5140), .A2(n5139), .ZN(n8940) );
  AOI21_X1 U5654 ( .B1(n5141), .B2(n5143), .A(n5090), .ZN(n5139) );
  NAND2_X1 U5655 ( .A1(n8919), .A2(n5141), .ZN(n5140) );
  AOI21_X1 U5656 ( .B1(n5142), .B2(n5146), .A(n5075), .ZN(n5141) );
  NOR2_X1 U5657 ( .A1(n5157), .A2(n5151), .ZN(n5150) );
  AND2_X1 U5658 ( .A1(n8963), .A2(n8962), .ZN(n5157) );
  INV_X1 U5659 ( .A(n8968), .ZN(n5151) );
  AND2_X1 U5660 ( .A1(n5212), .A2(n5211), .ZN(n5210) );
  NAND2_X1 U5661 ( .A1(n8653), .A2(n8652), .ZN(n5213) );
  NOR2_X1 U5662 ( .A1(n8651), .A2(n8758), .ZN(n5211) );
  NAND2_X1 U5663 ( .A1(n5284), .A2(n5282), .ZN(n10305) );
  INV_X1 U5664 ( .A(n10309), .ZN(n5277) );
  OAI21_X1 U5665 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_78), .A(n10308), 
        .ZN(n5276) );
  INV_X1 U5666 ( .A(n10520), .ZN(n5465) );
  INV_X1 U5667 ( .A(n10519), .ZN(n5464) );
  NOR2_X1 U5668 ( .A1(n10518), .A2(n5101), .ZN(n5463) );
  NOR2_X1 U5669 ( .A1(n10311), .A2(n5272), .ZN(n5271) );
  NOR2_X1 U5670 ( .A1(n10313), .A2(keyinput_81), .ZN(n5272) );
  INV_X1 U5671 ( .A(n5458), .ZN(n5457) );
  OAI22_X1 U5672 ( .A1(n10527), .A2(n10526), .B1(P2_DATAO_REG_11__SCAN_IN), 
        .B2(keyinput_213), .ZN(n5458) );
  AOI21_X1 U5673 ( .B1(n5155), .B2(n5156), .A(n5153), .ZN(n5152) );
  INV_X1 U5674 ( .A(n8974), .ZN(n5153) );
  NAND2_X1 U5675 ( .A1(n8967), .A2(n8968), .ZN(n5156) );
  OAI21_X1 U5676 ( .B1(n5068), .B2(n8669), .A(n8670), .ZN(n8671) );
  NAND2_X1 U5677 ( .A1(n5273), .A2(n5271), .ZN(n10314) );
  AND2_X1 U5678 ( .A1(n5314), .A2(n5313), .ZN(n5312) );
  NAND2_X1 U5679 ( .A1(n10317), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U5680 ( .A1(n10527), .A2(keyinput_85), .ZN(n5314) );
  AND2_X1 U5681 ( .A1(n10522), .A2(keyinput_82), .ZN(n5315) );
  NAND2_X1 U5682 ( .A1(n10535), .A2(n10319), .ZN(n5309) );
  NAND2_X1 U5683 ( .A1(keyinput_87), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n5308)
         );
  NAND2_X1 U5684 ( .A1(n5459), .A2(n5457), .ZN(n10532) );
  AOI21_X1 U5685 ( .B1(n5311), .B2(n5310), .A(n5307), .ZN(n10330) );
  AOI22_X1 U5686 ( .A1(n10318), .A2(n10528), .B1(keyinput_86), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U5687 ( .A1(n5309), .A2(n5308), .ZN(n5307) );
  OAI21_X1 U5688 ( .B1(n10316), .B2(n5315), .A(n5312), .ZN(n5311) );
  INV_X1 U5689 ( .A(n8644), .ZN(n8643) );
  INV_X1 U5690 ( .A(keyinput_104), .ZN(n5299) );
  NAND2_X1 U5691 ( .A1(n5442), .A2(n10562), .ZN(n5441) );
  NAND2_X1 U5692 ( .A1(n10550), .A2(n10549), .ZN(n5442) );
  AND2_X1 U5693 ( .A1(n5163), .A2(n5162), .ZN(n5161) );
  NAND2_X1 U5694 ( .A1(n5603), .A2(n10880), .ZN(n8579) );
  INV_X1 U5695 ( .A(SI_12_), .ZN(n10391) );
  INV_X1 U5696 ( .A(SI_10_), .ZN(n10228) );
  INV_X1 U5697 ( .A(SI_8_), .ZN(n10234) );
  NAND2_X1 U5698 ( .A1(n10344), .A2(n5297), .ZN(n5296) );
  AND2_X1 U5699 ( .A1(n10345), .A2(n5298), .ZN(n5297) );
  XNOR2_X1 U5700 ( .A(n5299), .B(P1_IR_REG_13__SCAN_IN), .ZN(n5298) );
  AOI22_X1 U5701 ( .A1(n10346), .A2(n10565), .B1(keyinput_107), .B2(
        P1_IR_REG_16__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U5702 ( .A1(n5440), .A2(n5438), .ZN(n10578) );
  NOR2_X1 U5703 ( .A1(n10564), .A2(n5439), .ZN(n5438) );
  NAND2_X1 U5704 ( .A1(n5441), .A2(n5102), .ZN(n5440) );
  XNOR2_X1 U5705 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_234), .ZN(n5439) );
  OAI22_X1 U5706 ( .A1(n10566), .A2(n10565), .B1(P1_IR_REG_16__SCAN_IN), .B2(
        keyinput_235), .ZN(n10567) );
  XNOR2_X1 U5707 ( .A(n5456), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5455) );
  INV_X1 U5708 ( .A(keyinput_243), .ZN(n5456) );
  INV_X1 U5709 ( .A(n9023), .ZN(n5399) );
  NOR2_X1 U5710 ( .A1(n5543), .A2(n5539), .ZN(n5538) );
  INV_X1 U5711 ( .A(n7214), .ZN(n5543) );
  INV_X1 U5712 ( .A(n7207), .ZN(n5539) );
  NAND2_X1 U5713 ( .A1(n7214), .A2(n5542), .ZN(n5541) );
  INV_X1 U5714 ( .A(n7212), .ZN(n5542) );
  INV_X1 U5715 ( .A(n5202), .ZN(n5204) );
  AND2_X1 U5716 ( .A1(n10053), .A2(n8455), .ZN(n8789) );
  INV_X1 U5717 ( .A(n8411), .ZN(n5630) );
  AND2_X1 U5718 ( .A1(n8436), .A2(n5504), .ZN(n5503) );
  NAND2_X1 U5719 ( .A1(n6249), .A2(n5751), .ZN(n5504) );
  INV_X1 U5720 ( .A(n5751), .ZN(n5501) );
  NOR2_X1 U5721 ( .A1(n6202), .A2(n5520), .ZN(n5519) );
  INV_X1 U5722 ( .A(n5730), .ZN(n5520) );
  INV_X1 U5723 ( .A(SI_21_), .ZN(n10407) );
  NAND2_X1 U5724 ( .A1(n5690), .A2(n10391), .ZN(n5693) );
  NOR2_X1 U5725 ( .A1(n5498), .A2(n5494), .ZN(n5493) );
  INV_X1 U5726 ( .A(n5680), .ZN(n5498) );
  NAND2_X1 U5727 ( .A1(n5497), .A2(n5680), .ZN(n5496) );
  INV_X1 U5728 ( .A(n5640), .ZN(n5497) );
  NOR2_X1 U5729 ( .A1(n5958), .A2(n5262), .ZN(n5261) );
  INV_X1 U5730 ( .A(n5671), .ZN(n5262) );
  NAND2_X1 U5731 ( .A1(n5932), .A2(n5881), .ZN(n5184) );
  INV_X1 U5732 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6059) );
  OR2_X1 U5733 ( .A1(n9611), .A2(n9442), .ZN(n9006) );
  NAND2_X1 U5734 ( .A1(n5330), .A2(n9501), .ZN(n5329) );
  INV_X1 U5735 ( .A(n6191), .ZN(n6190) );
  NOR2_X1 U5736 ( .A1(n9658), .A2(n9079), .ZN(n5320) );
  NOR2_X1 U5737 ( .A1(n5368), .A2(n5131), .ZN(n5130) );
  INV_X1 U5738 ( .A(n7868), .ZN(n5131) );
  NAND2_X1 U5739 ( .A1(n5370), .A2(n8027), .ZN(n5368) );
  INV_X1 U5740 ( .A(n8027), .ZN(n5367) );
  NAND2_X1 U5741 ( .A1(n5130), .A2(n5128), .ZN(n5127) );
  INV_X1 U5742 ( .A(n8866), .ZN(n5128) );
  NOR2_X1 U5743 ( .A1(n5334), .A2(n11065), .ZN(n5332) );
  NAND2_X1 U5744 ( .A1(n5335), .A2(n7819), .ZN(n5334) );
  NOR2_X1 U5745 ( .A1(n7820), .A2(n7768), .ZN(n5335) );
  OR2_X1 U5746 ( .A1(n8914), .A2(n7671), .ZN(n7714) );
  NAND2_X1 U5747 ( .A1(n5321), .A2(n10886), .ZN(n5323) );
  AND3_X1 U5748 ( .A1(n5077), .A2(n7258), .A3(n10852), .ZN(n5321) );
  NOR2_X1 U5749 ( .A1(n5323), .A2(n8916), .ZN(n7564) );
  NAND2_X1 U5750 ( .A1(n5779), .A2(n5437), .ZN(n5436) );
  INV_X1 U5751 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U5752 ( .A1(n5778), .A2(n5374), .ZN(n5373) );
  INV_X1 U5753 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5778) );
  INV_X1 U5754 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5374) );
  INV_X1 U5755 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6325) );
  NOR2_X1 U5756 ( .A1(n5777), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5428) );
  INV_X1 U5757 ( .A(n5776), .ZN(n5777) );
  INV_X1 U5758 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5766) );
  INV_X1 U5759 ( .A(n9717), .ZN(n5552) );
  AOI21_X1 U5760 ( .B1(n5202), .B2(n5203), .A(n8721), .ZN(n5201) );
  NOR2_X1 U5761 ( .A1(n5206), .A2(n8722), .ZN(n5203) );
  INV_X1 U5762 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U5763 ( .A1(n8473), .A2(n9801), .ZN(n8727) );
  NAND2_X1 U5764 ( .A1(n8471), .A2(n5220), .ZN(n5219) );
  NAND2_X1 U5765 ( .A1(n5044), .A2(n8384), .ZN(n5602) );
  NOR2_X1 U5766 ( .A1(n10082), .A2(n5230), .ZN(n5229) );
  INV_X1 U5767 ( .A(n5231), .ZN(n5230) );
  NOR2_X1 U5768 ( .A1(n10087), .A2(n10093), .ZN(n5231) );
  AND2_X1 U5769 ( .A1(n8681), .A2(n8680), .ZN(n8765) );
  INV_X1 U5770 ( .A(n5254), .ZN(n5253) );
  AOI21_X1 U5771 ( .B1(n5254), .B2(n5252), .A(n5251), .ZN(n5250) );
  NOR2_X1 U5772 ( .A1(n8656), .A2(n8561), .ZN(n5254) );
  NOR2_X1 U5773 ( .A1(n8657), .A2(n5257), .ZN(n5256) );
  INV_X1 U5774 ( .A(n8646), .ZN(n5257) );
  INV_X1 U5775 ( .A(n7531), .ZN(n5617) );
  INV_X1 U5776 ( .A(n5388), .ZN(n5387) );
  AOI21_X1 U5777 ( .B1(n5388), .B2(n5386), .A(n5385), .ZN(n5384) );
  INV_X1 U5778 ( .A(n10996), .ZN(n5385) );
  OAI21_X1 U5779 ( .B1(n7096), .B2(n5623), .A(n8754), .ZN(n5622) );
  INV_X1 U5780 ( .A(n8634), .ZN(n5623) );
  NOR2_X1 U5781 ( .A1(n7074), .A2(n7073), .ZN(n7217) );
  INV_X1 U5782 ( .A(n8586), .ZN(n5393) );
  INV_X1 U5783 ( .A(n8589), .ZN(n5391) );
  NAND2_X1 U5784 ( .A1(n7109), .A2(n5394), .ZN(n7160) );
  INV_X1 U5785 ( .A(n5392), .ZN(n5394) );
  INV_X1 U5786 ( .A(n5225), .ZN(n5223) );
  INV_X1 U5787 ( .A(n5607), .ZN(n5606) );
  OAI21_X1 U5788 ( .B1(n8447), .B2(n6886), .A(n6884), .ZN(n5607) );
  NOR2_X1 U5789 ( .A1(n6640), .A2(n7118), .ZN(n7189) );
  OAI21_X1 U5790 ( .B1(n6250), .B2(n5502), .A(n5499), .ZN(n8527) );
  INV_X1 U5791 ( .A(n5503), .ZN(n5502) );
  NOR2_X1 U5792 ( .A1(n5500), .A2(n5089), .ZN(n5499) );
  AND2_X1 U5793 ( .A1(n5503), .A2(n5501), .ZN(n5500) );
  AOI21_X1 U5794 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_21__SCAN_IN), .ZN(n5570) );
  INV_X1 U5795 ( .A(n6185), .ZN(n5521) );
  NAND2_X1 U5796 ( .A1(n5728), .A2(n5727), .ZN(n6186) );
  INV_X1 U5797 ( .A(n5508), .ZN(n5507) );
  OAI21_X1 U5798 ( .B1(n5510), .B2(n6132), .A(n5717), .ZN(n5508) );
  INV_X1 U5799 ( .A(n6057), .ZN(n5702) );
  INV_X1 U5800 ( .A(n6006), .ZN(n5687) );
  XNOR2_X1 U5801 ( .A(n5688), .B(n5686), .ZN(n6006) );
  INV_X1 U5802 ( .A(SI_11_), .ZN(n5686) );
  INV_X1 U5803 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5485) );
  AND2_X1 U5804 ( .A1(n6300), .A2(n6298), .ZN(n9206) );
  AND2_X1 U5805 ( .A1(n6265), .A2(n6264), .ZN(n9249) );
  NAND2_X1 U5806 ( .A1(n6246), .A2(n5060), .ZN(n9248) );
  NAND2_X1 U5807 ( .A1(n6102), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6122) );
  OR2_X1 U5808 ( .A1(n6234), .A2(n10480), .ZN(n6255) );
  AOI21_X1 U5809 ( .B1(n5453), .B2(n10592), .A(n5103), .ZN(n10594) );
  AND2_X1 U5810 ( .A1(n6213), .A2(n5584), .ZN(n5583) );
  NAND2_X1 U5811 ( .A1(n9239), .A2(n5585), .ZN(n5584) );
  INV_X1 U5812 ( .A(n6184), .ZN(n5585) );
  NAND2_X1 U5813 ( .A1(n9248), .A2(n9249), .ZN(n9308) );
  OR2_X1 U5814 ( .A1(n6085), .A2(n6084), .ZN(n6103) );
  OAI21_X1 U5815 ( .B1(n5168), .B2(n9032), .A(n9031), .ZN(n9036) );
  AOI21_X1 U5816 ( .B1(n5169), .B2(n9027), .A(n9026), .ZN(n5168) );
  AOI21_X1 U5817 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9368), .A(n9367), .ZN(
        n9371) );
  NAND2_X1 U5818 ( .A1(n8833), .A2(n8832), .ZN(n9400) );
  OR2_X1 U5819 ( .A1(n6302), .A2(n6301), .ZN(n9197) );
  NOR2_X1 U5820 ( .A1(n9406), .A2(n9589), .ZN(n9399) );
  NAND2_X1 U5821 ( .A1(n5325), .A2(n5324), .ZN(n9406) );
  OAI21_X1 U5822 ( .B1(n8821), .B2(n5432), .A(n5430), .ZN(n9462) );
  INV_X1 U5823 ( .A(n8823), .ZN(n5432) );
  AOI21_X1 U5824 ( .B1(n8823), .B2(n8995), .A(n5431), .ZN(n5430) );
  AND2_X1 U5825 ( .A1(n9455), .A2(n9460), .ZN(n9456) );
  NOR2_X1 U5826 ( .A1(n9551), .A2(n5328), .ZN(n9511) );
  INV_X1 U5827 ( .A(n5330), .ZN(n5328) );
  NAND2_X1 U5828 ( .A1(n9525), .A2(n9179), .ZN(n9510) );
  AOI21_X1 U5829 ( .B1(n5417), .B2(n5419), .A(n5415), .ZN(n5414) );
  INV_X1 U5830 ( .A(n8977), .ZN(n5415) );
  OR2_X1 U5831 ( .A1(n9562), .A2(n9642), .ZN(n9551) );
  NAND2_X1 U5832 ( .A1(n9526), .A2(n9531), .ZN(n9525) );
  NAND2_X1 U5833 ( .A1(n6157), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6173) );
  INV_X1 U5834 ( .A(n6159), .ZN(n6157) );
  OR2_X1 U5835 ( .A1(n6139), .A2(n6138), .ZN(n6159) );
  NOR2_X1 U5836 ( .A1(n9653), .A2(n5319), .ZN(n5318) );
  INV_X1 U5837 ( .A(n5320), .ZN(n5319) );
  AOI21_X1 U5838 ( .B1(n5352), .B2(n8963), .A(n5350), .ZN(n5349) );
  INV_X1 U5839 ( .A(n5352), .ZN(n5351) );
  INV_X1 U5840 ( .A(n9173), .ZN(n5350) );
  NAND2_X1 U5841 ( .A1(n8204), .A2(n5320), .ZN(n9189) );
  NAND2_X1 U5842 ( .A1(n8204), .A2(n11124), .ZN(n8293) );
  OAI21_X1 U5843 ( .B1(n7823), .B2(n5129), .A(n5126), .ZN(n8028) );
  INV_X1 U5844 ( .A(n5130), .ZN(n5129) );
  AND2_X1 U5845 ( .A1(n5366), .A2(n5127), .ZN(n5126) );
  OR2_X1 U5846 ( .A1(n5369), .A2(n5367), .ZN(n5366) );
  AND4_X1 U5847 ( .A1(n6071), .A2(n6070), .A3(n6069), .A4(n6068), .ZN(n9081)
         );
  AND4_X1 U5848 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n9068)
         );
  AND2_X1 U5849 ( .A1(n8946), .A2(n8025), .ZN(n5369) );
  NAND2_X1 U5850 ( .A1(n7869), .A2(n7868), .ZN(n7871) );
  AND4_X1 U5851 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n8518)
         );
  NAND2_X1 U5852 ( .A1(n7823), .A2(n8866), .ZN(n7869) );
  NAND2_X1 U5853 ( .A1(n5424), .A2(n5422), .ZN(n8029) );
  NOR2_X1 U5854 ( .A1(n7761), .A2(n5423), .ZN(n5422) );
  INV_X1 U5855 ( .A(n8933), .ZN(n5423) );
  OR2_X1 U5856 ( .A1(n5994), .A2(n5993), .ZN(n6013) );
  OAI21_X1 U5857 ( .B1(n7750), .B2(n8864), .A(n5069), .ZN(n7752) );
  NAND2_X1 U5858 ( .A1(n5138), .A2(n5078), .ZN(n7746) );
  INV_X1 U5859 ( .A(n7714), .ZN(n5138) );
  AND2_X1 U5860 ( .A1(n7670), .A2(n7569), .ZN(n7571) );
  NAND2_X1 U5861 ( .A1(n7571), .A2(n7570), .ZN(n7715) );
  NAND2_X1 U5862 ( .A1(n5406), .A2(n5407), .ZN(n5404) );
  NAND2_X1 U5863 ( .A1(n9330), .A2(n7683), .ZN(n8921) );
  INV_X1 U5864 ( .A(n5408), .ZN(n5407) );
  NAND2_X1 U5865 ( .A1(n8921), .A2(n8920), .ZN(n8860) );
  INV_X1 U5866 ( .A(n5354), .ZN(n5353) );
  NAND2_X1 U5867 ( .A1(n7466), .A2(n7465), .ZN(n7485) );
  NAND2_X1 U5868 ( .A1(n5322), .A2(n10886), .ZN(n7482) );
  INV_X1 U5869 ( .A(n7385), .ZN(n5322) );
  INV_X1 U5870 ( .A(n8862), .ZN(n8896) );
  NAND2_X1 U5871 ( .A1(n7258), .A2(n10852), .ZN(n7385) );
  AND4_X2 U5872 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n7254)
         );
  NAND2_X1 U5873 ( .A1(n7243), .A2(n7242), .ZN(n7262) );
  OR2_X1 U5874 ( .A1(n11125), .A2(n10922), .ZN(n7236) );
  INV_X1 U5875 ( .A(n5638), .ZN(n5347) );
  NAND2_X1 U5876 ( .A1(n9419), .A2(n9187), .ZN(n9405) );
  NAND2_X1 U5877 ( .A1(n9425), .A2(n9443), .ZN(n9187) );
  NAND2_X1 U5878 ( .A1(n6287), .A2(n6286), .ZN(n9600) );
  NAND2_X1 U5879 ( .A1(n6267), .A2(n6266), .ZN(n9607) );
  NAND2_X1 U5880 ( .A1(n6225), .A2(n6224), .ZN(n9615) );
  NAND2_X1 U5881 ( .A1(n6220), .A2(n6219), .ZN(n9620) );
  NAND2_X1 U5882 ( .A1(n6171), .A2(n6170), .ZN(n9635) );
  AND2_X1 U5883 ( .A1(n8026), .A2(n8025), .ZN(n8099) );
  NOR2_X1 U5884 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  INV_X1 U5885 ( .A(n11125), .ZN(n11067) );
  INV_X1 U5886 ( .A(n11066), .ZN(n11123) );
  AND2_X1 U5887 ( .A1(n6950), .A2(n6949), .ZN(n7234) );
  AND2_X1 U5888 ( .A1(n7236), .A2(n7231), .ZN(n6959) );
  XNOR2_X1 U5889 ( .A(n6321), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6329) );
  INV_X1 U5890 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5799) );
  INV_X1 U5891 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5795) );
  AND2_X1 U5892 ( .A1(n5988), .A2(n6008), .ZN(n7402) );
  INV_X1 U5893 ( .A(n5429), .ZN(n5955) );
  NOR2_X1 U5894 ( .A1(n5883), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U5895 ( .A1(n5764), .A2(n5765), .ZN(n5316) );
  NAND2_X1 U5896 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  INV_X1 U5897 ( .A(n9146), .ZN(n9147) );
  NAND2_X1 U5898 ( .A1(n5567), .A2(n9149), .ZN(n5566) );
  INV_X1 U5899 ( .A(n9695), .ZN(n5567) );
  NAND2_X1 U5900 ( .A1(n5523), .A2(n6698), .ZN(n6700) );
  NAND2_X1 U5901 ( .A1(n7548), .A2(n7547), .ZN(n5569) );
  NAND2_X1 U5902 ( .A1(n7441), .A2(n7440), .ZN(n7549) );
  AOI21_X1 U5903 ( .B1(n6640), .B2(n9159), .A(n6639), .ZN(n6645) );
  NOR2_X1 U5904 ( .A1(n8328), .A2(n9755), .ZN(n8337) );
  NAND2_X1 U5905 ( .A1(n5551), .A2(n5548), .ZN(n5556) );
  AND2_X1 U5906 ( .A1(n9777), .A2(n5552), .ZN(n5551) );
  AND2_X1 U5907 ( .A1(n7899), .A2(n7898), .ZN(n8006) );
  NAND2_X1 U5908 ( .A1(n7733), .A2(n7732), .ZN(n8003) );
  NAND2_X1 U5909 ( .A1(n8150), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6506) );
  BUF_X4 U5910 ( .A(n6825), .Z(n9160) );
  NAND2_X1 U5911 ( .A1(n8177), .A2(n8176), .ZN(n8180) );
  NOR2_X1 U5912 ( .A1(n5191), .A2(n5190), .ZN(n5189) );
  NAND2_X1 U5913 ( .A1(n8777), .A2(n8738), .ZN(n5190) );
  INV_X1 U5914 ( .A(n5196), .ZN(n5191) );
  AOI21_X1 U5915 ( .B1(n8743), .B2(n5053), .A(n8798), .ZN(n5195) );
  AOI22_X1 U5916 ( .A1(n6833), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n6834), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n6836) );
  AND2_X1 U5917 ( .A1(n5632), .A2(n6410), .ZN(n5214) );
  INV_X1 U5918 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U5919 ( .A1(n6986), .A2(n5396), .ZN(n6416) );
  AND2_X1 U5920 ( .A1(n6384), .A2(n5632), .ZN(n5396) );
  NAND2_X1 U5921 ( .A1(n5041), .A2(n9825), .ZN(n9824) );
  OR2_X1 U5922 ( .A1(n6547), .A2(n6546), .ZN(n6661) );
  NAND2_X1 U5923 ( .A1(n7327), .A2(n7328), .ZN(n7624) );
  XNOR2_X1 U5924 ( .A(n7794), .B(n7801), .ZN(n7626) );
  NAND2_X1 U5925 ( .A1(n7624), .A2(n5121), .ZN(n7794) );
  OR2_X1 U5926 ( .A1(n7960), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5121) );
  NOR2_X1 U5927 ( .A1(n7626), .A2(n7625), .ZN(n7795) );
  OR2_X1 U5928 ( .A1(n8109), .A2(n8108), .ZN(n5117) );
  AND2_X1 U5929 ( .A1(n5117), .A2(n5116), .ZN(n10722) );
  NAND2_X1 U5930 ( .A1(n9843), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5116) );
  INV_X1 U5931 ( .A(n8501), .ZN(n5270) );
  AND2_X1 U5932 ( .A1(n8718), .A2(n9867), .ZN(n9892) );
  INV_X1 U5933 ( .A(n8624), .ZN(n5380) );
  INV_X1 U5934 ( .A(n8707), .ZN(n5379) );
  AND2_X1 U5935 ( .A1(n9977), .A2(n5228), .ZN(n9924) );
  AND2_X1 U5936 ( .A1(n5229), .A2(n9916), .ZN(n5228) );
  NAND2_X1 U5937 ( .A1(n9977), .A2(n5229), .ZN(n9934) );
  AOI21_X1 U5938 ( .B1(n5610), .B2(n5612), .A(n5059), .ZN(n5608) );
  AND2_X1 U5939 ( .A1(n8556), .A2(n8700), .ZN(n9970) );
  NAND2_X1 U5940 ( .A1(n9977), .A2(n9967), .ZN(n9961) );
  AND2_X1 U5941 ( .A1(n8555), .A2(n8551), .ZN(n9984) );
  AND2_X1 U5942 ( .A1(n5244), .A2(n8458), .ZN(n5243) );
  NAND2_X1 U5943 ( .A1(n5246), .A2(n5249), .ZN(n5244) );
  OAI21_X1 U5944 ( .B1(n8457), .B2(n5249), .A(n5246), .ZN(n10013) );
  AND2_X1 U5945 ( .A1(n8067), .A2(n5081), .ZN(n10008) );
  NAND2_X1 U5946 ( .A1(n8067), .A2(n5235), .ZN(n10038) );
  NAND2_X1 U5947 ( .A1(n5245), .A2(n8680), .ZN(n10027) );
  NAND2_X1 U5948 ( .A1(n8457), .A2(n8681), .ZN(n5245) );
  NOR2_X1 U5949 ( .A1(n7968), .A2(n7967), .ZN(n8148) );
  NAND2_X1 U5950 ( .A1(n8067), .A2(n11110), .ZN(n8159) );
  AND2_X1 U5951 ( .A1(n8674), .A2(n8673), .ZN(n8763) );
  AND2_X1 U5952 ( .A1(n7992), .A2(n11094), .ZN(n8067) );
  NAND2_X1 U5953 ( .A1(n5225), .A2(n5227), .ZN(n5224) );
  INV_X1 U5954 ( .A(n11054), .ZN(n5227) );
  NOR2_X1 U5955 ( .A1(n7521), .A2(n6474), .ZN(n7645) );
  NAND2_X1 U5956 ( .A1(n5255), .A2(n7643), .ZN(n7964) );
  NAND2_X1 U5957 ( .A1(n7610), .A2(n5256), .ZN(n5255) );
  NAND2_X1 U5958 ( .A1(n7610), .A2(n8646), .ZN(n7642) );
  NOR2_X1 U5959 ( .A1(n10988), .A2(n5226), .ZN(n7613) );
  AND2_X1 U5960 ( .A1(n8649), .A2(n8646), .ZN(n8756) );
  NAND2_X1 U5961 ( .A1(n5383), .A2(n5388), .ZN(n10997) );
  NAND2_X1 U5962 ( .A1(n8780), .A2(n8639), .ZN(n5383) );
  NAND2_X1 U5963 ( .A1(n7532), .A2(n7531), .ZN(n10986) );
  OAI21_X1 U5964 ( .B1(n8780), .B2(n7301), .A(n8639), .ZN(n7494) );
  NAND2_X1 U5965 ( .A1(n5215), .A2(n10913), .ZN(n7154) );
  NOR2_X1 U5966 ( .A1(n7154), .A2(n10935), .ZN(n7338) );
  AND3_X1 U5967 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7045) );
  NAND2_X1 U5968 ( .A1(n7160), .A2(n8586), .ZN(n7111) );
  INV_X1 U5969 ( .A(n8750), .ZN(n7094) );
  NAND2_X1 U5970 ( .A1(n7109), .A2(n8583), .ZN(n7278) );
  INV_X1 U5971 ( .A(n10870), .ZN(n5216) );
  NOR2_X1 U5972 ( .A1(n7192), .A2(n7183), .ZN(n10868) );
  NAND2_X1 U5973 ( .A1(n10868), .A2(n10880), .ZN(n10870) );
  NAND2_X1 U5974 ( .A1(n7172), .A2(n8746), .ZN(n7088) );
  OAI22_X1 U5975 ( .A1(n7186), .A2(n7187), .B1(n7197), .B2(n7085), .ZN(n7172)
         );
  INV_X1 U5976 ( .A(n8746), .ZN(n7173) );
  NAND2_X1 U5977 ( .A1(n6680), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U5978 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  AND2_X1 U5979 ( .A1(n7103), .A2(n11057), .ZN(n10911) );
  INV_X1 U5980 ( .A(n7197), .ZN(n10824) );
  XNOR2_X1 U5981 ( .A(n8538), .B(n8537), .ZN(n9678) );
  NAND2_X1 U5982 ( .A1(n8535), .A2(n8534), .ZN(n8538) );
  XNOR2_X1 U5983 ( .A(n8527), .B(n8528), .ZN(n8443) );
  AND2_X1 U5984 ( .A1(n5762), .A2(n8438), .ZN(n5763) );
  NAND2_X1 U5985 ( .A1(n6388), .A2(n6389), .ZN(n6409) );
  INV_X1 U5986 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6385) );
  XNOR2_X1 U5987 ( .A(n6223), .B(n6222), .ZN(n8373) );
  AND2_X1 U5988 ( .A1(n6394), .A2(n6382), .ZN(n5572) );
  AND3_X1 U5989 ( .A1(n10565), .A2(n10571), .A3(n10572), .ZN(n6394) );
  NAND2_X1 U5990 ( .A1(n5513), .A2(n5510), .ZN(n6133) );
  NAND2_X1 U5991 ( .A1(n6097), .A2(n5514), .ZN(n5513) );
  NAND2_X1 U5992 ( .A1(n5509), .A2(n5710), .ZN(n6115) );
  AND2_X1 U5993 ( .A1(n6908), .A2(n6876), .ZN(n7878) );
  NAND2_X1 U5994 ( .A1(n5495), .A2(n5680), .ZN(n5982) );
  NAND2_X1 U5995 ( .A1(n5967), .A2(n5640), .ZN(n5495) );
  AND2_X1 U5996 ( .A1(n6502), .A2(n6501), .ZN(n7292) );
  NAND2_X1 U5997 ( .A1(n5263), .A2(n5671), .ZN(n5959) );
  NOR2_X1 U5998 ( .A1(n5185), .A2(n5181), .ZN(n5180) );
  INV_X1 U5999 ( .A(n5881), .ZN(n5181) );
  NAND2_X1 U6000 ( .A1(n6063), .A2(n6062), .ZN(n11101) );
  NAND2_X1 U6001 ( .A1(n7705), .A2(n5981), .ZN(n7688) );
  AND2_X1 U6002 ( .A1(n9043), .A2(n6354), .ZN(n9251) );
  NAND2_X1 U6003 ( .A1(n6109), .A2(n8215), .ZN(n8221) );
  AND3_X1 U6004 ( .A1(n6239), .A2(n6238), .A3(n6237), .ZN(n9284) );
  NOR3_X1 U6005 ( .A1(n10362), .A2(n10361), .A3(n10360), .ZN(n10375) );
  AND4_X1 U6006 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n7695)
         );
  AOI21_X1 U6007 ( .B1(n5577), .B2(n5579), .A(n5095), .ZN(n5575) );
  INV_X1 U6008 ( .A(n6036), .ZN(n5579) );
  OAI21_X1 U6009 ( .B1(n9238), .B2(n5586), .A(n5583), .ZN(n9279) );
  NAND2_X1 U6010 ( .A1(n9238), .A2(n6184), .ZN(n5582) );
  NAND2_X1 U6011 ( .A1(n5916), .A2(n5915), .ZN(n8491) );
  AND2_X1 U6012 ( .A1(n7014), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10616) );
  AND2_X1 U6013 ( .A1(n9305), .A2(n5592), .ZN(n5591) );
  INV_X1 U6014 ( .A(n6246), .ZN(n5587) );
  INV_X1 U6015 ( .A(n10616), .ZN(n9294) );
  INV_X1 U6016 ( .A(n7695), .ZN(n9329) );
  OR2_X1 U6017 ( .A1(n5922), .A2(n7474), .ZN(n5888) );
  OR2_X1 U6018 ( .A1(n6365), .A2(n10770), .ZN(n5176) );
  OR2_X1 U6019 ( .A1(n8842), .A2(n6738), .ZN(n5820) );
  AOI21_X1 U6020 ( .B1(n6735), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6753), .ZN(
        n6767) );
  AOI21_X1 U6021 ( .B1(n6733), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6765), .ZN(
        n6779) );
  AOI21_X1 U6022 ( .B1(n6804), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6803), .ZN(
        n6808) );
  NOR2_X1 U6023 ( .A1(n5968), .A2(n5792), .ZN(n6026) );
  AND2_X1 U6024 ( .A1(n6489), .A2(n6488), .ZN(n10787) );
  AOI21_X1 U6025 ( .B1(n9349), .B2(P2_REG2_REG_16__SCAN_IN), .A(n9348), .ZN(
        n9352) );
  INV_X1 U6026 ( .A(n9400), .ZN(n9588) );
  NAND2_X1 U6027 ( .A1(n9399), .A2(n9588), .ZN(n9585) );
  AND2_X1 U6028 ( .A1(n8828), .A2(n8827), .ZN(n9191) );
  AND2_X1 U6029 ( .A1(n9432), .A2(n9431), .ZN(n9603) );
  NAND2_X1 U6030 ( .A1(n9436), .A2(n5636), .ZN(n9421) );
  INV_X1 U6031 ( .A(n9607), .ZN(n9450) );
  AND2_X1 U6032 ( .A1(n8821), .A2(n8992), .ZN(n5645) );
  AND2_X1 U6033 ( .A1(n5363), .A2(n5361), .ZN(n9483) );
  NOR2_X1 U6034 ( .A1(n9509), .A2(n9180), .ZN(n9496) );
  NAND2_X1 U6035 ( .A1(n5416), .A2(n8816), .ZN(n9544) );
  NAND2_X1 U6036 ( .A1(n9570), .A2(n9561), .ZN(n5416) );
  NAND2_X1 U6037 ( .A1(n8290), .A2(n5352), .ZN(n9174) );
  NAND2_X1 U6038 ( .A1(n6043), .A2(n6042), .ZN(n9067) );
  AND2_X1 U6039 ( .A1(n5424), .A2(n7760), .ZN(n7813) );
  INV_X1 U6040 ( .A(n10959), .ZN(n7683) );
  NAND2_X1 U6041 ( .A1(n7466), .A2(n5411), .ZN(n5410) );
  INV_X1 U6042 ( .A(n7359), .ZN(n5357) );
  INV_X1 U6043 ( .A(n10832), .ZN(n7258) );
  INV_X1 U6044 ( .A(n9568), .ZN(n9542) );
  AND3_X2 U6045 ( .A1(n7234), .A2(n6959), .A3(n7232), .ZN(n11132) );
  AND2_X1 U6046 ( .A1(n6486), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10760) );
  OR2_X1 U6047 ( .A1(n5816), .A2(n9679), .ZN(n5814) );
  NAND2_X1 U6048 ( .A1(n5781), .A2(n5780), .ZN(n5783) );
  NAND2_X1 U6049 ( .A1(n5784), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5785) );
  INV_X1 U6050 ( .A(n6329), .ZN(n8089) );
  INV_X1 U6051 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7778) );
  INV_X1 U6052 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8305) );
  INV_X1 U6053 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7058) );
  INV_X1 U6054 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6676) );
  INV_X1 U6055 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6576) );
  INV_X1 U6056 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6514) );
  INV_X1 U6057 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6504) );
  INV_X1 U6058 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U6059 ( .A1(n7213), .A2(n7214), .ZN(n7438) );
  NAND2_X1 U6060 ( .A1(n5544), .A2(n7212), .ZN(n7213) );
  NAND2_X1 U6061 ( .A1(n7071), .A2(n7207), .ZN(n5544) );
  NAND2_X1 U6062 ( .A1(n9788), .A2(n9149), .ZN(n9697) );
  NAND2_X2 U6063 ( .A1(n8414), .A2(n8413), .ZN(n10062) );
  NAND2_X1 U6064 ( .A1(n7962), .A2(n7961), .ZN(n8046) );
  NAND2_X1 U6065 ( .A1(n5548), .A2(n9777), .ZN(n9715) );
  AND2_X1 U6066 ( .A1(n5564), .A2(n5563), .ZN(n5558) );
  OAI21_X1 U6067 ( .B1(n5564), .B2(n9163), .A(n5560), .ZN(n5559) );
  NAND2_X1 U6068 ( .A1(n5564), .A2(n5561), .ZN(n5560) );
  NAND2_X1 U6069 ( .A1(n5566), .A2(n5563), .ZN(n5561) );
  OR2_X1 U6070 ( .A1(n5566), .A2(n5563), .ZN(n5562) );
  NAND2_X1 U6071 ( .A1(n5524), .A2(n6697), .ZN(n6702) );
  NAND2_X1 U6072 ( .A1(n5546), .A2(n5549), .ZN(n9727) );
  NAND2_X1 U6073 ( .A1(n5550), .A2(n5554), .ZN(n5549) );
  NAND2_X1 U6074 ( .A1(n5076), .A2(n5555), .ZN(n5550) );
  NAND2_X1 U6075 ( .A1(n5526), .A2(n5525), .ZN(n9737) );
  INV_X1 U6076 ( .A(n5530), .ZN(n5525) );
  OAI21_X1 U6077 ( .B1(n5534), .B2(n5529), .A(n9132), .ZN(n5530) );
  NAND2_X1 U6078 ( .A1(n8147), .A2(n8146), .ZN(n10119) );
  NAND2_X1 U6079 ( .A1(n5533), .A2(n5532), .ZN(n9744) );
  AOI21_X1 U6080 ( .B1(n9704), .B2(n9707), .A(n5536), .ZN(n5532) );
  INV_X1 U6081 ( .A(n6934), .ZN(n6935) );
  NAND2_X1 U6082 ( .A1(n7498), .A2(n7497), .ZN(n10987) );
  AND2_X1 U6083 ( .A1(n6705), .A2(n10990), .ZN(n9791) );
  NAND2_X1 U6084 ( .A1(n8327), .A2(n8326), .ZN(n10097) );
  INV_X1 U6085 ( .A(n9802), .ZN(n10018) );
  CLKBUF_X1 U6086 ( .A(n7208), .Z(n7071) );
  INV_X1 U6087 ( .A(n9785), .ZN(n9787) );
  AND2_X1 U6088 ( .A1(n8428), .A2(n8405), .ZN(n9887) );
  INV_X1 U6089 ( .A(n9760), .ZN(n9796) );
  XNOR2_X1 U6090 ( .A(n6682), .B(n6524), .ZN(n6525) );
  NAND2_X1 U6091 ( .A1(n6525), .A2(n9813), .ZN(n6535) );
  INV_X1 U6092 ( .A(n5120), .ZN(n10732) );
  NAND2_X1 U6093 ( .A1(n10685), .A2(n10684), .ZN(n10683) );
  AND2_X1 U6094 ( .A1(n5120), .A2(n5119), .ZN(n10685) );
  NAND2_X1 U6095 ( .A1(n6559), .A2(n6541), .ZN(n5119) );
  NAND2_X1 U6096 ( .A1(n7003), .A2(n7004), .ZN(n10708) );
  NOR2_X1 U6097 ( .A1(n8106), .A2(n5118), .ZN(n8109) );
  AND2_X1 U6098 ( .A1(n8145), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5118) );
  INV_X1 U6099 ( .A(n5117), .ZN(n9842) );
  INV_X1 U6100 ( .A(n9852), .ZN(n10048) );
  NAND2_X1 U6101 ( .A1(n5222), .A2(n10053), .ZN(n5221) );
  XNOR2_X1 U6102 ( .A(n8456), .B(n8773), .ZN(n10056) );
  NAND2_X1 U6103 ( .A1(n8494), .A2(n5635), .ZN(n8456) );
  OR2_X1 U6104 ( .A1(n5220), .A2(n9700), .ZN(n5635) );
  AOI21_X1 U6105 ( .B1(n9874), .B2(n10998), .A(n9873), .ZN(n10065) );
  NAND2_X1 U6106 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  OAI21_X1 U6107 ( .B1(n9914), .B2(n5044), .A(n8384), .ZN(n9898) );
  NAND2_X1 U6108 ( .A1(n9918), .A2(n9919), .ZN(n9917) );
  NAND2_X1 U6109 ( .A1(n9959), .A2(n8347), .ZN(n9947) );
  AND2_X1 U6110 ( .A1(n8322), .A2(n8321), .ZN(n9998) );
  INV_X1 U6111 ( .A(n10879), .ZN(n11012) );
  NAND2_X1 U6112 ( .A1(n7983), .A2(n7958), .ZN(n8049) );
  AND2_X1 U6113 ( .A1(n7956), .A2(n7955), .ZN(n7984) );
  NAND2_X1 U6114 ( .A1(n7287), .A2(n8634), .ZN(n7334) );
  NAND2_X1 U6115 ( .A1(n5618), .A2(n7093), .ZN(n7148) );
  INV_X1 U6116 ( .A(n7118), .ZN(n7191) );
  INV_X1 U6117 ( .A(n11016), .ZN(n9863) );
  NAND2_X1 U6118 ( .A1(n8505), .A2(n11114), .ZN(n5268) );
  AND2_X1 U6119 ( .A1(n6879), .A2(n6424), .ZN(n10669) );
  INV_X1 U6120 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10139) );
  INV_X1 U6121 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6466) );
  INV_X1 U6122 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7777) );
  INV_X1 U6123 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10511) );
  INV_X1 U6124 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10516) );
  INV_X1 U6125 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10525) );
  INV_X1 U6126 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10528) );
  INV_X1 U6127 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10321) );
  INV_X1 U6128 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10543) );
  AND2_X1 U6129 ( .A1(n6462), .A2(n6459), .ZN(n10682) );
  NOR2_X1 U6130 ( .A1(n7941), .A2(n7940), .ZN(n10656) );
  NOR2_X1 U6131 ( .A1(n10654), .A2(n10653), .ZN(n7940) );
  OAI21_X1 U6132 ( .B1(n6350), .B2(n10611), .A(n5573), .ZN(n6372) );
  AND2_X1 U6133 ( .A1(n7009), .A2(n5836), .ZN(n6980) );
  INV_X1 U6134 ( .A(n5489), .ZN(n5488) );
  OAI211_X1 U6135 ( .C1(n9594), .C2(n5039), .A(n5348), .B(n5339), .ZN(P2_U3517) );
  NAND2_X1 U6136 ( .A1(n5340), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5348) );
  OR2_X1 U6137 ( .A1(n9593), .A2(n5340), .ZN(n5339) );
  OR2_X1 U6138 ( .A1(n8812), .A2(n8811), .ZN(n5104) );
  NAND2_X1 U6139 ( .A1(n5113), .A2(n5062), .ZN(P1_U3260) );
  OR2_X1 U6140 ( .A1(n5114), .A2(n10808), .ZN(n5113) );
  XNOR2_X1 U6141 ( .A(n9848), .B(n9847), .ZN(n5114) );
  NAND2_X1 U6142 ( .A1(n5266), .A2(n5264), .ZN(P1_U3551) );
  OR2_X1 U6143 ( .A1(n10847), .A2(n5265), .ZN(n5264) );
  NAND2_X1 U6144 ( .A1(n10125), .A2(n10847), .ZN(n5266) );
  INV_X1 U6145 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5265) );
  AND2_X1 U6146 ( .A1(n8761), .A2(n7955), .ZN(n5029) );
  OR2_X1 U6147 ( .A1(n10062), .A2(n9893), .ZN(n5030) );
  OR2_X1 U6148 ( .A1(n5792), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5031) );
  OR2_X1 U6149 ( .A1(n8048), .A2(n5626), .ZN(n5032) );
  AND2_X1 U6150 ( .A1(n5384), .A2(n5387), .ZN(n5033) );
  AND2_X1 U6151 ( .A1(n9331), .A2(n10943), .ZN(n5034) );
  INV_X1 U6152 ( .A(n8798), .ZN(n8777) );
  OR2_X2 U6153 ( .A1(n5031), .A2(n5067), .ZN(n5035) );
  AND2_X1 U6154 ( .A1(n9069), .A2(n6038), .ZN(n5036) );
  NAND2_X1 U6155 ( .A1(n5768), .A2(n5767), .ZN(n5883) );
  INV_X1 U6156 ( .A(n5146), .ZN(n5145) );
  OAI21_X1 U6157 ( .B1(n8917), .B2(n8918), .A(n8914), .ZN(n5146) );
  OR2_X1 U6158 ( .A1(n10062), .A2(n8419), .ZN(n8778) );
  INV_X1 U6159 ( .A(n5143), .ZN(n5142) );
  NAND2_X1 U6160 ( .A1(n5073), .A2(n5144), .ZN(n5143) );
  AND2_X1 U6161 ( .A1(n6216), .A2(n6215), .ZN(n5037) );
  AND2_X1 U6162 ( .A1(n7094), .A2(n7093), .ZN(n5038) );
  NAND2_X1 U6163 ( .A1(n9977), .A2(n5231), .ZN(n5232) );
  NAND2_X1 U6164 ( .A1(n6885), .A2(n5606), .ZN(n7089) );
  INV_X1 U6165 ( .A(n7089), .ZN(n10880) );
  OR2_X1 U6166 ( .A1(n5340), .A2(n11082), .ZN(n5039) );
  NAND2_X1 U6167 ( .A1(n7296), .A2(n8753), .ZN(n7532) );
  AND2_X1 U6168 ( .A1(n6348), .A2(n6354), .ZN(n10623) );
  OR2_X1 U6169 ( .A1(n10988), .A2(n5224), .ZN(n5040) );
  INV_X1 U6170 ( .A(n8421), .ZN(n7291) );
  AND2_X4 U6171 ( .A1(n6681), .A2(n6680), .ZN(n8421) );
  NOR2_X1 U6172 ( .A1(n5784), .A2(n5433), .ZN(n5816) );
  AND2_X1 U6173 ( .A1(n10745), .A2(n6538), .ZN(n5041) );
  AND4_X1 U6174 ( .A1(n5931), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n7559)
         );
  NAND2_X1 U6175 ( .A1(n5582), .A2(n9239), .ZN(n9241) );
  AND2_X1 U6176 ( .A1(n9859), .A2(n5221), .ZN(n5042) );
  AND2_X1 U6177 ( .A1(n6986), .A2(n6384), .ZN(n6388) );
  AND2_X1 U6178 ( .A1(n9490), .A2(n8992), .ZN(n5043) );
  NAND2_X1 U6179 ( .A1(n6252), .A2(n6251), .ZN(n9611) );
  AND2_X1 U6180 ( .A1(n8941), .A2(n8030), .ZN(n8939) );
  INV_X1 U6181 ( .A(n8939), .ZN(n5370) );
  AND2_X1 U6182 ( .A1(n10078), .A2(n9942), .ZN(n5044) );
  OR2_X1 U6183 ( .A1(n6681), .A2(n10810), .ZN(n5045) );
  NOR2_X1 U6184 ( .A1(n10097), .A2(n10001), .ZN(n5046) );
  AND2_X1 U6185 ( .A1(n8727), .A2(n8549), .ZN(n8791) );
  NAND2_X1 U6186 ( .A1(n8894), .A2(n8897), .ZN(n7353) );
  XOR2_X1 U6187 ( .A(n9040), .B(n10922), .Z(n5047) );
  XNOR2_X1 U6188 ( .A(n5814), .B(n5813), .ZN(n5819) );
  INV_X1 U6189 ( .A(n5819), .ZN(n5818) );
  AND2_X1 U6190 ( .A1(n5932), .A2(n5182), .ZN(n5048) );
  OR2_X1 U6191 ( .A1(n5664), .A2(n5663), .ZN(n5049) );
  AND2_X1 U6192 ( .A1(n5556), .A2(n5555), .ZN(n5050) );
  INV_X1 U6193 ( .A(n9595), .ZN(n5324) );
  INV_X1 U6194 ( .A(n10057), .ZN(n5220) );
  XNOR2_X1 U6195 ( .A(n9625), .B(n9519), .ZN(n9182) );
  XNOR2_X1 U6196 ( .A(n10863), .B(n7086), .ZN(n8746) );
  NAND2_X1 U6197 ( .A1(n5363), .A2(n5364), .ZN(n9482) );
  NOR2_X1 U6198 ( .A1(n8004), .A2(n8006), .ZN(n5051) );
  AND2_X1 U6199 ( .A1(n9015), .A2(n9016), .ZN(n9427) );
  NOR2_X1 U6200 ( .A1(n7758), .A2(n7759), .ZN(n5052) );
  INV_X1 U6201 ( .A(n5675), .ZN(n5494) );
  AND2_X1 U6202 ( .A1(n8449), .A2(n8448), .ZN(n8473) );
  INV_X1 U6203 ( .A(n8473), .ZN(n10053) );
  AND2_X1 U6204 ( .A1(n8804), .A2(n8744), .ZN(n5053) );
  NAND2_X1 U6205 ( .A1(n5429), .A2(n5428), .ZN(n5805) );
  OR3_X1 U6206 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .A3(
        P2_IR_REG_22__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6207 ( .A1(n8361), .A2(n8360), .ZN(n10082) );
  INV_X1 U6208 ( .A(n10886), .ZN(n8898) );
  AND3_X1 U6209 ( .A1(n5857), .A2(n5856), .A3(n5855), .ZN(n10886) );
  AND2_X1 U6210 ( .A1(n9868), .A2(n9867), .ZN(n5055) );
  NAND2_X1 U6211 ( .A1(n6188), .A2(n6187), .ZN(n9630) );
  AND2_X1 U6212 ( .A1(n10987), .A2(n9808), .ZN(n5056) );
  NOR2_X1 U6213 ( .A1(n9079), .A2(n9322), .ZN(n5057) );
  NAND2_X1 U6214 ( .A1(n8053), .A2(n8052), .ZN(n8191) );
  INV_X1 U6215 ( .A(n8963), .ZN(n8272) );
  AND2_X1 U6216 ( .A1(n8966), .A2(n8965), .ZN(n8963) );
  NAND2_X1 U6217 ( .A1(n6083), .A2(n6082), .ZN(n9079) );
  AND2_X1 U6218 ( .A1(n8917), .A2(n8915), .ZN(n5058) );
  AND2_X1 U6219 ( .A1(n10087), .A2(n9971), .ZN(n5059) );
  AND2_X1 U6220 ( .A1(n6248), .A2(n6247), .ZN(n5060) );
  INV_X1 U6221 ( .A(n9746), .ZN(n5536) );
  AND2_X1 U6222 ( .A1(n5821), .A2(n5822), .ZN(n5061) );
  AND2_X1 U6223 ( .A1(n5112), .A2(n5110), .ZN(n5062) );
  INV_X1 U6224 ( .A(n5325), .ZN(n9422) );
  NOR2_X1 U6225 ( .A1(n9444), .A2(n9600), .ZN(n5325) );
  INV_X1 U6226 ( .A(n8771), .ZN(n8496) );
  AND2_X1 U6227 ( .A1(n8549), .A2(n8725), .ZN(n8771) );
  NAND2_X1 U6228 ( .A1(n8637), .A2(n8645), .ZN(n10995) );
  OR2_X1 U6229 ( .A1(n11094), .A2(n8047), .ZN(n5063) );
  INV_X1 U6230 ( .A(n5122), .ZN(n10804) );
  NAND2_X1 U6231 ( .A1(n6534), .A2(n6535), .ZN(n5122) );
  NOR2_X1 U6232 ( .A1(n7289), .A2(n9809), .ZN(n5064) );
  AND2_X1 U6233 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n5065) );
  NOR2_X1 U6234 ( .A1(n9595), .A2(n9213), .ZN(n5066) );
  INV_X1 U6235 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6389) );
  NAND3_X1 U6236 ( .A1(n6078), .A2(n6059), .A3(n5794), .ZN(n5067) );
  OR2_X1 U6237 ( .A1(n8667), .A2(n8668), .ZN(n5068) );
  OR2_X1 U6238 ( .A1(n9630), .A2(n9533), .ZN(n8988) );
  NAND2_X1 U6239 ( .A1(n7749), .A2(n11024), .ZN(n5069) );
  OR2_X1 U6240 ( .A1(n5955), .A2(n5777), .ZN(n5070) );
  INV_X1 U6241 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5793) );
  AND2_X1 U6242 ( .A1(n8666), .A2(n8660), .ZN(n5071) );
  AND2_X1 U6243 ( .A1(n5213), .A2(n5210), .ZN(n5072) );
  AND2_X1 U6244 ( .A1(n8923), .A2(n8922), .ZN(n5073) );
  OR2_X1 U6245 ( .A1(n9868), .A2(n5630), .ZN(n5074) );
  INV_X1 U6246 ( .A(n9331), .ZN(n9052) );
  NAND4_X1 U6247 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n9331)
         );
  NAND2_X1 U6248 ( .A1(n8316), .A2(n8315), .ZN(n10107) );
  OR2_X1 U6249 ( .A1(n5148), .A2(n5147), .ZN(n5075) );
  NAND2_X1 U6250 ( .A1(n9105), .A2(n9752), .ZN(n5076) );
  NAND2_X1 U6251 ( .A1(n8375), .A2(n8374), .ZN(n10078) );
  AND2_X1 U6252 ( .A1(n10904), .A2(n7473), .ZN(n5077) );
  NAND2_X1 U6253 ( .A1(n9329), .A2(n7713), .ZN(n5078) );
  AND2_X1 U6254 ( .A1(n5554), .A2(n5552), .ZN(n5079) );
  NOR2_X1 U6255 ( .A1(n9427), .A2(n5132), .ZN(n5080) );
  AND2_X1 U6256 ( .A1(n10011), .A2(n5233), .ZN(n5081) );
  INV_X1 U6257 ( .A(n8410), .ZN(n5631) );
  AND2_X1 U6258 ( .A1(n5641), .A2(n5496), .ZN(n5082) );
  AND2_X1 U6259 ( .A1(n9569), .A2(n5318), .ZN(n5083) );
  AND2_X1 U6260 ( .A1(n5137), .A2(n11129), .ZN(n5084) );
  INV_X1 U6261 ( .A(n5206), .ZN(n5205) );
  NAND2_X1 U6262 ( .A1(n8771), .A2(n5207), .ZN(n5206) );
  AND2_X1 U6263 ( .A1(n6935), .A2(n6924), .ZN(n5085) );
  AND2_X1 U6264 ( .A1(n5205), .A2(n5198), .ZN(n5086) );
  AND2_X1 U6265 ( .A1(n5364), .A2(n5362), .ZN(n5361) );
  INV_X1 U6266 ( .A(n9005), .ZN(n5166) );
  INV_X1 U6267 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9679) );
  INV_X1 U6268 ( .A(n9123), .ZN(n5529) );
  NAND2_X1 U6269 ( .A1(n8155), .A2(n8673), .ZN(n8457) );
  NAND2_X1 U6270 ( .A1(n8179), .A2(n8180), .ZN(n8227) );
  NAND2_X1 U6271 ( .A1(n8026), .A2(n5369), .ZN(n8100) );
  NAND2_X1 U6272 ( .A1(n7783), .A2(n6036), .ZN(n8081) );
  NAND2_X1 U6273 ( .A1(n8221), .A2(n6113), .ZN(n8260) );
  INV_X1 U6274 ( .A(n8903), .ZN(n5356) );
  NAND2_X1 U6275 ( .A1(n7289), .A2(n7288), .ZN(n8639) );
  INV_X1 U6276 ( .A(n8639), .ZN(n5386) );
  INV_X1 U6277 ( .A(n9239), .ZN(n5586) );
  NAND2_X1 U6278 ( .A1(n8291), .A2(n8272), .ZN(n8290) );
  NAND2_X1 U6279 ( .A1(n7514), .A2(n7513), .ZN(n7738) );
  NOR3_X1 U6280 ( .A1(n9551), .A2(n9620), .A3(n5329), .ZN(n5326) );
  NAND2_X1 U6281 ( .A1(n8067), .A2(n5233), .ZN(n5236) );
  OR2_X1 U6282 ( .A1(n6849), .A2(n6662), .ZN(n5087) );
  NAND2_X1 U6283 ( .A1(n8204), .A2(n5318), .ZN(n5088) );
  OR2_X1 U6284 ( .A1(n5644), .A2(n5637), .ZN(n5089) );
  INV_X1 U6285 ( .A(n5327), .ZN(n9497) );
  NOR2_X1 U6286 ( .A1(n9551), .A2(n5329), .ZN(n5327) );
  NAND2_X1 U6287 ( .A1(n5371), .A2(n5370), .ZN(n8026) );
  NAND2_X1 U6288 ( .A1(n8929), .A2(n8933), .ZN(n5090) );
  INV_X1 U6289 ( .A(n5106), .ZN(n6116) );
  NAND2_X1 U6290 ( .A1(n5108), .A2(n5107), .ZN(n5106) );
  NAND2_X1 U6291 ( .A1(n7503), .A2(n7502), .ZN(n7614) );
  AND2_X1 U6292 ( .A1(n5467), .A2(n5466), .ZN(n5091) );
  AND2_X1 U6293 ( .A1(n8290), .A2(n8273), .ZN(n5092) );
  OR2_X1 U6294 ( .A1(n5968), .A2(n5035), .ZN(n5093) );
  NAND2_X1 U6295 ( .A1(n5783), .A2(n5812), .ZN(n6355) );
  NAND2_X1 U6296 ( .A1(n6023), .A2(n7781), .ZN(n7783) );
  NAND2_X1 U6297 ( .A1(n5357), .A2(n7360), .ZN(n7469) );
  AND3_X2 U6298 ( .A1(n7234), .A2(n6959), .A3(n6951), .ZN(n11135) );
  INV_X1 U6299 ( .A(n11135), .ZN(n5340) );
  AOI21_X1 U6300 ( .B1(n7301), .B2(n8639), .A(n5389), .ZN(n5388) );
  OR2_X1 U6301 ( .A1(n10988), .A2(n10987), .ZN(n5094) );
  NAND2_X1 U6302 ( .A1(n5576), .A2(n5575), .ZN(n8516) );
  NAND2_X1 U6303 ( .A1(n8805), .A2(n9850), .ZN(n8735) );
  NAND2_X1 U6304 ( .A1(n5569), .A2(n7549), .ZN(n7575) );
  NAND2_X1 U6305 ( .A1(n7581), .A2(n7580), .ZN(n7731) );
  NAND2_X1 U6306 ( .A1(n5410), .A2(n8910), .ZN(n7558) );
  XOR2_X1 U6307 ( .A(n8519), .B(n6054), .Z(n5095) );
  INV_X1 U6308 ( .A(n5603), .ZN(n7175) );
  AND2_X1 U6309 ( .A1(n6357), .A2(n6353), .ZN(n10611) );
  OR2_X1 U6310 ( .A1(n7769), .A2(n5334), .ZN(n5096) );
  OR2_X1 U6311 ( .A1(n10988), .A2(n5223), .ZN(n5097) );
  NAND2_X1 U6312 ( .A1(n6925), .A2(n6924), .ZN(n6933) );
  INV_X1 U6313 ( .A(n7781), .ZN(n5578) );
  NAND2_X1 U6314 ( .A1(n5427), .A2(n5429), .ZN(n6322) );
  NOR2_X1 U6315 ( .A1(n7717), .A2(n8864), .ZN(n5098) );
  INV_X1 U6316 ( .A(n5115), .ZN(n6848) );
  NOR2_X1 U6317 ( .A1(n6664), .A2(n6663), .ZN(n5115) );
  NAND2_X1 U6318 ( .A1(n5216), .A2(n10894), .ZN(n7273) );
  INV_X1 U6319 ( .A(n7273), .ZN(n5215) );
  NAND2_X1 U6320 ( .A1(n7669), .A2(n7571), .ZN(n5099) );
  OR2_X1 U6321 ( .A1(n6322), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n5100) );
  INV_X1 U6322 ( .A(n5425), .ZN(n7762) );
  NAND2_X1 U6323 ( .A1(n7720), .A2(n8924), .ZN(n5425) );
  OR2_X1 U6324 ( .A1(n6647), .A2(n8524), .ZN(n6689) );
  INV_X1 U6325 ( .A(n10967), .ZN(n5187) );
  NAND2_X1 U6326 ( .A1(n6702), .A2(n6704), .ZN(n6701) );
  AND2_X1 U6327 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_209), .ZN(n5101)
         );
  AND4_X1 U6328 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n9332)
         );
  XNOR2_X1 U6329 ( .A(n5804), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8891) );
  INV_X1 U6330 ( .A(n8891), .ZN(n8843) );
  AND2_X1 U6331 ( .A1(n10561), .A2(n10560), .ZN(n5102) );
  OR2_X1 U6332 ( .A1(n10591), .A2(n10590), .ZN(n5103) );
  INV_X1 U6333 ( .A(n9047), .ZN(n5490) );
  NAND2_X1 U6334 ( .A1(n6826), .A2(n6827), .ZN(n6828) );
  NAND2_X1 U6335 ( .A1(n5105), .A2(n5104), .ZN(P1_U3240) );
  XNOR2_X1 U6336 ( .A(n6392), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6431) );
  NAND3_X1 U6337 ( .A1(n8179), .A2(n8180), .A3(n5545), .ZN(n8246) );
  NAND2_X1 U6338 ( .A1(n5179), .A2(n5652), .ZN(n5842) );
  NAND2_X1 U6339 ( .A1(n7033), .A2(n7032), .ZN(n7043) );
  OAI21_X1 U6340 ( .B1(n6007), .B2(n5687), .A(n5689), .ZN(n6025) );
  NAND2_X1 U6341 ( .A1(n6218), .A2(n6217), .ZN(n5743) );
  NAND2_X1 U6342 ( .A1(n5263), .A2(n5261), .ZN(n5676) );
  NAND2_X1 U6343 ( .A1(n5505), .A2(n5507), .ZN(n6151) );
  NAND2_X1 U6344 ( .A1(n5492), .A2(n5082), .ZN(n5685) );
  OAI21_X1 U6345 ( .B1(n5195), .B2(n9926), .A(n5196), .ZN(n5192) );
  NAND3_X1 U6346 ( .A1(n7009), .A2(n6979), .A3(n5836), .ZN(n6978) );
  NAND2_X1 U6347 ( .A1(n5833), .A2(n5832), .ZN(n7009) );
  INV_X1 U6348 ( .A(n5622), .ZN(n5621) );
  INV_X4 U6349 ( .A(n5650), .ZN(n6422) );
  NAND2_X1 U6350 ( .A1(n10060), .A2(n5267), .ZN(n10125) );
  INV_X1 U6351 ( .A(n6415), .ZN(n6412) );
  NAND2_X1 U6352 ( .A1(n7607), .A2(n7536), .ZN(n7631) );
  NAND2_X1 U6353 ( .A1(n6248), .A2(n5589), .ZN(n5588) );
  NAND2_X1 U6354 ( .A1(n5620), .A2(n5619), .ZN(n7297) );
  NOR2_X2 U6355 ( .A1(n5035), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5107) );
  NOR2_X2 U6356 ( .A1(n5955), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6357 ( .A1(n10994), .A2(n8645), .ZN(n7611) );
  NAND2_X2 U6358 ( .A1(n7611), .A2(n8756), .ZN(n7610) );
  AND2_X2 U6359 ( .A1(n10014), .A2(n8553), .ZN(n5646) );
  NAND2_X1 U6360 ( .A1(n9952), .A2(n9953), .ZN(n9951) );
  NAND2_X1 U6361 ( .A1(n7985), .A2(n7986), .ZN(n8056) );
  NAND2_X1 U6362 ( .A1(n5123), .A2(n5659), .ZN(n5899) );
  NAND2_X1 U6363 ( .A1(n5180), .A2(n5186), .ZN(n5133) );
  INV_X1 U6364 ( .A(n9824), .ZN(n6539) );
  OAI21_X1 U6365 ( .B1(n10697), .B2(n9849), .A(n9841), .ZN(n5111) );
  XNOR2_X1 U6366 ( .A(n5123), .B(n5872), .ZN(n6926) );
  NAND2_X1 U6367 ( .A1(n5658), .A2(n5657), .ZN(n5123) );
  MUX2_X1 U6368 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5650), .Z(n5807) );
  AND2_X2 U6369 ( .A1(n5125), .A2(n5124), .ZN(n5650) );
  NAND3_X1 U6370 ( .A1(n5485), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5124) );
  NAND3_X1 U6371 ( .A1(n5487), .A2(n9849), .A3(n5486), .ZN(n5125) );
  NAND2_X1 U6372 ( .A1(n8028), .A2(n8036), .ZN(n8200) );
  NAND2_X1 U6373 ( .A1(n9436), .A2(n5080), .ZN(n9419) );
  NAND3_X1 U6374 ( .A1(n5135), .A2(n5137), .A3(n5134), .ZN(n9594) );
  NAND3_X1 U6375 ( .A1(n5135), .A2(n5084), .A3(n5134), .ZN(n5136) );
  NAND2_X1 U6376 ( .A1(n5136), .A2(n9593), .ZN(n9664) );
  NAND2_X1 U6377 ( .A1(n5341), .A2(n5342), .ZN(n5137) );
  NAND2_X1 U6378 ( .A1(n8964), .A2(n5155), .ZN(n5154) );
  NAND2_X1 U6379 ( .A1(n5154), .A2(n5152), .ZN(n8975) );
  AND2_X2 U6380 ( .A1(n5768), .A2(n5597), .ZN(n5429) );
  NAND2_X1 U6381 ( .A1(n5160), .A2(n5161), .ZN(n9009) );
  NAND3_X1 U6382 ( .A1(n8991), .A2(n5165), .A3(n8990), .ZN(n5160) );
  NAND3_X2 U6383 ( .A1(n5820), .A2(n5176), .A3(n5061), .ZN(n7229) );
  NAND4_X1 U6384 ( .A1(n5177), .A2(n9041), .A3(n5421), .A4(n5490), .ZN(n5420)
         );
  NAND2_X1 U6385 ( .A1(n5178), .A2(n5654), .ZN(n5853) );
  NAND2_X1 U6386 ( .A1(n5842), .A2(n5843), .ZN(n5178) );
  NAND2_X1 U6387 ( .A1(n5807), .A2(n5808), .ZN(n5179) );
  NAND2_X1 U6388 ( .A1(n5899), .A2(n5665), .ZN(n5186) );
  NAND2_X1 U6389 ( .A1(n5187), .A2(n10992), .ZN(n8638) );
  NAND2_X1 U6390 ( .A1(n8739), .A2(n5189), .ZN(n5193) );
  NAND2_X1 U6391 ( .A1(n8739), .A2(n8738), .ZN(n5194) );
  NAND3_X1 U6392 ( .A1(n5203), .A2(n5198), .A3(n8717), .ZN(n5200) );
  AND2_X1 U6393 ( .A1(n5199), .A2(n5197), .ZN(n8724) );
  NAND2_X1 U6394 ( .A1(n8717), .A2(n5086), .ZN(n5197) );
  OR2_X1 U6395 ( .A1(n5206), .A2(n5204), .ZN(n5199) );
  NAND2_X1 U6396 ( .A1(n5201), .A2(n5200), .ZN(n8723) );
  INV_X1 U6397 ( .A(n8778), .ZN(n5208) );
  NAND3_X1 U6398 ( .A1(n6986), .A2(n6384), .A3(n5214), .ZN(n6415) );
  AND2_X2 U6399 ( .A1(n6447), .A2(n6380), .ZN(n6986) );
  NOR2_X2 U6400 ( .A1(n6377), .A2(n6376), .ZN(n6380) );
  AND2_X2 U6401 ( .A1(n6445), .A2(n10544), .ZN(n6447) );
  NAND2_X1 U6402 ( .A1(n9875), .A2(n8471), .ZN(n9877) );
  NAND2_X1 U6403 ( .A1(n9875), .A2(n5217), .ZN(n5222) );
  INV_X1 U6404 ( .A(n5232), .ZN(n9933) );
  INV_X1 U6405 ( .A(n5236), .ZN(n10037) );
  OAI21_X1 U6406 ( .B1(n6684), .B2(n6680), .A(n5239), .ZN(n5238) );
  NAND2_X4 U6407 ( .A1(n9816), .A2(n10675), .ZN(n6681) );
  NAND2_X1 U6408 ( .A1(n5238), .A2(n6681), .ZN(n5237) );
  MUX2_X1 U6409 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5650), .Z(n5653) );
  NAND2_X1 U6410 ( .A1(n8457), .A2(n5246), .ZN(n5242) );
  NAND2_X1 U6411 ( .A1(n5242), .A2(n5243), .ZN(n10014) );
  OAI21_X2 U6412 ( .B1(n7610), .B2(n5253), .A(n5250), .ZN(n7985) );
  AND2_X2 U6413 ( .A1(n6743), .A2(n6422), .ZN(n5934) );
  NAND3_X1 U6414 ( .A1(n5764), .A2(n5765), .A3(n5766), .ZN(n5902) );
  NAND2_X1 U6415 ( .A1(n5316), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5873) );
  NOR2_X2 U6416 ( .A1(n5054), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6417 ( .A1(n8204), .A2(n5083), .ZN(n9562) );
  INV_X1 U6418 ( .A(n5323), .ZN(n7481) );
  NAND2_X1 U6419 ( .A1(n6317), .A2(n5784), .ZN(n8240) );
  INV_X1 U6420 ( .A(n5326), .ZN(n9485) );
  INV_X1 U6421 ( .A(n7769), .ZN(n5331) );
  NAND2_X1 U6422 ( .A1(n5331), .A2(n5332), .ZN(n5642) );
  OR2_X4 U6423 ( .A1(n9686), .A2(n5818), .ZN(n8842) );
  INV_X1 U6424 ( .A(n9686), .ZN(n5336) );
  NAND2_X1 U6425 ( .A1(n7354), .A2(n7353), .ZN(n7356) );
  NAND2_X1 U6426 ( .A1(n5338), .A2(n10852), .ZN(n8894) );
  INV_X1 U6427 ( .A(n9332), .ZN(n5338) );
  OAI21_X1 U6428 ( .B1(n8291), .B2(n5351), .A(n5349), .ZN(n9560) );
  NAND2_X1 U6429 ( .A1(n7359), .A2(n8903), .ZN(n5355) );
  OAI21_X1 U6430 ( .B1(n7360), .B2(n5356), .A(n7470), .ZN(n5354) );
  NAND2_X1 U6431 ( .A1(n5355), .A2(n5353), .ZN(n7472) );
  AOI21_X1 U6432 ( .B1(n5358), .B2(n5361), .A(n5359), .ZN(n9469) );
  INV_X1 U6433 ( .A(n7871), .ZN(n5371) );
  NAND3_X1 U6434 ( .A1(n5427), .A2(n5429), .A3(n5372), .ZN(n5812) );
  AOI21_X1 U6435 ( .B1(n9454), .B2(n9461), .A(n9186), .ZN(n9438) );
  AOI21_X1 U6436 ( .B1(n8271), .B2(n8270), .A(n5057), .ZN(n8291) );
  NAND2_X1 U6437 ( .A1(n7755), .A2(n7754), .ZN(n7822) );
  NAND2_X1 U6438 ( .A1(n9470), .A2(n9185), .ZN(n9454) );
  NOR2_X2 U6439 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5770) );
  AOI21_X1 U6441 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(n10262) );
  NAND2_X1 U6442 ( .A1(n10236), .A2(n10235), .ZN(n10240) );
  INV_X1 U6443 ( .A(n10214), .ZN(n10220) );
  NAND2_X1 U6444 ( .A1(n8057), .A2(n8763), .ZN(n8155) );
  AOI21_X2 U6445 ( .B1(n8056), .B2(n8055), .A(n8054), .ZN(n8057) );
  INV_X1 U6446 ( .A(n5375), .ZN(n9905) );
  NAND2_X1 U6447 ( .A1(n8581), .A2(n7173), .ZN(n7107) );
  NAND2_X1 U6448 ( .A1(n8780), .A2(n5384), .ZN(n5382) );
  INV_X1 U6449 ( .A(n8638), .ZN(n5389) );
  NAND2_X1 U6450 ( .A1(n5382), .A2(n5381), .ZN(n10994) );
  NOR2_X1 U6451 ( .A1(n10995), .A2(n5033), .ZN(n5381) );
  OAI21_X2 U6452 ( .B1(n7109), .B2(n5393), .A(n5390), .ZN(n8628) );
  AOI21_X1 U6453 ( .B1(n5392), .B2(n8586), .A(n5391), .ZN(n5390) );
  OR2_X1 U6454 ( .A1(n5395), .A2(n8582), .ZN(n5392) );
  NAND4_X1 U6455 ( .A1(n6395), .A2(n6381), .A3(n10571), .A4(n10568), .ZN(n5397) );
  AND2_X1 U6456 ( .A1(n7262), .A2(n8890), .ZN(n7264) );
  NAND2_X1 U6457 ( .A1(n5400), .A2(n5398), .ZN(n8830) );
  AOI21_X1 U6458 ( .B1(n5401), .B2(n9188), .A(n5399), .ZN(n5398) );
  NAND2_X1 U6459 ( .A1(n9426), .A2(n5401), .ZN(n5400) );
  NAND2_X1 U6460 ( .A1(n7466), .A2(n5406), .ZN(n5405) );
  OAI21_X1 U6461 ( .B1(n7466), .B2(n5407), .A(n5406), .ZN(n7676) );
  NAND3_X1 U6462 ( .A1(n5405), .A2(n8920), .A3(n5404), .ZN(n7719) );
  NAND2_X1 U6463 ( .A1(n9570), .A2(n5417), .ZN(n5413) );
  NAND2_X1 U6464 ( .A1(n5413), .A2(n5414), .ZN(n9532) );
  NAND2_X1 U6465 ( .A1(n5488), .A2(n5420), .ZN(P2_U3244) );
  NAND2_X1 U6466 ( .A1(n7720), .A2(n5426), .ZN(n5424) );
  NOR2_X1 U6467 ( .A1(n5784), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5782) );
  NAND3_X1 U6468 ( .A1(n10499), .A2(n10497), .A3(n10498), .ZN(n5483) );
  XNOR2_X1 U6469 ( .A(n5484), .B(n8545), .ZN(n9171) );
  NAND2_X1 U6470 ( .A1(n5676), .A2(n5493), .ZN(n5492) );
  OAI21_X2 U6471 ( .B1(n6250), .B2(n6249), .A(n5751), .ZN(n8437) );
  NAND2_X1 U6472 ( .A1(n6097), .A2(n5506), .ZN(n5505) );
  OR2_X1 U6473 ( .A1(n6097), .A2(n6096), .ZN(n5509) );
  NAND2_X1 U6474 ( .A1(n6186), .A2(n5519), .ZN(n5516) );
  OAI21_X1 U6475 ( .B1(n6186), .B2(n5521), .A(n5730), .ZN(n6203) );
  NAND2_X1 U6476 ( .A1(n5516), .A2(n5517), .ZN(n6218) );
  INV_X1 U6477 ( .A(n5524), .ZN(n5523) );
  NAND2_X1 U6478 ( .A1(n9124), .A2(n5527), .ZN(n5526) );
  OAI21_X1 U6479 ( .B1(n9706), .B2(n9707), .A(n9704), .ZN(n9745) );
  NAND2_X1 U6480 ( .A1(n7208), .A2(n5538), .ZN(n5537) );
  NAND2_X1 U6481 ( .A1(n8178), .A2(n8182), .ZN(n8179) );
  NAND2_X1 U6482 ( .A1(n8246), .A2(n8245), .ZN(n9094) );
  NAND2_X1 U6483 ( .A1(n5553), .A2(n5547), .ZN(n5546) );
  CLKBUF_X1 U6484 ( .A(n5553), .Z(n5548) );
  INV_X1 U6485 ( .A(n5556), .ZN(n9716) );
  NAND2_X1 U6486 ( .A1(n9753), .A2(n9106), .ZN(n5554) );
  NAND2_X1 U6487 ( .A1(n9790), .A2(n5558), .ZN(n5557) );
  OAI211_X1 U6488 ( .C1(n9790), .C2(n5562), .A(n5559), .B(n5557), .ZN(n9170)
         );
  NAND2_X1 U6489 ( .A1(n9790), .A2(n9789), .ZN(n9788) );
  NAND2_X1 U6490 ( .A1(n6925), .A2(n5085), .ZN(n7033) );
  NAND2_X1 U6491 ( .A1(n8015), .A2(n8012), .ZN(n8011) );
  NAND3_X1 U6492 ( .A1(n5569), .A2(n7577), .A3(n7549), .ZN(n7581) );
  OAI21_X1 U6493 ( .B1(n6402), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U6494 ( .A1(n6402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U6495 ( .A1(n6402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6606) );
  NAND3_X1 U6496 ( .A1(n6380), .A2(n6447), .A3(n6382), .ZN(n6989) );
  NAND3_X1 U6497 ( .A1(n6380), .A2(n6447), .A3(n5572), .ZN(n6400) );
  XNOR2_X1 U6498 ( .A(n6314), .B(n6313), .ZN(n6350) );
  NAND2_X1 U6499 ( .A1(n6023), .A2(n5577), .ZN(n5576) );
  NAND2_X1 U6500 ( .A1(n9238), .A2(n5583), .ZN(n5580) );
  NAND2_X1 U6501 ( .A1(n5580), .A2(n5581), .ZN(n6243) );
  NAND2_X1 U6502 ( .A1(n8491), .A2(n5595), .ZN(n7367) );
  NAND2_X1 U6503 ( .A1(n7705), .A2(n5596), .ZN(n7689) );
  NAND2_X2 U6504 ( .A1(n7456), .A2(n5977), .ZN(n7705) );
  NAND2_X1 U6505 ( .A1(n6978), .A2(n5851), .ZN(n5866) );
  OAI21_X2 U6506 ( .B1(n8260), .B2(n8261), .A(n8262), .ZN(n9295) );
  NAND2_X1 U6507 ( .A1(n5600), .A2(n5601), .ZN(n8397) );
  NAND2_X1 U6508 ( .A1(n9913), .A2(n8384), .ZN(n5600) );
  NAND2_X1 U6509 ( .A1(n7175), .A2(n7089), .ZN(n8583) );
  NAND2_X1 U6510 ( .A1(n5603), .A2(n7089), .ZN(n5604) );
  NAND2_X1 U6511 ( .A1(n5605), .A2(n5604), .ZN(n7108) );
  NAND2_X1 U6512 ( .A1(n9960), .A2(n5610), .ZN(n5609) );
  NAND2_X1 U6513 ( .A1(n5613), .A2(n5614), .ZN(n7609) );
  NAND2_X1 U6514 ( .A1(n7296), .A2(n5615), .ZN(n5613) );
  NAND2_X1 U6515 ( .A1(n5618), .A2(n5038), .ZN(n7146) );
  NAND2_X1 U6516 ( .A1(n7097), .A2(n5621), .ZN(n5620) );
  AOI21_X1 U6517 ( .B1(n5621), .B2(n5623), .A(n5064), .ZN(n5619) );
  NAND2_X1 U6518 ( .A1(n6412), .A2(n6411), .ZN(n6468) );
  OAI21_X1 U6519 ( .B1(n9885), .B2(n8410), .A(n8411), .ZN(n9881) );
  OAI21_X2 U6520 ( .B1(n9885), .B2(n5629), .A(n5628), .ZN(n8492) );
  INV_X1 U6521 ( .A(n7443), .ZN(n7441) );
  OR2_X1 U6522 ( .A1(n6681), .A2(n6553), .ZN(n6683) );
  NAND2_X1 U6523 ( .A1(n10440), .A2(n10439), .ZN(n10443) );
  CLKBUF_X1 U6524 ( .A(n6640), .Z(n9812) );
  INV_X1 U6525 ( .A(n6636), .ZN(n8795) );
  NAND2_X1 U6526 ( .A1(n6690), .A2(n9157), .ZN(n6692) );
  INV_X1 U6527 ( .A(n6697), .ZN(n6698) );
  NAND2_X1 U6528 ( .A1(n8200), .A2(n8199), .ZN(n8271) );
  NAND2_X1 U6529 ( .A1(n8443), .A2(SI_29_), .ZN(n8531) );
  NAND2_X1 U6530 ( .A1(n9332), .A2(n7255), .ZN(n8897) );
  MUX2_X1 U6531 ( .A(n10674), .B(n10148), .S(n6681), .Z(n7118) );
  XNOR2_X1 U6532 ( .A(n6250), .B(n6249), .ZN(n8385) );
  OAI21_X1 U6533 ( .B1(n9295), .B2(n9296), .A(n9297), .ZN(n9232) );
  OR2_X1 U6534 ( .A1(n6365), .A2(n10485), .ZN(n5824) );
  NAND2_X1 U6535 ( .A1(n6833), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U6536 ( .A1(n5026), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U6537 ( .A1(n5026), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6602) );
  INV_X1 U6538 ( .A(n8505), .ZN(n10061) );
  NAND2_X1 U6539 ( .A1(n7265), .A2(n7253), .ZN(n7242) );
  OR2_X1 U6540 ( .A1(n8842), .A2(n10762), .ZN(n5826) );
  INV_X1 U6541 ( .A(n10062), .ZN(n8471) );
  INV_X1 U6542 ( .A(n9875), .ZN(n9886) );
  INV_X1 U6543 ( .A(n9615), .ZN(n9184) );
  NAND2_X2 U6544 ( .A1(n7238), .A2(n9554), .ZN(n10933) );
  NAND2_X1 U6545 ( .A1(n8015), .A2(n8014), .ZN(n8166) );
  XOR2_X1 U6546 ( .A(n10394), .B(keyinput_6), .Z(n5633) );
  AND2_X1 U6547 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_162), .ZN(n5634) );
  OR2_X1 U6548 ( .A1(n9450), .A2(n9250), .ZN(n5636) );
  AND2_X1 U6549 ( .A1(n8442), .A2(n8441), .ZN(n5637) );
  AND2_X1 U6550 ( .A1(n5324), .A2(n9213), .ZN(n5638) );
  INV_X1 U6551 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5779) );
  AND2_X1 U6552 ( .A1(n6836), .A2(n6835), .ZN(n5639) );
  AND2_X1 U6553 ( .A1(n5680), .A2(n5679), .ZN(n5640) );
  AND2_X1 U6554 ( .A1(n5684), .A2(n5683), .ZN(n5641) );
  AND2_X1 U6555 ( .A1(n6293), .A2(n6292), .ZN(n9443) );
  OR2_X1 U6556 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5643) );
  AND4_X1 U6557 ( .A1(n6165), .A2(n6164), .A3(n6163), .A4(n6162), .ZN(n9273)
         );
  INV_X1 U6558 ( .A(n9273), .ZN(n9177) );
  AND3_X1 U6559 ( .A1(n6231), .A2(n6230), .A3(n6229), .ZN(n9261) );
  INV_X1 U6560 ( .A(n9992), .ZN(n8460) );
  NOR2_X1 U6561 ( .A1(n8439), .A2(n8438), .ZN(n5644) );
  OR2_X1 U6562 ( .A1(n6819), .A2(n10666), .ZN(n11120) );
  INV_X1 U6563 ( .A(n10900), .ZN(n11118) );
  NAND2_X1 U6564 ( .A1(n9172), .A2(n6472), .ZN(n6600) );
  INV_X1 U6565 ( .A(keyinput_144), .ZN(n10417) );
  XNOR2_X1 U6566 ( .A(n10417), .B(SI_16_), .ZN(n10418) );
  XNOR2_X1 U6567 ( .A(n10217), .B(keyinput_16), .ZN(n10218) );
  INV_X1 U6568 ( .A(keyinput_23), .ZN(n10229) );
  NOR2_X1 U6569 ( .A1(keyinput_162), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10441) );
  NOR2_X1 U6570 ( .A1(n5634), .A2(n10441), .ZN(n10442) );
  INV_X1 U6571 ( .A(keyinput_165), .ZN(n10448) );
  XNOR2_X1 U6572 ( .A(n10449), .B(n10448), .ZN(n10450) );
  OAI22_X1 U6573 ( .A1(n10455), .A2(n10454), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(keyinput_167), .ZN(n10456) );
  OAI22_X1 U6574 ( .A1(n6158), .A2(keyinput_169), .B1(n10459), .B2(
        P2_REG3_REG_19__SCAN_IN), .ZN(n10460) );
  INV_X1 U6575 ( .A(n10460), .ZN(n10461) );
  INV_X1 U6576 ( .A(keyinput_172), .ZN(n10466) );
  XNOR2_X1 U6577 ( .A(n10770), .B(n10466), .ZN(n10467) );
  XNOR2_X1 U6578 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n10275) );
  INV_X1 U6579 ( .A(keyinput_189), .ZN(n10496) );
  NOR2_X1 U6580 ( .A1(n10276), .A2(n10275), .ZN(n10277) );
  XNOR2_X1 U6581 ( .A(n10496), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n10497) );
  XNOR2_X1 U6582 ( .A(n5923), .B(keyinput_61), .ZN(n10286) );
  NAND2_X1 U6583 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  INV_X1 U6584 ( .A(n10292), .ZN(n10293) );
  AOI21_X1 U6585 ( .B1(n10305), .B2(n10304), .A(n10303), .ZN(n10306) );
  AND2_X1 U6586 ( .A1(n10313), .A2(keyinput_81), .ZN(n10311) );
  OAI22_X1 U6587 ( .A1(n10529), .A2(n10528), .B1(P2_DATAO_REG_10__SCAN_IN), 
        .B2(keyinput_214), .ZN(n10530) );
  INV_X1 U6588 ( .A(n10530), .ZN(n10531) );
  NAND2_X1 U6589 ( .A1(n10572), .A2(keyinput_236), .ZN(n10573) );
  NAND2_X1 U6590 ( .A1(n10334), .A2(n10333), .ZN(n10335) );
  NOR2_X1 U6591 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  INV_X1 U6592 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U6593 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_110), .ZN(n10348) );
  NOR2_X1 U6594 ( .A1(n10349), .A2(n10348), .ZN(n10350) );
  INV_X1 U6595 ( .A(n6066), .ZN(n6065) );
  INV_X1 U6596 ( .A(n6103), .ZN(n6102) );
  NAND2_X1 U6597 ( .A1(n10351), .A2(n10350), .ZN(n10359) );
  INV_X1 U6598 ( .A(n8883), .ZN(n8852) );
  AND2_X1 U6599 ( .A1(n9620), .A2(n9504), .ZN(n9183) );
  INV_X1 U6600 ( .A(n8858), .ZN(n7360) );
  INV_X1 U6601 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7302) );
  OR2_X1 U6602 ( .A1(n7646), .A2(n6475), .ZN(n7968) );
  INV_X1 U6603 ( .A(n8756), .ZN(n7534) );
  AND2_X1 U6604 ( .A1(n6281), .A2(n5757), .ZN(n8435) );
  INV_X1 U6605 ( .A(SI_19_), .ZN(n10208) );
  INV_X1 U6606 ( .A(n7365), .ZN(n5944) );
  NAND2_X1 U6607 ( .A1(n6065), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6085) );
  INV_X1 U6608 ( .A(n7687), .ZN(n6004) );
  NAND2_X1 U6609 ( .A1(n6227), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6234) );
  OR2_X1 U6610 ( .A1(n6173), .A2(n10488), .ZN(n6191) );
  OR2_X1 U6611 ( .A1(n6013), .A2(n9339), .ZN(n6047) );
  AOI21_X1 U6612 ( .B1(n8853), .B2(n8852), .A(n8854), .ZN(n9040) );
  OR2_X1 U6613 ( .A1(n9312), .A2(n6365), .ZN(n6275) );
  NAND2_X2 U6614 ( .A1(n5818), .A2(n9686), .ZN(n5922) );
  OR2_X1 U6615 ( .A1(n10146), .A2(n8826), .ZN(n8828) );
  AND2_X1 U6616 ( .A1(n6303), .A2(n9197), .ZN(n9408) );
  NAND2_X1 U6617 ( .A1(n6190), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6206) );
  OR2_X1 U6618 ( .A1(n6047), .A2(n6044), .ZN(n6066) );
  AND2_X1 U6619 ( .A1(n9045), .A2(n8891), .ZN(n6954) );
  NAND2_X1 U6620 ( .A1(n5779), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5780) );
  INV_X1 U6621 ( .A(n9157), .ZN(n6696) );
  INV_X1 U6622 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7504) );
  AND2_X1 U6623 ( .A1(n8148), .A2(n6490), .ZN(n8150) );
  INV_X1 U6624 ( .A(n8362), .ZN(n8364) );
  OR2_X1 U6625 ( .A1(n7303), .A2(n7302), .ZN(n7505) );
  INV_X1 U6626 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6411) );
  INV_X1 U6627 ( .A(n8751), .ZN(n7096) );
  INV_X1 U6628 ( .A(n7183), .ZN(n7086) );
  INV_X1 U6629 ( .A(n8046), .ZN(n11094) );
  NAND2_X1 U6630 ( .A1(n7535), .A2(n7534), .ZN(n7607) );
  NAND2_X1 U6631 ( .A1(n6468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U6632 ( .A1(n5695), .A2(n5694), .ZN(n5698) );
  NOR2_X1 U6633 ( .A1(n10598), .A2(P1_D_REG_4__SCAN_IN), .ZN(n10599) );
  NAND2_X2 U6634 ( .A1(n6743), .A2(n6680), .ZN(n8826) );
  NOR2_X1 U6635 ( .A1(n9037), .A2(n8307), .ZN(n8879) );
  AND2_X1 U6636 ( .A1(n6275), .A2(n6274), .ZN(n9250) );
  INV_X1 U6637 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U6638 ( .A1(n9184), .A2(n9261), .ZN(n9185) );
  NAND2_X1 U6639 ( .A1(n9642), .A2(n9177), .ZN(n9178) );
  NAND2_X1 U6640 ( .A1(n7715), .A2(n5078), .ZN(n7750) );
  NAND2_X1 U6641 ( .A1(n8918), .A2(n8860), .ZN(n7670) );
  INV_X1 U6642 ( .A(n10185), .ZN(n7235) );
  NAND2_X1 U6643 ( .A1(n10836), .A2(n7239), .ZN(n10832) );
  AND2_X1 U6644 ( .A1(n6315), .A2(n8880), .ZN(n11066) );
  INV_X1 U6645 ( .A(n9572), .ZN(n9548) );
  OR2_X1 U6646 ( .A1(n6506), .A2(n6505), .ZN(n8328) );
  INV_X1 U6647 ( .A(n8187), .ZN(n8047) );
  OR2_X1 U6648 ( .A1(n7505), .A2(n7504), .ZN(n7521) );
  INV_X1 U6649 ( .A(n9791), .ZN(n9756) );
  AND3_X1 U6650 ( .A1(n6510), .A2(n6509), .A3(n6508), .ZN(n10019) );
  INV_X1 U6651 ( .A(n9970), .ZN(n8346) );
  AND2_X1 U6652 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  NOR2_X1 U6653 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10640), .ZN(n7920) );
  INV_X1 U6654 ( .A(n8240), .ZN(n6332) );
  AND3_X1 U6655 ( .A1(n6260), .A2(n6259), .A3(n6258), .ZN(n9442) );
  AND4_X1 U6656 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n9074)
         );
  INV_X1 U6657 ( .A(n10788), .ZN(n10761) );
  AND2_X1 U6658 ( .A1(n6745), .A2(n6744), .ZN(n10796) );
  INV_X1 U6659 ( .A(n9182), .ZN(n9503) );
  OR2_X1 U6660 ( .A1(n7236), .A2(n7235), .ZN(n9554) );
  INV_X1 U6661 ( .A(n9550), .ZN(n9574) );
  AND2_X1 U6662 ( .A1(n6335), .A2(n10756), .ZN(n7232) );
  AND2_X1 U6663 ( .A1(n8275), .A2(n10850), .ZN(n11082) );
  INV_X1 U6664 ( .A(n11082), .ZN(n11129) );
  AND2_X1 U6665 ( .A1(n6705), .A2(n10993), .ZN(n9758) );
  AND3_X1 U6666 ( .A1(n8544), .A2(n8543), .A3(n8542), .ZN(n9856) );
  INV_X1 U6667 ( .A(n10019), .ZN(n9985) );
  INV_X1 U6668 ( .A(n10808), .ZN(n10746) );
  OR2_X1 U6669 ( .A1(n10693), .A2(n9821), .ZN(n10809) );
  INV_X1 U6670 ( .A(n10697), .ZN(n10813) );
  INV_X1 U6671 ( .A(n8769), .ZN(n9907) );
  INV_X1 U6672 ( .A(n8765), .ZN(n8683) );
  OR2_X1 U6673 ( .A1(n7153), .A2(n6877), .ZN(n11109) );
  OR2_X1 U6674 ( .A1(n7153), .A2(n8801), .ZN(n11111) );
  OR2_X1 U6675 ( .A1(n8735), .A2(n8801), .ZN(n11057) );
  OR3_X1 U6676 ( .A1(n6625), .A2(n6624), .A3(n6634), .ZN(n6819) );
  AND2_X1 U6677 ( .A1(n6627), .A2(n6626), .ZN(n10666) );
  AND2_X1 U6678 ( .A1(n7128), .A2(n7412), .ZN(n9843) );
  AND2_X1 U6679 ( .A1(n6578), .A2(n6573), .ZN(n7501) );
  NOR2_X1 U6680 ( .A1(n10641), .A2(n7920), .ZN(n7921) );
  NOR2_X1 U6681 ( .A1(n10652), .A2(n10651), .ZN(n7937) );
  INV_X1 U6682 ( .A(n10760), .ZN(n6421) );
  INV_X1 U6683 ( .A(n10611), .ZN(n9319) );
  AND4_X1 U6684 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n9547)
         );
  NAND2_X1 U6685 ( .A1(n6729), .A2(n6726), .ZN(n10788) );
  NAND2_X1 U6686 ( .A1(n10933), .A2(n10924), .ZN(n9568) );
  INV_X1 U6687 ( .A(n10933), .ZN(n9541) );
  NAND2_X1 U6688 ( .A1(n10933), .A2(n10919), .ZN(n9581) );
  INV_X1 U6689 ( .A(n11132), .ZN(n11131) );
  AND3_X1 U6690 ( .A1(n11051), .A2(n11050), .A3(n11049), .ZN(n11052) );
  AND2_X1 U6691 ( .A1(n10984), .A2(n10983), .ZN(n10985) );
  NAND2_X1 U6692 ( .A1(n10185), .A2(n10184), .ZN(n10757) );
  INV_X1 U6693 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6906) );
  OR2_X1 U6694 ( .A1(n6879), .A2(n6407), .ZN(n6515) );
  INV_X1 U6695 ( .A(n9773), .ZN(n9799) );
  OR2_X1 U6696 ( .A1(n10671), .A2(n6518), .ZN(n10702) );
  NAND2_X1 U6697 ( .A1(n11019), .A2(n7120), .ZN(n11016) );
  NAND2_X1 U6698 ( .A1(n11019), .A2(n7150), .ZN(n10025) );
  NOR2_X1 U6699 ( .A1(n6819), .A2(n6628), .ZN(n10900) );
  AND2_X1 U6700 ( .A1(n11098), .A2(n11097), .ZN(n11100) );
  CLKBUF_X1 U6701 ( .A(n10181), .Z(n10169) );
  INV_X1 U6702 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7416) );
  INV_X1 U6703 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10523) );
  INV_X1 U6704 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10535) );
  CLKBUF_X1 U6705 ( .A(n8024), .Z(n10147) );
  INV_X1 U6706 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10771) );
  NOR2_X1 U6707 ( .A1(n7938), .A2(n7937), .ZN(n10654) );
  INV_X1 U6708 ( .A(SI_2_), .ZN(n5647) );
  XNOR2_X1 U6709 ( .A(n5653), .B(n5647), .ZN(n5843) );
  AND2_X1 U6710 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6711 ( .A1(n5650), .A2(n5648), .ZN(n5829) );
  NAND2_X1 U6712 ( .A1(n5651), .A2(SI_1_), .ZN(n5652) );
  NAND2_X1 U6713 ( .A1(n5653), .A2(SI_2_), .ZN(n5654) );
  MUX2_X1 U6714 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6422), .Z(n5656) );
  XNOR2_X1 U6715 ( .A(n5656), .B(SI_3_), .ZN(n5852) );
  INV_X1 U6716 ( .A(n5852), .ZN(n5655) );
  NAND2_X1 U6717 ( .A1(n5853), .A2(n5655), .ZN(n5658) );
  NAND2_X1 U6718 ( .A1(n5656), .A2(SI_3_), .ZN(n5657) );
  MUX2_X1 U6719 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6422), .Z(n5660) );
  XNOR2_X1 U6720 ( .A(n5660), .B(SI_4_), .ZN(n5872) );
  INV_X1 U6721 ( .A(n5872), .ZN(n5659) );
  NAND2_X1 U6722 ( .A1(n5660), .A2(SI_4_), .ZN(n5898) );
  MUX2_X1 U6723 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6422), .Z(n5662) );
  NAND2_X1 U6724 ( .A1(n5662), .A2(SI_5_), .ZN(n5661) );
  AND2_X1 U6725 ( .A1(n5898), .A2(n5661), .ZN(n5665) );
  INV_X1 U6726 ( .A(n5661), .ZN(n5664) );
  XNOR2_X1 U6727 ( .A(n5662), .B(SI_5_), .ZN(n5900) );
  INV_X1 U6728 ( .A(n5900), .ZN(n5663) );
  MUX2_X1 U6729 ( .A(n6461), .B(n10543), .S(n6422), .Z(n5666) );
  XNOR2_X1 U6730 ( .A(n5666), .B(SI_6_), .ZN(n5881) );
  INV_X1 U6731 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U6732 ( .A1(n5667), .A2(SI_6_), .ZN(n5668) );
  MUX2_X1 U6733 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6422), .Z(n5670) );
  INV_X1 U6734 ( .A(SI_7_), .ZN(n5669) );
  XNOR2_X1 U6735 ( .A(n5670), .B(n5669), .ZN(n5932) );
  NAND2_X1 U6736 ( .A1(n5670), .A2(SI_7_), .ZN(n5671) );
  MUX2_X1 U6737 ( .A(n6504), .B(n10321), .S(n6422), .Z(n5672) );
  NAND2_X1 U6738 ( .A1(n5672), .A2(n10234), .ZN(n5675) );
  INV_X1 U6739 ( .A(n5672), .ZN(n5673) );
  NAND2_X1 U6740 ( .A1(n5673), .A2(SI_8_), .ZN(n5674) );
  NAND2_X1 U6741 ( .A1(n5675), .A2(n5674), .ZN(n5958) );
  MUX2_X1 U6742 ( .A(n6514), .B(n10535), .S(n6422), .Z(n5677) );
  NAND2_X1 U6743 ( .A1(n5677), .A2(n10425), .ZN(n5680) );
  INV_X1 U6744 ( .A(n5677), .ZN(n5678) );
  NAND2_X1 U6745 ( .A1(n5678), .A2(SI_9_), .ZN(n5679) );
  INV_X1 U6746 ( .A(n6422), .ZN(n6680) );
  MUX2_X1 U6747 ( .A(n6576), .B(n10528), .S(n5752), .Z(n5681) );
  INV_X1 U6748 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U6749 ( .A1(n5682), .A2(SI_10_), .ZN(n5683) );
  NAND2_X1 U6750 ( .A1(n5685), .A2(n5684), .ZN(n6007) );
  MUX2_X1 U6751 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5752), .Z(n5688) );
  NAND2_X1 U6752 ( .A1(n5688), .A2(SI_11_), .ZN(n5689) );
  MUX2_X1 U6753 ( .A(n6676), .B(n10525), .S(n5752), .Z(n5690) );
  INV_X1 U6754 ( .A(n5690), .ZN(n5691) );
  NAND2_X1 U6755 ( .A1(n5691), .A2(SI_12_), .ZN(n5692) );
  NAND2_X1 U6756 ( .A1(n5693), .A2(n5692), .ZN(n6024) );
  MUX2_X1 U6757 ( .A(n6906), .B(n10523), .S(n5752), .Z(n5695) );
  INV_X1 U6758 ( .A(n5695), .ZN(n5696) );
  NAND2_X1 U6759 ( .A1(n5696), .A2(SI_13_), .ZN(n5697) );
  NAND2_X1 U6760 ( .A1(n6040), .A2(n6039), .ZN(n5699) );
  MUX2_X1 U6761 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5752), .Z(n5700) );
  NAND2_X1 U6762 ( .A1(n5700), .A2(SI_14_), .ZN(n5701) );
  MUX2_X1 U6763 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5752), .Z(n5704) );
  XNOR2_X1 U6764 ( .A(n5704), .B(SI_15_), .ZN(n6076) );
  INV_X1 U6765 ( .A(n6076), .ZN(n5703) );
  NAND2_X1 U6766 ( .A1(n6077), .A2(n5703), .ZN(n5706) );
  NAND2_X1 U6767 ( .A1(n5704), .A2(SI_15_), .ZN(n5705) );
  MUX2_X1 U6768 ( .A(n7058), .B(n10516), .S(n5752), .Z(n5707) );
  NAND2_X1 U6769 ( .A1(n5707), .A2(n10217), .ZN(n5710) );
  INV_X1 U6770 ( .A(n5707), .ZN(n5708) );
  NAND2_X1 U6771 ( .A1(n5708), .A2(SI_16_), .ZN(n5709) );
  NAND2_X1 U6772 ( .A1(n5710), .A2(n5709), .ZN(n6096) );
  MUX2_X1 U6773 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5752), .Z(n5712) );
  INV_X1 U6774 ( .A(SI_17_), .ZN(n5711) );
  XNOR2_X1 U6775 ( .A(n5712), .B(n5711), .ZN(n6114) );
  INV_X1 U6776 ( .A(n6114), .ZN(n5714) );
  NAND2_X1 U6777 ( .A1(n5712), .A2(SI_17_), .ZN(n5713) );
  MUX2_X1 U6778 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5752), .Z(n5716) );
  XNOR2_X1 U6779 ( .A(n5716), .B(SI_18_), .ZN(n6132) );
  INV_X1 U6780 ( .A(n6132), .ZN(n5715) );
  NAND2_X1 U6781 ( .A1(n5716), .A2(SI_18_), .ZN(n5717) );
  INV_X1 U6782 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n5718) );
  MUX2_X1 U6783 ( .A(n5718), .B(n7416), .S(n5752), .Z(n5719) );
  NAND2_X1 U6784 ( .A1(n5719), .A2(n10208), .ZN(n5722) );
  INV_X1 U6785 ( .A(n5719), .ZN(n5720) );
  NAND2_X1 U6786 ( .A1(n5720), .A2(SI_19_), .ZN(n5721) );
  NAND2_X1 U6787 ( .A1(n5722), .A2(n5721), .ZN(n6150) );
  MUX2_X1 U6788 ( .A(n8305), .B(n10511), .S(n5752), .Z(n5724) );
  INV_X1 U6789 ( .A(SI_20_), .ZN(n5723) );
  NAND2_X1 U6790 ( .A1(n5724), .A2(n5723), .ZN(n5727) );
  INV_X1 U6791 ( .A(n5724), .ZN(n5725) );
  NAND2_X1 U6792 ( .A1(n5725), .A2(SI_20_), .ZN(n5726) );
  NAND2_X1 U6793 ( .A1(n6169), .A2(n6168), .ZN(n5728) );
  MUX2_X1 U6794 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5752), .Z(n5729) );
  XNOR2_X1 U6795 ( .A(n5729), .B(n10407), .ZN(n6185) );
  NAND2_X1 U6796 ( .A1(n5729), .A2(SI_21_), .ZN(n5730) );
  MUX2_X1 U6797 ( .A(n7778), .B(n7777), .S(n5752), .Z(n5732) );
  INV_X1 U6798 ( .A(SI_22_), .ZN(n5731) );
  NAND2_X1 U6799 ( .A1(n5732), .A2(n5731), .ZN(n5735) );
  INV_X1 U6800 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U6801 ( .A1(n5733), .A2(SI_22_), .ZN(n5734) );
  NAND2_X1 U6802 ( .A1(n5735), .A2(n5734), .ZN(n6202) );
  INV_X1 U6803 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5737) );
  INV_X1 U6804 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5736) );
  MUX2_X1 U6805 ( .A(n5737), .B(n5736), .S(n5752), .Z(n5739) );
  INV_X1 U6806 ( .A(SI_23_), .ZN(n5738) );
  NAND2_X1 U6807 ( .A1(n5739), .A2(n5738), .ZN(n5742) );
  INV_X1 U6808 ( .A(n5739), .ZN(n5740) );
  NAND2_X1 U6809 ( .A1(n5740), .A2(SI_23_), .ZN(n5741) );
  MUX2_X1 U6810 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n5752), .Z(n5745) );
  INV_X1 U6811 ( .A(SI_24_), .ZN(n5744) );
  XNOR2_X1 U6812 ( .A(n5745), .B(n5744), .ZN(n6222) );
  INV_X1 U6813 ( .A(n6222), .ZN(n5747) );
  NAND2_X1 U6814 ( .A1(n5745), .A2(SI_24_), .ZN(n5746) );
  OAI21_X2 U6815 ( .B1(n6223), .B2(n5747), .A(n5746), .ZN(n6250) );
  INV_X1 U6816 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8194) );
  INV_X1 U6817 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8198) );
  MUX2_X1 U6818 ( .A(n8194), .B(n8198), .S(n5752), .Z(n5748) );
  NAND2_X1 U6819 ( .A1(n5748), .A2(n10395), .ZN(n5751) );
  INV_X1 U6820 ( .A(n5748), .ZN(n5749) );
  NAND2_X1 U6821 ( .A1(n5749), .A2(SI_25_), .ZN(n5750) );
  NAND2_X1 U6822 ( .A1(n5751), .A2(n5750), .ZN(n6249) );
  INV_X1 U6823 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8238) );
  INV_X1 U6824 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5753) );
  MUX2_X1 U6825 ( .A(n8238), .B(n5753), .S(n5752), .Z(n5754) );
  INV_X1 U6826 ( .A(SI_26_), .ZN(n10394) );
  NAND2_X1 U6827 ( .A1(n5754), .A2(n10394), .ZN(n6282) );
  INV_X1 U6828 ( .A(n5754), .ZN(n5755) );
  NAND2_X1 U6829 ( .A1(n5755), .A2(SI_26_), .ZN(n5756) );
  MUX2_X1 U6830 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n5752), .Z(n5759) );
  NAND2_X1 U6831 ( .A1(n5759), .A2(SI_27_), .ZN(n5757) );
  NAND2_X1 U6832 ( .A1(n8437), .A2(n8435), .ZN(n5762) );
  INV_X1 U6833 ( .A(n5757), .ZN(n5761) );
  INV_X1 U6834 ( .A(SI_27_), .ZN(n5758) );
  XNOR2_X1 U6835 ( .A(n5759), .B(n5758), .ZN(n6284) );
  AND2_X1 U6836 ( .A1(n6282), .A2(n6284), .ZN(n5760) );
  MUX2_X1 U6837 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5752), .Z(n8440) );
  XNOR2_X1 U6838 ( .A(n8440), .B(SI_28_), .ZN(n8439) );
  NOR2_X2 U6839 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5765) );
  NOR2_X2 U6840 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5764) );
  NOR2_X1 U6841 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5772) );
  NAND4_X1 U6842 ( .A1(n5791), .A2(n5772), .A3(n5771), .A4(n5770), .ZN(n5775)
         );
  NAND4_X1 U6843 ( .A1(n5773), .A2(n5797), .A3(n5793), .A4(n6078), .ZN(n5774)
         );
  NOR2_X1 U6844 ( .A1(n5775), .A2(n5774), .ZN(n5776) );
  OAI21_X1 U6845 ( .B1(n5782), .B2(n9679), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n5781) );
  INV_X1 U6846 ( .A(n5782), .ZN(n5786) );
  NAND2_X1 U6847 ( .A1(n8420), .A2(n8848), .ZN(n5789) );
  NAND2_X1 U6848 ( .A1(n5934), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U6849 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  INV_X1 U6850 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5794) );
  AOI21_X1 U6851 ( .B1(n6116), .B2(n5795), .A(n9679), .ZN(n5796) );
  INV_X2 U6852 ( .A(n5796), .ZN(n6134) );
  NAND2_X1 U6853 ( .A1(n6134), .A2(n5797), .ZN(n5798) );
  XNOR2_X2 U6854 ( .A(n5800), .B(n5799), .ZN(n10922) );
  NAND2_X1 U6855 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  INV_X1 U6856 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5802) );
  XNOR2_X2 U6857 ( .A(n5803), .B(n5802), .ZN(n8307) );
  NAND2_X1 U6858 ( .A1(n5070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5804) );
  MUX2_X2 U6859 ( .A(n10922), .B(n8307), .S(n8891), .Z(n5806) );
  NAND2_X1 U6860 ( .A1(n5805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6319) );
  INV_X1 U6861 ( .A(n9045), .ZN(n7780) );
  XNOR2_X1 U6862 ( .A(n5808), .B(n5807), .ZN(n6684) );
  INV_X2 U6863 ( .A(n6743), .ZN(n5937) );
  NAND2_X1 U6864 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5809) );
  NAND2_X1 U6865 ( .A1(n5937), .A2(n10778), .ZN(n5810) );
  OAI211_X2 U6866 ( .C1(n8826), .C2(n6684), .A(n5811), .B(n5810), .ZN(n7253)
         );
  XNOR2_X1 U6867 ( .A(n5028), .B(n7253), .ZN(n5835) );
  INV_X1 U6868 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U6869 ( .A1(n5812), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5815) );
  INV_X1 U6870 ( .A(n5816), .ZN(n9680) );
  INV_X1 U6871 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10770) );
  INV_X1 U6872 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7250) );
  OR2_X1 U6873 ( .A1(n5922), .A2(n7250), .ZN(n5822) );
  INV_X1 U6874 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6738) );
  XNOR2_X1 U6875 ( .A(n5835), .B(n5834), .ZN(n7012) );
  INV_X1 U6876 ( .A(n7012), .ZN(n5833) );
  INV_X1 U6877 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10762) );
  INV_X1 U6878 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7373) );
  OR2_X1 U6879 ( .A1(n5922), .A2(n7373), .ZN(n5825) );
  INV_X1 U6880 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10485) );
  NAND2_X1 U6881 ( .A1(n5921), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U6882 ( .A1(n6680), .A2(SI_0_), .ZN(n5828) );
  INV_X1 U6883 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U6884 ( .A1(n5828), .A2(n5827), .ZN(n5830) );
  AND2_X1 U6885 ( .A1(n5830), .A2(n5829), .ZN(n9692) );
  MUX2_X1 U6886 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9692), .S(n6743), .Z(n7375) );
  INV_X1 U6887 ( .A(n7375), .ZN(n7239) );
  NOR2_X1 U6888 ( .A1(n7254), .A2(n7239), .ZN(n7230) );
  NAND2_X1 U6889 ( .A1(n7230), .A2(n7237), .ZN(n6914) );
  NAND2_X1 U6890 ( .A1(n7239), .A2(n6226), .ZN(n5831) );
  NAND2_X1 U6891 ( .A1(n6914), .A2(n5831), .ZN(n7011) );
  NAND2_X1 U6892 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  INV_X1 U6893 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7259) );
  OR2_X1 U6894 ( .A1(n6365), .A2(n7259), .ZN(n5841) );
  NAND2_X1 U6895 ( .A1(n5921), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5840) );
  INV_X1 U6896 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6737) );
  OR2_X1 U6897 ( .A1(n8842), .A2(n6737), .ZN(n5839) );
  INV_X1 U6898 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5837) );
  OR2_X1 U6899 ( .A1(n5922), .A2(n5837), .ZN(n5838) );
  NOR2_X1 U6900 ( .A1(n9332), .A2(n5027), .ZN(n5847) );
  XNOR2_X1 U6901 ( .A(n5842), .B(n5843), .ZN(n6824) );
  NAND2_X1 U6902 ( .A1(n5934), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U6903 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5643), .ZN(n5844) );
  XNOR2_X1 U6904 ( .A(n5844), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10793) );
  NAND2_X1 U6905 ( .A1(n5937), .A2(n10793), .ZN(n5845) );
  OAI211_X1 U6906 ( .C1(n8826), .C2(n6824), .A(n5846), .B(n5845), .ZN(n7255)
         );
  XNOR2_X1 U6907 ( .A(n10852), .B(n5028), .ZN(n5848) );
  NAND2_X1 U6908 ( .A1(n5847), .A2(n5848), .ZN(n5851) );
  INV_X1 U6909 ( .A(n5847), .ZN(n5849) );
  INV_X1 U6910 ( .A(n5848), .ZN(n7020) );
  NAND2_X1 U6911 ( .A1(n5849), .A2(n7020), .ZN(n5850) );
  AND2_X1 U6912 ( .A1(n5851), .A2(n5850), .ZN(n6979) );
  CLKBUF_X3 U6913 ( .A(n5934), .Z(n8831) );
  NAND2_X1 U6914 ( .A1(n8831), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5857) );
  XNOR2_X1 U6915 ( .A(n5852), .B(n5853), .ZN(n6435) );
  NAND2_X1 U6916 ( .A1(n8848), .A2(n6435), .ZN(n5856) );
  OAI21_X1 U6917 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(n5643), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U6918 ( .A(n5854), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U6919 ( .A1(n5937), .A2(n6735), .ZN(n5855) );
  XNOR2_X1 U6920 ( .A(n10886), .B(n6226), .ZN(n5862) );
  NAND2_X1 U6921 ( .A1(n5921), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5861) );
  OR2_X1 U6922 ( .A1(n6365), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5860) );
  INV_X1 U6923 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6736) );
  OR2_X1 U6924 ( .A1(n8842), .A2(n6736), .ZN(n5859) );
  INV_X1 U6925 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6717) );
  OR2_X1 U6926 ( .A1(n5922), .A2(n6717), .ZN(n5858) );
  NAND4_X1 U6927 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n7347)
         );
  AND2_X1 U6928 ( .A1(n7347), .A2(n7237), .ZN(n5863) );
  NAND2_X1 U6929 ( .A1(n5862), .A2(n5863), .ZN(n5877) );
  INV_X1 U6930 ( .A(n5862), .ZN(n10606) );
  INV_X1 U6931 ( .A(n5863), .ZN(n5864) );
  NAND2_X1 U6932 ( .A1(n10606), .A2(n5864), .ZN(n5865) );
  AND2_X1 U6933 ( .A1(n5877), .A2(n5865), .ZN(n7018) );
  NAND2_X1 U6934 ( .A1(n5866), .A2(n7018), .ZN(n7021) );
  NAND2_X1 U6935 ( .A1(n5921), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5871) );
  INV_X1 U6936 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6734) );
  OR2_X1 U6937 ( .A1(n8842), .A2(n6734), .ZN(n5870) );
  INV_X1 U6938 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5867) );
  OR2_X1 U6939 ( .A1(n5922), .A2(n5867), .ZN(n5869) );
  NAND2_X1 U6940 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5892) );
  OAI21_X1 U6941 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5892), .ZN(n10614) );
  OR2_X1 U6942 ( .A1(n6365), .A2(n10614), .ZN(n5868) );
  OR2_X1 U6943 ( .A1(n7381), .A2(n9039), .ZN(n5880) );
  NAND2_X1 U6944 ( .A1(n8848), .A2(n6926), .ZN(n5876) );
  NAND2_X1 U6945 ( .A1(n8831), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5875) );
  XNOR2_X1 U6946 ( .A(n5873), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U6947 ( .A1(n5937), .A2(n6733), .ZN(n5874) );
  XNOR2_X1 U6948 ( .A(n10904), .B(n6226), .ZN(n9053) );
  XNOR2_X1 U6949 ( .A(n5880), .B(n9053), .ZN(n10626) );
  AND2_X1 U6950 ( .A1(n10626), .A2(n5877), .ZN(n5878) );
  NAND2_X1 U6951 ( .A1(n7021), .A2(n5878), .ZN(n8482) );
  INV_X1 U6952 ( .A(n9053), .ZN(n5879) );
  NAND2_X1 U6953 ( .A1(n5880), .A2(n5879), .ZN(n8483) );
  NAND2_X1 U6954 ( .A1(n5934), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U6955 ( .A1(n5883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5884) );
  XNOR2_X1 U6956 ( .A(n5884), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U6957 ( .A1(n5937), .A2(n6793), .ZN(n5885) );
  XNOR2_X1 U6958 ( .A(n6226), .B(n8916), .ZN(n5919) );
  NAND2_X1 U6959 ( .A1(n5921), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5891) );
  INV_X1 U6960 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6742) );
  OR2_X1 U6961 ( .A1(n8842), .A2(n6742), .ZN(n5890) );
  INV_X1 U6962 ( .A(n5892), .ZN(n5887) );
  NAND2_X1 U6963 ( .A1(n5887), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5924) );
  INV_X1 U6964 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5923) );
  XNOR2_X1 U6965 ( .A(n5924), .B(n5923), .ZN(n8479) );
  OR2_X1 U6966 ( .A1(n6365), .A2(n8479), .ZN(n5889) );
  INV_X1 U6967 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7474) );
  AND2_X1 U6968 ( .A1(n9331), .A2(n7237), .ZN(n5917) );
  XNOR2_X1 U6969 ( .A(n5919), .B(n5917), .ZN(n8485) );
  INV_X1 U6970 ( .A(n8485), .ZN(n5908) );
  NAND2_X1 U6971 ( .A1(n5921), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5897) );
  INV_X1 U6972 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6719) );
  OR2_X1 U6973 ( .A1(n5922), .A2(n6719), .ZN(n5896) );
  INV_X1 U6974 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U6975 ( .A1(n5892), .A2(n10473), .ZN(n5893) );
  NAND2_X1 U6976 ( .A1(n5924), .A2(n5893), .ZN(n9048) );
  OR2_X1 U6977 ( .A1(n6365), .A2(n9048), .ZN(n5895) );
  INV_X1 U6978 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6732) );
  OR2_X1 U6979 ( .A1(n8842), .A2(n6732), .ZN(n5894) );
  OR2_X1 U6980 ( .A1(n8486), .A2(n9039), .ZN(n5912) );
  NAND2_X1 U6981 ( .A1(n5899), .A2(n5898), .ZN(n5901) );
  XNOR2_X1 U6982 ( .A(n5901), .B(n5900), .ZN(n7034) );
  NAND2_X1 U6983 ( .A1(n8848), .A2(n7034), .ZN(n5906) );
  NAND2_X1 U6984 ( .A1(n8831), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U6985 ( .A1(n5902), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5903) );
  XNOR2_X1 U6986 ( .A(n5903), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U6987 ( .A1(n5937), .A2(n6731), .ZN(n5904) );
  XNOR2_X1 U6988 ( .A(n7473), .B(n6226), .ZN(n5911) );
  INV_X1 U6989 ( .A(n5911), .ZN(n8487) );
  NAND2_X1 U6990 ( .A1(n5912), .A2(n8487), .ZN(n5907) );
  OR2_X1 U6991 ( .A1(n5908), .A2(n5907), .ZN(n5910) );
  AND2_X1 U6992 ( .A1(n8483), .A2(n5910), .ZN(n5909) );
  NAND2_X1 U6993 ( .A1(n8482), .A2(n5909), .ZN(n5916) );
  INV_X1 U6994 ( .A(n5910), .ZN(n5914) );
  XNOR2_X1 U6995 ( .A(n5912), .B(n5911), .ZN(n9057) );
  AND2_X1 U6996 ( .A1(n9057), .A2(n8485), .ZN(n5913) );
  OR2_X1 U6997 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  INV_X1 U6998 ( .A(n5917), .ZN(n5918) );
  NAND2_X1 U6999 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  NAND2_X1 U7000 ( .A1(n5921), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5931) );
  INV_X1 U7001 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7678) );
  OR2_X1 U7002 ( .A1(n5922), .A2(n7678), .ZN(n5930) );
  OAI21_X1 U7003 ( .B1(n5924), .B2(n5923), .A(n10445), .ZN(n5927) );
  INV_X1 U7004 ( .A(n5924), .ZN(n5926) );
  AND2_X1 U7005 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n5925) );
  NAND2_X1 U7006 ( .A1(n5926), .A2(n5925), .ZN(n5949) );
  NAND2_X1 U7007 ( .A1(n5927), .A2(n5949), .ZN(n7682) );
  OR2_X1 U7008 ( .A1(n6365), .A2(n7682), .ZN(n5929) );
  INV_X1 U7009 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6796) );
  OR2_X1 U7010 ( .A1(n8842), .A2(n6796), .ZN(n5928) );
  NOR2_X1 U7011 ( .A1(n7559), .A2(n9039), .ZN(n5940) );
  NAND2_X1 U7012 ( .A1(n5934), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5939) );
  OR2_X1 U7013 ( .A1(n5935), .A2(n9679), .ZN(n5936) );
  XNOR2_X1 U7014 ( .A(n5936), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U7015 ( .A1(n5937), .A2(n6804), .ZN(n5938) );
  XNOR2_X1 U7016 ( .A(n7683), .B(n6226), .ZN(n5941) );
  NAND2_X1 U7017 ( .A1(n5940), .A2(n5941), .ZN(n5945) );
  INV_X1 U7018 ( .A(n5940), .ZN(n5942) );
  INV_X1 U7019 ( .A(n5941), .ZN(n7455) );
  NAND2_X1 U7020 ( .A1(n5942), .A2(n7455), .ZN(n5943) );
  NAND2_X1 U7021 ( .A1(n5945), .A2(n5943), .ZN(n7365) );
  NAND2_X1 U7022 ( .A1(n7367), .A2(n5945), .ZN(n5966) );
  NAND2_X1 U7023 ( .A1(n8834), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5954) );
  INV_X1 U7024 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5946) );
  OR2_X1 U7025 ( .A1(n5947), .A2(n5946), .ZN(n5953) );
  INV_X1 U7026 ( .A(n5949), .ZN(n5948) );
  INV_X1 U7027 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U7028 ( .A1(n5949), .A2(n10258), .ZN(n5950) );
  NAND2_X1 U7029 ( .A1(n5994), .A2(n5950), .ZN(n7563) );
  OR2_X1 U7030 ( .A1(n6365), .A2(n7563), .ZN(n5952) );
  INV_X1 U7031 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6812) );
  OR2_X1 U7032 ( .A1(n8842), .A2(n6812), .ZN(n5951) );
  NOR2_X1 U7033 ( .A1(n7695), .A2(n9039), .ZN(n5962) );
  NAND2_X1 U7034 ( .A1(n5955), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5957) );
  INV_X1 U7035 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7036 ( .A(n5957), .B(n5956), .ZN(n6865) );
  NAND2_X1 U7037 ( .A1(n7290), .A2(n8848), .ZN(n5961) );
  NAND2_X1 U7038 ( .A1(n8831), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n5960) );
  OAI211_X1 U7039 ( .C1(n6743), .C2(n6865), .A(n5961), .B(n5960), .ZN(n7713)
         );
  XNOR2_X1 U7040 ( .A(n6311), .B(n7713), .ZN(n5963) );
  NAND2_X1 U7041 ( .A1(n5962), .A2(n5963), .ZN(n5976) );
  INV_X1 U7042 ( .A(n5962), .ZN(n5964) );
  INV_X1 U7043 ( .A(n5963), .ZN(n7696) );
  NAND2_X1 U7044 ( .A1(n5964), .A2(n7696), .ZN(n5965) );
  AND2_X1 U7045 ( .A1(n5976), .A2(n5965), .ZN(n7453) );
  NAND2_X1 U7046 ( .A1(n5966), .A2(n7453), .ZN(n7456) );
  NAND2_X1 U7047 ( .A1(n7495), .A2(n8848), .ZN(n5970) );
  NAND2_X1 U7048 ( .A1(n5968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5984) );
  XNOR2_X1 U7049 ( .A(n5984), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6963) );
  AOI22_X1 U7050 ( .A1(n8831), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5937), .B2(
        n6963), .ZN(n5969) );
  XNOR2_X1 U7051 ( .A(n7768), .B(n6311), .ZN(n5978) );
  NAND2_X1 U7052 ( .A1(n8834), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5975) );
  INV_X1 U7053 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5971) );
  INV_X1 U7054 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7055 ( .A(n5994), .B(n5992), .ZN(n7723) );
  OR2_X1 U7056 ( .A1(n6365), .A2(n7723), .ZN(n5973) );
  INV_X1 U7057 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6866) );
  OR2_X1 U7058 ( .A1(n8842), .A2(n6866), .ZN(n5972) );
  OR2_X1 U7059 ( .A1(n7749), .A2(n9039), .ZN(n5979) );
  XNOR2_X1 U7060 ( .A(n5978), .B(n5979), .ZN(n7710) );
  AND2_X1 U7061 ( .A1(n7710), .A2(n5976), .ZN(n5977) );
  INV_X1 U7062 ( .A(n5978), .ZN(n5980) );
  NAND2_X1 U7063 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  XNOR2_X1 U7064 ( .A(n5982), .B(n5641), .ZN(n7500) );
  NAND2_X1 U7065 ( .A1(n7500), .A2(n8848), .ZN(n5990) );
  INV_X1 U7066 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7067 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  NAND2_X1 U7068 ( .A1(n5985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5987) );
  INV_X1 U7069 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5986) );
  OR2_X1 U7070 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7071 ( .A1(n5987), .A2(n5986), .ZN(n6008) );
  AOI22_X1 U7072 ( .A1(n8831), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5937), .B2(
        n7402), .ZN(n5989) );
  NAND2_X1 U7073 ( .A1(n5990), .A2(n5989), .ZN(n7820) );
  XNOR2_X1 U7074 ( .A(n7820), .B(n6311), .ZN(n6000) );
  NAND2_X1 U7075 ( .A1(n8834), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5999) );
  INV_X1 U7076 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5991) );
  OR2_X1 U7077 ( .A1(n5947), .A2(n5991), .ZN(n5998) );
  OAI21_X1 U7078 ( .B1(n5994), .B2(n5992), .A(n10455), .ZN(n5995) );
  NAND2_X1 U7079 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n5993) );
  NAND2_X1 U7080 ( .A1(n5995), .A2(n6013), .ZN(n7766) );
  OR2_X1 U7081 ( .A1(n6365), .A2(n7766), .ZN(n5997) );
  INV_X1 U7082 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6970) );
  OR2_X1 U7083 ( .A1(n8842), .A2(n6970), .ZN(n5996) );
  NOR2_X1 U7084 ( .A1(n7788), .A2(n9039), .ZN(n6001) );
  NAND2_X1 U7085 ( .A1(n6000), .A2(n6001), .ZN(n6005) );
  INV_X1 U7086 ( .A(n6000), .ZN(n7782) );
  INV_X1 U7087 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7088 ( .A1(n7782), .A2(n6002), .ZN(n6003) );
  NAND2_X1 U7089 ( .A1(n6005), .A2(n6003), .ZN(n7687) );
  NAND2_X1 U7090 ( .A1(n7689), .A2(n6005), .ZN(n6023) );
  XNOR2_X1 U7091 ( .A(n6007), .B(n6006), .ZN(n7512) );
  NAND2_X1 U7092 ( .A1(n7512), .A2(n8848), .ZN(n6011) );
  NAND2_X1 U7093 ( .A1(n6008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6009) );
  XNOR2_X1 U7094 ( .A(n6009), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9338) );
  AOI22_X1 U7095 ( .A1(n8831), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5937), .B2(
        n9338), .ZN(n6010) );
  NAND2_X1 U7096 ( .A1(n6011), .A2(n6010), .ZN(n11045) );
  XNOR2_X1 U7097 ( .A(n11045), .B(n6311), .ZN(n6019) );
  NAND2_X1 U7098 ( .A1(n8834), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6018) );
  INV_X1 U7099 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6012) );
  OR2_X1 U7100 ( .A1(n5947), .A2(n6012), .ZN(n6017) );
  NAND2_X1 U7101 ( .A1(n6013), .A2(n9339), .ZN(n6014) );
  NAND2_X1 U7102 ( .A1(n6047), .A2(n6014), .ZN(n7786) );
  OR2_X1 U7103 ( .A1(n6365), .A2(n7786), .ZN(n6016) );
  INV_X1 U7104 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7391) );
  OR2_X1 U7105 ( .A1(n8842), .A2(n7391), .ZN(n6015) );
  NOR2_X1 U7106 ( .A1(n8073), .A2(n9039), .ZN(n6020) );
  NAND2_X1 U7107 ( .A1(n6019), .A2(n6020), .ZN(n6035) );
  INV_X1 U7108 ( .A(n6019), .ZN(n8074) );
  INV_X1 U7109 ( .A(n6020), .ZN(n6021) );
  NAND2_X1 U7110 ( .A1(n8074), .A2(n6021), .ZN(n6022) );
  AND2_X1 U7111 ( .A1(n6035), .A2(n6022), .ZN(n7781) );
  XNOR2_X1 U7112 ( .A(n6025), .B(n6024), .ZN(n7634) );
  NAND2_X1 U7113 ( .A1(n7634), .A2(n8848), .ZN(n6029) );
  OR2_X1 U7114 ( .A1(n6026), .A2(n9679), .ZN(n6027) );
  XNOR2_X1 U7115 ( .A(n6027), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7423) );
  AOI22_X1 U7116 ( .A1(n8831), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5937), .B2(
        n7423), .ZN(n6028) );
  XNOR2_X1 U7117 ( .A(n11065), .B(n6226), .ZN(n9069) );
  NAND2_X1 U7118 ( .A1(n5921), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6034) );
  INV_X1 U7119 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6030) );
  OR2_X1 U7120 ( .A1(n5922), .A2(n6030), .ZN(n6033) );
  INV_X1 U7121 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6046) );
  XNOR2_X1 U7122 ( .A(n6047), .B(n6046), .ZN(n8080) );
  OR2_X1 U7123 ( .A1(n6365), .A2(n8080), .ZN(n6032) );
  INV_X1 U7124 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7395) );
  OR2_X1 U7125 ( .A1(n8842), .A2(n7395), .ZN(n6031) );
  NOR2_X1 U7126 ( .A1(n9068), .A2(n9039), .ZN(n6037) );
  XNOR2_X1 U7127 ( .A(n9069), .B(n6037), .ZN(n8086) );
  AND2_X1 U7128 ( .A1(n8086), .A2(n6035), .ZN(n6036) );
  INV_X1 U7129 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7130 ( .A1(n7877), .A2(n8848), .ZN(n6043) );
  OR2_X1 U7131 ( .A1(n6041), .A2(n9679), .ZN(n6060) );
  XNOR2_X1 U7132 ( .A(n6060), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7599) );
  AOI22_X1 U7133 ( .A1(n8831), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5937), .B2(
        n7599), .ZN(n6042) );
  XNOR2_X1 U7134 ( .A(n9067), .B(n6226), .ZN(n8519) );
  NAND2_X1 U7135 ( .A1(n5921), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6053) );
  INV_X1 U7136 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8095) );
  OR2_X1 U7137 ( .A1(n5922), .A2(n8095), .ZN(n6052) );
  NAND2_X1 U7138 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .ZN(n6044) );
  INV_X1 U7139 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6045) );
  OAI21_X1 U7140 ( .B1(n6047), .B2(n6046), .A(n6045), .ZN(n6048) );
  NAND2_X1 U7141 ( .A1(n6066), .A2(n6048), .ZN(n9065) );
  OR2_X1 U7142 ( .A1(n6365), .A2(n9065), .ZN(n6051) );
  INV_X1 U7143 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6049) );
  OR2_X1 U7144 ( .A1(n8842), .A2(n6049), .ZN(n6050) );
  NOR2_X1 U7145 ( .A1(n8518), .A2(n9039), .ZN(n6054) );
  INV_X1 U7146 ( .A(n6054), .ZN(n6055) );
  NAND2_X1 U7147 ( .A1(n8519), .A2(n6055), .ZN(n6056) );
  NAND2_X1 U7148 ( .A1(n8516), .A2(n6056), .ZN(n6072) );
  XNOR2_X1 U7149 ( .A(n6058), .B(n6057), .ZN(n7959) );
  NAND2_X1 U7150 ( .A1(n7959), .A2(n8848), .ZN(n6063) );
  NAND2_X1 U7151 ( .A1(n6060), .A2(n6059), .ZN(n6061) );
  NAND2_X1 U7152 ( .A1(n6061), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6079) );
  XNOR2_X1 U7153 ( .A(n6079), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7848) );
  AOI22_X1 U7154 ( .A1(n8831), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5937), .B2(
        n7848), .ZN(n6062) );
  XNOR2_X1 U7155 ( .A(n11101), .B(n6226), .ZN(n9082) );
  NAND2_X1 U7156 ( .A1(n5921), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6071) );
  INV_X1 U7157 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6064) );
  OR2_X1 U7158 ( .A1(n8842), .A2(n6064), .ZN(n6070) );
  INV_X1 U7159 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10449) );
  NAND2_X1 U7160 ( .A1(n6066), .A2(n10449), .ZN(n6067) );
  NAND2_X1 U7161 ( .A1(n6085), .A2(n6067), .ZN(n8514) );
  OR2_X1 U7162 ( .A1(n6365), .A2(n8514), .ZN(n6069) );
  INV_X1 U7163 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8040) );
  OR2_X1 U7164 ( .A1(n5922), .A2(n8040), .ZN(n6068) );
  NOR2_X1 U7165 ( .A1(n9081), .A2(n9039), .ZN(n6073) );
  XNOR2_X1 U7166 ( .A(n9082), .B(n6073), .ZN(n8517) );
  NAND2_X1 U7167 ( .A1(n6072), .A2(n8517), .ZN(n8509) );
  INV_X1 U7168 ( .A(n6073), .ZN(n6074) );
  NAND2_X1 U7169 ( .A1(n9082), .A2(n6074), .ZN(n6075) );
  NAND2_X1 U7170 ( .A1(n8509), .A2(n6075), .ZN(n6092) );
  XNOR2_X1 U7171 ( .A(n6077), .B(n6076), .ZN(n8050) );
  NAND2_X1 U7172 ( .A1(n8050), .A2(n8848), .ZN(n6083) );
  NAND2_X1 U7173 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  NAND2_X1 U7174 ( .A1(n6080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6081) );
  XNOR2_X1 U7175 ( .A(n6081), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8121) );
  AOI22_X1 U7176 ( .A1(n8831), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5937), .B2(
        n8121), .ZN(n6082) );
  XNOR2_X1 U7177 ( .A(n9079), .B(n6226), .ZN(n8216) );
  NAND2_X1 U7178 ( .A1(n5921), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6091) );
  INV_X1 U7179 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8205) );
  OR2_X1 U7180 ( .A1(n5922), .A2(n8205), .ZN(n6090) );
  INV_X1 U7181 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7182 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  NAND2_X1 U7183 ( .A1(n6103), .A2(n6086), .ZN(n9077) );
  OR2_X1 U7184 ( .A1(n6365), .A2(n9077), .ZN(n6089) );
  INV_X1 U7185 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6087) );
  OR2_X1 U7186 ( .A1(n8842), .A2(n6087), .ZN(n6088) );
  NOR2_X1 U7187 ( .A1(n8511), .A2(n9039), .ZN(n6093) );
  XNOR2_X1 U7188 ( .A(n8216), .B(n6093), .ZN(n9080) );
  NAND2_X1 U7189 ( .A1(n6092), .A2(n9080), .ZN(n8214) );
  INV_X1 U7190 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7191 ( .A1(n8216), .A2(n6094), .ZN(n6095) );
  NAND2_X1 U7192 ( .A1(n8214), .A2(n6095), .ZN(n6109) );
  XNOR2_X1 U7193 ( .A(n6097), .B(n6096), .ZN(n8144) );
  NAND2_X1 U7194 ( .A1(n8144), .A2(n8848), .ZN(n6100) );
  NAND2_X1 U7195 ( .A1(n5093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6098) );
  XNOR2_X1 U7196 ( .A(n6098), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9349) );
  AOI22_X1 U7197 ( .A1(n8831), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5937), .B2(
        n9349), .ZN(n6099) );
  XNOR2_X1 U7198 ( .A(n9658), .B(n6226), .ZN(n6112) );
  NAND2_X1 U7199 ( .A1(n5921), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6108) );
  INV_X1 U7200 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6101) );
  OR2_X1 U7201 ( .A1(n5922), .A2(n6101), .ZN(n6107) );
  INV_X1 U7202 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10474) );
  NAND2_X1 U7203 ( .A1(n6103), .A2(n10474), .ZN(n6104) );
  NAND2_X1 U7204 ( .A1(n6122), .A2(n6104), .ZN(n8294) );
  OR2_X1 U7205 ( .A1(n6365), .A2(n8294), .ZN(n6106) );
  INV_X1 U7206 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9356) );
  OR2_X1 U7207 ( .A1(n8842), .A2(n9356), .ZN(n6105) );
  NOR2_X1 U7208 ( .A1(n9074), .A2(n9039), .ZN(n6110) );
  XNOR2_X1 U7209 ( .A(n6112), .B(n6110), .ZN(n8215) );
  INV_X1 U7210 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7211 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  XNOR2_X1 U7212 ( .A(n6115), .B(n6114), .ZN(n8247) );
  NAND2_X1 U7213 ( .A1(n8247), .A2(n8848), .ZN(n6119) );
  NAND2_X1 U7214 ( .A1(n5106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6117) );
  XNOR2_X1 U7215 ( .A(n6117), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9368) );
  AOI22_X1 U7216 ( .A1(n8831), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5937), .B2(
        n9368), .ZN(n6118) );
  XNOR2_X1 U7217 ( .A(n9653), .B(n6226), .ZN(n6128) );
  NAND2_X1 U7218 ( .A1(n5921), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6127) );
  INV_X1 U7219 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8284) );
  OR2_X1 U7220 ( .A1(n5922), .A2(n8284), .ZN(n6126) );
  INV_X1 U7221 ( .A(n6122), .ZN(n6120) );
  NAND2_X1 U7222 ( .A1(n6120), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6139) );
  INV_X1 U7223 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7224 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  NAND2_X1 U7225 ( .A1(n6139), .A2(n6123), .ZN(n8283) );
  OR2_X1 U7226 ( .A1(n6365), .A2(n8283), .ZN(n6125) );
  INV_X1 U7227 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9374) );
  OR2_X1 U7228 ( .A1(n8842), .A2(n9374), .ZN(n6124) );
  NAND4_X1 U7229 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n9573)
         );
  NAND2_X1 U7230 ( .A1(n9573), .A2(n7237), .ZN(n6129) );
  AND2_X1 U7231 ( .A1(n6128), .A2(n6129), .ZN(n8261) );
  INV_X1 U7232 ( .A(n6128), .ZN(n6131) );
  INV_X1 U7233 ( .A(n6129), .ZN(n6130) );
  NAND2_X1 U7234 ( .A1(n6131), .A2(n6130), .ZN(n8262) );
  XNOR2_X1 U7235 ( .A(n6133), .B(n6132), .ZN(n8314) );
  NAND2_X1 U7236 ( .A1(n8314), .A2(n8848), .ZN(n6136) );
  XNOR2_X1 U7237 ( .A(n6134), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9382) );
  AOI22_X1 U7238 ( .A1(n8831), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5937), .B2(
        n9382), .ZN(n6135) );
  XNOR2_X1 U7239 ( .A(n9645), .B(n6311), .ZN(n6146) );
  NAND2_X1 U7240 ( .A1(n5921), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6145) );
  INV_X1 U7241 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6137) );
  OR2_X1 U7242 ( .A1(n8842), .A2(n6137), .ZN(n6144) );
  INV_X1 U7243 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7244 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  NAND2_X1 U7245 ( .A1(n6159), .A2(n6140), .ZN(n9564) );
  OR2_X1 U7246 ( .A1(n6365), .A2(n9564), .ZN(n6143) );
  INV_X1 U7247 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7248 ( .A1(n5922), .A2(n6141), .ZN(n6142) );
  NOR2_X1 U7249 ( .A1(n9547), .A2(n9039), .ZN(n6147) );
  AND2_X1 U7250 ( .A1(n6146), .A2(n6147), .ZN(n9296) );
  INV_X1 U7251 ( .A(n6146), .ZN(n6149) );
  INV_X1 U7252 ( .A(n6147), .ZN(n6148) );
  NAND2_X1 U7253 ( .A1(n6149), .A2(n6148), .ZN(n9297) );
  NAND2_X1 U7254 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  NAND2_X1 U7255 ( .A1(n6153), .A2(n6152), .ZN(n8319) );
  NAND2_X1 U7256 ( .A1(n8319), .A2(n8848), .ZN(n6155) );
  INV_X1 U7257 ( .A(n10922), .ZN(n9555) );
  AOI22_X1 U7258 ( .A1(n8831), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5937), .B2(
        n9555), .ZN(n6154) );
  XNOR2_X1 U7259 ( .A(n9642), .B(n6226), .ZN(n9230) );
  NAND2_X1 U7260 ( .A1(n5921), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6165) );
  INV_X1 U7261 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6156) );
  OR2_X1 U7262 ( .A1(n5922), .A2(n6156), .ZN(n6164) );
  INV_X1 U7263 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7264 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  NAND2_X1 U7265 ( .A1(n6173), .A2(n6160), .ZN(n9553) );
  OR2_X1 U7266 ( .A1(n6365), .A2(n9553), .ZN(n6163) );
  INV_X1 U7267 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n6161) );
  OR2_X1 U7268 ( .A1(n8842), .A2(n6161), .ZN(n6162) );
  OR2_X1 U7269 ( .A1(n9273), .A2(n9039), .ZN(n9229) );
  OAI21_X1 U7270 ( .B1(n9232), .B2(n9230), .A(n9229), .ZN(n6167) );
  NAND2_X1 U7271 ( .A1(n9232), .A2(n9230), .ZN(n6166) );
  NAND2_X1 U7272 ( .A1(n6167), .A2(n6166), .ZN(n9270) );
  XNOR2_X1 U7273 ( .A(n6169), .B(n6168), .ZN(n8325) );
  NAND2_X1 U7274 ( .A1(n8325), .A2(n8848), .ZN(n6171) );
  NAND2_X1 U7275 ( .A1(n8831), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6170) );
  XNOR2_X1 U7276 ( .A(n9635), .B(n6311), .ZN(n6180) );
  NAND2_X1 U7277 ( .A1(n8834), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6179) );
  INV_X1 U7278 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6172) );
  OR2_X1 U7279 ( .A1(n5947), .A2(n6172), .ZN(n6178) );
  INV_X1 U7280 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U7281 ( .A1(n6173), .A2(n10488), .ZN(n6174) );
  NAND2_X1 U7282 ( .A1(n6191), .A2(n6174), .ZN(n9272) );
  OR2_X1 U7283 ( .A1(n6365), .A2(n9272), .ZN(n6177) );
  INV_X1 U7284 ( .A(n8842), .ZN(n6257) );
  INV_X1 U7285 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6175) );
  OR2_X1 U7286 ( .A1(n8842), .A2(n6175), .ZN(n6176) );
  NOR2_X1 U7287 ( .A1(n9549), .A2(n9039), .ZN(n6181) );
  NAND2_X1 U7288 ( .A1(n6180), .A2(n6181), .ZN(n6184) );
  INV_X1 U7289 ( .A(n6180), .ZN(n9240) );
  INV_X1 U7290 ( .A(n6181), .ZN(n6182) );
  NAND2_X1 U7291 ( .A1(n9240), .A2(n6182), .ZN(n6183) );
  NAND2_X1 U7292 ( .A1(n6184), .A2(n6183), .ZN(n9269) );
  OR2_X2 U7293 ( .A1(n9270), .A2(n9269), .ZN(n9238) );
  XNOR2_X1 U7294 ( .A(n6186), .B(n6185), .ZN(n8334) );
  NAND2_X1 U7295 ( .A1(n8334), .A2(n8848), .ZN(n6188) );
  NAND2_X1 U7296 ( .A1(n5934), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6187) );
  XNOR2_X1 U7297 ( .A(n9630), .B(n6311), .ZN(n6198) );
  NAND2_X1 U7298 ( .A1(n8834), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6197) );
  INV_X1 U7299 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6189) );
  OR2_X1 U7300 ( .A1(n5947), .A2(n6189), .ZN(n6196) );
  INV_X1 U7301 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10471) );
  NAND2_X1 U7302 ( .A1(n6191), .A2(n10471), .ZN(n6192) );
  NAND2_X1 U7303 ( .A1(n6206), .A2(n6192), .ZN(n9521) );
  OR2_X1 U7304 ( .A1(n6365), .A2(n9521), .ZN(n6195) );
  INV_X1 U7305 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6193) );
  OR2_X1 U7306 ( .A1(n8842), .A2(n6193), .ZN(n6194) );
  NAND4_X1 U7307 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n9533)
         );
  AND2_X1 U7308 ( .A1(n9533), .A2(n7237), .ZN(n6199) );
  NAND2_X1 U7309 ( .A1(n6198), .A2(n6199), .ZN(n6212) );
  INV_X1 U7310 ( .A(n6198), .ZN(n9280) );
  INV_X1 U7311 ( .A(n6199), .ZN(n6200) );
  NAND2_X1 U7312 ( .A1(n9280), .A2(n6200), .ZN(n6201) );
  AND2_X1 U7313 ( .A1(n6212), .A2(n6201), .ZN(n9239) );
  XNOR2_X1 U7314 ( .A(n6203), .B(n6202), .ZN(n8348) );
  NAND2_X1 U7315 ( .A1(n8348), .A2(n8848), .ZN(n6205) );
  NAND2_X1 U7316 ( .A1(n8831), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6204) );
  XNOR2_X1 U7317 ( .A(n9625), .B(n6311), .ZN(n6214) );
  INV_X1 U7318 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U7319 ( .A1(n6206), .A2(n10490), .ZN(n6207) );
  NAND2_X1 U7320 ( .A1(n6232), .A2(n6207), .ZN(n9283) );
  OR2_X1 U7321 ( .A1(n9283), .A2(n6365), .ZN(n6211) );
  NAND2_X1 U7322 ( .A1(n5921), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7323 ( .A1(n8834), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7324 ( .A1(n6257), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6208) );
  NAND4_X1 U7325 ( .A1(n6211), .A2(n6210), .A3(n6209), .A4(n6208), .ZN(n9519)
         );
  NAND2_X1 U7326 ( .A1(n9519), .A2(n7237), .ZN(n6215) );
  XNOR2_X1 U7327 ( .A(n6214), .B(n6215), .ZN(n9281) );
  AND2_X1 U7328 ( .A1(n9281), .A2(n6212), .ZN(n6213) );
  INV_X1 U7329 ( .A(n6214), .ZN(n6216) );
  XNOR2_X1 U7330 ( .A(n6218), .B(n6217), .ZN(n8359) );
  NAND2_X1 U7331 ( .A1(n8359), .A2(n8848), .ZN(n6220) );
  NAND2_X1 U7332 ( .A1(n5934), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6219) );
  XNOR2_X1 U7333 ( .A(n9620), .B(n6226), .ZN(n6242) );
  INV_X1 U7334 ( .A(n6242), .ZN(n6221) );
  NAND2_X1 U7335 ( .A1(n8373), .A2(n8848), .ZN(n6225) );
  NAND2_X1 U7336 ( .A1(n5934), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6224) );
  XNOR2_X1 U7337 ( .A(n9615), .B(n6226), .ZN(n6244) );
  INV_X1 U7338 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10480) );
  NAND2_X1 U7339 ( .A1(n6234), .A2(n10480), .ZN(n6228) );
  AND2_X1 U7340 ( .A1(n6255), .A2(n6228), .ZN(n9472) );
  INV_X1 U7341 ( .A(n6365), .ZN(n6304) );
  NAND2_X1 U7342 ( .A1(n9472), .A2(n6304), .ZN(n6231) );
  AOI22_X1 U7343 ( .A1(n8834), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n5921), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7344 ( .A1(n6257), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6229) );
  INV_X1 U7345 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U7346 ( .A1(n6232), .A2(n10452), .ZN(n6233) );
  NAND2_X1 U7347 ( .A1(n6234), .A2(n6233), .ZN(n9223) );
  OR2_X1 U7348 ( .A1(n9223), .A2(n6365), .ZN(n6239) );
  NAND2_X1 U7349 ( .A1(n8834), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7350 ( .A1(n5921), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6235) );
  AND2_X1 U7351 ( .A1(n6236), .A2(n6235), .ZN(n6238) );
  NAND2_X1 U7352 ( .A1(n6257), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6237) );
  OR2_X1 U7353 ( .A1(n9284), .A2(n9039), .ZN(n9219) );
  AOI21_X1 U7354 ( .B1(n6244), .B2(n9261), .A(n9219), .ZN(n6240) );
  NAND2_X1 U7355 ( .A1(n9221), .A2(n6240), .ZN(n6248) );
  INV_X1 U7356 ( .A(n6244), .ZN(n9259) );
  OR2_X1 U7357 ( .A1(n9261), .A2(n9039), .ZN(n9263) );
  INV_X1 U7358 ( .A(n9263), .ZN(n6241) );
  NAND2_X1 U7359 ( .A1(n9259), .A2(n6241), .ZN(n6247) );
  AND2_X1 U7360 ( .A1(n6244), .A2(n9263), .ZN(n6245) );
  OR2_X2 U7361 ( .A1(n9257), .A2(n6245), .ZN(n6246) );
  NAND2_X1 U7362 ( .A1(n8385), .A2(n8848), .ZN(n6252) );
  NAND2_X1 U7363 ( .A1(n5934), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6251) );
  XNOR2_X1 U7364 ( .A(n9611), .B(n6311), .ZN(n6261) );
  INV_X1 U7365 ( .A(n6255), .ZN(n6253) );
  NAND2_X1 U7366 ( .A1(n6253), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6268) );
  INV_X1 U7367 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7368 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  NAND2_X1 U7369 ( .A1(n6268), .A2(n6256), .ZN(n9252) );
  OR2_X1 U7370 ( .A1(n9252), .A2(n6365), .ZN(n6260) );
  AOI22_X1 U7371 ( .A1(n8834), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n5921), .B2(
        P2_REG0_REG_25__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7372 ( .A1(n6257), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6258) );
  NOR2_X1 U7373 ( .A1(n9442), .A2(n9039), .ZN(n6262) );
  NAND2_X1 U7374 ( .A1(n6261), .A2(n6262), .ZN(n6265) );
  INV_X1 U7375 ( .A(n6261), .ZN(n9309) );
  INV_X1 U7376 ( .A(n6262), .ZN(n6263) );
  NAND2_X1 U7377 ( .A1(n9309), .A2(n6263), .ZN(n6264) );
  XNOR2_X1 U7378 ( .A(n8437), .B(n6281), .ZN(n8398) );
  NAND2_X1 U7379 ( .A1(n8398), .A2(n8848), .ZN(n6267) );
  NAND2_X1 U7380 ( .A1(n5934), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6266) );
  XNOR2_X1 U7381 ( .A(n9607), .B(n6311), .ZN(n6276) );
  INV_X1 U7382 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10284) );
  NAND2_X1 U7383 ( .A1(n6268), .A2(n10284), .ZN(n6269) );
  NAND2_X1 U7384 ( .A1(n6302), .A2(n6269), .ZN(n9312) );
  INV_X1 U7385 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7386 ( .A1(n8834), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7387 ( .A1(n5921), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6270) );
  OAI211_X1 U7388 ( .C1(n6272), .C2(n8842), .A(n6271), .B(n6270), .ZN(n6273)
         );
  INV_X1 U7389 ( .A(n6273), .ZN(n6274) );
  NOR2_X1 U7390 ( .A1(n9250), .A2(n9039), .ZN(n6277) );
  NAND2_X1 U7391 ( .A1(n6276), .A2(n6277), .ZN(n6280) );
  INV_X1 U7392 ( .A(n6276), .ZN(n9208) );
  INV_X1 U7393 ( .A(n6277), .ZN(n6278) );
  NAND2_X1 U7394 ( .A1(n9208), .A2(n6278), .ZN(n6279) );
  NAND2_X1 U7395 ( .A1(n9205), .A2(n6280), .ZN(n6299) );
  NAND2_X1 U7396 ( .A1(n8437), .A2(n6281), .ZN(n6283) );
  NAND2_X1 U7397 ( .A1(n6283), .A2(n6282), .ZN(n6285) );
  NAND2_X1 U7398 ( .A1(n8412), .A2(n8848), .ZN(n6287) );
  NAND2_X1 U7399 ( .A1(n5934), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6286) );
  XNOR2_X1 U7400 ( .A(n9600), .B(n6311), .ZN(n6294) );
  XNOR2_X1 U7401 ( .A(n6302), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U7402 ( .A1(n9423), .A2(n6304), .ZN(n6293) );
  INV_X1 U7403 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7404 ( .A1(n8834), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7405 ( .A1(n5921), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6288) );
  OAI211_X1 U7406 ( .C1(n6290), .C2(n8842), .A(n6289), .B(n6288), .ZN(n6291)
         );
  INV_X1 U7407 ( .A(n6291), .ZN(n6292) );
  NOR2_X1 U7408 ( .A1(n9443), .A2(n9039), .ZN(n6295) );
  NAND2_X1 U7409 ( .A1(n6294), .A2(n6295), .ZN(n6300) );
  INV_X1 U7410 ( .A(n6294), .ZN(n6297) );
  INV_X1 U7411 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U7412 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  NAND2_X1 U7413 ( .A1(n6299), .A2(n9206), .ZN(n9209) );
  NAND2_X1 U7414 ( .A1(n9209), .A2(n6300), .ZN(n6314) );
  INV_X1 U7415 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9212) );
  INV_X1 U7416 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6366) );
  OAI21_X1 U7417 ( .B1(n6302), .B2(n9212), .A(n6366), .ZN(n6303) );
  NAND2_X1 U7418 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6301) );
  NAND2_X1 U7419 ( .A1(n9408), .A2(n6304), .ZN(n6310) );
  INV_X1 U7420 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U7421 ( .A1(n8834), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7422 ( .A1(n5921), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6305) );
  OAI211_X1 U7423 ( .C1(n6307), .C2(n8842), .A(n6306), .B(n6305), .ZN(n6308)
         );
  INV_X1 U7424 ( .A(n6308), .ZN(n6309) );
  NAND2_X1 U7425 ( .A1(n9430), .A2(n7237), .ZN(n6312) );
  MUX2_X1 U7426 ( .A(n6312), .B(n9430), .S(n6311), .Z(n6313) );
  INV_X1 U7427 ( .A(n6350), .ZN(n6349) );
  NAND2_X1 U7428 ( .A1(n5100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6316) );
  MUX2_X1 U7429 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6316), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6317) );
  INV_X1 U7430 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U7431 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  NAND2_X1 U7432 ( .A1(n6328), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U7433 ( .A1(n6322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6323) );
  MUX2_X1 U7434 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6323), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6324) );
  AND2_X1 U7435 ( .A1(n6324), .A2(n5100), .ZN(n6333) );
  NAND3_X1 U7436 ( .A1(n6332), .A2(n6329), .A3(n6333), .ZN(n6721) );
  OR2_X1 U7437 ( .A1(n6326), .A2(n6325), .ZN(n6327) );
  NAND2_X1 U7438 ( .A1(n6328), .A2(n6327), .ZN(n6486) );
  INV_X1 U7439 ( .A(n6954), .ZN(n6356) );
  NAND2_X1 U7440 ( .A1(n10185), .A2(n6356), .ZN(n6724) );
  NOR2_X1 U7441 ( .A1(n11066), .A2(n6724), .ZN(n6348) );
  INV_X1 U7442 ( .A(P2_B_REG_SCAN_IN), .ZN(n10500) );
  AOI22_X1 U7443 ( .A1(P2_B_REG_SCAN_IN), .A2(n8089), .B1(n6329), .B2(n10500), 
        .ZN(n6330) );
  OR2_X1 U7444 ( .A1(n6333), .A2(n6330), .ZN(n6331) );
  INV_X1 U7445 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U7446 ( .A1(n10183), .A2(n10186), .ZN(n6334) );
  INV_X1 U7447 ( .A(n6333), .ZN(n8195) );
  NAND2_X1 U7448 ( .A1(n8195), .A2(n8240), .ZN(n10182) );
  NAND2_X1 U7449 ( .A1(n6334), .A2(n10182), .ZN(n7231) );
  INV_X1 U7450 ( .A(n7231), .ZN(n6336) );
  INV_X1 U7451 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10758) );
  NAND2_X1 U7452 ( .A1(n10183), .A2(n10758), .ZN(n6335) );
  NAND2_X1 U7453 ( .A1(n8089), .A2(n8240), .ZN(n10756) );
  AND2_X1 U7454 ( .A1(n6336), .A2(n7232), .ZN(n6347) );
  NOR4_X1 U7455 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6340) );
  NOR4_X1 U7456 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6339) );
  NOR4_X1 U7457 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6338) );
  NOR4_X1 U7458 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6337) );
  NAND4_X1 U7459 ( .A1(n6340), .A2(n6339), .A3(n6338), .A4(n6337), .ZN(n6346)
         );
  NOR2_X1 U7460 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6344) );
  NOR4_X1 U7461 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6343) );
  NOR4_X1 U7462 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6342) );
  NOR4_X1 U7463 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6341) );
  NAND4_X1 U7464 ( .A1(n6344), .A2(n6343), .A3(n6342), .A4(n6341), .ZN(n6345)
         );
  OAI21_X1 U7465 ( .B1(n6346), .B2(n6345), .A(n10183), .ZN(n6948) );
  NAND2_X1 U7466 ( .A1(n6347), .A2(n6948), .ZN(n6352) );
  INV_X1 U7467 ( .A(n6352), .ZN(n6354) );
  NAND2_X1 U7468 ( .A1(n6349), .A2(n10623), .ZN(n6373) );
  INV_X1 U7469 ( .A(n8307), .ZN(n8877) );
  NAND2_X1 U7470 ( .A1(n8307), .A2(n8880), .ZN(n11125) );
  INV_X1 U7471 ( .A(n6721), .ZN(n6351) );
  AOI21_X1 U7472 ( .B1(n7236), .B2(n6352), .A(n6351), .ZN(n6357) );
  AND2_X1 U7473 ( .A1(n11066), .A2(n10760), .ZN(n6353) );
  NOR2_X1 U7474 ( .A1(n6315), .A2(n7235), .ZN(n9043) );
  NOR2_X2 U7475 ( .A1(n6355), .A2(n6356), .ZN(n9572) );
  NAND2_X1 U7476 ( .A1(n9251), .A2(n9572), .ZN(n9313) );
  NOR2_X1 U7477 ( .A1(n9443), .A2(n9313), .ZN(n6370) );
  INV_X1 U7478 ( .A(n6357), .ZN(n6359) );
  NAND2_X1 U7479 ( .A1(n6315), .A2(n6954), .ZN(n6949) );
  NAND2_X1 U7480 ( .A1(n6949), .A2(n6486), .ZN(n6358) );
  INV_X1 U7481 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U7482 ( .A1(n8834), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U7483 ( .A1(n5921), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6360) );
  OAI211_X1 U7484 ( .C1(n6362), .C2(n8842), .A(n6361), .B(n6360), .ZN(n6363)
         );
  INV_X1 U7485 ( .A(n6363), .ZN(n6364) );
  OAI21_X1 U7486 ( .B1(n9197), .B2(n6365), .A(n6364), .ZN(n9412) );
  INV_X1 U7487 ( .A(n9412), .ZN(n8829) );
  NAND2_X1 U7488 ( .A1(n6355), .A2(n6954), .ZN(n9550) );
  NAND2_X1 U7489 ( .A1(n9251), .A2(n9574), .ZN(n9314) );
  OAI22_X1 U7490 ( .A1(n8829), .A2(n9314), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6366), .ZN(n6367) );
  AOI21_X1 U7491 ( .B1(n9408), .B2(n10616), .A(n6367), .ZN(n6368) );
  INV_X1 U7492 ( .A(n6368), .ZN(n6369) );
  NOR2_X1 U7493 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  OAI211_X1 U7494 ( .C1(n9595), .C2(n6373), .A(n6372), .B(n6371), .ZN(P2_U3222) );
  NAND4_X1 U7495 ( .A1(n6497), .A2(n6375), .A3(n6374), .A4(n10552), .ZN(n6377)
         );
  INV_X2 U7496 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6874) );
  INV_X2 U7497 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6457) );
  NAND4_X1 U7498 ( .A1(n6874), .A2(n10190), .A3(n6457), .A4(n6570), .ZN(n6376)
         );
  NOR2_X1 U7499 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6395) );
  NAND4_X1 U7500 ( .A1(n10353), .A2(n6382), .A3(n10565), .A4(n10572), .ZN(
        n6383) );
  NAND2_X1 U7501 ( .A1(n6409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7502 ( .A1(n6386), .A2(n6385), .ZN(n6391) );
  OR2_X1 U7503 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  NAND2_X1 U7504 ( .A1(n6391), .A2(n6387), .ZN(n8196) );
  INV_X1 U7505 ( .A(n6388), .ZN(n6398) );
  NAND2_X1 U7506 ( .A1(n6398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6390) );
  NOR2_X1 U7507 ( .A1(n8196), .A2(n8023), .ZN(n6393) );
  NAND2_X1 U7508 ( .A1(n6391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6392) );
  NAND3_X1 U7509 ( .A1(n6395), .A2(n10353), .A3(n10568), .ZN(n6396) );
  OAI21_X1 U7510 ( .B1(n6400), .B2(n6396), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6397) );
  MUX2_X1 U7511 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6397), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6399) );
  NAND2_X1 U7512 ( .A1(n6399), .A2(n6398), .ZN(n7859) );
  INV_X1 U7513 ( .A(n7859), .ZN(n6407) );
  NOR2_X2 U7514 ( .A1(n6515), .A2(P1_U3084), .ZN(P1_U4006) );
  INV_X1 U7515 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U7516 ( .A1(n6401), .A2(n10568), .ZN(n6402) );
  INV_X1 U7517 ( .A(n6595), .ZN(n8525) );
  OR2_X1 U7518 ( .A1(n6647), .A2(n6407), .ZN(n6408) );
  NAND2_X1 U7519 ( .A1(n6408), .A2(n6515), .ZN(n10671) );
  NAND2_X1 U7520 ( .A1(n6415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U7521 ( .A1(n6416), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6417) );
  MUX2_X1 U7522 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6417), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n6418) );
  OR2_X1 U7523 ( .A1(n10671), .A2(n8320), .ZN(n6420) );
  NAND2_X1 U7524 ( .A1(n6420), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X2 U7525 ( .A1(n6721), .A2(n6421), .ZN(P2_U3966) );
  INV_X1 U7526 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AND2_X1 U7527 ( .A1(n6422), .A2(n9691), .ZN(n9682) );
  AOI22_X1 U7528 ( .A1(n9682), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n10793), .ZN(n6423) );
  OAI21_X1 U7529 ( .B1(n6824), .B2(n9684), .A(n6423), .ZN(P2_U3356) );
  AND2_X1 U7530 ( .A1(n7859), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6424) );
  INV_X1 U7531 ( .A(n10669), .ZN(n10151) );
  NAND3_X1 U7532 ( .A1(n8196), .A2(P1_B_REG_SCAN_IN), .A3(n8023), .ZN(n6428)
         );
  INV_X1 U7533 ( .A(n8023), .ZN(n6426) );
  INV_X1 U7534 ( .A(P1_B_REG_SCAN_IN), .ZN(n6425) );
  NAND2_X1 U7535 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  INV_X1 U7536 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U7537 ( .A1(n10150), .A2(n6430), .ZN(n6433) );
  INV_X1 U7538 ( .A(n6431), .ZN(n8222) );
  NAND2_X1 U7539 ( .A1(n8222), .A2(n8196), .ZN(n6432) );
  NAND2_X1 U7540 ( .A1(n6433), .A2(n6432), .ZN(n6631) );
  NAND2_X1 U7541 ( .A1(n10151), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6434) );
  OAI21_X1 U7542 ( .B1(n10151), .B2(n6631), .A(n6434), .ZN(P1_U3441) );
  INV_X2 U7543 ( .A(n9682), .ZN(n9687) );
  INV_X1 U7544 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6436) );
  INV_X1 U7545 ( .A(n6435), .ZN(n6886) );
  INV_X1 U7546 ( .A(n6735), .ZN(n6762) );
  INV_X1 U7547 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n9691) );
  OAI222_X1 U7548 ( .A1(n9687), .A2(n6436), .B1(n9684), .B2(n6886), .C1(n6762), 
        .C2(n9691), .ZN(P2_U3355) );
  INV_X1 U7549 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6437) );
  INV_X1 U7550 ( .A(n10778), .ZN(n6739) );
  OAI222_X1 U7551 ( .A1(n9687), .A2(n6437), .B1(n9684), .B2(n6684), .C1(n6739), 
        .C2(n9691), .ZN(P2_U3357) );
  NAND2_X1 U7552 ( .A1(n5752), .A2(P1_U3084), .ZN(n8024) );
  NOR2_X1 U7553 ( .A1(n5752), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10141) );
  OAI21_X1 U7554 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(P1_IR_REG_0__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6443) );
  INV_X1 U7555 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U7556 ( .A1(n6443), .A2(n10540), .ZN(n6438) );
  NAND2_X1 U7557 ( .A1(n6438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6439) );
  XNOR2_X1 U7558 ( .A(n6439), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U7559 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n10141), .B1(n10743), 
        .B2(P1_STATE_REG_SCAN_IN), .ZN(n6440) );
  OAI21_X1 U7560 ( .B1(n6886), .B2(n10147), .A(n6440), .ZN(P1_U3350) );
  INV_X1 U7561 ( .A(n10141), .ZN(n10144) );
  INV_X1 U7562 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U7563 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6441) );
  INV_X1 U7564 ( .A(n6682), .ZN(n6553) );
  OAI222_X1 U7565 ( .A1(n10144), .A2(n6442), .B1(n10147), .B2(n6684), .C1(
        P1_U3084), .C2(n6553), .ZN(P1_U3352) );
  INV_X1 U7566 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6444) );
  XNOR2_X1 U7567 ( .A(n6443), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10802) );
  INV_X1 U7568 ( .A(n10802), .ZN(n10810) );
  OAI222_X1 U7569 ( .A1(n10144), .A2(n6444), .B1(n10147), .B2(n6824), .C1(
        P1_U3084), .C2(n10810), .ZN(P1_U3351) );
  NOR2_X1 U7570 ( .A1(n6445), .A2(n10139), .ZN(n6446) );
  MUX2_X1 U7571 ( .A(n10139), .B(n6446), .S(P1_IR_REG_4__SCAN_IN), .Z(n6448)
         );
  NOR2_X1 U7572 ( .A1(n6448), .A2(n6447), .ZN(n9833) );
  INV_X1 U7573 ( .A(n9833), .ZN(n6558) );
  INV_X1 U7574 ( .A(n6926), .ZN(n6450) );
  INV_X1 U7575 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6658) );
  OAI222_X1 U7576 ( .A1(n6558), .A2(P1_U3084), .B1(n10147), .B2(n6450), .C1(
        n10144), .C2(n6658), .ZN(P1_U3349) );
  INV_X1 U7577 ( .A(n6733), .ZN(n6774) );
  INV_X1 U7578 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6449) );
  OAI222_X1 U7579 ( .A1(n6774), .A2(n9691), .B1(n9684), .B2(n6450), .C1(n6449), 
        .C2(n9687), .ZN(P2_U3354) );
  INV_X1 U7580 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6451) );
  INV_X1 U7581 ( .A(n7034), .ZN(n6453) );
  INV_X1 U7582 ( .A(n6731), .ZN(n6785) );
  OAI222_X1 U7583 ( .A1(n9687), .A2(n6451), .B1(n9684), .B2(n6453), .C1(n6785), 
        .C2(n9691), .ZN(P2_U3353) );
  INV_X1 U7584 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6454) );
  OR2_X1 U7585 ( .A1(n6447), .A2(n10139), .ZN(n6452) );
  XNOR2_X1 U7586 ( .A(n6452), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10731) );
  INV_X1 U7587 ( .A(n10731), .ZN(n6559) );
  OAI222_X1 U7588 ( .A1(n10144), .A2(n6454), .B1(n10147), .B2(n6453), .C1(
        P1_U3084), .C2(n6559), .ZN(P1_U3348) );
  INV_X1 U7589 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U7590 ( .A1(n6447), .A2(n6455), .ZN(n6456) );
  NAND2_X1 U7591 ( .A1(n6456), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U7592 ( .A1(n6458), .A2(n6457), .ZN(n6462) );
  OR2_X1 U7593 ( .A1(n6458), .A2(n6457), .ZN(n6459) );
  INV_X1 U7594 ( .A(n10682), .ZN(n6460) );
  INV_X1 U7595 ( .A(n6793), .ZN(n6750) );
  INV_X1 U7596 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U7597 ( .A1(n6462), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6463) );
  XNOR2_X1 U7598 ( .A(n6463), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7201) );
  INV_X1 U7599 ( .A(n7201), .ZN(n6562) );
  OAI222_X1 U7600 ( .A1(n10144), .A2(n6464), .B1(n10147), .B2(n7200), .C1(
        P1_U3084), .C2(n6562), .ZN(P1_U3346) );
  INV_X1 U7601 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6465) );
  INV_X1 U7602 ( .A(n6804), .ZN(n6811) );
  OAI222_X1 U7603 ( .A1(n9687), .A2(n6465), .B1(n9684), .B2(n7200), .C1(n6811), 
        .C2(n9691), .ZN(P2_U3351) );
  INV_X1 U7604 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6912) );
  XNOR2_X2 U7605 ( .A(n6467), .B(n6466), .ZN(n9172) );
  BUF_X4 U7606 ( .A(n6833), .Z(n8401) );
  NAND2_X1 U7607 ( .A1(n8401), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U7608 ( .A1(n8541), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U7609 ( .A1(n7045), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U7610 ( .A1(n7217), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7303) );
  NAND2_X1 U7611 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n6474) );
  NAND2_X1 U7612 ( .A1(n7645), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7646) );
  INV_X1 U7613 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7614 ( .A1(n7646), .A2(n6475), .ZN(n6476) );
  AND2_X1 U7615 ( .A1(n7968), .A2(n6476), .ZN(n8017) );
  NAND2_X1 U7616 ( .A1(n5026), .A2(n8017), .ZN(n6478) );
  NAND2_X1 U7617 ( .A1(n6834), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6477) );
  NAND4_X1 U7618 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n8187)
         );
  NAND2_X1 U7619 ( .A1(n8187), .A2(P1_U4006), .ZN(n6481) );
  OAI21_X1 U7620 ( .B1(n6912), .B2(P1_U4006), .A(n6481), .ZN(P1_U3569) );
  INV_X1 U7621 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U7622 ( .A1(n8541), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U7623 ( .A1(n8401), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U7624 ( .A1(n6834), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6482) );
  AND3_X1 U7625 ( .A1(n6484), .A2(n6483), .A3(n6482), .ZN(n8614) );
  INV_X1 U7626 ( .A(n8614), .ZN(n8464) );
  NAND2_X1 U7627 ( .A1(n8464), .A2(P1_U4006), .ZN(n6485) );
  OAI21_X1 U7628 ( .B1(n9203), .B2(P1_U4006), .A(n6485), .ZN(P1_U3585) );
  OR2_X1 U7629 ( .A1(n6486), .A2(n9691), .ZN(n9047) );
  NAND2_X1 U7630 ( .A1(n7235), .A2(n9047), .ZN(n6489) );
  NAND2_X1 U7631 ( .A1(n10185), .A2(n6954), .ZN(n6487) );
  NAND2_X1 U7632 ( .A1(n6487), .A2(n6743), .ZN(n6488) );
  NOR2_X1 U7633 ( .A1(n10787), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7634 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7410) );
  INV_X1 U7635 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7967) );
  AND2_X1 U7636 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n6490) );
  OR2_X1 U7637 ( .A1(n8150), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6491) );
  AND2_X1 U7638 ( .A1(n6506), .A2(n6491), .ZN(n10009) );
  NAND2_X1 U7639 ( .A1(n10009), .A2(n5026), .ZN(n6495) );
  NAND2_X1 U7640 ( .A1(n8401), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U7641 ( .A1(n8541), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U7642 ( .A1(n6834), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6492) );
  NAND4_X1 U7643 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n10000)
         );
  NAND2_X1 U7644 ( .A1(n10000), .A2(P1_U4006), .ZN(n6496) );
  OAI21_X1 U7645 ( .B1(n7410), .B2(P1_U4006), .A(n6496), .ZN(P1_U3573) );
  INV_X1 U7646 ( .A(n7290), .ZN(n6503) );
  AND2_X1 U7647 ( .A1(n6497), .A2(n6457), .ZN(n6498) );
  NAND2_X1 U7648 ( .A1(n6447), .A2(n6498), .ZN(n6499) );
  INV_X1 U7649 ( .A(n6571), .ZN(n6502) );
  NAND2_X1 U7650 ( .A1(n6499), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6500) );
  MUX2_X1 U7651 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6500), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6501) );
  INV_X1 U7652 ( .A(n7292), .ZN(n6667) );
  OAI222_X1 U7653 ( .A1(n10144), .A2(n10321), .B1(n10147), .B2(n6503), .C1(
        P1_U3084), .C2(n6667), .ZN(P1_U3345) );
  OAI222_X1 U7654 ( .A1(n9687), .A2(n6504), .B1(n9684), .B2(n6503), .C1(n6865), 
        .C2(n9691), .ZN(P2_U3350) );
  INV_X1 U7655 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U7656 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  AND2_X1 U7657 ( .A1(n8328), .A2(n6507), .ZN(n9996) );
  NAND2_X1 U7658 ( .A1(n9996), .A2(n5026), .ZN(n6510) );
  AOI22_X1 U7659 ( .A1(n8401), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n6834), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U7660 ( .A1(n8541), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U7661 ( .A1(n9985), .A2(P1_U4006), .ZN(n6511) );
  OAI21_X1 U7662 ( .B1(n5718), .B2(P1_U4006), .A(n6511), .ZN(P1_U3574) );
  INV_X1 U7663 ( .A(n7495), .ZN(n6513) );
  OR2_X1 U7664 ( .A1(n6571), .A2(n10139), .ZN(n6512) );
  XNOR2_X1 U7665 ( .A(n6512), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7496) );
  INV_X1 U7666 ( .A(n7496), .ZN(n6849) );
  OAI222_X1 U7667 ( .A1(n10147), .A2(n6513), .B1(n6849), .B2(P1_U3084), .C1(
        n10535), .C2(n10144), .ZN(P1_U3344) );
  INV_X1 U7668 ( .A(n6963), .ZN(n6969) );
  OAI222_X1 U7669 ( .A1(n9687), .A2(n6514), .B1(n9684), .B2(n6513), .C1(n9691), 
        .C2(n6969), .ZN(P2_U3349) );
  INV_X1 U7670 ( .A(n6515), .ZN(n6516) );
  OR2_X1 U7671 ( .A1(P1_U3083), .A2(n6516), .ZN(n10697) );
  INV_X1 U7672 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6528) );
  NOR2_X1 U7673 ( .A1(n10675), .A2(P1_U3084), .ZN(n8236) );
  INV_X1 U7674 ( .A(n8236), .ZN(n6517) );
  OR2_X1 U7675 ( .A1(n10671), .A2(n6517), .ZN(n10693) );
  INV_X1 U7676 ( .A(n9816), .ZN(n9821) );
  INV_X1 U7677 ( .A(n10809), .ZN(n10744) );
  INV_X1 U7678 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7194) );
  INV_X1 U7679 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10674) );
  INV_X1 U7680 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10673) );
  NOR2_X1 U7681 ( .A1(n10674), .A2(n10673), .ZN(n6521) );
  INV_X1 U7682 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6554) );
  MUX2_X1 U7683 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6554), .S(n6682), .Z(n6520)
         );
  NOR2_X1 U7684 ( .A1(n9816), .A2(P1_U3084), .ZN(n8241) );
  NAND2_X1 U7685 ( .A1(n8241), .A2(n10675), .ZN(n6518) );
  INV_X1 U7686 ( .A(n10702), .ZN(n10815) );
  MUX2_X1 U7687 ( .A(n6554), .B(P1_REG1_REG_1__SCAN_IN), .S(n6682), .Z(n6519)
         );
  OR3_X1 U7688 ( .A1(n6519), .A2(n10673), .A3(n10674), .ZN(n6552) );
  OAI211_X1 U7689 ( .C1(n6521), .C2(n6520), .A(n10815), .B(n6552), .ZN(n6522)
         );
  OAI21_X1 U7690 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7194), .A(n6522), .ZN(n6523) );
  AOI21_X1 U7691 ( .B1(n6682), .B2(n10744), .A(n6523), .ZN(n6527) );
  INV_X1 U7692 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6524) );
  AND2_X1 U7693 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9813) );
  OR2_X1 U7694 ( .A1(n10693), .A2(n9816), .ZN(n10808) );
  OAI211_X1 U7695 ( .C1(n6525), .C2(n9813), .A(n10746), .B(n6535), .ZN(n6526)
         );
  OAI211_X1 U7696 ( .C1(n10697), .C2(n6528), .A(n6527), .B(n6526), .ZN(
        P1_U3242) );
  NOR2_X1 U7697 ( .A1(n7201), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U7698 ( .A1(n10682), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6542) );
  INV_X1 U7699 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6529) );
  MUX2_X1 U7700 ( .A(n6529), .B(P1_REG2_REG_6__SCAN_IN), .S(n10682), .Z(n6530)
         );
  INV_X1 U7701 ( .A(n6530), .ZN(n10684) );
  INV_X1 U7702 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6541) );
  INV_X1 U7703 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U7704 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n10743), .ZN(n6538) );
  INV_X1 U7705 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6531) );
  MUX2_X1 U7706 ( .A(n6531), .B(P1_REG2_REG_3__SCAN_IN), .S(n10743), .Z(n6532)
         );
  INV_X1 U7707 ( .A(n6532), .ZN(n10747) );
  INV_X1 U7708 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6533) );
  MUX2_X1 U7709 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6533), .S(n10802), .Z(n6536)
         );
  NAND2_X1 U7710 ( .A1(n6682), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U7711 ( .A1(n6536), .A2(n5122), .ZN(n10805) );
  NAND2_X1 U7712 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n10802), .ZN(n6537) );
  NAND2_X1 U7713 ( .A1(n10805), .A2(n6537), .ZN(n10748) );
  NAND2_X1 U7714 ( .A1(n10747), .A2(n10748), .ZN(n10745) );
  MUX2_X1 U7715 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6540), .S(n9833), .Z(n9825)
         );
  AOI21_X1 U7716 ( .B1(n6540), .B2(n6558), .A(n6539), .ZN(n10734) );
  MUX2_X1 U7717 ( .A(n6541), .B(P1_REG2_REG_5__SCAN_IN), .S(n10731), .Z(n10733) );
  INV_X1 U7718 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7336) );
  MUX2_X1 U7719 ( .A(n7336), .B(P1_REG2_REG_7__SCAN_IN), .S(n7201), .Z(n6585)
         );
  NOR2_X1 U7720 ( .A1(n6586), .A2(n6585), .ZN(n6584) );
  NOR2_X1 U7721 ( .A1(n6543), .A2(n6584), .ZN(n6547) );
  INV_X1 U7722 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6544) );
  MUX2_X1 U7723 ( .A(n6544), .B(P1_REG2_REG_8__SCAN_IN), .S(n7292), .Z(n6546)
         );
  INV_X1 U7724 ( .A(n6661), .ZN(n6545) );
  AOI21_X1 U7725 ( .B1(n6547), .B2(n6546), .A(n6545), .ZN(n6569) );
  INV_X1 U7726 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6548) );
  NOR2_X1 U7727 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6548), .ZN(n7446) );
  NOR2_X1 U7728 ( .A1(n10809), .A2(n6667), .ZN(n6549) );
  AOI211_X1 U7729 ( .C1(n10813), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n7446), .B(
        n6549), .ZN(n6568) );
  INV_X1 U7730 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10974) );
  MUX2_X1 U7731 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10974), .S(n7292), .Z(n6565)
         );
  NOR2_X1 U7732 ( .A1(n7201), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7733 ( .A1(n10682), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6561) );
  INV_X1 U7734 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6550) );
  MUX2_X1 U7735 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6550), .S(n10682), .Z(n10687) );
  INV_X1 U7736 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6560) );
  INV_X1 U7737 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U7738 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n10743), .ZN(n6557) );
  INV_X1 U7739 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6551) );
  MUX2_X1 U7740 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6551), .S(n10743), .Z(n10750) );
  NAND2_X1 U7741 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(n10802), .ZN(n6556) );
  OAI21_X1 U7742 ( .B1(n6554), .B2(n6553), .A(n6552), .ZN(n10817) );
  INV_X1 U7743 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6555) );
  MUX2_X1 U7744 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6555), .S(n10802), .Z(n10816) );
  NAND2_X1 U7745 ( .A1(n10817), .A2(n10816), .ZN(n10814) );
  NAND2_X1 U7746 ( .A1(n6556), .A2(n10814), .ZN(n10751) );
  NAND2_X1 U7747 ( .A1(n10750), .A2(n10751), .ZN(n10749) );
  NAND2_X1 U7748 ( .A1(n6557), .A2(n10749), .ZN(n9828) );
  MUX2_X1 U7749 ( .A(n10899), .B(P1_REG1_REG_4__SCAN_IN), .S(n9833), .Z(n9827)
         );
  NOR2_X1 U7750 ( .A1(n9828), .A2(n9827), .ZN(n9826) );
  AOI21_X1 U7751 ( .B1(n10899), .B2(n6558), .A(n9826), .ZN(n10738) );
  MUX2_X1 U7752 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6560), .S(n10731), .Z(n10737) );
  NAND2_X1 U7753 ( .A1(n10738), .A2(n10737), .ZN(n10736) );
  OAI21_X1 U7754 ( .B1(n6560), .B2(n6559), .A(n10736), .ZN(n10688) );
  NAND2_X1 U7755 ( .A1(n10687), .A2(n10688), .ZN(n10686) );
  NAND2_X1 U7756 ( .A1(n6561), .A2(n10686), .ZN(n6583) );
  INV_X1 U7757 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U7758 ( .A1(n7201), .A2(n10956), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6562), .ZN(n6582) );
  NOR2_X1 U7759 ( .A1(n6583), .A2(n6582), .ZN(n6581) );
  OR2_X1 U7760 ( .A1(n6563), .A2(n6581), .ZN(n6564) );
  NAND2_X1 U7761 ( .A1(n6564), .A2(n6565), .ZN(n6671) );
  OAI21_X1 U7762 ( .B1(n6565), .B2(n6564), .A(n6671), .ZN(n6566) );
  NAND2_X1 U7763 ( .A1(n6566), .A2(n10815), .ZN(n6567) );
  OAI211_X1 U7764 ( .C1(n6569), .C2(n10808), .A(n6568), .B(n6567), .ZN(
        P1_U3249) );
  INV_X1 U7765 ( .A(n7500), .ZN(n6575) );
  NAND2_X1 U7766 ( .A1(n6571), .A2(n6570), .ZN(n6677) );
  NAND2_X1 U7767 ( .A1(n6677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U7768 ( .A1(n6572), .A2(n10552), .ZN(n6578) );
  OR2_X1 U7769 ( .A1(n6572), .A2(n10552), .ZN(n6573) );
  INV_X1 U7770 ( .A(n7501), .ZN(n6847) );
  OAI222_X1 U7771 ( .A1(n8024), .A2(n6575), .B1(n6847), .B2(P1_U3084), .C1(
        n10528), .C2(n10144), .ZN(P1_U3343) );
  INV_X1 U7772 ( .A(n7512), .ZN(n6580) );
  AOI22_X1 U7773 ( .A1(n9338), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9682), .ZN(n6574) );
  OAI21_X1 U7774 ( .B1(n6580), .B2(n9684), .A(n6574), .ZN(P2_U3347) );
  INV_X1 U7775 ( .A(n7402), .ZN(n7393) );
  OAI222_X1 U7776 ( .A1(n9687), .A2(n6576), .B1(n9684), .B2(n6575), .C1(n9691), 
        .C2(n7393), .ZN(P2_U3348) );
  INV_X2 U7777 ( .A(P2_U3966), .ZN(n9333) );
  NAND2_X1 U7778 ( .A1(n9333), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n6577) );
  OAI21_X1 U7779 ( .B1(n9547), .B2(n9333), .A(n6577), .ZN(P2_U3570) );
  NAND2_X1 U7780 ( .A1(n6578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6579) );
  XNOR2_X1 U7781 ( .A(n6579), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10703) );
  INV_X1 U7782 ( .A(n10703), .ZN(n10710) );
  INV_X1 U7783 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10527) );
  OAI222_X1 U7784 ( .A1(n8024), .A2(n6580), .B1(n10710), .B2(P1_U3084), .C1(
        n10527), .C2(n10144), .ZN(P1_U3342) );
  AOI21_X1 U7785 ( .B1(n6583), .B2(n6582), .A(n6581), .ZN(n6592) );
  AOI21_X1 U7786 ( .B1(n6586), .B2(n6585), .A(n6584), .ZN(n6589) );
  AND2_X1 U7787 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7216) );
  AOI21_X1 U7788 ( .B1(n10744), .B2(n7201), .A(n7216), .ZN(n6588) );
  NAND2_X1 U7789 ( .A1(n10813), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6587) );
  OAI211_X1 U7790 ( .C1(n6589), .C2(n10808), .A(n6588), .B(n6587), .ZN(n6590)
         );
  INV_X1 U7791 ( .A(n6590), .ZN(n6591) );
  OAI21_X1 U7792 ( .B1(n6592), .B2(n10702), .A(n6591), .ZN(P1_U3248) );
  NAND2_X1 U7793 ( .A1(n5752), .A2(SI_0_), .ZN(n6594) );
  INV_X1 U7794 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6593) );
  XNOR2_X1 U7795 ( .A(n6594), .B(n6593), .ZN(n10148) );
  INV_X1 U7796 ( .A(n7153), .ZN(n6609) );
  NAND2_X1 U7797 ( .A1(n5026), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U7798 ( .A1(n5024), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6596) );
  INV_X1 U7799 ( .A(n7085), .ZN(n7174) );
  INV_X1 U7800 ( .A(n6647), .ZN(n8744) );
  INV_X1 U7801 ( .A(n10990), .ZN(n10030) );
  NAND2_X1 U7802 ( .A1(n6833), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7803 ( .A1(n5024), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7804 ( .A1(n6834), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6601) );
  NAND4_X1 U7805 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n6640)
         );
  INV_X1 U7806 ( .A(n7189), .ZN(n6605) );
  NAND2_X1 U7807 ( .A1(n9812), .A2(n7118), .ZN(n8575) );
  NAND2_X1 U7808 ( .A1(n6605), .A2(n8575), .ZN(n8747) );
  NAND2_X1 U7809 ( .A1(n6400), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6607) );
  INV_X1 U7810 ( .A(n6877), .ZN(n8524) );
  NAND3_X1 U7811 ( .A1(n8747), .A2(n6689), .A3(n7153), .ZN(n6608) );
  OAI21_X1 U7812 ( .B1(n7174), .B2(n10030), .A(n6608), .ZN(n7169) );
  AOI21_X1 U7813 ( .B1(n7191), .B2(n6609), .A(n7169), .ZN(n6822) );
  NOR2_X1 U7814 ( .A1(n11057), .A2(n6636), .ZN(n6625) );
  INV_X1 U7815 ( .A(n10150), .ZN(n6621) );
  NOR4_X1 U7816 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6613) );
  NOR4_X1 U7817 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6612) );
  NOR4_X1 U7818 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6611) );
  NOR4_X1 U7819 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6610) );
  NAND4_X1 U7820 ( .A1(n6613), .A2(n6612), .A3(n6611), .A4(n6610), .ZN(n6619)
         );
  NOR2_X1 U7821 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6617) );
  NOR4_X1 U7822 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6616) );
  NOR4_X1 U7823 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6615) );
  NOR4_X1 U7824 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6614) );
  NAND4_X1 U7825 ( .A1(n6617), .A2(n6616), .A3(n6615), .A4(n6614), .ZN(n6618)
         );
  NOR2_X1 U7826 ( .A1(n6619), .A2(n6618), .ZN(n6620) );
  NOR2_X1 U7827 ( .A1(n6621), .A2(n6620), .ZN(n6630) );
  INV_X1 U7828 ( .A(n6630), .ZN(n6622) );
  NAND2_X1 U7829 ( .A1(n6622), .A2(n6631), .ZN(n6624) );
  OR2_X1 U7830 ( .A1(n6647), .A2(n6877), .ZN(n6623) );
  NAND2_X1 U7831 ( .A1(n6623), .A2(n10669), .ZN(n6634) );
  INV_X1 U7832 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U7833 ( .A1(n10150), .A2(n10668), .ZN(n6627) );
  NAND2_X1 U7834 ( .A1(n8222), .A2(n8023), .ZN(n6626) );
  INV_X1 U7835 ( .A(n10666), .ZN(n6628) );
  NAND2_X1 U7836 ( .A1(n11118), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6629) );
  OAI21_X1 U7837 ( .B1(n6822), .B2(n11118), .A(n6629), .ZN(P1_U3523) );
  OR2_X1 U7838 ( .A1(n6631), .A2(n6630), .ZN(n7098) );
  INV_X1 U7839 ( .A(n7098), .ZN(n6632) );
  NAND2_X1 U7840 ( .A1(n6632), .A2(n10666), .ZN(n6646) );
  OR2_X1 U7841 ( .A1(n7153), .A2(n7593), .ZN(n6650) );
  NAND2_X1 U7842 ( .A1(n6689), .A2(n6650), .ZN(n6633) );
  AND3_X1 U7843 ( .A1(n6646), .A2(n10669), .A3(n6633), .ZN(n6882) );
  NAND2_X1 U7844 ( .A1(n6646), .A2(n11109), .ZN(n6878) );
  INV_X1 U7845 ( .A(n6634), .ZN(n7100) );
  NAND2_X1 U7846 ( .A1(n6878), .A2(n7100), .ZN(n6635) );
  NOR2_X1 U7847 ( .A1(n6882), .A2(n6635), .ZN(n6838) );
  INV_X1 U7848 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U7849 ( .A1(n7101), .A2(n6879), .ZN(n9087) );
  INV_X1 U7850 ( .A(n9087), .ZN(n6642) );
  NAND2_X1 U7851 ( .A1(n8805), .A2(n6877), .ZN(n6637) );
  INV_X1 U7852 ( .A(n6879), .ZN(n6638) );
  OAI22_X1 U7853 ( .A1(n7118), .A2(n9128), .B1(n6879), .B2(n10674), .ZN(n6639)
         );
  NAND2_X1 U7854 ( .A1(n6640), .A2(n6825), .ZN(n6644) );
  NOR2_X1 U7855 ( .A1(n6879), .A2(n10673), .ZN(n6641) );
  AOI21_X1 U7856 ( .B1(n7191), .B2(n6642), .A(n6641), .ZN(n6643) );
  NAND2_X1 U7857 ( .A1(n6644), .A2(n6643), .ZN(n6687) );
  NAND2_X1 U7858 ( .A1(n6645), .A2(n6687), .ZN(n6691) );
  OAI21_X1 U7859 ( .B1(n6645), .B2(n6687), .A(n6691), .ZN(n9814) );
  INV_X1 U7860 ( .A(n6646), .ZN(n6651) );
  AND3_X1 U7861 ( .A1(n11109), .A2(n10669), .A3(n6647), .ZN(n6648) );
  NAND2_X1 U7862 ( .A1(n9814), .A2(n9787), .ZN(n6655) );
  AND2_X1 U7863 ( .A1(n10669), .A2(n6877), .ZN(n6649) );
  AND2_X1 U7864 ( .A1(n6651), .A2(n6649), .ZN(n6705) );
  INV_X1 U7865 ( .A(n6650), .ZN(n7120) );
  NAND3_X1 U7866 ( .A1(n6651), .A2(n10669), .A3(n7120), .ZN(n6653) );
  NAND2_X1 U7867 ( .A1(n10669), .A2(n8795), .ZN(n6652) );
  AOI22_X1 U7868 ( .A1(n9791), .A2(n7085), .B1(n7191), .B2(n9773), .ZN(n6654)
         );
  OAI211_X1 U7869 ( .C1(n6838), .C2(n6656), .A(n6655), .B(n6654), .ZN(P1_U3230) );
  NAND2_X1 U7870 ( .A1(n9054), .A2(P2_U3966), .ZN(n6657) );
  OAI21_X1 U7871 ( .B1(P2_U3966), .B2(n6658), .A(n6657), .ZN(P2_U3556) );
  NOR2_X1 U7872 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7302), .ZN(n7550) );
  INV_X1 U7873 ( .A(n7550), .ZN(n6659) );
  OAI21_X1 U7874 ( .B1(n10809), .B2(n6849), .A(n6659), .ZN(n6666) );
  NAND2_X1 U7875 ( .A1(n6667), .A2(n6544), .ZN(n6660) );
  NAND2_X1 U7876 ( .A1(n6661), .A2(n6660), .ZN(n6664) );
  INV_X1 U7877 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6662) );
  MUX2_X1 U7878 ( .A(n6662), .B(P1_REG2_REG_9__SCAN_IN), .S(n7496), .Z(n6663)
         );
  AOI211_X1 U7879 ( .C1(n6664), .C2(n6663), .A(n10808), .B(n5115), .ZN(n6665)
         );
  AOI211_X1 U7880 ( .C1(n10813), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n6666), .B(
        n6665), .ZN(n6674) );
  NAND2_X1 U7881 ( .A1(n6667), .A2(n10974), .ZN(n6669) );
  INV_X1 U7882 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6668) );
  MUX2_X1 U7883 ( .A(n6668), .B(P1_REG1_REG_9__SCAN_IN), .S(n7496), .Z(n6670)
         );
  AOI21_X1 U7884 ( .B1(n6671), .B2(n6669), .A(n6670), .ZN(n6843) );
  AND3_X1 U7885 ( .A1(n6671), .A2(n6670), .A3(n6669), .ZN(n6672) );
  OAI21_X1 U7886 ( .B1(n6843), .B2(n6672), .A(n10815), .ZN(n6673) );
  NAND2_X1 U7887 ( .A1(n6674), .A2(n6673), .ZN(P1_U3250) );
  INV_X1 U7888 ( .A(n7254), .ZN(n6913) );
  NAND2_X1 U7889 ( .A1(n6913), .A2(P2_U3966), .ZN(n6675) );
  OAI21_X1 U7890 ( .B1(P2_U3966), .B2(n6593), .A(n6675), .ZN(P2_U3552) );
  INV_X1 U7891 ( .A(n7423), .ZN(n7419) );
  INV_X1 U7892 ( .A(n7634), .ZN(n6679) );
  OAI222_X1 U7893 ( .A1(n7419), .A2(P2_U3152), .B1(n9684), .B2(n6679), .C1(
        n6676), .C2(n9687), .ZN(P2_U3346) );
  NAND2_X1 U7894 ( .A1(n6873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6678) );
  XNOR2_X1 U7895 ( .A(n6678), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7635) );
  INV_X1 U7896 ( .A(n7635), .ZN(n7002) );
  OAI222_X1 U7897 ( .A1(n10144), .A2(n10525), .B1(n8024), .B2(n6679), .C1(
        P1_U3084), .C2(n7002), .ZN(P1_U3341) );
  NAND2_X1 U7898 ( .A1(n7085), .A2(n9159), .ZN(n6686) );
  NAND2_X1 U7899 ( .A1(n7197), .A2(n9160), .ZN(n6685) );
  NAND2_X1 U7900 ( .A1(n6686), .A2(n6685), .ZN(n6704) );
  INV_X1 U7901 ( .A(n6687), .ZN(n6690) );
  AOI21_X1 U7902 ( .B1(n8805), .B2(n8801), .A(n9850), .ZN(n6688) );
  NAND2_X4 U7903 ( .A1(n7103), .A2(n7101), .ZN(n9157) );
  NAND2_X1 U7904 ( .A1(n6692), .A2(n6691), .ZN(n6697) );
  NAND2_X1 U7905 ( .A1(n7085), .A2(n6825), .ZN(n6694) );
  NAND2_X1 U7906 ( .A1(n7197), .A2(n9133), .ZN(n6693) );
  NAND2_X1 U7907 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  INV_X1 U7908 ( .A(n6701), .ZN(n6699) );
  NAND2_X1 U7909 ( .A1(n6699), .A2(n6700), .ZN(n6703) );
  AOI22_X1 U7910 ( .A1(n6704), .A2(n6703), .B1(n6830), .B2(n6702), .ZN(n6713)
         );
  AND2_X2 U7911 ( .A1(n8744), .A2(n9821), .ZN(n10993) );
  AOI22_X1 U7912 ( .A1(n9758), .A2(n9812), .B1(n7197), .B2(n9773), .ZN(n6712)
         );
  INV_X1 U7913 ( .A(n6838), .ZN(n6710) );
  NAND2_X1 U7914 ( .A1(n6833), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U7915 ( .A1(n5024), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U7916 ( .A1(n6834), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6706) );
  AOI22_X1 U7917 ( .A1(n6710), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9791), .B2(
        n10863), .ZN(n6711) );
  OAI211_X1 U7918 ( .C1(n6713), .C2(n9785), .A(n6712), .B(n6711), .ZN(P1_U3220) );
  INV_X1 U7919 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10779) );
  MUX2_X1 U7920 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7250), .S(n10778), .Z(n6714)
         );
  INV_X1 U7921 ( .A(n6714), .ZN(n10774) );
  NOR3_X1 U7922 ( .A1(n10779), .A2(n7373), .A3(n10774), .ZN(n10773) );
  AND2_X1 U7923 ( .A1(n10778), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U7924 ( .A1(n10793), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6716) );
  OAI21_X1 U7925 ( .B1(n10793), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6716), .ZN(
        n10790) );
  NOR2_X1 U7926 ( .A1(n10791), .A2(n10790), .ZN(n10789) );
  AOI21_X1 U7927 ( .B1(n10793), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10789), .ZN(
        n6755) );
  MUX2_X1 U7928 ( .A(n6717), .B(P2_REG2_REG_3__SCAN_IN), .S(n6735), .Z(n6754)
         );
  NOR2_X1 U7929 ( .A1(n6755), .A2(n6754), .ZN(n6753) );
  NAND2_X1 U7930 ( .A1(n6733), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6718) );
  OAI21_X1 U7931 ( .B1(n6733), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6718), .ZN(
        n6766) );
  NOR2_X1 U7932 ( .A1(n6767), .A2(n6766), .ZN(n6765) );
  MUX2_X1 U7933 ( .A(n6719), .B(P2_REG2_REG_5__SCAN_IN), .S(n6731), .Z(n6778)
         );
  NOR2_X1 U7934 ( .A1(n6779), .A2(n6778), .ZN(n6777) );
  AOI21_X1 U7935 ( .B1(n6731), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6777), .ZN(
        n6728) );
  NAND2_X1 U7936 ( .A1(n6793), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6720) );
  OAI21_X1 U7937 ( .B1(n6793), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6720), .ZN(
        n6727) );
  NOR2_X1 U7938 ( .A1(n6728), .A2(n6727), .ZN(n6788) );
  OAI21_X1 U7939 ( .B1(n6721), .B2(P2_U3152), .A(n9047), .ZN(n6722) );
  INV_X1 U7940 ( .A(n6722), .ZN(n6723) );
  NAND2_X1 U7941 ( .A1(n6724), .A2(n6723), .ZN(n6745) );
  NAND2_X1 U7942 ( .A1(n6745), .A2(n6743), .ZN(n6725) );
  NAND2_X1 U7943 ( .A1(n6725), .A2(n9333), .ZN(n6729) );
  NOR2_X1 U7944 ( .A1(n6355), .A2(n9690), .ZN(n6726) );
  AOI211_X1 U7945 ( .C1(n6728), .C2(n6727), .A(n6788), .B(n10788), .ZN(n6752)
         );
  NAND2_X1 U7946 ( .A1(n6729), .A2(n6355), .ZN(n10763) );
  NAND2_X1 U7947 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8477) );
  INV_X1 U7948 ( .A(n8477), .ZN(n6730) );
  AOI21_X1 U7949 ( .B1(n10787), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6730), .ZN(
        n6749) );
  MUX2_X1 U7950 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6732), .S(n6731), .Z(n6781)
         );
  NAND2_X1 U7951 ( .A1(n6733), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6741) );
  MUX2_X1 U7952 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6734), .S(n6733), .Z(n6770)
         );
  MUX2_X1 U7953 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6736), .S(n6735), .Z(n6758)
         );
  NAND2_X1 U7954 ( .A1(n10793), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6740) );
  MUX2_X1 U7955 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6737), .S(n10793), .Z(n10797) );
  MUX2_X1 U7956 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6738), .S(n10778), .Z(n10781) );
  NAND3_X1 U7957 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10781), .ZN(n10780) );
  OAI21_X1 U7958 ( .B1(n6739), .B2(n6738), .A(n10780), .ZN(n10798) );
  NAND2_X1 U7959 ( .A1(n10797), .A2(n10798), .ZN(n10795) );
  NAND2_X1 U7960 ( .A1(n6740), .A2(n10795), .ZN(n6759) );
  NAND2_X1 U7961 ( .A1(n6758), .A2(n6759), .ZN(n6757) );
  OAI21_X1 U7962 ( .B1(n6762), .B2(n6736), .A(n6757), .ZN(n6771) );
  NAND2_X1 U7963 ( .A1(n6770), .A2(n6771), .ZN(n6769) );
  NAND2_X1 U7964 ( .A1(n6741), .A2(n6769), .ZN(n6782) );
  NAND2_X1 U7965 ( .A1(n6781), .A2(n6782), .ZN(n6780) );
  OAI21_X1 U7966 ( .B1(n6785), .B2(n6732), .A(n6780), .ZN(n6747) );
  MUX2_X1 U7967 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6742), .S(n6793), .Z(n6746)
         );
  AND2_X1 U7968 ( .A1(n6743), .A2(n9690), .ZN(n6744) );
  NAND2_X1 U7969 ( .A1(n6746), .A2(n6747), .ZN(n6794) );
  OAI211_X1 U7970 ( .C1(n6747), .C2(n6746), .A(n10796), .B(n6794), .ZN(n6748)
         );
  OAI211_X1 U7971 ( .C1(n10763), .C2(n6750), .A(n6749), .B(n6748), .ZN(n6751)
         );
  OR2_X1 U7972 ( .A1(n6752), .A2(n6751), .ZN(P2_U3251) );
  AOI211_X1 U7973 ( .C1(n6755), .C2(n6754), .A(n6753), .B(n10788), .ZN(n6764)
         );
  INV_X1 U7974 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10458) );
  NOR2_X1 U7975 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10458), .ZN(n6756) );
  AOI21_X1 U7976 ( .B1(n10787), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6756), .ZN(
        n6761) );
  OAI211_X1 U7977 ( .C1(n6759), .C2(n6758), .A(n10796), .B(n6757), .ZN(n6760)
         );
  OAI211_X1 U7978 ( .C1(n10763), .C2(n6762), .A(n6761), .B(n6760), .ZN(n6763)
         );
  OR2_X1 U7979 ( .A1(n6764), .A2(n6763), .ZN(P2_U3248) );
  AOI211_X1 U7980 ( .C1(n6767), .C2(n6766), .A(n6765), .B(n10788), .ZN(n6776)
         );
  INV_X1 U7981 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10483) );
  NOR2_X1 U7982 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10483), .ZN(n6768) );
  AOI21_X1 U7983 ( .B1(n10787), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6768), .ZN(
        n6773) );
  OAI211_X1 U7984 ( .C1(n6771), .C2(n6770), .A(n10796), .B(n6769), .ZN(n6772)
         );
  OAI211_X1 U7985 ( .C1(n10763), .C2(n6774), .A(n6773), .B(n6772), .ZN(n6775)
         );
  OR2_X1 U7986 ( .A1(n6776), .A2(n6775), .ZN(P2_U3249) );
  AOI211_X1 U7987 ( .C1(n6779), .C2(n6778), .A(n6777), .B(n10788), .ZN(n6787)
         );
  NOR2_X1 U7988 ( .A1(n10473), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9049) );
  AOI21_X1 U7989 ( .B1(n10787), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9049), .ZN(
        n6784) );
  OAI211_X1 U7990 ( .C1(n6782), .C2(n6781), .A(n10796), .B(n6780), .ZN(n6783)
         );
  OAI211_X1 U7991 ( .C1(n10763), .C2(n6785), .A(n6784), .B(n6783), .ZN(n6786)
         );
  OR2_X1 U7992 ( .A1(n6787), .A2(n6786), .ZN(P2_U3250) );
  AOI21_X1 U7993 ( .B1(n6793), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6788), .ZN(
        n6791) );
  MUX2_X1 U7994 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7678), .S(n6804), .Z(n6789)
         );
  INV_X1 U7995 ( .A(n6789), .ZN(n6790) );
  NOR2_X1 U7996 ( .A1(n6791), .A2(n6790), .ZN(n6803) );
  AOI211_X1 U7997 ( .C1(n6791), .C2(n6790), .A(n6803), .B(n10788), .ZN(n6802)
         );
  INV_X1 U7998 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10445) );
  NOR2_X1 U7999 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10445), .ZN(n6792) );
  AOI21_X1 U8000 ( .B1(n10787), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6792), .ZN(
        n6800) );
  NAND2_X1 U8001 ( .A1(n6793), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U8002 ( .A1(n6795), .A2(n6794), .ZN(n6798) );
  MUX2_X1 U8003 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6796), .S(n6804), .Z(n6797)
         );
  NAND2_X1 U8004 ( .A1(n6797), .A2(n6798), .ZN(n6810) );
  OAI211_X1 U8005 ( .C1(n6798), .C2(n6797), .A(n10796), .B(n6810), .ZN(n6799)
         );
  OAI211_X1 U8006 ( .C1(n10763), .C2(n6811), .A(n6800), .B(n6799), .ZN(n6801)
         );
  OR2_X1 U8007 ( .A1(n6802), .A2(n6801), .ZN(P2_U3252) );
  INV_X1 U8008 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6805) );
  MUX2_X1 U8009 ( .A(n6805), .B(P2_REG2_REG_8__SCAN_IN), .S(n6865), .Z(n6806)
         );
  INV_X1 U8010 ( .A(n6806), .ZN(n6807) );
  NOR2_X1 U8011 ( .A1(n6808), .A2(n6807), .ZN(n6859) );
  AOI211_X1 U8012 ( .C1(n6808), .C2(n6807), .A(n6859), .B(n10788), .ZN(n6818)
         );
  NOR2_X1 U8013 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10258), .ZN(n6809) );
  AOI21_X1 U8014 ( .B1(n10787), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6809), .ZN(
        n6816) );
  OAI21_X1 U8015 ( .B1(n6811), .B2(n6796), .A(n6810), .ZN(n6814) );
  MUX2_X1 U8016 ( .A(n6812), .B(P2_REG1_REG_8__SCAN_IN), .S(n6865), .Z(n6813)
         );
  NAND2_X1 U8017 ( .A1(n6813), .A2(n6814), .ZN(n6864) );
  OAI211_X1 U8018 ( .C1(n6814), .C2(n6813), .A(n10796), .B(n6864), .ZN(n6815)
         );
  OAI211_X1 U8019 ( .C1(n10763), .C2(n6865), .A(n6816), .B(n6815), .ZN(n6817)
         );
  OR2_X1 U8020 ( .A1(n6818), .A2(n6817), .ZN(P2_U3253) );
  INV_X2 U8021 ( .A(n11120), .ZN(n10137) );
  INV_X1 U8022 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6820) );
  OR2_X1 U8023 ( .A1(n10137), .A2(n6820), .ZN(n6821) );
  OAI21_X1 U8024 ( .B1(n6822), .B2(n11120), .A(n6821), .ZN(P1_U3454) );
  NAND2_X1 U8025 ( .A1(n8421), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6823) );
  INV_X2 U8026 ( .A(n9087), .ZN(n9133) );
  NAND2_X1 U8027 ( .A1(n7183), .A2(n9133), .ZN(n6827) );
  NAND2_X1 U8028 ( .A1(n10863), .A2(n9143), .ZN(n6826) );
  XNOR2_X1 U8029 ( .A(n6828), .B(n9157), .ZN(n6891) );
  AND2_X1 U8030 ( .A1(n7183), .A2(n9160), .ZN(n6829) );
  AOI21_X1 U8031 ( .B1(n10863), .B2(n9159), .A(n6829), .ZN(n6892) );
  XNOR2_X1 U8032 ( .A(n6891), .B(n6892), .ZN(n6831) );
  NAND2_X1 U8033 ( .A1(n6830), .A2(n6831), .ZN(n6895) );
  OAI21_X1 U8034 ( .B1(n6831), .B2(n6830), .A(n6895), .ZN(n6841) );
  INV_X1 U8035 ( .A(n9758), .ZN(n9793) );
  INV_X1 U8036 ( .A(n7183), .ZN(n10842) );
  OAI22_X1 U8037 ( .A1(n9793), .A2(n7174), .B1(n10842), .B2(n9799), .ZN(n6840)
         );
  INV_X1 U8038 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8039 ( .A1(n5026), .A2(n6832), .ZN(n6837) );
  NAND2_X1 U8040 ( .A1(n5024), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6835) );
  INV_X1 U8041 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10820) );
  OAI22_X1 U8042 ( .A1(n7175), .A2(n9756), .B1(n6838), .B2(n10820), .ZN(n6839)
         );
  AOI211_X1 U8043 ( .C1(n6841), .C2(n9787), .A(n6840), .B(n6839), .ZN(n6842)
         );
  INV_X1 U8044 ( .A(n6842), .ZN(P1_U3235) );
  AOI21_X1 U8045 ( .B1(n6668), .B2(n6849), .A(n6843), .ZN(n6845) );
  INV_X1 U8046 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7620) );
  AOI22_X1 U8047 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6847), .B1(n7501), .B2(
        n7620), .ZN(n6844) );
  NOR2_X1 U8048 ( .A1(n6845), .A2(n6844), .ZN(n6993) );
  AOI21_X1 U8049 ( .B1(n6845), .B2(n6844), .A(n6993), .ZN(n6858) );
  NAND2_X1 U8050 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n6846) );
  OAI21_X1 U8051 ( .B1(n10809), .B2(n6847), .A(n6846), .ZN(n6856) );
  INV_X1 U8052 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6850) );
  MUX2_X1 U8053 ( .A(n6850), .B(P1_REG2_REG_10__SCAN_IN), .S(n7501), .Z(n6851)
         );
  INV_X1 U8054 ( .A(n6851), .ZN(n6852) );
  OAI211_X1 U8055 ( .C1(n6853), .C2(n6852), .A(n10746), .B(n7003), .ZN(n6854)
         );
  INV_X1 U8056 ( .A(n6854), .ZN(n6855) );
  AOI211_X1 U8057 ( .C1(n10813), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n6856), .B(
        n6855), .ZN(n6857) );
  OAI21_X1 U8058 ( .B1(n6858), .B2(n10702), .A(n6857), .ZN(P1_U3251) );
  INV_X1 U8059 ( .A(n6865), .ZN(n6860) );
  AOI21_X1 U8060 ( .B1(n6860), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6859), .ZN(
        n6863) );
  NAND2_X1 U8061 ( .A1(n6963), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6861) );
  OAI21_X1 U8062 ( .B1(n6963), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6861), .ZN(
        n6862) );
  NOR2_X1 U8063 ( .A1(n6863), .A2(n6862), .ZN(n6962) );
  AOI211_X1 U8064 ( .C1(n6863), .C2(n6862), .A(n6962), .B(n10788), .ZN(n6872)
         );
  NOR2_X1 U8065 ( .A1(n5992), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7700) );
  AOI21_X1 U8066 ( .B1(n10787), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7700), .ZN(
        n6870) );
  OAI21_X1 U8067 ( .B1(n6865), .B2(n6812), .A(n6864), .ZN(n6868) );
  MUX2_X1 U8068 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6866), .S(n6963), .Z(n6867)
         );
  NAND2_X1 U8069 ( .A1(n6867), .A2(n6868), .ZN(n6968) );
  OAI211_X1 U8070 ( .C1(n6868), .C2(n6867), .A(n10796), .B(n6968), .ZN(n6869)
         );
  OAI211_X1 U8071 ( .C1(n10763), .C2(n6969), .A(n6870), .B(n6869), .ZN(n6871)
         );
  OR2_X1 U8072 ( .A1(n6872), .A2(n6871), .ZN(P2_U3254) );
  INV_X1 U8073 ( .A(n7877), .ZN(n6907) );
  OAI21_X1 U8074 ( .B1(n6873), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U8075 ( .A1(n6875), .A2(n6874), .ZN(n6908) );
  OR2_X1 U8076 ( .A1(n6875), .A2(n6874), .ZN(n6876) );
  INV_X1 U8077 ( .A(n7878), .ZN(n7138) );
  OAI222_X1 U8078 ( .A1(n8024), .A2(n6907), .B1(n7138), .B2(P1_U3084), .C1(
        n10523), .C2(n10144), .ZN(P1_U3340) );
  MUX2_X1 U8079 ( .A(n6878), .B(n6877), .S(n8744), .Z(n6881) );
  AND2_X1 U8080 ( .A1(n6879), .A2(n7859), .ZN(n6880) );
  NAND2_X1 U8081 ( .A1(n6881), .A2(n6880), .ZN(n6883) );
  AOI21_X2 U8082 ( .B1(n6883), .B2(P1_STATE_REG_SCAN_IN), .A(n6882), .ZN(n9760) );
  NAND2_X1 U8083 ( .A1(n5603), .A2(n9160), .ZN(n6888) );
  NAND2_X1 U8084 ( .A1(n8421), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U8085 ( .A1(n8320), .A2(n10743), .ZN(n6884) );
  NAND2_X1 U8086 ( .A1(n7089), .A2(n9133), .ZN(n6887) );
  NAND2_X1 U8087 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  XNOR2_X1 U8088 ( .A(n6889), .B(n9157), .ZN(n6921) );
  AND2_X1 U8089 ( .A1(n7089), .A2(n9160), .ZN(n6890) );
  AOI21_X1 U8090 ( .B1(n5603), .B2(n9159), .A(n6890), .ZN(n6922) );
  XNOR2_X1 U8091 ( .A(n6921), .B(n6922), .ZN(n6919) );
  INV_X1 U8092 ( .A(n6891), .ZN(n6893) );
  NAND2_X1 U8093 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  NAND2_X1 U8094 ( .A1(n6895), .A2(n6894), .ZN(n6920) );
  XNOR2_X1 U8095 ( .A(n6919), .B(n6920), .ZN(n6896) );
  NAND2_X1 U8096 ( .A1(n6896), .A2(n9787), .ZN(n6905) );
  NAND2_X1 U8097 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10754) );
  INV_X1 U8098 ( .A(n10754), .ZN(n6903) );
  NAND2_X1 U8099 ( .A1(n5024), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U8100 ( .A1(n8401), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6900) );
  INV_X1 U8101 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6897) );
  XNOR2_X1 U8102 ( .A(n6897), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7274) );
  NAND2_X1 U8103 ( .A1(n5026), .A2(n7274), .ZN(n6899) );
  NAND2_X1 U8104 ( .A1(n6834), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6898) );
  INV_X1 U8105 ( .A(n10862), .ZN(n7092) );
  OAI22_X1 U8106 ( .A1(n9756), .A2(n7092), .B1(n10880), .B2(n9799), .ZN(n6902)
         );
  AOI211_X1 U8107 ( .C1(n9758), .C2(n10863), .A(n6903), .B(n6902), .ZN(n6904)
         );
  OAI211_X1 U8108 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9760), .A(n6905), .B(
        n6904), .ZN(P1_U3216) );
  INV_X1 U8109 ( .A(n7599), .ZN(n7595) );
  OAI222_X1 U8110 ( .A1(n9691), .A2(n7595), .B1(n9684), .B2(n6907), .C1(n6906), 
        .C2(n9687), .ZN(P2_U3345) );
  INV_X1 U8111 ( .A(n7959), .ZN(n6911) );
  NAND2_X1 U8112 ( .A1(n6908), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6909) );
  XNOR2_X1 U8113 ( .A(n6909), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7960) );
  INV_X1 U8114 ( .A(n7960), .ZN(n6910) );
  INV_X1 U8115 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10522) );
  OAI222_X1 U8116 ( .A1(n8024), .A2(n6911), .B1(n6910), .B2(P1_U3084), .C1(
        n10522), .C2(n10144), .ZN(P1_U3339) );
  INV_X1 U8117 ( .A(n7848), .ZN(n7854) );
  OAI222_X1 U8118 ( .A1(n7854), .A2(P2_U3152), .B1(n9687), .B2(n6912), .C1(
        n6911), .C2(n9684), .ZN(P2_U3344) );
  NAND2_X1 U8119 ( .A1(n10623), .A2(n7237), .ZN(n10607) );
  INV_X1 U8120 ( .A(n10607), .ZN(n9055) );
  AOI22_X1 U8121 ( .A1(n9055), .A2(n6913), .B1(n7375), .B2(n10623), .ZN(n6918)
         );
  INV_X1 U8122 ( .A(n6914), .ZN(n6917) );
  INV_X1 U8123 ( .A(n9314), .ZN(n10613) );
  NOR2_X1 U8124 ( .A1(n10485), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10766) );
  AOI21_X1 U8125 ( .B1(n10613), .B2(n7229), .A(n10766), .ZN(n6916) );
  AOI22_X1 U8126 ( .A1(n10611), .A2(n7375), .B1(n7014), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n6915) );
  OAI211_X1 U8127 ( .C1(n6918), .C2(n6917), .A(n6916), .B(n6915), .ZN(P2_U3234) );
  INV_X1 U8128 ( .A(n7274), .ZN(n6947) );
  NAND2_X1 U8129 ( .A1(n6920), .A2(n6919), .ZN(n6925) );
  INV_X1 U8130 ( .A(n6921), .ZN(n6923) );
  NAND2_X1 U8131 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  NAND2_X1 U8132 ( .A1(n10862), .A2(n9160), .ZN(n6930) );
  NAND2_X1 U8133 ( .A1(n8546), .A2(n6926), .ZN(n6928) );
  NAND2_X1 U8134 ( .A1(n8320), .A2(n9833), .ZN(n6927) );
  NAND2_X1 U8135 ( .A1(n7275), .A2(n9133), .ZN(n6929) );
  NAND2_X1 U8136 ( .A1(n6930), .A2(n6929), .ZN(n6931) );
  XNOR2_X1 U8137 ( .A(n6931), .B(n9152), .ZN(n7028) );
  AND2_X1 U8138 ( .A1(n7275), .A2(n9160), .ZN(n6932) );
  AOI21_X1 U8139 ( .B1(n10862), .B2(n9159), .A(n6932), .ZN(n7029) );
  XNOR2_X1 U8140 ( .A(n7028), .B(n7029), .ZN(n6934) );
  AOI21_X1 U8141 ( .B1(n6933), .B2(n6934), .A(n9785), .ZN(n6936) );
  NAND2_X1 U8142 ( .A1(n6936), .A2(n7033), .ZN(n6946) );
  NAND2_X1 U8143 ( .A1(n5024), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U8144 ( .A1(n8401), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6940) );
  AOI21_X1 U8145 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6937) );
  NOR2_X1 U8146 ( .A1(n6937), .A2(n7045), .ZN(n7151) );
  NAND2_X1 U8147 ( .A1(n5026), .A2(n7151), .ZN(n6939) );
  NAND2_X1 U8148 ( .A1(n6834), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U8149 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9829) );
  INV_X1 U8150 ( .A(n9829), .ZN(n6942) );
  AOI21_X1 U8151 ( .B1(n9758), .B2(n5603), .A(n6942), .ZN(n6943) );
  OAI21_X1 U8152 ( .B1(n9756), .B2(n7104), .A(n6943), .ZN(n6944) );
  AOI21_X1 U8153 ( .B1(n7275), .B2(n9773), .A(n6944), .ZN(n6945) );
  OAI211_X1 U8154 ( .C1(n9760), .C2(n6947), .A(n6946), .B(n6945), .ZN(P1_U3228) );
  AND2_X1 U8155 ( .A1(n6948), .A2(n10185), .ZN(n6950) );
  INV_X1 U8156 ( .A(n7232), .ZN(n6951) );
  INV_X1 U8157 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6958) );
  OR2_X1 U8158 ( .A1(n7254), .A2(n7375), .ZN(n8892) );
  NAND2_X1 U8159 ( .A1(n7254), .A2(n7375), .ZN(n7243) );
  NAND2_X1 U8160 ( .A1(n8892), .A2(n7243), .ZN(n8884) );
  NAND2_X1 U8161 ( .A1(n8877), .A2(n8891), .ZN(n6952) );
  NAND2_X1 U8162 ( .A1(n9555), .A2(n9045), .ZN(n9033) );
  NAND2_X2 U8163 ( .A1(n6952), .A2(n9033), .ZN(n9576) );
  AOI22_X1 U8164 ( .A1(n8884), .A2(n9576), .B1(n9574), .B2(n7229), .ZN(n7378)
         );
  NAND3_X1 U8165 ( .A1(n8877), .A2(n9045), .A3(n10922), .ZN(n6953) );
  OAI21_X1 U8166 ( .B1(n6315), .B2(n6954), .A(n6953), .ZN(n6955) );
  NAND2_X1 U8167 ( .A1(n6955), .A2(n9034), .ZN(n8275) );
  OR3_X1 U8168 ( .A1(n8877), .A2(n9045), .A3(n10922), .ZN(n10850) );
  AOI22_X1 U8169 ( .A1(n8884), .A2(n11129), .B1(n8880), .B2(n7375), .ZN(n6956)
         );
  NAND2_X1 U8170 ( .A1(n7378), .A2(n6956), .ZN(n6960) );
  NAND2_X1 U8171 ( .A1(n6960), .A2(n11135), .ZN(n6957) );
  OAI21_X1 U8172 ( .B1(n11135), .B2(n6958), .A(n6957), .ZN(P2_U3451) );
  NAND2_X1 U8173 ( .A1(n6960), .A2(n11132), .ZN(n6961) );
  OAI21_X1 U8174 ( .B1(n11132), .B2(n10762), .A(n6961), .ZN(P2_U3520) );
  AOI21_X1 U8175 ( .B1(n6963), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6962), .ZN(
        n6966) );
  NAND2_X1 U8176 ( .A1(n7402), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6964) );
  OAI21_X1 U8177 ( .B1(n7402), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6964), .ZN(
        n6965) );
  NOR2_X1 U8178 ( .A1(n6966), .A2(n6965), .ZN(n7401) );
  AOI211_X1 U8179 ( .C1(n6966), .C2(n6965), .A(n7401), .B(n10788), .ZN(n6976)
         );
  INV_X1 U8180 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10455) );
  NOR2_X1 U8181 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10455), .ZN(n6967) );
  AOI21_X1 U8182 ( .B1(n10787), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6967), .ZN(
        n6974) );
  OAI21_X1 U8183 ( .B1(n6969), .B2(n6866), .A(n6968), .ZN(n6972) );
  MUX2_X1 U8184 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6970), .S(n7402), .Z(n6971)
         );
  NAND2_X1 U8185 ( .A1(n6971), .A2(n6972), .ZN(n7392) );
  OAI211_X1 U8186 ( .C1(n6972), .C2(n6971), .A(n10796), .B(n7392), .ZN(n6973)
         );
  OAI211_X1 U8187 ( .C1(n10763), .C2(n7393), .A(n6974), .B(n6973), .ZN(n6975)
         );
  OR2_X1 U8188 ( .A1(n6976), .A2(n6975), .ZN(P2_U3255) );
  INV_X1 U8189 ( .A(n9250), .ZN(n9429) );
  NAND2_X1 U8190 ( .A1(n9429), .A2(P2_U3966), .ZN(n6977) );
  OAI21_X1 U8191 ( .B1(n5753), .B2(P2_U3966), .A(n6977), .ZN(P2_U3578) );
  OAI211_X1 U8192 ( .C1(n6980), .C2(n6979), .A(n6978), .B(n10623), .ZN(n6984)
         );
  NAND2_X1 U8193 ( .A1(n9691), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n10785) );
  OAI21_X1 U8194 ( .B1(n9313), .B2(n7265), .A(n10785), .ZN(n6982) );
  INV_X1 U8195 ( .A(n7347), .ZN(n10605) );
  OAI22_X1 U8196 ( .A1(n9319), .A2(n10852), .B1(n10605), .B2(n9314), .ZN(n6981) );
  AOI211_X1 U8197 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n7014), .A(n6982), .B(
        n6981), .ZN(n6983) );
  NAND2_X1 U8198 ( .A1(n6984), .A2(n6983), .ZN(P2_U3239) );
  INV_X1 U8199 ( .A(n8121), .ZN(n8127) );
  INV_X1 U8200 ( .A(n8050), .ZN(n6991) );
  INV_X1 U8201 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6985) );
  OAI222_X1 U8202 ( .A1(n8127), .A2(P2_U3152), .B1(n9684), .B2(n6991), .C1(
        n6985), .C2(n9687), .ZN(P2_U3343) );
  INV_X1 U8203 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10313) );
  INV_X1 U8204 ( .A(n6986), .ZN(n6987) );
  NAND2_X1 U8205 ( .A1(n6987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6988) );
  MUX2_X1 U8206 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6988), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6990) );
  NAND2_X1 U8207 ( .A1(n6990), .A2(n6989), .ZN(n7801) );
  OAI222_X1 U8208 ( .A1(n10144), .A2(n10313), .B1(n8024), .B2(n6991), .C1(
        P1_U3084), .C2(n7801), .ZN(P1_U3338) );
  NAND2_X1 U8209 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7839) );
  INV_X1 U8210 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6992) );
  MUX2_X1 U8211 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6992), .S(n7635), .Z(n6999)
         );
  NAND2_X1 U8212 ( .A1(n10703), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6996) );
  OR2_X1 U8213 ( .A1(n7501), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6995) );
  INV_X1 U8214 ( .A(n6993), .ZN(n6994) );
  NAND2_X1 U8215 ( .A1(n6995), .A2(n6994), .ZN(n10709) );
  NAND2_X1 U8216 ( .A1(n6996), .A2(n10709), .ZN(n6998) );
  OR2_X1 U8217 ( .A1(n10703), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6997) );
  NAND2_X1 U8218 ( .A1(n6998), .A2(n6997), .ZN(n10712) );
  NAND2_X1 U8219 ( .A1(n10712), .A2(n6999), .ZN(n7133) );
  OAI21_X1 U8220 ( .B1(n6999), .B2(n10712), .A(n7133), .ZN(n7000) );
  NAND2_X1 U8221 ( .A1(n10815), .A2(n7000), .ZN(n7001) );
  OAI211_X1 U8222 ( .C1(n10809), .C2(n7002), .A(n7839), .B(n7001), .ZN(n7007)
         );
  XNOR2_X1 U8223 ( .A(n7635), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U8224 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7501), .ZN(n7004) );
  AND2_X1 U8225 ( .A1(n10708), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10700) );
  OAI22_X1 U8226 ( .A1(n10700), .A2(n10703), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n10708), .ZN(n10706) );
  NOR2_X1 U8227 ( .A1(n10706), .A2(n7005), .ZN(n7139) );
  AOI211_X1 U8228 ( .C1(n7005), .C2(n10706), .A(n10808), .B(n7139), .ZN(n7006)
         );
  AOI211_X1 U8229 ( .C1(n10813), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7007), .B(
        n7006), .ZN(n7008) );
  INV_X1 U8230 ( .A(n7008), .ZN(P1_U3253) );
  INV_X1 U8231 ( .A(n7009), .ZN(n7010) );
  AOI21_X1 U8232 ( .B1(n7012), .B2(n7011), .A(n7010), .ZN(n7017) );
  INV_X2 U8233 ( .A(n10623), .ZN(n9306) );
  OAI22_X1 U8234 ( .A1(n7254), .A2(n9313), .B1(n9314), .B2(n9332), .ZN(n7013)
         );
  AOI21_X1 U8235 ( .B1(n10611), .B2(n7253), .A(n7013), .ZN(n7016) );
  OAI21_X1 U8236 ( .B1(n7014), .B2(P2_U3152), .A(P2_REG3_REG_1__SCAN_IN), .ZN(
        n7015) );
  OAI211_X1 U8237 ( .C1(n7017), .C2(n9306), .A(n7016), .B(n7015), .ZN(P2_U3224) );
  INV_X1 U8238 ( .A(n7018), .ZN(n7019) );
  AOI21_X1 U8239 ( .B1(n6978), .B2(n7019), .A(n9306), .ZN(n7023) );
  NOR3_X1 U8240 ( .A1(n10607), .A2(n7020), .A3(n9332), .ZN(n7022) );
  OAI21_X1 U8241 ( .B1(n7023), .B2(n7022), .A(n7021), .ZN(n7027) );
  OAI22_X1 U8242 ( .A1(n9319), .A2(n10886), .B1(n7381), .B2(n9314), .ZN(n7025)
         );
  OAI22_X1 U8243 ( .A1(n9313), .A2(n9332), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10458), .ZN(n7024) );
  NOR2_X1 U8244 ( .A1(n7025), .A2(n7024), .ZN(n7026) );
  OAI211_X1 U8245 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9294), .A(n7027), .B(
        n7026), .ZN(P2_U3220) );
  INV_X1 U8246 ( .A(n7028), .ZN(n7031) );
  INV_X1 U8247 ( .A(n7029), .ZN(n7030) );
  NAND2_X1 U8248 ( .A1(n7031), .A2(n7030), .ZN(n7032) );
  INV_X1 U8249 ( .A(n7043), .ZN(n7041) );
  NAND2_X1 U8250 ( .A1(n9811), .A2(n9160), .ZN(n7038) );
  AOI22_X1 U8251 ( .A1(n8421), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8320), .B2(
        n10731), .ZN(n7036) );
  NAND2_X1 U8252 ( .A1(n7034), .A2(n8546), .ZN(n7035) );
  NAND2_X1 U8253 ( .A1(n7036), .A2(n7035), .ZN(n7158) );
  NAND2_X1 U8254 ( .A1(n7158), .A2(n9133), .ZN(n7037) );
  NAND2_X1 U8255 ( .A1(n7038), .A2(n7037), .ZN(n7039) );
  XNOR2_X1 U8256 ( .A(n7039), .B(n9157), .ZN(n7042) );
  INV_X1 U8257 ( .A(n7042), .ZN(n7040) );
  NAND2_X1 U8258 ( .A1(n7041), .A2(n7040), .ZN(n7061) );
  NAND2_X1 U8259 ( .A1(n7043), .A2(n7042), .ZN(n7060) );
  NAND2_X1 U8260 ( .A1(n7061), .A2(n7060), .ZN(n7044) );
  AOI22_X1 U8261 ( .A1(n9811), .A2(n9159), .B1(n9143), .B2(n7158), .ZN(n7059)
         );
  XNOR2_X1 U8262 ( .A(n7044), .B(n7059), .ZN(n7056) );
  INV_X1 U8263 ( .A(n7158), .ZN(n10913) );
  NAND2_X1 U8264 ( .A1(n8401), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U8265 ( .A1(n6834), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7049) );
  OAI21_X1 U8266 ( .B1(n7045), .B2(P1_REG3_REG_6__SCAN_IN), .A(n7074), .ZN(
        n7121) );
  INV_X1 U8267 ( .A(n7121), .ZN(n7046) );
  NAND2_X1 U8268 ( .A1(n5026), .A2(n7046), .ZN(n7048) );
  NAND2_X1 U8269 ( .A1(n5024), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7047) );
  NAND4_X1 U8270 ( .A1(n7050), .A2(n7049), .A3(n7048), .A4(n7047), .ZN(n9810)
         );
  NAND2_X1 U8271 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10741) );
  INV_X1 U8272 ( .A(n10741), .ZN(n7052) );
  NOR2_X1 U8273 ( .A1(n9793), .A2(n7092), .ZN(n7051) );
  AOI211_X1 U8274 ( .C1(n9791), .C2(n9810), .A(n7052), .B(n7051), .ZN(n7053)
         );
  OAI21_X1 U8275 ( .B1(n10913), .B2(n9799), .A(n7053), .ZN(n7054) );
  AOI21_X1 U8276 ( .B1(n7151), .B2(n9796), .A(n7054), .ZN(n7055) );
  OAI21_X1 U8277 ( .B1(n7056), .B2(n9785), .A(n7055), .ZN(P1_U3225) );
  INV_X1 U8278 ( .A(n8144), .ZN(n7057) );
  NAND2_X1 U8279 ( .A1(n6989), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7125) );
  XNOR2_X1 U8280 ( .A(n7125), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8145) );
  INV_X1 U8281 ( .A(n8145), .ZN(n7809) );
  OAI222_X1 U8282 ( .A1(n10144), .A2(n10516), .B1(n8024), .B2(n7057), .C1(
        P1_U3084), .C2(n7809), .ZN(P1_U3337) );
  INV_X1 U8283 ( .A(n9349), .ZN(n9357) );
  OAI222_X1 U8284 ( .A1(n9687), .A2(n7058), .B1(n9684), .B2(n7057), .C1(n9357), 
        .C2(n9691), .ZN(P2_U3342) );
  NAND2_X1 U8285 ( .A1(n7060), .A2(n7059), .ZN(n7062) );
  NAND2_X1 U8286 ( .A1(n7062), .A2(n7061), .ZN(n7208) );
  AOI22_X1 U8287 ( .A1(n8421), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8320), .B2(
        n10682), .ZN(n7064) );
  NAND2_X1 U8288 ( .A1(n10935), .A2(n9133), .ZN(n7067) );
  NAND2_X1 U8289 ( .A1(n9810), .A2(n9160), .ZN(n7066) );
  NAND2_X1 U8290 ( .A1(n7067), .A2(n7066), .ZN(n7068) );
  XNOR2_X1 U8291 ( .A(n7068), .B(n9152), .ZN(n7211) );
  NAND2_X1 U8292 ( .A1(n10935), .A2(n9160), .ZN(n7070) );
  NAND2_X1 U8293 ( .A1(n9810), .A2(n9159), .ZN(n7069) );
  NAND2_X1 U8294 ( .A1(n7070), .A2(n7069), .ZN(n7209) );
  XNOR2_X1 U8295 ( .A(n7211), .B(n7209), .ZN(n7207) );
  XOR2_X1 U8296 ( .A(n7071), .B(n7207), .Z(n7084) );
  NAND2_X1 U8297 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10691) );
  INV_X1 U8298 ( .A(n10691), .ZN(n7072) );
  AOI21_X1 U8299 ( .B1(n9758), .B2(n9811), .A(n7072), .ZN(n7081) );
  NAND2_X1 U8300 ( .A1(n8401), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7079) );
  NAND2_X1 U8301 ( .A1(n5024), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7078) );
  AND2_X1 U8302 ( .A1(n7074), .A2(n7073), .ZN(n7075) );
  NOR2_X1 U8303 ( .A1(n7217), .A2(n7075), .ZN(n7215) );
  NAND2_X1 U8304 ( .A1(n5026), .A2(n7215), .ZN(n7077) );
  NAND2_X1 U8305 ( .A1(n6834), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7076) );
  NAND4_X1 U8306 ( .A1(n7079), .A2(n7078), .A3(n7077), .A4(n7076), .ZN(n9809)
         );
  NAND2_X1 U8307 ( .A1(n9791), .A2(n9809), .ZN(n7080) );
  OAI211_X1 U8308 ( .C1(n9760), .C2(n7121), .A(n7081), .B(n7080), .ZN(n7082)
         );
  AOI21_X1 U8309 ( .B1(n10935), .B2(n9773), .A(n7082), .ZN(n7083) );
  OAI21_X1 U8310 ( .B1(n7084), .B2(n9785), .A(n7083), .ZN(P1_U3237) );
  AND2_X1 U8311 ( .A1(n6640), .A2(n7191), .ZN(n7187) );
  INV_X1 U8312 ( .A(n10863), .ZN(n7106) );
  NAND2_X1 U8313 ( .A1(n7106), .A2(n10842), .ZN(n7087) );
  NAND2_X1 U8314 ( .A1(n7088), .A2(n7087), .ZN(n10861) );
  INV_X1 U8315 ( .A(n7108), .ZN(n10860) );
  NAND2_X1 U8316 ( .A1(n10861), .A2(n10860), .ZN(n7091) );
  NAND2_X1 U8317 ( .A1(n7175), .A2(n10880), .ZN(n7090) );
  NAND2_X1 U8318 ( .A1(n7091), .A2(n7090), .ZN(n7271) );
  XNOR2_X1 U8319 ( .A(n10862), .B(n7275), .ZN(n8749) );
  INV_X1 U8320 ( .A(n8749), .ZN(n7277) );
  NAND2_X1 U8321 ( .A1(n7092), .A2(n10894), .ZN(n7093) );
  NAND2_X1 U8322 ( .A1(n7104), .A2(n7158), .ZN(n8589) );
  NAND2_X1 U8323 ( .A1(n9811), .A2(n10913), .ZN(n7110) );
  NAND2_X1 U8324 ( .A1(n9811), .A2(n7158), .ZN(n7095) );
  INV_X1 U8325 ( .A(n9810), .ZN(n7285) );
  NAND2_X1 U8326 ( .A1(n7285), .A2(n10935), .ZN(n8588) );
  INV_X1 U8327 ( .A(n10935), .ZN(n7286) );
  NAND2_X1 U8328 ( .A1(n7286), .A2(n9810), .ZN(n8591) );
  OAI21_X1 U8329 ( .B1(n7097), .B2(n7096), .A(n7287), .ZN(n7117) );
  INV_X1 U8330 ( .A(n7117), .ZN(n10939) );
  NOR2_X1 U8331 ( .A1(n7098), .A2(n10666), .ZN(n7099) );
  NAND2_X1 U8332 ( .A1(n7100), .A2(n7099), .ZN(n7155) );
  NAND2_X2 U8333 ( .A1(n7155), .A2(n10879), .ZN(n11019) );
  OR2_X1 U8334 ( .A1(n7101), .A2(n9926), .ZN(n7149) );
  INV_X1 U8335 ( .A(n7149), .ZN(n7102) );
  NAND2_X1 U8336 ( .A1(n11019), .A2(n7102), .ZN(n10042) );
  INV_X1 U8337 ( .A(n7103), .ZN(n11062) );
  INV_X1 U8338 ( .A(n9809), .ZN(n7288) );
  INV_X1 U8339 ( .A(n10993), .ZN(n10028) );
  OAI22_X1 U8340 ( .A1(n7288), .A2(n10030), .B1(n7104), .B2(n10028), .ZN(n7116) );
  NAND2_X1 U8341 ( .A1(n7174), .A2(n7197), .ZN(n7105) );
  NAND2_X1 U8342 ( .A1(n7106), .A2(n7183), .ZN(n8577) );
  NOR2_X1 U8343 ( .A1(n10862), .A2(n10894), .ZN(n8582) );
  NAND2_X1 U8344 ( .A1(n10862), .A2(n10894), .ZN(n7159) );
  AND2_X1 U8345 ( .A1(n7110), .A2(n7159), .ZN(n8586) );
  NAND2_X1 U8346 ( .A1(n8628), .A2(n8751), .ZN(n7300) );
  NAND3_X1 U8347 ( .A1(n7111), .A2(n8589), .A3(n7096), .ZN(n7114) );
  AND2_X1 U8348 ( .A1(n6636), .A2(n8801), .ZN(n8806) );
  INV_X1 U8349 ( .A(n8806), .ZN(n7113) );
  OR2_X1 U8350 ( .A1(n8805), .A2(n9926), .ZN(n7112) );
  INV_X1 U8351 ( .A(n10998), .ZN(n10867) );
  AOI21_X1 U8352 ( .B1(n7300), .B2(n7114), .A(n10867), .ZN(n7115) );
  AOI211_X1 U8353 ( .C1(n7117), .C2(n11062), .A(n7116), .B(n7115), .ZN(n10938)
         );
  MUX2_X1 U8354 ( .A(n6529), .B(n10938), .S(n11019), .Z(n7124) );
  NAND2_X1 U8355 ( .A1(n10824), .A2(n7118), .ZN(n7192) );
  AOI21_X1 U8356 ( .B1(n10935), .B2(n7154), .A(n7338), .ZN(n10936) );
  NOR2_X1 U8357 ( .A1(n7153), .A2(n8524), .ZN(n7119) );
  OAI22_X1 U8358 ( .A1(n11016), .A2(n7286), .B1(n7121), .B2(n10879), .ZN(n7122) );
  AOI21_X1 U8359 ( .B1(n10936), .B2(n11009), .A(n7122), .ZN(n7123) );
  OAI211_X1 U8360 ( .C1(n10939), .C2(n10042), .A(n7124), .B(n7123), .ZN(
        P1_U3285) );
  INV_X1 U8361 ( .A(n8247), .ZN(n7130) );
  NAND2_X1 U8362 ( .A1(n7125), .A2(n10565), .ZN(n7126) );
  NAND2_X1 U8363 ( .A1(n7126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7127) );
  OR2_X1 U8364 ( .A1(n7127), .A2(n10572), .ZN(n7128) );
  NAND2_X1 U8365 ( .A1(n7127), .A2(n10572), .ZN(n7412) );
  INV_X1 U8366 ( .A(n9843), .ZN(n8116) );
  INV_X1 U8367 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10517) );
  OAI222_X1 U8368 ( .A1(n8024), .A2(n7130), .B1(n8116), .B2(P1_U3084), .C1(
        n10517), .C2(n10144), .ZN(P1_U3336) );
  INV_X1 U8369 ( .A(n9368), .ZN(n9373) );
  INV_X1 U8370 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7129) );
  OAI222_X1 U8371 ( .A1(P2_U3152), .A2(n9373), .B1(n9684), .B2(n7130), .C1(
        n7129), .C2(n9687), .ZN(P2_U3341) );
  NAND2_X1 U8372 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7907) );
  INV_X1 U8373 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7131) );
  MUX2_X1 U8374 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7131), .S(n7878), .Z(n7135)
         );
  OR2_X1 U8375 ( .A1(n7635), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U8376 ( .A1(n7133), .A2(n7132), .ZN(n7134) );
  NAND2_X1 U8377 ( .A1(n7134), .A2(n7135), .ZN(n7318) );
  OAI21_X1 U8378 ( .B1(n7135), .B2(n7134), .A(n7318), .ZN(n7136) );
  NAND2_X1 U8379 ( .A1(n10815), .A2(n7136), .ZN(n7137) );
  OAI211_X1 U8380 ( .C1(n10809), .C2(n7138), .A(n7907), .B(n7137), .ZN(n7144)
         );
  AOI21_X1 U8381 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7635), .A(n7139), .ZN(
        n7142) );
  NAND2_X1 U8382 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7878), .ZN(n7140) );
  OAI21_X1 U8383 ( .B1(n7878), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7140), .ZN(
        n7141) );
  NOR2_X1 U8384 ( .A1(n7142), .A2(n7141), .ZN(n7325) );
  AOI211_X1 U8385 ( .C1(n7142), .C2(n7141), .A(n10808), .B(n7325), .ZN(n7143)
         );
  AOI211_X1 U8386 ( .C1(n10813), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7144), .B(
        n7143), .ZN(n7145) );
  INV_X1 U8387 ( .A(n7145), .ZN(P1_U3254) );
  INV_X1 U8388 ( .A(n7146), .ZN(n7147) );
  AOI21_X1 U8389 ( .B1(n8750), .B2(n7148), .A(n7147), .ZN(n10916) );
  INV_X1 U8390 ( .A(n10916), .ZN(n7167) );
  NAND2_X1 U8391 ( .A1(n7103), .A2(n7149), .ZN(n7150) );
  INV_X1 U8392 ( .A(n7151), .ZN(n7152) );
  OAI22_X1 U8393 ( .A1(n11019), .A2(n6541), .B1(n7152), .B2(n10879), .ZN(n7157) );
  OAI211_X1 U8394 ( .C1(n5215), .C2(n10913), .A(n10968), .B(n7154), .ZN(n10912) );
  NOR2_X1 U8395 ( .A1(n7155), .A2(n9850), .ZN(n10005) );
  INV_X1 U8396 ( .A(n10005), .ZN(n7979) );
  NOR2_X1 U8397 ( .A1(n10912), .A2(n7979), .ZN(n7156) );
  AOI211_X1 U8398 ( .C1(n9863), .C2(n7158), .A(n7157), .B(n7156), .ZN(n7166)
         );
  NAND2_X1 U8399 ( .A1(n7160), .A2(n7159), .ZN(n7161) );
  XNOR2_X1 U8400 ( .A(n7161), .B(n7094), .ZN(n7162) );
  NAND2_X1 U8401 ( .A1(n7162), .A2(n10998), .ZN(n7164) );
  AOI22_X1 U8402 ( .A1(n10993), .A2(n10862), .B1(n9810), .B2(n10990), .ZN(
        n7163) );
  NAND2_X1 U8403 ( .A1(n7164), .A2(n7163), .ZN(n10914) );
  NAND2_X1 U8404 ( .A1(n10914), .A2(n11019), .ZN(n7165) );
  OAI211_X1 U8405 ( .C1(n7167), .C2(n10025), .A(n7166), .B(n7165), .ZN(
        P1_U3286) );
  INV_X1 U8406 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U8407 ( .A1(n10879), .A2(n6656), .ZN(n7168) );
  OAI21_X1 U8408 ( .B1(n7169), .B2(n7168), .A(n11019), .ZN(n7171) );
  OAI21_X1 U8409 ( .B1(n9863), .B2(n11009), .A(n7191), .ZN(n7170) );
  OAI211_X1 U8410 ( .C1(n9818), .C2(n11019), .A(n7171), .B(n7170), .ZN(
        P1_U3291) );
  XNOR2_X1 U8411 ( .A(n7173), .B(n7172), .ZN(n10841) );
  XNOR2_X1 U8412 ( .A(n8581), .B(n7173), .ZN(n7177) );
  OAI22_X1 U8413 ( .A1(n7175), .A2(n10030), .B1(n7174), .B2(n10028), .ZN(n7176) );
  AOI21_X1 U8414 ( .B1(n7177), .B2(n10998), .A(n7176), .ZN(n7178) );
  OAI21_X1 U8415 ( .B1(n10841), .B2(n7103), .A(n7178), .ZN(n10844) );
  NAND2_X1 U8416 ( .A1(n10844), .A2(n11019), .ZN(n7185) );
  OAI22_X1 U8417 ( .A1(n11019), .A2(n6533), .B1(n10820), .B2(n10879), .ZN(
        n7182) );
  INV_X1 U8418 ( .A(n7192), .ZN(n7180) );
  INV_X1 U8419 ( .A(n10868), .ZN(n7179) );
  OAI21_X1 U8420 ( .B1(n10842), .B2(n7180), .A(n7179), .ZN(n10843) );
  INV_X1 U8421 ( .A(n11009), .ZN(n9866) );
  NOR2_X1 U8422 ( .A1(n10843), .A2(n9866), .ZN(n7181) );
  AOI211_X1 U8423 ( .C1(n9863), .C2(n7183), .A(n7182), .B(n7181), .ZN(n7184)
         );
  OAI211_X1 U8424 ( .C1(n10841), .C2(n10042), .A(n7185), .B(n7184), .ZN(
        P1_U3289) );
  INV_X1 U8425 ( .A(n7186), .ZN(n8748) );
  XNOR2_X1 U8426 ( .A(n8748), .B(n7187), .ZN(n10821) );
  OAI21_X1 U8427 ( .B1(n7189), .B2(n7186), .A(n7188), .ZN(n7190) );
  INV_X1 U8428 ( .A(n10823), .ZN(n7196) );
  AOI21_X1 U8429 ( .B1(n7191), .B2(n7197), .A(n11111), .ZN(n7193) );
  NAND2_X1 U8430 ( .A1(n7193), .A2(n7192), .ZN(n10822) );
  OAI22_X1 U8431 ( .A1(n10822), .A2(n9850), .B1(n7194), .B2(n10879), .ZN(n7195) );
  OAI21_X1 U8432 ( .B1(n7196), .B2(n7195), .A(n11019), .ZN(n7199) );
  AOI22_X1 U8433 ( .A1(n9863), .A2(n7197), .B1(n11014), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7198) );
  OAI211_X1 U8434 ( .C1(n10025), .C2(n10821), .A(n7199), .B(n7198), .ZN(
        P1_U3290) );
  OR2_X1 U8435 ( .A1(n7200), .A2(n8447), .ZN(n7203) );
  AOI22_X1 U8436 ( .A1(n8421), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8320), .B2(
        n7201), .ZN(n7202) );
  NAND2_X1 U8437 ( .A1(n7289), .A2(n9133), .ZN(n7205) );
  NAND2_X1 U8438 ( .A1(n9809), .A2(n9143), .ZN(n7204) );
  NAND2_X1 U8439 ( .A1(n7205), .A2(n7204), .ZN(n7206) );
  XNOR2_X1 U8440 ( .A(n7206), .B(n9157), .ZN(n7434) );
  AOI22_X1 U8441 ( .A1(n7289), .A2(n9160), .B1(n9159), .B2(n9809), .ZN(n7435)
         );
  XNOR2_X1 U8442 ( .A(n7434), .B(n7435), .ZN(n7214) );
  INV_X1 U8443 ( .A(n7209), .ZN(n7210) );
  NAND2_X1 U8444 ( .A1(n7211), .A2(n7210), .ZN(n7212) );
  OAI21_X1 U8445 ( .B1(n7214), .B2(n7213), .A(n7438), .ZN(n7227) );
  INV_X1 U8446 ( .A(n7289), .ZN(n10952) );
  NOR2_X1 U8447 ( .A1(n10952), .A2(n9799), .ZN(n7226) );
  INV_X1 U8448 ( .A(n7215), .ZN(n7339) );
  AOI21_X1 U8449 ( .B1(n9758), .B2(n9810), .A(n7216), .ZN(n7224) );
  NAND2_X1 U8450 ( .A1(n5024), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7222) );
  NAND2_X1 U8451 ( .A1(n8401), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7221) );
  OR2_X1 U8452 ( .A1(n7217), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7218) );
  AND2_X1 U8453 ( .A1(n7303), .A2(n7218), .ZN(n7445) );
  NAND2_X1 U8454 ( .A1(n5026), .A2(n7445), .ZN(n7220) );
  NAND2_X1 U8455 ( .A1(n6834), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7219) );
  NAND2_X1 U8456 ( .A1(n9791), .A2(n10992), .ZN(n7223) );
  OAI211_X1 U8457 ( .C1(n9760), .C2(n7339), .A(n7224), .B(n7223), .ZN(n7225)
         );
  AOI211_X1 U8458 ( .C1(n7227), .C2(n9787), .A(n7226), .B(n7225), .ZN(n7228)
         );
  INV_X1 U8459 ( .A(n7228), .ZN(P1_U3211) );
  INV_X1 U8460 ( .A(n7253), .ZN(n10836) );
  NAND2_X1 U8461 ( .A1(n7242), .A2(n8890), .ZN(n8885) );
  XNOR2_X1 U8462 ( .A(n7230), .B(n8885), .ZN(n10830) );
  NOR2_X1 U8463 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  NAND2_X1 U8464 ( .A1(n7234), .A2(n7233), .ZN(n7238) );
  NAND3_X1 U8465 ( .A1(n8307), .A2(n9555), .A3(n8891), .ZN(n7256) );
  NAND2_X1 U8466 ( .A1(n8275), .A2(n7256), .ZN(n10919) );
  INV_X1 U8467 ( .A(n9554), .ZN(n10927) );
  NOR2_X1 U8468 ( .A1(n8307), .A2(n9034), .ZN(n10924) );
  NOR2_X1 U8469 ( .A1(n9568), .A2(n10836), .ZN(n7241) );
  NOR2_X2 U8470 ( .A1(n7238), .A2(n7237), .ZN(n9579) );
  INV_X1 U8471 ( .A(n9579), .ZN(n9398) );
  AND2_X1 U8472 ( .A1(n7375), .A2(n7253), .ZN(n10831) );
  NOR3_X1 U8473 ( .A1(n9398), .A2(n7258), .A3(n10831), .ZN(n7240) );
  AOI211_X1 U8474 ( .C1(n10927), .C2(P2_REG3_REG_1__SCAN_IN), .A(n7241), .B(
        n7240), .ZN(n7252) );
  INV_X1 U8475 ( .A(n8890), .ZN(n7246) );
  INV_X1 U8476 ( .A(n7243), .ZN(n7244) );
  NAND2_X1 U8477 ( .A1(n8885), .A2(n7244), .ZN(n7245) );
  OAI211_X1 U8478 ( .C1(n7262), .C2(n7246), .A(n7245), .B(n9576), .ZN(n7249)
         );
  OAI22_X1 U8479 ( .A1(n7254), .A2(n9548), .B1(n9332), .B2(n9550), .ZN(n7247)
         );
  INV_X1 U8480 ( .A(n7247), .ZN(n7248) );
  AND2_X1 U8481 ( .A1(n7249), .A2(n7248), .ZN(n10835) );
  MUX2_X1 U8482 ( .A(n10835), .B(n7250), .S(n9566), .Z(n7251) );
  OAI211_X1 U8483 ( .C1(n10830), .C2(n9581), .A(n7252), .B(n7251), .ZN(
        P2_U3295) );
  XNOR2_X1 U8484 ( .A(n7354), .B(n7263), .ZN(n10851) );
  INV_X1 U8485 ( .A(n7256), .ZN(n7257) );
  AND2_X1 U8486 ( .A1(n10933), .A2(n7257), .ZN(n8286) );
  INV_X1 U8487 ( .A(n8286), .ZN(n7776) );
  NOR2_X1 U8488 ( .A1(n9568), .A2(n10852), .ZN(n7261) );
  OAI21_X1 U8489 ( .B1(n7258), .B2(n10852), .A(n7385), .ZN(n10853) );
  OAI22_X1 U8490 ( .A1(n9398), .A2(n10853), .B1(n7259), .B2(n9554), .ZN(n7260)
         );
  AOI211_X1 U8491 ( .C1(n9541), .C2(P2_REG2_REG_2__SCAN_IN), .A(n7261), .B(
        n7260), .ZN(n7270) );
  INV_X1 U8492 ( .A(n7353), .ZN(n7263) );
  OAI21_X1 U8493 ( .B1(n7264), .B2(n7263), .A(n8889), .ZN(n7267) );
  OAI22_X1 U8494 ( .A1(n10605), .A2(n9550), .B1(n7265), .B2(n9548), .ZN(n7266)
         );
  AOI21_X1 U8495 ( .B1(n7267), .B2(n9576), .A(n7266), .ZN(n7268) );
  OAI21_X1 U8496 ( .B1(n10851), .B2(n8275), .A(n7268), .ZN(n10854) );
  NAND2_X1 U8497 ( .A1(n10854), .A2(n10933), .ZN(n7269) );
  OAI211_X1 U8498 ( .C1(n10851), .C2(n7776), .A(n7270), .B(n7269), .ZN(
        P2_U3294) );
  XNOR2_X1 U8499 ( .A(n7271), .B(n7277), .ZN(n10893) );
  INV_X1 U8500 ( .A(n10042), .ZN(n11010) );
  NAND2_X1 U8501 ( .A1(n10870), .A2(n7275), .ZN(n7272) );
  NAND2_X1 U8502 ( .A1(n7273), .A2(n7272), .ZN(n10895) );
  AOI22_X1 U8503 ( .A1(n9863), .A2(n7275), .B1(n11012), .B2(n7274), .ZN(n7276)
         );
  OAI21_X1 U8504 ( .B1(n10895), .B2(n9866), .A(n7276), .ZN(n7283) );
  XNOR2_X1 U8505 ( .A(n7278), .B(n7277), .ZN(n7281) );
  NAND2_X1 U8506 ( .A1(n10893), .A2(n11062), .ZN(n7280) );
  AOI22_X1 U8507 ( .A1(n10993), .A2(n5603), .B1(n9811), .B2(n10990), .ZN(n7279) );
  OAI211_X1 U8508 ( .C1(n10867), .C2(n7281), .A(n7280), .B(n7279), .ZN(n10898)
         );
  MUX2_X1 U8509 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10898), .S(n11019), .Z(n7282) );
  AOI211_X1 U8510 ( .C1(n10893), .C2(n11010), .A(n7283), .B(n7282), .ZN(n7284)
         );
  INV_X1 U8511 ( .A(n7284), .ZN(P1_U3287) );
  NAND2_X1 U8512 ( .A1(n7286), .A2(n7285), .ZN(n8634) );
  OR2_X1 U8513 ( .A1(n7288), .A2(n7289), .ZN(n8632) );
  NAND2_X1 U8514 ( .A1(n8632), .A2(n8639), .ZN(n8754) );
  INV_X1 U8515 ( .A(n7297), .ZN(n7296) );
  NAND2_X1 U8516 ( .A1(n7290), .A2(n8546), .ZN(n7294) );
  AOI22_X1 U8517 ( .A1(n8421), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8320), .B2(
        n7292), .ZN(n7293) );
  INV_X1 U8518 ( .A(n10992), .ZN(n7295) );
  NAND2_X1 U8519 ( .A1(n10967), .A2(n7295), .ZN(n10996) );
  NAND2_X1 U8520 ( .A1(n8638), .A2(n10996), .ZN(n8753) );
  INV_X1 U8521 ( .A(n8753), .ZN(n7298) );
  NAND2_X1 U8522 ( .A1(n7297), .A2(n7298), .ZN(n7299) );
  NAND2_X1 U8523 ( .A1(n7532), .A2(n7299), .ZN(n10971) );
  AND2_X2 U8524 ( .A1(n7300), .A2(n8588), .ZN(n8780) );
  INV_X1 U8525 ( .A(n8632), .ZN(n7301) );
  XNOR2_X1 U8526 ( .A(n7494), .B(n8753), .ZN(n7311) );
  OR2_X1 U8527 ( .A1(n10971), .A2(n7103), .ZN(n7310) );
  NAND2_X1 U8528 ( .A1(n8401), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7308) );
  NAND2_X1 U8529 ( .A1(n6834), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7307) );
  NAND2_X1 U8530 ( .A1(n7303), .A2(n7302), .ZN(n7304) );
  AND2_X1 U8531 ( .A1(n7505), .A2(n7304), .ZN(n11013) );
  NAND2_X1 U8532 ( .A1(n5026), .A2(n11013), .ZN(n7306) );
  NAND2_X1 U8533 ( .A1(n5024), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7305) );
  NAND4_X1 U8534 ( .A1(n7308), .A2(n7307), .A3(n7306), .A4(n7305), .ZN(n9808)
         );
  AOI22_X1 U8535 ( .A1(n10993), .A2(n9809), .B1(n9808), .B2(n10990), .ZN(n7309) );
  OAI211_X1 U8536 ( .C1(n10867), .C2(n7311), .A(n7310), .B(n7309), .ZN(n10973)
         );
  NAND2_X1 U8537 ( .A1(n10973), .A2(n11019), .ZN(n7316) );
  NAND2_X1 U8538 ( .A1(n7338), .A2(n10952), .ZN(n7337) );
  OR2_X1 U8539 ( .A1(n7337), .A2(n10967), .ZN(n10988) );
  NAND2_X1 U8540 ( .A1(n7337), .A2(n10967), .ZN(n7312) );
  AND2_X1 U8541 ( .A1(n10988), .A2(n7312), .ZN(n10969) );
  AOI22_X1 U8542 ( .A1(n11014), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7445), .B2(
        n11012), .ZN(n7313) );
  OAI21_X1 U8543 ( .B1(n5187), .B2(n11016), .A(n7313), .ZN(n7314) );
  AOI21_X1 U8544 ( .B1(n10969), .B2(n11009), .A(n7314), .ZN(n7315) );
  OAI211_X1 U8545 ( .C1(n10971), .C2(n10042), .A(n7316), .B(n7315), .ZN(
        P1_U3283) );
  OR2_X1 U8546 ( .A1(n7878), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7317) );
  NAND2_X1 U8547 ( .A1(n7318), .A2(n7317), .ZN(n7321) );
  INV_X1 U8548 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7319) );
  MUX2_X1 U8549 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7319), .S(n7960), .Z(n7320)
         );
  NAND2_X1 U8550 ( .A1(n7320), .A2(n7321), .ZN(n7621) );
  OAI21_X1 U8551 ( .B1(n7321), .B2(n7320), .A(n7621), .ZN(n7332) );
  INV_X1 U8552 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U8553 ( .A1(n10744), .A2(n7960), .ZN(n7323) );
  NAND2_X1 U8554 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7322) );
  OAI211_X1 U8555 ( .C1(n10697), .C2(n7324), .A(n7323), .B(n7322), .ZN(n7331)
         );
  AOI21_X1 U8556 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7878), .A(n7325), .ZN(
        n7327) );
  NOR2_X1 U8557 ( .A1(n7960), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7326) );
  AOI21_X1 U8558 ( .B1(n7960), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7326), .ZN(
        n7328) );
  OR2_X1 U8559 ( .A1(n7327), .A2(n7328), .ZN(n7329) );
  AOI21_X1 U8560 ( .B1(n7329), .B2(n7624), .A(n10808), .ZN(n7330) );
  AOI211_X1 U8561 ( .C1(n10815), .C2(n7332), .A(n7331), .B(n7330), .ZN(n7333)
         );
  INV_X1 U8562 ( .A(n7333), .ZN(P1_U3255) );
  XOR2_X1 U8563 ( .A(n7334), .B(n8754), .Z(n10953) );
  XNOR2_X1 U8564 ( .A(n8780), .B(n8754), .ZN(n7335) );
  MUX2_X1 U8565 ( .A(n7336), .B(n10951), .S(n11019), .Z(n7343) );
  OAI211_X1 U8566 ( .C1(n7338), .C2(n10952), .A(n7337), .B(n10968), .ZN(n10950) );
  INV_X1 U8567 ( .A(n10950), .ZN(n7341) );
  OAI22_X1 U8568 ( .A1(n10952), .A2(n11016), .B1(n7339), .B2(n10879), .ZN(
        n7340) );
  AOI21_X1 U8569 ( .B1(n7341), .B2(n10005), .A(n7340), .ZN(n7342) );
  OAI211_X1 U8570 ( .C1(n10025), .C2(n10953), .A(n7343), .B(n7342), .ZN(
        P1_U3284) );
  NAND2_X1 U8571 ( .A1(n8889), .A2(n8897), .ZN(n7380) );
  XNOR2_X1 U8572 ( .A(n7347), .B(n10886), .ZN(n8862) );
  NAND2_X1 U8573 ( .A1(n7380), .A2(n8896), .ZN(n7345) );
  NAND2_X1 U8574 ( .A1(n7381), .A2(n10904), .ZN(n8908) );
  INV_X2 U8575 ( .A(n10904), .ZN(n10610) );
  NAND2_X1 U8576 ( .A1(n9054), .A2(n10610), .ZN(n8903) );
  NAND2_X1 U8577 ( .A1(n8908), .A2(n8903), .ZN(n8858) );
  NAND2_X1 U8578 ( .A1(n10605), .A2(n8898), .ZN(n7346) );
  AND2_X1 U8579 ( .A1(n8858), .A2(n7346), .ZN(n7344) );
  NAND2_X1 U8580 ( .A1(n7345), .A2(n7344), .ZN(n7466) );
  NAND2_X1 U8581 ( .A1(n7466), .A2(n9576), .ZN(n7350) );
  AOI21_X1 U8582 ( .B1(n7345), .B2(n7346), .A(n8858), .ZN(n7349) );
  INV_X1 U8583 ( .A(n8486), .ZN(n10612) );
  AOI22_X1 U8584 ( .A1(n10612), .A2(n9574), .B1(n9572), .B2(n7347), .ZN(n7348)
         );
  OAI21_X1 U8585 ( .B1(n7350), .B2(n7349), .A(n7348), .ZN(n10906) );
  INV_X1 U8586 ( .A(n10906), .ZN(n7364) );
  OAI22_X1 U8587 ( .A1(n10933), .A2(n5867), .B1(n10614), .B2(n9554), .ZN(n7352) );
  XNOR2_X1 U8588 ( .A(n7482), .B(n10610), .ZN(n10905) );
  NOR2_X1 U8589 ( .A1(n10905), .A2(n9398), .ZN(n7351) );
  AOI211_X1 U8590 ( .C1(n9542), .C2(n10610), .A(n7352), .B(n7351), .ZN(n7363)
         );
  NAND2_X1 U8591 ( .A1(n9332), .A2(n10852), .ZN(n7355) );
  NAND2_X1 U8592 ( .A1(n7356), .A2(n7355), .ZN(n7379) );
  NAND2_X1 U8593 ( .A1(n7379), .A2(n8862), .ZN(n7358) );
  NAND2_X1 U8594 ( .A1(n10605), .A2(n10886), .ZN(n7357) );
  NAND2_X1 U8595 ( .A1(n7358), .A2(n7357), .ZN(n7359) );
  AND2_X1 U8596 ( .A1(n7359), .A2(n8858), .ZN(n10903) );
  INV_X1 U8597 ( .A(n10903), .ZN(n7361) );
  INV_X1 U8598 ( .A(n9581), .ZN(n8101) );
  NAND3_X1 U8599 ( .A1(n7361), .A2(n8101), .A3(n7469), .ZN(n7362) );
  OAI211_X1 U8600 ( .C1(n7364), .C2(n9566), .A(n7363), .B(n7362), .ZN(P2_U3292) );
  AOI21_X1 U8601 ( .B1(n7366), .B2(n7365), .A(n9306), .ZN(n7368) );
  NAND2_X1 U8602 ( .A1(n7368), .A2(n7367), .ZN(n7372) );
  OAI22_X1 U8603 ( .A1(n9313), .A2(n9052), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10445), .ZN(n7370) );
  NOR2_X1 U8604 ( .A1(n9294), .A2(n7682), .ZN(n7369) );
  AOI211_X1 U8605 ( .C1(n10613), .C2(n9329), .A(n7370), .B(n7369), .ZN(n7371)
         );
  OAI211_X1 U8606 ( .C1(n7683), .C2(n9319), .A(n7372), .B(n7371), .ZN(P2_U3215) );
  OAI22_X1 U8607 ( .A1(n10933), .A2(n7373), .B1(n10485), .B2(n9554), .ZN(n7374) );
  AOI21_X1 U8608 ( .B1(n8101), .B2(n8884), .A(n7374), .ZN(n7377) );
  OAI21_X1 U8609 ( .B1(n9542), .B2(n9579), .A(n7375), .ZN(n7376) );
  OAI211_X1 U8610 ( .C1(n7378), .C2(n9541), .A(n7377), .B(n7376), .ZN(P2_U3296) );
  XNOR2_X1 U8611 ( .A(n7379), .B(n8896), .ZN(n10885) );
  OAI21_X1 U8612 ( .B1(n7380), .B2(n8896), .A(n7345), .ZN(n7383) );
  OAI22_X1 U8613 ( .A1(n7381), .A2(n9550), .B1(n9332), .B2(n9548), .ZN(n7382)
         );
  AOI21_X1 U8614 ( .B1(n7383), .B2(n9576), .A(n7382), .ZN(n7384) );
  OAI21_X1 U8615 ( .B1(n8275), .B2(n10885), .A(n7384), .ZN(n10888) );
  NAND2_X1 U8616 ( .A1(n10888), .A2(n10933), .ZN(n7390) );
  OAI22_X1 U8617 ( .A1(n10933), .A2(n6717), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9554), .ZN(n7388) );
  NAND2_X1 U8618 ( .A1(n7385), .A2(n8898), .ZN(n7386) );
  NAND2_X1 U8619 ( .A1(n7482), .A2(n7386), .ZN(n10887) );
  NOR2_X1 U8620 ( .A1(n9398), .A2(n10887), .ZN(n7387) );
  AOI211_X1 U8621 ( .C1(n9542), .C2(n8898), .A(n7388), .B(n7387), .ZN(n7389)
         );
  OAI211_X1 U8622 ( .C1(n10885), .C2(n7776), .A(n7390), .B(n7389), .ZN(
        P2_U3293) );
  INV_X1 U8623 ( .A(n10763), .ZN(n10794) );
  INV_X1 U8624 ( .A(n10796), .ZN(n8138) );
  INV_X1 U8625 ( .A(n9338), .ZN(n7394) );
  MUX2_X1 U8626 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7391), .S(n9338), .Z(n9342)
         );
  OAI21_X1 U8627 ( .B1(n7393), .B2(n6970), .A(n7392), .ZN(n9343) );
  NAND2_X1 U8628 ( .A1(n9342), .A2(n9343), .ZN(n9341) );
  OAI21_X1 U8629 ( .B1(n7394), .B2(n7391), .A(n9341), .ZN(n7397) );
  MUX2_X1 U8630 ( .A(n7395), .B(P2_REG1_REG_12__SCAN_IN), .S(n7423), .Z(n7396)
         );
  NOR2_X1 U8631 ( .A1(n7396), .A2(n7397), .ZN(n7418) );
  AOI21_X1 U8632 ( .B1(n7397), .B2(n7396), .A(n7418), .ZN(n7400) );
  NAND2_X1 U8633 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8077) );
  INV_X1 U8634 ( .A(n8077), .ZN(n7398) );
  AOI21_X1 U8635 ( .B1(n10787), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7398), .ZN(
        n7399) );
  OAI21_X1 U8636 ( .B1(n8138), .B2(n7400), .A(n7399), .ZN(n7408) );
  NOR2_X1 U8637 ( .A1(n9338), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7403) );
  AOI21_X1 U8638 ( .B1(n9338), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7403), .ZN(
        n9336) );
  NAND2_X1 U8639 ( .A1(n9335), .A2(n9336), .ZN(n9334) );
  OAI21_X1 U8640 ( .B1(n9338), .B2(P2_REG2_REG_11__SCAN_IN), .A(n9334), .ZN(
        n7406) );
  NAND2_X1 U8641 ( .A1(n7423), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7404) );
  OAI21_X1 U8642 ( .B1(n7423), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7404), .ZN(
        n7405) );
  NOR2_X1 U8643 ( .A1(n7405), .A2(n7406), .ZN(n7422) );
  AOI211_X1 U8644 ( .C1(n7406), .C2(n7405), .A(n7422), .B(n10788), .ZN(n7407)
         );
  AOI211_X1 U8645 ( .C1(n10794), .C2(n7423), .A(n7408), .B(n7407), .ZN(n7409)
         );
  INV_X1 U8646 ( .A(n7409), .ZN(P2_U3257) );
  INV_X1 U8647 ( .A(n9382), .ZN(n7411) );
  INV_X1 U8648 ( .A(n8314), .ZN(n7414) );
  OAI222_X1 U8649 ( .A1(n7411), .A2(P2_U3152), .B1(n9684), .B2(n7414), .C1(
        n9687), .C2(n7410), .ZN(P2_U3340) );
  INV_X1 U8650 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7415) );
  NAND2_X1 U8651 ( .A1(n7412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7413) );
  XNOR2_X1 U8652 ( .A(n7413), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9846) );
  INV_X1 U8653 ( .A(n9846), .ZN(n10727) );
  OAI222_X1 U8654 ( .A1(n10144), .A2(n7415), .B1(n10147), .B2(n7414), .C1(
        P1_U3084), .C2(n10727), .ZN(P1_U3335) );
  INV_X1 U8655 ( .A(n8319), .ZN(n7417) );
  OAI222_X1 U8656 ( .A1(n10144), .A2(n7416), .B1(n10147), .B2(n7417), .C1(
        P1_U3084), .C2(n9926), .ZN(P1_U3334) );
  OAI222_X1 U8657 ( .A1(P2_U3152), .A2(n10922), .B1(n9684), .B2(n7417), .C1(
        n9687), .C2(n5718), .ZN(P2_U3339) );
  AOI21_X1 U8658 ( .B1(n7419), .B2(n7395), .A(n7418), .ZN(n7421) );
  AOI22_X1 U8659 ( .A1(n7599), .A2(n6049), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7595), .ZN(n7420) );
  NOR2_X1 U8660 ( .A1(n7421), .A2(n7420), .ZN(n7594) );
  AOI21_X1 U8661 ( .B1(n7421), .B2(n7420), .A(n7594), .ZN(n7430) );
  AOI22_X1 U8662 ( .A1(n7599), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8095), .B2(
        n7595), .ZN(n7424) );
  NAND2_X1 U8663 ( .A1(n7425), .A2(n7424), .ZN(n7598) );
  OAI21_X1 U8664 ( .B1(n7425), .B2(n7424), .A(n7598), .ZN(n7426) );
  NAND2_X1 U8665 ( .A1(n7426), .A2(n10761), .ZN(n7429) );
  INV_X1 U8666 ( .A(n10787), .ZN(n10772) );
  INV_X1 U8667 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U8668 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(n9691), .ZN(n9062) );
  OAI21_X1 U8669 ( .B1(n10772), .B2(n7939), .A(n9062), .ZN(n7427) );
  AOI21_X1 U8670 ( .B1(n7599), .B2(n10794), .A(n7427), .ZN(n7428) );
  OAI211_X1 U8671 ( .C1(n7430), .C2(n8138), .A(n7429), .B(n7428), .ZN(P2_U3258) );
  NAND2_X1 U8672 ( .A1(n10967), .A2(n9133), .ZN(n7432) );
  NAND2_X1 U8673 ( .A1(n10992), .A2(n9160), .ZN(n7431) );
  NAND2_X1 U8674 ( .A1(n7432), .A2(n7431), .ZN(n7433) );
  XNOR2_X1 U8675 ( .A(n7433), .B(n9157), .ZN(n7547) );
  INV_X1 U8676 ( .A(n7434), .ZN(n7436) );
  NAND2_X1 U8677 ( .A1(n7436), .A2(n7435), .ZN(n7437) );
  AND2_X1 U8678 ( .A1(n10992), .A2(n9159), .ZN(n7439) );
  AOI21_X1 U8679 ( .B1(n10967), .B2(n9143), .A(n7439), .ZN(n7442) );
  INV_X1 U8680 ( .A(n7442), .ZN(n7440) );
  NAND2_X1 U8681 ( .A1(n7443), .A2(n7442), .ZN(n7548) );
  NAND2_X1 U8682 ( .A1(n7549), .A2(n7548), .ZN(n7444) );
  XOR2_X1 U8683 ( .A(n7547), .B(n7444), .Z(n7452) );
  INV_X1 U8684 ( .A(n7445), .ZN(n7449) );
  AOI21_X1 U8685 ( .B1(n9758), .B2(n9809), .A(n7446), .ZN(n7448) );
  NAND2_X1 U8686 ( .A1(n9791), .A2(n9808), .ZN(n7447) );
  OAI211_X1 U8687 ( .C1(n9760), .C2(n7449), .A(n7448), .B(n7447), .ZN(n7450)
         );
  AOI21_X1 U8688 ( .B1(n10967), .B2(n9773), .A(n7450), .ZN(n7451) );
  OAI21_X1 U8689 ( .B1(n7452), .B2(n9785), .A(n7451), .ZN(P1_U3219) );
  INV_X1 U8690 ( .A(n7713), .ZN(n10981) );
  INV_X1 U8691 ( .A(n7453), .ZN(n7454) );
  AOI21_X1 U8692 ( .B1(n7367), .B2(n7454), .A(n9306), .ZN(n7458) );
  NOR3_X1 U8693 ( .A1(n10607), .A2(n7455), .A3(n7559), .ZN(n7457) );
  OAI21_X1 U8694 ( .B1(n7458), .B2(n7457), .A(n7456), .ZN(n7464) );
  INV_X1 U8695 ( .A(n7563), .ZN(n7462) );
  OR2_X1 U8696 ( .A1(n7559), .A2(n9548), .ZN(n7459) );
  OAI21_X1 U8697 ( .B1(n7749), .B2(n9550), .A(n7459), .ZN(n7561) );
  INV_X1 U8698 ( .A(n7561), .ZN(n7460) );
  INV_X1 U8699 ( .A(n9251), .ZN(n7789) );
  OAI22_X1 U8700 ( .A1(n7460), .A2(n7789), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10258), .ZN(n7461) );
  AOI21_X1 U8701 ( .B1(n7462), .B2(n10616), .A(n7461), .ZN(n7463) );
  OAI211_X1 U8702 ( .C1(n10981), .C2(n9319), .A(n7464), .B(n7463), .ZN(
        P2_U3223) );
  INV_X1 U8703 ( .A(n9576), .ZN(n9546) );
  NAND2_X1 U8704 ( .A1(n9054), .A2(n10904), .ZN(n7465) );
  NAND2_X1 U8705 ( .A1(n10612), .A2(n7473), .ZN(n8911) );
  INV_X1 U8706 ( .A(n8911), .ZN(n7467) );
  NAND2_X1 U8707 ( .A1(n8486), .A2(n10925), .ZN(n8910) );
  INV_X1 U8708 ( .A(n8916), .ZN(n10943) );
  NAND2_X1 U8709 ( .A1(n9052), .A2(n10943), .ZN(n7672) );
  AND2_X1 U8710 ( .A1(n9331), .A2(n8916), .ZN(n7671) );
  INV_X1 U8711 ( .A(n7671), .ZN(n8915) );
  AND2_X1 U8712 ( .A1(n7672), .A2(n8915), .ZN(n8861) );
  XNOR2_X1 U8713 ( .A(n7558), .B(n8861), .ZN(n7468) );
  OAI222_X1 U8714 ( .A1(n9550), .A2(n7559), .B1(n9548), .B2(n8486), .C1(n9546), 
        .C2(n7468), .ZN(n10945) );
  INV_X1 U8715 ( .A(n10945), .ZN(n7479) );
  NAND2_X1 U8716 ( .A1(n8486), .A2(n7473), .ZN(n7470) );
  NAND2_X1 U8717 ( .A1(n8910), .A2(n8911), .ZN(n8857) );
  OR2_X1 U8718 ( .A1(n8857), .A2(n8486), .ZN(n7471) );
  NAND2_X1 U8719 ( .A1(n7472), .A2(n7471), .ZN(n7745) );
  XOR2_X1 U8720 ( .A(n7745), .B(n8861), .Z(n10947) );
  INV_X1 U8721 ( .A(n7564), .ZN(n7681) );
  OAI21_X1 U8722 ( .B1(n10943), .B2(n7481), .A(n7681), .ZN(n10944) );
  OAI22_X1 U8723 ( .A1(n10933), .A2(n7474), .B1(n8479), .B2(n9554), .ZN(n7475)
         );
  AOI21_X1 U8724 ( .B1(n9542), .B2(n8916), .A(n7475), .ZN(n7476) );
  OAI21_X1 U8725 ( .B1(n10944), .B2(n9398), .A(n7476), .ZN(n7477) );
  AOI21_X1 U8726 ( .B1(n10947), .B2(n8101), .A(n7477), .ZN(n7478) );
  OAI21_X1 U8727 ( .B1(n7479), .B2(n9541), .A(n7478), .ZN(P2_U3290) );
  XNOR2_X1 U8728 ( .A(n7480), .B(n8857), .ZN(n10921) );
  NOR2_X1 U8729 ( .A1(n7481), .A2(n11125), .ZN(n7484) );
  OAI21_X1 U8730 ( .B1(n7482), .B2(n10610), .A(n10925), .ZN(n7483) );
  AND2_X1 U8731 ( .A1(n7484), .A2(n7483), .ZN(n10923) );
  XNOR2_X1 U8732 ( .A(n7485), .B(n8857), .ZN(n7486) );
  NAND2_X1 U8733 ( .A1(n7486), .A2(n9576), .ZN(n7488) );
  AOI22_X1 U8734 ( .A1(n9054), .A2(n9572), .B1(n9574), .B2(n9331), .ZN(n7487)
         );
  NAND2_X1 U8735 ( .A1(n7488), .A2(n7487), .ZN(n10931) );
  AOI211_X1 U8736 ( .C1(n11066), .C2(n10925), .A(n10923), .B(n10931), .ZN(
        n7489) );
  OAI21_X1 U8737 ( .B1(n11082), .B2(n10921), .A(n7489), .ZN(n7491) );
  NAND2_X1 U8738 ( .A1(n7491), .A2(n11132), .ZN(n7490) );
  OAI21_X1 U8739 ( .B1(n11132), .B2(n6732), .A(n7490), .ZN(P2_U3525) );
  INV_X1 U8740 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7493) );
  NAND2_X1 U8741 ( .A1(n7491), .A2(n11135), .ZN(n7492) );
  OAI21_X1 U8742 ( .B1(n11135), .B2(n7493), .A(n7492), .ZN(P2_U3466) );
  NAND2_X1 U8743 ( .A1(n7495), .A2(n8546), .ZN(n7498) );
  AOI22_X1 U8744 ( .A1(n8421), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8320), .B2(
        n7496), .ZN(n7497) );
  INV_X1 U8745 ( .A(n9808), .ZN(n7499) );
  OR2_X1 U8746 ( .A1(n10987), .A2(n7499), .ZN(n8637) );
  NAND2_X1 U8747 ( .A1(n7500), .A2(n8546), .ZN(n7503) );
  AOI22_X1 U8748 ( .A1(n8421), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8320), .B2(
        n7501), .ZN(n7502) );
  NAND2_X1 U8749 ( .A1(n8401), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U8750 ( .A1(n6834), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U8751 ( .A1(n7505), .A2(n7504), .ZN(n7506) );
  AND2_X1 U8752 ( .A1(n7521), .A2(n7506), .ZN(n7660) );
  NAND2_X1 U8753 ( .A1(n5026), .A2(n7660), .ZN(n7508) );
  NAND2_X1 U8754 ( .A1(n5024), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7507) );
  NAND4_X1 U8755 ( .A1(n7510), .A2(n7509), .A3(n7508), .A4(n7507), .ZN(n10991)
         );
  INV_X1 U8756 ( .A(n10991), .ZN(n7511) );
  OR2_X1 U8757 ( .A1(n7614), .A2(n7511), .ZN(n8649) );
  NAND2_X1 U8758 ( .A1(n7614), .A2(n7511), .ZN(n8646) );
  NAND2_X1 U8759 ( .A1(n7512), .A2(n8546), .ZN(n7514) );
  AOI22_X1 U8760 ( .A1(n8421), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8320), .B2(
        n10703), .ZN(n7513) );
  NAND2_X1 U8761 ( .A1(n8541), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U8762 ( .A1(n8401), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7517) );
  XNOR2_X1 U8763 ( .A(n7521), .B(P1_REG3_REG_11__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U8764 ( .A1(n5026), .A2(n7742), .ZN(n7516) );
  NAND2_X1 U8765 ( .A1(n6834), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7515) );
  NAND4_X1 U8766 ( .A1(n7518), .A2(n7517), .A3(n7516), .A4(n7515), .ZN(n9807)
         );
  INV_X1 U8767 ( .A(n9807), .ZN(n7589) );
  NOR2_X1 U8768 ( .A1(n7738), .A2(n7589), .ZN(n8656) );
  INV_X1 U8769 ( .A(n8656), .ZN(n7643) );
  NAND2_X1 U8770 ( .A1(n7738), .A2(n7589), .ZN(n8562) );
  NAND2_X1 U8771 ( .A1(n7643), .A2(n8562), .ZN(n8758) );
  INV_X1 U8772 ( .A(n8758), .ZN(n7519) );
  XNOR2_X1 U8773 ( .A(n7642), .B(n7519), .ZN(n7520) );
  NAND2_X1 U8774 ( .A1(n7520), .A2(n10998), .ZN(n7530) );
  NAND2_X1 U8775 ( .A1(n8401), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U8776 ( .A1(n6834), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7527) );
  INV_X1 U8777 ( .A(n7521), .ZN(n7522) );
  AOI21_X1 U8778 ( .B1(n7522), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n7523) );
  OR2_X1 U8779 ( .A1(n7523), .A2(n7645), .ZN(n7843) );
  INV_X1 U8780 ( .A(n7843), .ZN(n7524) );
  NAND2_X1 U8781 ( .A1(n5026), .A2(n7524), .ZN(n7526) );
  NAND2_X1 U8782 ( .A1(n8541), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7525) );
  NAND4_X1 U8783 ( .A1(n7528), .A2(n7527), .A3(n7526), .A4(n7525), .ZN(n9806)
         );
  AOI22_X1 U8784 ( .A1(n10993), .A2(n10991), .B1(n9806), .B2(n10990), .ZN(
        n7529) );
  NAND2_X1 U8785 ( .A1(n7530), .A2(n7529), .ZN(n11040) );
  INV_X1 U8786 ( .A(n11040), .ZN(n7542) );
  NAND2_X1 U8787 ( .A1(n10967), .A2(n10992), .ZN(n7531) );
  OR2_X1 U8788 ( .A1(n10987), .A2(n9808), .ZN(n7533) );
  INV_X1 U8789 ( .A(n7609), .ZN(n7535) );
  OR2_X1 U8790 ( .A1(n7614), .A2(n10991), .ZN(n7536) );
  XNOR2_X1 U8791 ( .A(n7631), .B(n8758), .ZN(n11042) );
  INV_X1 U8792 ( .A(n10025), .ZN(n7540) );
  INV_X1 U8793 ( .A(n7614), .ZN(n7662) );
  INV_X1 U8794 ( .A(n7738), .ZN(n11038) );
  OAI21_X1 U8795 ( .B1(n7613), .B2(n11038), .A(n5097), .ZN(n11039) );
  AOI22_X1 U8796 ( .A1(n11014), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7742), .B2(
        n11012), .ZN(n7538) );
  NAND2_X1 U8797 ( .A1(n7738), .A2(n9863), .ZN(n7537) );
  OAI211_X1 U8798 ( .C1(n11039), .C2(n9866), .A(n7538), .B(n7537), .ZN(n7539)
         );
  AOI21_X1 U8799 ( .B1(n11042), .B2(n7540), .A(n7539), .ZN(n7541) );
  OAI21_X1 U8800 ( .B1(n7542), .B2(n11014), .A(n7541), .ZN(P1_U3280) );
  NAND2_X1 U8801 ( .A1(n10987), .A2(n9133), .ZN(n7544) );
  NAND2_X1 U8802 ( .A1(n9808), .A2(n9160), .ZN(n7543) );
  NAND2_X1 U8803 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  XNOR2_X1 U8804 ( .A(n7545), .B(n9152), .ZN(n7579) );
  AND2_X1 U8805 ( .A1(n9808), .A2(n9159), .ZN(n7546) );
  AOI21_X1 U8806 ( .B1(n10987), .B2(n9143), .A(n7546), .ZN(n7578) );
  XNOR2_X1 U8807 ( .A(n7579), .B(n7578), .ZN(n7576) );
  XOR2_X1 U8808 ( .A(n7576), .B(n7575), .Z(n7556) );
  INV_X1 U8809 ( .A(n11013), .ZN(n7553) );
  AOI21_X1 U8810 ( .B1(n9758), .B2(n10992), .A(n7550), .ZN(n7552) );
  NAND2_X1 U8811 ( .A1(n9791), .A2(n10991), .ZN(n7551) );
  OAI211_X1 U8812 ( .C1(n9760), .C2(n7553), .A(n7552), .B(n7551), .ZN(n7554)
         );
  AOI21_X1 U8813 ( .B1(n10987), .B2(n9773), .A(n7554), .ZN(n7555) );
  OAI21_X1 U8814 ( .B1(n7556), .B2(n9785), .A(n7555), .ZN(P1_U3229) );
  NOR2_X1 U8815 ( .A1(n9331), .A2(n10943), .ZN(n7557) );
  NAND2_X1 U8816 ( .A1(n7559), .A2(n10959), .ZN(n8920) );
  INV_X1 U8817 ( .A(n7559), .ZN(n9330) );
  NAND2_X1 U8818 ( .A1(n7719), .A2(n8921), .ZN(n7560) );
  NAND2_X1 U8819 ( .A1(n7695), .A2(n7713), .ZN(n8924) );
  NAND2_X1 U8820 ( .A1(n9329), .A2(n10981), .ZN(n8925) );
  NAND2_X1 U8821 ( .A1(n8924), .A2(n8925), .ZN(n7570) );
  XNOR2_X1 U8822 ( .A(n7560), .B(n7570), .ZN(n7562) );
  AOI21_X1 U8823 ( .B1(n7562), .B2(n9576), .A(n7561), .ZN(n10983) );
  OAI22_X1 U8824 ( .A1(n10933), .A2(n6805), .B1(n7563), .B2(n9554), .ZN(n7568)
         );
  NAND2_X1 U8825 ( .A1(n7564), .A2(n7683), .ZN(n7679) );
  AOI21_X1 U8826 ( .B1(n7679), .B2(n7713), .A(n11125), .ZN(n7565) );
  OR2_X1 U8827 ( .A1(n7679), .A2(n7713), .ZN(n7769) );
  NAND2_X1 U8828 ( .A1(n7565), .A2(n7769), .ZN(n10979) );
  AND2_X1 U8829 ( .A1(n10933), .A2(n10922), .ZN(n9467) );
  INV_X1 U8830 ( .A(n9467), .ZN(n7566) );
  NOR2_X1 U8831 ( .A1(n10979), .A2(n7566), .ZN(n7567) );
  AOI211_X1 U8832 ( .C1(n9542), .C2(n7713), .A(n7568), .B(n7567), .ZN(n7574)
         );
  INV_X1 U8833 ( .A(n8860), .ZN(n8914) );
  OR2_X1 U8834 ( .A1(n7745), .A2(n7714), .ZN(n7669) );
  INV_X1 U8835 ( .A(n7672), .ZN(n8918) );
  NAND2_X1 U8836 ( .A1(n7559), .A2(n7683), .ZN(n7569) );
  INV_X1 U8837 ( .A(n7570), .ZN(n8923) );
  NAND2_X1 U8838 ( .A1(n5099), .A2(n8923), .ZN(n10978) );
  INV_X1 U8839 ( .A(n7715), .ZN(n7572) );
  NAND2_X1 U8840 ( .A1(n7669), .A2(n7572), .ZN(n10977) );
  NAND3_X1 U8841 ( .A1(n10978), .A2(n8101), .A3(n10977), .ZN(n7573) );
  OAI211_X1 U8842 ( .C1(n10983), .C2(n9566), .A(n7574), .B(n7573), .ZN(
        P2_U3288) );
  INV_X1 U8843 ( .A(n7576), .ZN(n7577) );
  NAND2_X1 U8844 ( .A1(n7579), .A2(n7578), .ZN(n7580) );
  NAND2_X1 U8845 ( .A1(n7614), .A2(n9133), .ZN(n7583) );
  NAND2_X1 U8846 ( .A1(n10991), .A2(n9160), .ZN(n7582) );
  NAND2_X1 U8847 ( .A1(n7583), .A2(n7582), .ZN(n7584) );
  XNOR2_X1 U8848 ( .A(n7584), .B(n9152), .ZN(n7730) );
  AND2_X1 U8849 ( .A1(n10991), .A2(n9159), .ZN(n7585) );
  AOI21_X1 U8850 ( .B1(n7614), .B2(n9143), .A(n7585), .ZN(n7729) );
  XNOR2_X1 U8851 ( .A(n7730), .B(n7729), .ZN(n7586) );
  XNOR2_X1 U8852 ( .A(n7731), .B(n7586), .ZN(n7592) );
  NAND2_X1 U8853 ( .A1(n9796), .A2(n7660), .ZN(n7588) );
  AOI22_X1 U8854 ( .A1(n9758), .A2(n9808), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3084), .ZN(n7587) );
  OAI211_X1 U8855 ( .C1(n7589), .C2(n9756), .A(n7588), .B(n7587), .ZN(n7590)
         );
  AOI21_X1 U8856 ( .B1(n7614), .B2(n9773), .A(n7590), .ZN(n7591) );
  OAI21_X1 U8857 ( .B1(n7592), .B2(n9785), .A(n7591), .ZN(P1_U3215) );
  INV_X1 U8858 ( .A(n8325), .ZN(n8306) );
  OAI222_X1 U8859 ( .A1(n10147), .A2(n8306), .B1(n7593), .B2(P1_U3084), .C1(
        n10511), .C2(n10144), .ZN(P1_U3333) );
  AOI21_X1 U8860 ( .B1(n7595), .B2(n6049), .A(n7594), .ZN(n7597) );
  AOI22_X1 U8861 ( .A1(n7848), .A2(n6064), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7854), .ZN(n7596) );
  NOR2_X1 U8862 ( .A1(n7597), .A2(n7596), .ZN(n7853) );
  AOI21_X1 U8863 ( .B1(n7597), .B2(n7596), .A(n7853), .ZN(n7606) );
  AOI22_X1 U8864 ( .A1(n7848), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8040), .B2(
        n7854), .ZN(n7601) );
  OAI21_X1 U8865 ( .B1(n7599), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7598), .ZN(
        n7600) );
  NAND2_X1 U8866 ( .A1(n7601), .A2(n7600), .ZN(n7847) );
  OAI21_X1 U8867 ( .B1(n7601), .B2(n7600), .A(n7847), .ZN(n7602) );
  NAND2_X1 U8868 ( .A1(n7602), .A2(n10761), .ZN(n7605) );
  INV_X1 U8869 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U8870 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8510) );
  OAI21_X1 U8871 ( .B1(n10772), .B2(n7942), .A(n8510), .ZN(n7603) );
  AOI21_X1 U8872 ( .B1(n7848), .B2(n10794), .A(n7603), .ZN(n7604) );
  OAI211_X1 U8873 ( .C1(n7606), .C2(n8138), .A(n7605), .B(n7604), .ZN(P2_U3259) );
  INV_X1 U8874 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7617) );
  INV_X1 U8875 ( .A(n7607), .ZN(n7608) );
  AOI21_X1 U8876 ( .B1(n8756), .B2(n7609), .A(n7608), .ZN(n7663) );
  OAI21_X1 U8877 ( .B1(n8756), .B2(n7611), .A(n7610), .ZN(n7612) );
  AOI222_X1 U8878 ( .A1(n10998), .A2(n7612), .B1(n9807), .B2(n10990), .C1(
        n9808), .C2(n10993), .ZN(n7668) );
  AOI211_X1 U8879 ( .C1(n7614), .C2(n5094), .A(n11111), .B(n7613), .ZN(n7666)
         );
  AOI21_X1 U8880 ( .B1(n11053), .B2(n7614), .A(n7666), .ZN(n7615) );
  OAI211_X1 U8881 ( .C1(n7663), .C2(n10911), .A(n7668), .B(n7615), .ZN(n7618)
         );
  NAND2_X1 U8882 ( .A1(n7618), .A2(n10137), .ZN(n7616) );
  OAI21_X1 U8883 ( .B1(n10137), .B2(n7617), .A(n7616), .ZN(P1_U3484) );
  INV_X2 U8884 ( .A(n11118), .ZN(n10847) );
  NAND2_X1 U8885 ( .A1(n7618), .A2(n10847), .ZN(n7619) );
  OAI21_X1 U8886 ( .B1(n10847), .B2(n7620), .A(n7619), .ZN(P1_U3533) );
  INV_X1 U8887 ( .A(n7801), .ZN(n8051) );
  AND2_X1 U8888 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8186) );
  OAI21_X1 U8889 ( .B1(n7960), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7621), .ZN(
        n7800) );
  XNOR2_X1 U8890 ( .A(n7801), .B(n7800), .ZN(n7622) );
  INV_X1 U8891 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11119) );
  NOR2_X1 U8892 ( .A1(n11119), .A2(n7622), .ZN(n7802) );
  AOI211_X1 U8893 ( .C1(n7622), .C2(n11119), .A(n7802), .B(n10702), .ZN(n7623)
         );
  AOI211_X1 U8894 ( .C1(n10744), .C2(n8051), .A(n8186), .B(n7623), .ZN(n7629)
         );
  INV_X1 U8895 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7625) );
  AOI211_X1 U8896 ( .C1(n7626), .C2(n7625), .A(n7795), .B(n10808), .ZN(n7627)
         );
  AOI21_X1 U8897 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n10813), .A(n7627), .ZN(
        n7628) );
  NAND2_X1 U8898 ( .A1(n7629), .A2(n7628), .ZN(P1_U3256) );
  NAND2_X1 U8899 ( .A1(n7738), .A2(n9807), .ZN(n7630) );
  NAND2_X1 U8900 ( .A1(n7631), .A2(n7630), .ZN(n7633) );
  OR2_X1 U8901 ( .A1(n7738), .A2(n9807), .ZN(n7632) );
  NAND2_X1 U8902 ( .A1(n7633), .A2(n7632), .ZN(n7639) );
  INV_X1 U8903 ( .A(n7639), .ZN(n7638) );
  NAND2_X1 U8904 ( .A1(n7634), .A2(n8546), .ZN(n7637) );
  AOI22_X1 U8905 ( .A1(n8421), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8320), .B2(
        n7635), .ZN(n7636) );
  INV_X1 U8906 ( .A(n9806), .ZN(n7987) );
  NOR2_X1 U8907 ( .A1(n11054), .A2(n7987), .ZN(n8561) );
  INV_X1 U8908 ( .A(n8561), .ZN(n8665) );
  NAND2_X1 U8909 ( .A1(n11054), .A2(n7987), .ZN(n8563) );
  NAND2_X1 U8910 ( .A1(n8665), .A2(n8563), .ZN(n8760) );
  INV_X1 U8911 ( .A(n8760), .ZN(n7640) );
  NAND2_X1 U8912 ( .A1(n7638), .A2(n8760), .ZN(n7956) );
  NAND2_X1 U8913 ( .A1(n7639), .A2(n7640), .ZN(n7641) );
  NAND2_X1 U8914 ( .A1(n7956), .A2(n7641), .ZN(n11058) );
  INV_X1 U8915 ( .A(n8562), .ZN(n8657) );
  XNOR2_X1 U8916 ( .A(n7964), .B(n8760), .ZN(n7644) );
  NAND2_X1 U8917 ( .A1(n7644), .A2(n10998), .ZN(n7653) );
  NAND2_X1 U8918 ( .A1(n8401), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U8919 ( .A1(n6834), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7650) );
  OR2_X1 U8920 ( .A1(n7645), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7647) );
  AND2_X1 U8921 ( .A1(n7647), .A2(n7646), .ZN(n7994) );
  NAND2_X1 U8922 ( .A1(n5026), .A2(n7994), .ZN(n7649) );
  NAND2_X1 U8923 ( .A1(n8541), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7648) );
  NAND4_X1 U8924 ( .A1(n7651), .A2(n7650), .A3(n7649), .A4(n7648), .ZN(n9805)
         );
  AOI22_X1 U8925 ( .A1(n10993), .A2(n9807), .B1(n9805), .B2(n10990), .ZN(n7652) );
  NAND2_X1 U8926 ( .A1(n7653), .A2(n7652), .ZN(n11060) );
  NAND2_X1 U8927 ( .A1(n11060), .A2(n11019), .ZN(n7659) );
  INV_X1 U8928 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7654) );
  OAI22_X1 U8929 ( .A1(n11019), .A2(n7654), .B1(n7843), .B2(n10879), .ZN(n7657) );
  AOI21_X1 U8930 ( .B1(n5097), .B2(n11054), .A(n11111), .ZN(n7655) );
  NAND2_X1 U8931 ( .A1(n7655), .A2(n5040), .ZN(n11056) );
  NOR2_X1 U8932 ( .A1(n11056), .A2(n7979), .ZN(n7656) );
  AOI211_X1 U8933 ( .C1(n9863), .C2(n11054), .A(n7657), .B(n7656), .ZN(n7658)
         );
  OAI211_X1 U8934 ( .C1(n10025), .C2(n11058), .A(n7659), .B(n7658), .ZN(
        P1_U3279) );
  AOI22_X1 U8935 ( .A1(n11014), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7660), .B2(
        n11012), .ZN(n7661) );
  OAI21_X1 U8936 ( .B1(n7662), .B2(n11016), .A(n7661), .ZN(n7665) );
  NOR2_X1 U8937 ( .A1(n7663), .A2(n10025), .ZN(n7664) );
  AOI211_X1 U8938 ( .C1(n7666), .C2(n10005), .A(n7665), .B(n7664), .ZN(n7667)
         );
  OAI21_X1 U8939 ( .B1(n11014), .B2(n7668), .A(n7667), .ZN(P1_U3281) );
  AND2_X1 U8940 ( .A1(n7670), .A2(n7669), .ZN(n7675) );
  OR2_X1 U8941 ( .A1(n7745), .A2(n7671), .ZN(n7673) );
  NAND3_X1 U8942 ( .A1(n7673), .A2(n8914), .A3(n7672), .ZN(n7674) );
  AND2_X1 U8943 ( .A1(n7675), .A2(n7674), .ZN(n10963) );
  XNOR2_X1 U8944 ( .A(n7676), .B(n8860), .ZN(n7677) );
  AOI222_X1 U8945 ( .A1(n9576), .A2(n7677), .B1(n9331), .B2(n9572), .C1(n9329), 
        .C2(n9574), .ZN(n10962) );
  MUX2_X1 U8946 ( .A(n7678), .B(n10962), .S(n10933), .Z(n7686) );
  INV_X1 U8947 ( .A(n7679), .ZN(n7680) );
  AOI21_X1 U8948 ( .B1(n10959), .B2(n7681), .A(n7680), .ZN(n10960) );
  OAI22_X1 U8949 ( .A1(n9568), .A2(n7683), .B1(n9554), .B2(n7682), .ZN(n7684)
         );
  AOI21_X1 U8950 ( .B1(n10960), .B2(n9579), .A(n7684), .ZN(n7685) );
  OAI211_X1 U8951 ( .C1(n10963), .C2(n9581), .A(n7686), .B(n7685), .ZN(
        P2_U3289) );
  INV_X1 U8952 ( .A(n7820), .ZN(n11031) );
  AOI21_X1 U8953 ( .B1(n7688), .B2(n7687), .A(n9306), .ZN(n7690) );
  NAND2_X1 U8954 ( .A1(n7690), .A2(n7689), .ZN(n7694) );
  INV_X1 U8955 ( .A(n8073), .ZN(n9326) );
  OAI22_X1 U8956 ( .A1(n9313), .A2(n7749), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10455), .ZN(n7692) );
  NOR2_X1 U8957 ( .A1(n9294), .A2(n7766), .ZN(n7691) );
  AOI211_X1 U8958 ( .C1(n10613), .C2(n9326), .A(n7692), .B(n7691), .ZN(n7693)
         );
  OAI211_X1 U8959 ( .C1(n11031), .C2(n9319), .A(n7694), .B(n7693), .ZN(
        P2_U3219) );
  INV_X1 U8960 ( .A(n8334), .ZN(n7712) );
  INV_X1 U8961 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10510) );
  OAI222_X1 U8962 ( .A1(n8024), .A2(n7712), .B1(P1_U3084), .B2(n8795), .C1(
        n10510), .C2(n10144), .ZN(P1_U3332) );
  INV_X1 U8963 ( .A(n7456), .ZN(n7698) );
  NOR3_X1 U8964 ( .A1(n10607), .A2(n7696), .A3(n7695), .ZN(n7697) );
  AOI21_X1 U8965 ( .B1(n7698), .B2(n10623), .A(n7697), .ZN(n7709) );
  INV_X1 U8966 ( .A(n7723), .ZN(n7699) );
  NAND2_X1 U8967 ( .A1(n10616), .A2(n7699), .ZN(n7704) );
  INV_X1 U8968 ( .A(n9313), .ZN(n10617) );
  NAND2_X1 U8969 ( .A1(n10617), .A2(n9329), .ZN(n7703) );
  INV_X1 U8970 ( .A(n7788), .ZN(n9327) );
  NAND2_X1 U8971 ( .A1(n10613), .A2(n9327), .ZN(n7702) );
  INV_X1 U8972 ( .A(n7700), .ZN(n7701) );
  NAND4_X1 U8973 ( .A1(n7704), .A2(n7703), .A3(n7702), .A4(n7701), .ZN(n7707)
         );
  NOR2_X1 U8974 ( .A1(n7705), .A2(n9306), .ZN(n7706) );
  AOI211_X1 U8975 ( .C1(n10611), .C2(n7768), .A(n7707), .B(n7706), .ZN(n7708)
         );
  OAI21_X1 U8976 ( .B1(n7710), .B2(n7709), .A(n7708), .ZN(P2_U3233) );
  INV_X1 U8977 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7711) );
  OAI222_X1 U8978 ( .A1(n8843), .A2(n9691), .B1(n9684), .B2(n7712), .C1(n7711), 
        .C2(n9687), .ZN(P2_U3337) );
  NAND2_X1 U8979 ( .A1(n7749), .A2(n7768), .ZN(n8932) );
  INV_X1 U8980 ( .A(n7768), .ZN(n11024) );
  OR2_X1 U8981 ( .A1(n7745), .A2(n7746), .ZN(n7716) );
  AND2_X1 U8982 ( .A1(n7716), .A2(n7750), .ZN(n7717) );
  AOI21_X1 U8983 ( .B1(n8864), .B2(n7717), .A(n5098), .ZN(n11023) );
  AOI22_X1 U8984 ( .A1(n9572), .A2(n9329), .B1(n9327), .B2(n9574), .ZN(n7722)
         );
  AND2_X1 U8985 ( .A1(n8921), .A2(n8923), .ZN(n7718) );
  NAND2_X1 U8986 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  INV_X1 U8987 ( .A(n8864), .ZN(n7758) );
  OR2_X1 U8988 ( .A1(n5425), .A2(n7758), .ZN(n7757) );
  OAI211_X1 U8989 ( .C1(n7762), .C2(n8864), .A(n9576), .B(n7757), .ZN(n7721)
         );
  OAI211_X1 U8990 ( .C1(n11023), .C2(n8275), .A(n7722), .B(n7721), .ZN(n11026)
         );
  NAND2_X1 U8991 ( .A1(n11026), .A2(n10933), .ZN(n7728) );
  INV_X1 U8992 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7724) );
  OAI22_X1 U8993 ( .A1(n10933), .A2(n7724), .B1(n7723), .B2(n9554), .ZN(n7726)
         );
  XNOR2_X1 U8994 ( .A(n7769), .B(n7768), .ZN(n11025) );
  NOR2_X1 U8995 ( .A1(n11025), .A2(n9398), .ZN(n7725) );
  AOI211_X1 U8996 ( .C1(n9542), .C2(n7768), .A(n7726), .B(n7725), .ZN(n7727)
         );
  OAI211_X1 U8997 ( .C1(n11023), .C2(n7776), .A(n7728), .B(n7727), .ZN(
        P2_U3287) );
  OAI21_X1 U8998 ( .B1(n7731), .B2(n7730), .A(n7729), .ZN(n7733) );
  NAND2_X1 U8999 ( .A1(n7731), .A2(n7730), .ZN(n7732) );
  NAND2_X1 U9000 ( .A1(n7738), .A2(n9133), .ZN(n7735) );
  NAND2_X1 U9001 ( .A1(n9807), .A2(n9160), .ZN(n7734) );
  NAND2_X1 U9002 ( .A1(n7735), .A2(n7734), .ZN(n7736) );
  XNOR2_X1 U9003 ( .A(n7736), .B(n9152), .ZN(n7828) );
  AND2_X1 U9004 ( .A1(n9807), .A2(n9159), .ZN(n7737) );
  AOI21_X1 U9005 ( .B1(n7738), .B2(n9143), .A(n7737), .ZN(n7829) );
  XNOR2_X1 U9006 ( .A(n7828), .B(n7829), .ZN(n7882) );
  AOI21_X1 U9007 ( .B1(n8003), .B2(n7882), .A(n9785), .ZN(n7739) );
  OR2_X1 U9008 ( .A1(n8003), .A2(n7882), .ZN(n7832) );
  NAND2_X1 U9009 ( .A1(n7739), .A2(n7832), .ZN(n7744) );
  AND2_X1 U9010 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10694) );
  AOI21_X1 U9011 ( .B1(n9758), .B2(n10991), .A(n10694), .ZN(n7740) );
  OAI21_X1 U9012 ( .B1(n9756), .B2(n7987), .A(n7740), .ZN(n7741) );
  AOI21_X1 U9013 ( .B1(n9796), .B2(n7742), .A(n7741), .ZN(n7743) );
  OAI211_X1 U9014 ( .C1(n11038), .C2(n9799), .A(n7744), .B(n7743), .ZN(
        P1_U3234) );
  INV_X1 U9015 ( .A(n7745), .ZN(n7748) );
  NAND2_X1 U9016 ( .A1(n7748), .A2(n7747), .ZN(n7755) );
  INV_X1 U9017 ( .A(n7752), .ZN(n7751) );
  AND2_X1 U9018 ( .A1(n7755), .A2(n7751), .ZN(n7756) );
  NAND2_X1 U9019 ( .A1(n7820), .A2(n7788), .ZN(n8931) );
  NAND2_X1 U9020 ( .A1(n8933), .A2(n8931), .ZN(n7759) );
  INV_X1 U9021 ( .A(n7759), .ZN(n7753) );
  NOR2_X1 U9022 ( .A1(n7753), .A2(n7752), .ZN(n7754) );
  OAI21_X1 U9023 ( .B1(n7756), .B2(n7759), .A(n7822), .ZN(n11030) );
  AOI22_X1 U9024 ( .A1(n9574), .A2(n9326), .B1(n9328), .B2(n9572), .ZN(n7765)
         );
  NAND2_X1 U9025 ( .A1(n7757), .A2(n8928), .ZN(n7763) );
  OR2_X1 U9026 ( .A1(n7759), .A2(n8928), .ZN(n7760) );
  INV_X1 U9027 ( .A(n7760), .ZN(n7761) );
  OAI211_X1 U9028 ( .C1(n7763), .C2(n7753), .A(n7813), .B(n9576), .ZN(n7764)
         );
  OAI211_X1 U9029 ( .C1(n11030), .C2(n8275), .A(n7765), .B(n7764), .ZN(n11033)
         );
  NAND2_X1 U9030 ( .A1(n11033), .A2(n10933), .ZN(n7775) );
  INV_X1 U9031 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7767) );
  OAI22_X1 U9032 ( .A1(n10933), .A2(n7767), .B1(n7766), .B2(n9554), .ZN(n7773)
         );
  NOR2_X1 U9033 ( .A1(n7770), .A2(n11031), .ZN(n7771) );
  OR2_X1 U9034 ( .A1(n7816), .A2(n7771), .ZN(n11032) );
  NOR2_X1 U9035 ( .A1(n11032), .A2(n9398), .ZN(n7772) );
  AOI211_X1 U9036 ( .C1(n9542), .C2(n7820), .A(n7773), .B(n7772), .ZN(n7774)
         );
  OAI211_X1 U9037 ( .C1(n11030), .C2(n7776), .A(n7775), .B(n7774), .ZN(
        P2_U3286) );
  INV_X1 U9038 ( .A(n8348), .ZN(n7779) );
  OAI222_X1 U9039 ( .A1(n10144), .A2(n7777), .B1(n10147), .B2(n7779), .C1(
        n8805), .C2(P1_U3084), .ZN(P1_U3331) );
  OAI222_X1 U9040 ( .A1(n9691), .A2(n7780), .B1(n9684), .B2(n7779), .C1(n7778), 
        .C2(n9687), .ZN(P2_U3336) );
  INV_X1 U9041 ( .A(n11045), .ZN(n7819) );
  AOI21_X1 U9042 ( .B1(n7689), .B2(n5578), .A(n9306), .ZN(n7785) );
  NOR3_X1 U9043 ( .A1(n7782), .A2(n7788), .A3(n10607), .ZN(n7784) );
  OAI21_X1 U9044 ( .B1(n7785), .B2(n7784), .A(n7783), .ZN(n7793) );
  INV_X1 U9045 ( .A(n7786), .ZN(n7817) );
  OR2_X1 U9046 ( .A1(n9068), .A2(n9550), .ZN(n7787) );
  OAI21_X1 U9047 ( .B1(n7788), .B2(n9548), .A(n7787), .ZN(n7814) );
  INV_X1 U9048 ( .A(n7814), .ZN(n7790) );
  OAI22_X1 U9049 ( .A1(n7790), .A2(n7789), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9339), .ZN(n7791) );
  AOI21_X1 U9050 ( .B1(n7817), .B2(n10616), .A(n7791), .ZN(n7792) );
  OAI211_X1 U9051 ( .C1(n7819), .C2(n9319), .A(n7793), .B(n7792), .ZN(P2_U3238) );
  NOR2_X1 U9052 ( .A1(n7801), .A2(n7794), .ZN(n7796) );
  NOR2_X1 U9053 ( .A1(n7796), .A2(n7795), .ZN(n7799) );
  NAND2_X1 U9054 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8145), .ZN(n7797) );
  OAI21_X1 U9055 ( .B1(n8145), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7797), .ZN(
        n7798) );
  NOR2_X1 U9056 ( .A1(n7799), .A2(n7798), .ZN(n8106) );
  AOI211_X1 U9057 ( .C1(n7799), .C2(n7798), .A(n8106), .B(n10808), .ZN(n7812)
         );
  NOR2_X1 U9058 ( .A1(n7801), .A2(n7800), .ZN(n7803) );
  NOR2_X1 U9059 ( .A1(n7803), .A2(n7802), .ZN(n7806) );
  NOR2_X1 U9060 ( .A1(n7809), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7804) );
  AOI21_X1 U9061 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n7809), .A(n7804), .ZN(
        n7805) );
  NOR2_X1 U9062 ( .A1(n7806), .A2(n7805), .ZN(n8110) );
  AOI211_X1 U9063 ( .C1(n7806), .C2(n7805), .A(n8110), .B(n10702), .ZN(n7811)
         );
  NAND2_X1 U9064 ( .A1(n10813), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U9065 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7807) );
  OAI211_X1 U9066 ( .C1(n10809), .C2(n7809), .A(n7808), .B(n7807), .ZN(n7810)
         );
  OR3_X1 U9067 ( .A1(n7812), .A2(n7811), .A3(n7810), .ZN(P1_U3257) );
  OR2_X1 U9068 ( .A1(n11045), .A2(n8073), .ZN(n8934) );
  NAND2_X1 U9069 ( .A1(n11045), .A2(n8073), .ZN(n8930) );
  NAND2_X1 U9070 ( .A1(n8934), .A2(n8930), .ZN(n8866) );
  XNOR2_X1 U9071 ( .A(n8029), .B(n8866), .ZN(n7815) );
  AOI21_X1 U9072 ( .B1(n7815), .B2(n9576), .A(n7814), .ZN(n11051) );
  OAI211_X1 U9073 ( .C1(n7816), .C2(n7819), .A(n11067), .B(n5096), .ZN(n11047)
         );
  INV_X1 U9074 ( .A(n11047), .ZN(n7826) );
  INV_X1 U9075 ( .A(n10933), .ZN(n9566) );
  AOI22_X1 U9076 ( .A1(n9566), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7817), .B2(
        n10927), .ZN(n7818) );
  OAI21_X1 U9077 ( .B1(n7819), .B2(n9568), .A(n7818), .ZN(n7825) );
  NAND2_X1 U9078 ( .A1(n7820), .A2(n9327), .ZN(n7821) );
  NAND2_X1 U9079 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  OAI21_X1 U9080 ( .B1(n7823), .B2(n8866), .A(n7869), .ZN(n11048) );
  NOR2_X1 U9081 ( .A1(n11048), .A2(n9581), .ZN(n7824) );
  AOI211_X1 U9082 ( .C1(n9467), .C2(n7826), .A(n7825), .B(n7824), .ZN(n7827)
         );
  OAI21_X1 U9083 ( .B1(n9541), .B2(n11051), .A(n7827), .ZN(P2_U3285) );
  INV_X1 U9084 ( .A(n7828), .ZN(n7831) );
  INV_X1 U9085 ( .A(n7829), .ZN(n7830) );
  NAND2_X1 U9086 ( .A1(n7831), .A2(n7830), .ZN(n7892) );
  NAND2_X1 U9087 ( .A1(n7832), .A2(n7892), .ZN(n7838) );
  NAND2_X1 U9088 ( .A1(n11054), .A2(n9133), .ZN(n7834) );
  NAND2_X1 U9089 ( .A1(n9806), .A2(n9160), .ZN(n7833) );
  NAND2_X1 U9090 ( .A1(n7834), .A2(n7833), .ZN(n7835) );
  XNOR2_X1 U9091 ( .A(n7835), .B(n9152), .ZN(n7888) );
  AND2_X1 U9092 ( .A1(n9806), .A2(n9159), .ZN(n7836) );
  AOI21_X1 U9093 ( .B1(n11054), .B2(n9143), .A(n7836), .ZN(n7881) );
  INV_X1 U9094 ( .A(n7881), .ZN(n7889) );
  XNOR2_X1 U9095 ( .A(n7888), .B(n7889), .ZN(n7837) );
  XNOR2_X1 U9096 ( .A(n7838), .B(n7837), .ZN(n7846) );
  INV_X1 U9097 ( .A(n7839), .ZN(n7841) );
  INV_X1 U9098 ( .A(n9805), .ZN(n7957) );
  NOR2_X1 U9099 ( .A1(n9756), .A2(n7957), .ZN(n7840) );
  AOI211_X1 U9100 ( .C1(n9758), .C2(n9807), .A(n7841), .B(n7840), .ZN(n7842)
         );
  OAI21_X1 U9101 ( .B1(n9760), .B2(n7843), .A(n7842), .ZN(n7844) );
  AOI21_X1 U9102 ( .B1(n11054), .B2(n9773), .A(n7844), .ZN(n7845) );
  OAI21_X1 U9103 ( .B1(n7846), .B2(n9785), .A(n7845), .ZN(P1_U3222) );
  OAI21_X1 U9104 ( .B1(n7848), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7847), .ZN(
        n8126) );
  XNOR2_X1 U9105 ( .A(n8126), .B(n8121), .ZN(n7849) );
  NAND2_X1 U9106 ( .A1(n7849), .A2(n8205), .ZN(n8128) );
  OAI21_X1 U9107 ( .B1(n7849), .B2(n8205), .A(n8128), .ZN(n7850) );
  INV_X1 U9108 ( .A(n7850), .ZN(n7858) );
  NAND2_X1 U9109 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n9073) );
  INV_X1 U9110 ( .A(n9073), .ZN(n7852) );
  NOR2_X1 U9111 ( .A1(n10763), .A2(n8127), .ZN(n7851) );
  AOI211_X1 U9112 ( .C1(n10787), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7852), .B(
        n7851), .ZN(n7857) );
  AOI21_X1 U9113 ( .B1(n7854), .B2(n6064), .A(n7853), .ZN(n8120) );
  XNOR2_X1 U9114 ( .A(n8120), .B(n8127), .ZN(n7855) );
  NAND2_X1 U9115 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7855), .ZN(n8122) );
  OAI211_X1 U9116 ( .C1(n7855), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10796), .B(
        n8122), .ZN(n7856) );
  OAI211_X1 U9117 ( .C1(n7858), .C2(n10788), .A(n7857), .B(n7856), .ZN(
        P2_U3260) );
  INV_X1 U9118 ( .A(n8359), .ZN(n7876) );
  NOR2_X1 U9119 ( .A1(n7859), .A2(P1_U3084), .ZN(n8808) );
  AOI21_X1 U9120 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10141), .A(n8808), .ZN(
        n7860) );
  OAI21_X1 U9121 ( .B1(n7876), .B2(n10147), .A(n7860), .ZN(P1_U3330) );
  NAND2_X1 U9122 ( .A1(n8029), .A2(n8930), .ZN(n7861) );
  NAND2_X1 U9123 ( .A1(n7861), .A2(n8934), .ZN(n7862) );
  OR2_X1 U9124 ( .A1(n11065), .A2(n9068), .ZN(n8941) );
  NAND2_X1 U9125 ( .A1(n11065), .A2(n9068), .ZN(n8030) );
  XNOR2_X1 U9126 ( .A(n7862), .B(n5370), .ZN(n7864) );
  OAI22_X1 U9127 ( .A1(n8518), .A2(n9550), .B1(n8073), .B2(n9548), .ZN(n7863)
         );
  AOI21_X1 U9128 ( .B1(n7864), .B2(n9576), .A(n7863), .ZN(n11070) );
  INV_X1 U9129 ( .A(n5642), .ZN(n8096) );
  AOI21_X1 U9130 ( .B1(n11065), .B2(n5096), .A(n8096), .ZN(n11068) );
  INV_X1 U9131 ( .A(n11065), .ZN(n7867) );
  INV_X1 U9132 ( .A(n8080), .ZN(n7865) );
  AOI22_X1 U9133 ( .A1(n9566), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7865), .B2(
        n10927), .ZN(n7866) );
  OAI21_X1 U9134 ( .B1(n7867), .B2(n9568), .A(n7866), .ZN(n7873) );
  NAND2_X1 U9135 ( .A1(n11045), .A2(n9326), .ZN(n7868) );
  INV_X1 U9136 ( .A(n8026), .ZN(n7870) );
  AOI21_X1 U9137 ( .B1(n8939), .B2(n7871), .A(n7870), .ZN(n11071) );
  NOR2_X1 U9138 ( .A1(n11071), .A2(n9581), .ZN(n7872) );
  AOI211_X1 U9139 ( .C1(n9579), .C2(n11068), .A(n7873), .B(n7872), .ZN(n7874)
         );
  OAI21_X1 U9140 ( .B1(n9566), .B2(n11070), .A(n7874), .ZN(P2_U3284) );
  NAND2_X1 U9141 ( .A1(n9682), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7875) );
  OAI211_X1 U9142 ( .C1(n7876), .C2(n9684), .A(n9047), .B(n7875), .ZN(P2_U3335) );
  NAND2_X1 U9143 ( .A1(n7877), .A2(n8546), .ZN(n7880) );
  AOI22_X1 U9144 ( .A1(n8421), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8320), .B2(
        n7878), .ZN(n7879) );
  INV_X1 U9145 ( .A(n7995), .ZN(n11075) );
  AND2_X1 U9146 ( .A1(n7888), .A2(n7881), .ZN(n7894) );
  OR2_X1 U9147 ( .A1(n7882), .A2(n7894), .ZN(n8004) );
  OR2_X1 U9148 ( .A1(n8003), .A2(n8004), .ZN(n7901) );
  NAND2_X1 U9149 ( .A1(n7995), .A2(n9133), .ZN(n7884) );
  NAND2_X1 U9150 ( .A1(n9805), .A2(n9160), .ZN(n7883) );
  NAND2_X1 U9151 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  XNOR2_X1 U9152 ( .A(n7885), .B(n9157), .ZN(n7896) );
  NAND2_X1 U9153 ( .A1(n7995), .A2(n9160), .ZN(n7887) );
  NAND2_X1 U9154 ( .A1(n9805), .A2(n9159), .ZN(n7886) );
  NAND2_X1 U9155 ( .A1(n7887), .A2(n7886), .ZN(n7897) );
  AND2_X1 U9156 ( .A1(n7896), .A2(n7897), .ZN(n7903) );
  INV_X1 U9157 ( .A(n7903), .ZN(n7895) );
  INV_X1 U9158 ( .A(n7888), .ZN(n7890) );
  NAND2_X1 U9159 ( .A1(n7890), .A2(n7889), .ZN(n7891) );
  AND2_X1 U9160 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  OR2_X1 U9161 ( .A1(n7894), .A2(n7893), .ZN(n7900) );
  AND2_X1 U9162 ( .A1(n7895), .A2(n7900), .ZN(n8005) );
  NAND2_X1 U9163 ( .A1(n7901), .A2(n8005), .ZN(n7905) );
  INV_X1 U9164 ( .A(n7896), .ZN(n7899) );
  INV_X1 U9165 ( .A(n7897), .ZN(n7898) );
  NAND2_X1 U9166 ( .A1(n7901), .A2(n7900), .ZN(n7902) );
  OAI21_X1 U9167 ( .B1(n8006), .B2(n7903), .A(n7902), .ZN(n7904) );
  OAI21_X1 U9168 ( .B1(n7905), .B2(n8006), .A(n7904), .ZN(n7906) );
  NAND2_X1 U9169 ( .A1(n7906), .A2(n9787), .ZN(n7912) );
  INV_X1 U9170 ( .A(n7907), .ZN(n7908) );
  AOI21_X1 U9171 ( .B1(n9758), .B2(n9806), .A(n7908), .ZN(n7909) );
  OAI21_X1 U9172 ( .B1(n9756), .B2(n8047), .A(n7909), .ZN(n7910) );
  AOI21_X1 U9173 ( .B1(n9796), .B2(n7994), .A(n7910), .ZN(n7911) );
  OAI211_X1 U9174 ( .C1(n11075), .C2(n9799), .A(n7912), .B(n7911), .ZN(
        P1_U3232) );
  NOR2_X1 U9175 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7950) );
  NOR2_X1 U9176 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7948) );
  NOR2_X1 U9177 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7946) );
  NOR2_X1 U9178 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7944) );
  NOR2_X1 U9179 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7941) );
  NOR2_X1 U9180 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7938) );
  NAND2_X1 U9181 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7936) );
  XOR2_X1 U9182 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10650) );
  NAND2_X1 U9183 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7934) );
  XOR2_X1 U9184 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10648) );
  NOR2_X1 U9185 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7918) );
  XNOR2_X1 U9186 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10639) );
  NAND2_X1 U9187 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7916) );
  XOR2_X1 U9188 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10637) );
  NAND2_X1 U9189 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7914) );
  XOR2_X1 U9190 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10635) );
  AOI21_X1 U9191 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10630) );
  NAND3_X1 U9192 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10632) );
  OAI21_X1 U9193 ( .B1(n10630), .B2(n10771), .A(n10632), .ZN(n10634) );
  NAND2_X1 U9194 ( .A1(n10635), .A2(n10634), .ZN(n7913) );
  NAND2_X1 U9195 ( .A1(n7914), .A2(n7913), .ZN(n10636) );
  NAND2_X1 U9196 ( .A1(n10637), .A2(n10636), .ZN(n7915) );
  NAND2_X1 U9197 ( .A1(n7916), .A2(n7915), .ZN(n10638) );
  NOR2_X1 U9198 ( .A1(n10639), .A2(n10638), .ZN(n7917) );
  NOR2_X1 U9199 ( .A1(n7918), .A2(n7917), .ZN(n7919) );
  NOR2_X1 U9200 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7919), .ZN(n10641) );
  AND2_X1 U9201 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7919), .ZN(n10640) );
  NAND2_X1 U9202 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7921), .ZN(n7923) );
  XOR2_X1 U9203 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7921), .Z(n10643) );
  NAND2_X1 U9204 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10643), .ZN(n7922) );
  NAND2_X1 U9205 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  NAND2_X1 U9206 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7924), .ZN(n7926) );
  XOR2_X1 U9207 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7924), .Z(n10644) );
  NAND2_X1 U9208 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10644), .ZN(n7925) );
  NAND2_X1 U9209 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  NAND2_X1 U9210 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7927), .ZN(n7929) );
  XOR2_X1 U9211 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7927), .Z(n10645) );
  NAND2_X1 U9212 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10645), .ZN(n7928) );
  NAND2_X1 U9213 ( .A1(n7929), .A2(n7928), .ZN(n7930) );
  NAND2_X1 U9214 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7930), .ZN(n7932) );
  XOR2_X1 U9215 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7930), .Z(n10646) );
  NAND2_X1 U9216 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10646), .ZN(n7931) );
  NAND2_X1 U9217 ( .A1(n7932), .A2(n7931), .ZN(n10647) );
  NAND2_X1 U9218 ( .A1(n10648), .A2(n10647), .ZN(n7933) );
  NAND2_X1 U9219 ( .A1(n7934), .A2(n7933), .ZN(n10649) );
  NAND2_X1 U9220 ( .A1(n10650), .A2(n10649), .ZN(n7935) );
  NAND2_X1 U9221 ( .A1(n7936), .A2(n7935), .ZN(n10652) );
  XNOR2_X1 U9222 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10651) );
  XOR2_X1 U9223 ( .A(n7939), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10653) );
  XOR2_X1 U9224 ( .A(n7942), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n10655) );
  NOR2_X1 U9225 ( .A1(n10656), .A2(n10655), .ZN(n7943) );
  NOR2_X1 U9226 ( .A1(n7944), .A2(n7943), .ZN(n10658) );
  XNOR2_X1 U9227 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10657) );
  NOR2_X1 U9228 ( .A1(n10658), .A2(n10657), .ZN(n7945) );
  NOR2_X1 U9229 ( .A1(n7946), .A2(n7945), .ZN(n10660) );
  XNOR2_X1 U9230 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10659) );
  NOR2_X1 U9231 ( .A1(n10660), .A2(n10659), .ZN(n7947) );
  NOR2_X1 U9232 ( .A1(n7948), .A2(n7947), .ZN(n10662) );
  XNOR2_X1 U9233 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10661) );
  NOR2_X1 U9234 ( .A1(n10662), .A2(n10661), .ZN(n7949) );
  NOR2_X1 U9235 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  AND2_X1 U9236 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7951), .ZN(n10663) );
  NOR2_X1 U9237 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10663), .ZN(n7952) );
  NOR2_X1 U9238 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7951), .ZN(n10664) );
  NOR2_X1 U9239 ( .A1(n7952), .A2(n10664), .ZN(n7954) );
  XNOR2_X1 U9240 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7953) );
  XNOR2_X1 U9241 ( .A(n7954), .B(n7953), .ZN(ADD_1071_U4) );
  NAND2_X1 U9242 ( .A1(n11054), .A2(n9806), .ZN(n7955) );
  OR2_X1 U9243 ( .A1(n7995), .A2(n7957), .ZN(n8662) );
  NAND2_X1 U9244 ( .A1(n7995), .A2(n7957), .ZN(n8663) );
  NAND2_X1 U9245 ( .A1(n8662), .A2(n8663), .ZN(n8761) );
  OR2_X1 U9246 ( .A1(n7995), .A2(n9805), .ZN(n7958) );
  NAND2_X1 U9247 ( .A1(n7959), .A2(n8546), .ZN(n7962) );
  AOI22_X1 U9248 ( .A1(n8421), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8320), .B2(
        n7960), .ZN(n7961) );
  OR2_X1 U9249 ( .A1(n8046), .A2(n8047), .ZN(n8661) );
  NAND2_X1 U9250 ( .A1(n8046), .A2(n8047), .ZN(n8670) );
  INV_X1 U9251 ( .A(n8764), .ZN(n7963) );
  XNOR2_X1 U9252 ( .A(n8049), .B(n7963), .ZN(n11092) );
  INV_X1 U9253 ( .A(n11092), .ZN(n7982) );
  INV_X1 U9254 ( .A(n8761), .ZN(n7986) );
  NAND2_X1 U9255 ( .A1(n8056), .A2(n8663), .ZN(n7965) );
  XNOR2_X1 U9256 ( .A(n7965), .B(n8764), .ZN(n7966) );
  NAND2_X1 U9257 ( .A1(n7966), .A2(n10998), .ZN(n7975) );
  NAND2_X1 U9258 ( .A1(n8401), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U9259 ( .A1(n6834), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7972) );
  AND2_X1 U9260 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  NOR2_X1 U9261 ( .A1(n8148), .A2(n7969), .ZN(n8185) );
  NAND2_X1 U9262 ( .A1(n5026), .A2(n8185), .ZN(n7971) );
  NAND2_X1 U9263 ( .A1(n8541), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7970) );
  NAND4_X1 U9264 ( .A1(n7973), .A2(n7972), .A3(n7971), .A4(n7970), .ZN(n9804)
         );
  AOI22_X1 U9265 ( .A1(n10993), .A2(n9805), .B1(n9804), .B2(n10990), .ZN(n7974) );
  NAND2_X1 U9266 ( .A1(n7975), .A2(n7974), .ZN(n11096) );
  OAI21_X1 U9267 ( .B1(n7992), .B2(n11094), .A(n10968), .ZN(n7976) );
  OR2_X1 U9268 ( .A1(n7976), .A2(n8067), .ZN(n11093) );
  AOI22_X1 U9269 ( .A1(n11014), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8017), .B2(
        n11012), .ZN(n7978) );
  NAND2_X1 U9270 ( .A1(n8046), .A2(n9863), .ZN(n7977) );
  OAI211_X1 U9271 ( .C1(n11093), .C2(n7979), .A(n7978), .B(n7977), .ZN(n7980)
         );
  AOI21_X1 U9272 ( .B1(n11096), .B2(n11019), .A(n7980), .ZN(n7981) );
  OAI21_X1 U9273 ( .B1(n7982), .B2(n10025), .A(n7981), .ZN(P1_U3277) );
  OAI21_X1 U9274 ( .B1(n7984), .B2(n8761), .A(n7983), .ZN(n11079) );
  INV_X1 U9275 ( .A(n11079), .ZN(n7991) );
  OAI21_X1 U9276 ( .B1(n7986), .B2(n7985), .A(n8056), .ZN(n7989) );
  OAI22_X1 U9277 ( .A1(n8047), .A2(n10030), .B1(n7987), .B2(n10028), .ZN(n7988) );
  AOI21_X1 U9278 ( .B1(n7989), .B2(n10998), .A(n7988), .ZN(n7990) );
  OAI21_X1 U9279 ( .B1(n7991), .B2(n7103), .A(n7990), .ZN(n11077) );
  INV_X1 U9280 ( .A(n11077), .ZN(n8000) );
  AND2_X1 U9281 ( .A1(n5040), .A2(n7995), .ZN(n7993) );
  OR2_X1 U9282 ( .A1(n7993), .A2(n7992), .ZN(n11076) );
  AOI22_X1 U9283 ( .A1(n11014), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7994), .B2(
        n11012), .ZN(n7997) );
  NAND2_X1 U9284 ( .A1(n7995), .A2(n9863), .ZN(n7996) );
  OAI211_X1 U9285 ( .C1(n11076), .C2(n9866), .A(n7997), .B(n7996), .ZN(n7998)
         );
  AOI21_X1 U9286 ( .B1(n11079), .B2(n11010), .A(n7998), .ZN(n7999) );
  OAI21_X1 U9287 ( .B1(n8000), .B2(n11014), .A(n7999), .ZN(P1_U3278) );
  NAND2_X1 U9288 ( .A1(n8046), .A2(n9160), .ZN(n8002) );
  NAND2_X1 U9289 ( .A1(n8187), .A2(n9159), .ZN(n8001) );
  NAND2_X1 U9290 ( .A1(n8002), .A2(n8001), .ZN(n8165) );
  OR2_X1 U9291 ( .A1(n8006), .A2(n8005), .ZN(n8012) );
  NAND2_X1 U9292 ( .A1(n8046), .A2(n9133), .ZN(n8008) );
  NAND2_X1 U9293 ( .A1(n8187), .A2(n9160), .ZN(n8007) );
  NAND2_X1 U9294 ( .A1(n8008), .A2(n8007), .ZN(n8009) );
  XNOR2_X1 U9295 ( .A(n8009), .B(n9152), .ZN(n8013) );
  INV_X1 U9296 ( .A(n8013), .ZN(n8010) );
  NAND2_X1 U9297 ( .A1(n8011), .A2(n8010), .ZN(n8167) );
  AND2_X1 U9298 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  NAND2_X1 U9299 ( .A1(n8167), .A2(n8166), .ZN(n8016) );
  XOR2_X1 U9300 ( .A(n8165), .B(n8016), .Z(n8022) );
  INV_X1 U9301 ( .A(n9804), .ZN(n8156) );
  NAND2_X1 U9302 ( .A1(n9796), .A2(n8017), .ZN(n8019) );
  AOI22_X1 U9303 ( .A1(n9758), .A2(n9805), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3084), .ZN(n8018) );
  OAI211_X1 U9304 ( .C1(n8156), .C2(n9756), .A(n8019), .B(n8018), .ZN(n8020)
         );
  AOI21_X1 U9305 ( .B1(n8046), .B2(n9773), .A(n8020), .ZN(n8021) );
  OAI21_X1 U9306 ( .B1(n8022), .B2(n9785), .A(n8021), .ZN(P1_U3213) );
  INV_X1 U9307 ( .A(n8373), .ZN(n8088) );
  INV_X1 U9308 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10382) );
  OAI222_X1 U9309 ( .A1(n8024), .A2(n8088), .B1(P1_U3084), .B2(n8023), .C1(
        n10382), .C2(n10144), .ZN(P1_U3329) );
  INV_X1 U9310 ( .A(n9068), .ZN(n9325) );
  OR2_X1 U9311 ( .A1(n11065), .A2(n9325), .ZN(n8025) );
  OR2_X1 U9312 ( .A1(n9067), .A2(n8518), .ZN(n8951) );
  NAND2_X1 U9313 ( .A1(n9067), .A2(n8518), .ZN(n8950) );
  NAND2_X1 U9314 ( .A1(n8951), .A2(n8950), .ZN(n8946) );
  INV_X1 U9315 ( .A(n8518), .ZN(n9324) );
  NAND2_X1 U9316 ( .A1(n9067), .A2(n9324), .ZN(n8027) );
  OR2_X1 U9317 ( .A1(n11101), .A2(n9081), .ZN(n8956) );
  NAND2_X1 U9318 ( .A1(n11101), .A2(n9081), .ZN(n8955) );
  NAND2_X1 U9319 ( .A1(n8956), .A2(n8955), .ZN(n8036) );
  OAI21_X1 U9320 ( .B1(n8028), .B2(n8036), .A(n8200), .ZN(n11106) );
  INV_X1 U9321 ( .A(n11106), .ZN(n8045) );
  AND2_X1 U9322 ( .A1(n8030), .A2(n8930), .ZN(n8943) );
  NAND2_X1 U9323 ( .A1(n8029), .A2(n8943), .ZN(n8090) );
  NAND2_X1 U9324 ( .A1(n8941), .A2(n8934), .ZN(n8031) );
  AND2_X1 U9325 ( .A1(n8031), .A2(n8030), .ZN(n8945) );
  NOR2_X1 U9326 ( .A1(n8946), .A2(n8945), .ZN(n8032) );
  NAND2_X1 U9327 ( .A1(n8090), .A2(n8032), .ZN(n8035) );
  INV_X1 U9328 ( .A(n8950), .ZN(n8033) );
  NOR2_X1 U9329 ( .A1(n8036), .A2(n8033), .ZN(n8034) );
  NAND2_X1 U9330 ( .A1(n8035), .A2(n8034), .ZN(n8201) );
  NAND2_X1 U9331 ( .A1(n8201), .A2(n9576), .ZN(n8039) );
  INV_X1 U9332 ( .A(n8036), .ZN(n8953) );
  AOI21_X1 U9333 ( .B1(n8035), .B2(n8950), .A(n8953), .ZN(n8038) );
  INV_X1 U9334 ( .A(n8511), .ZN(n9322) );
  AOI22_X1 U9335 ( .A1(n9574), .A2(n9322), .B1(n9324), .B2(n9572), .ZN(n8037)
         );
  OAI21_X1 U9336 ( .B1(n8039), .B2(n8038), .A(n8037), .ZN(n11105) );
  XNOR2_X1 U9337 ( .A(n8203), .B(n11101), .ZN(n11103) );
  OAI22_X1 U9338 ( .A1(n10933), .A2(n8040), .B1(n8514), .B2(n9554), .ZN(n8041)
         );
  AOI21_X1 U9339 ( .B1(n11101), .B2(n9542), .A(n8041), .ZN(n8042) );
  OAI21_X1 U9340 ( .B1(n11103), .B2(n9398), .A(n8042), .ZN(n8043) );
  AOI21_X1 U9341 ( .B1(n11105), .B2(n10933), .A(n8043), .ZN(n8044) );
  OAI21_X1 U9342 ( .B1(n8045), .B2(n9581), .A(n8044), .ZN(P2_U3282) );
  NOR2_X1 U9343 ( .A1(n8046), .A2(n8187), .ZN(n8048) );
  NAND2_X1 U9344 ( .A1(n8050), .A2(n8546), .ZN(n8053) );
  AOI22_X1 U9345 ( .A1(n8421), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8320), .B2(
        n8051), .ZN(n8052) );
  OR2_X1 U9346 ( .A1(n8191), .A2(n8156), .ZN(n8674) );
  NAND2_X1 U9347 ( .A1(n8191), .A2(n8156), .ZN(n8673) );
  XNOR2_X1 U9348 ( .A(n8141), .B(n8763), .ZN(n11115) );
  AND2_X1 U9349 ( .A1(n8764), .A2(n8663), .ZN(n8055) );
  INV_X1 U9350 ( .A(n8661), .ZN(n8054) );
  OAI21_X1 U9351 ( .B1(n8763), .B2(n8057), .A(n8155), .ZN(n8058) );
  NAND2_X1 U9352 ( .A1(n8058), .A2(n10998), .ZN(n8065) );
  NAND2_X1 U9353 ( .A1(n8401), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U9354 ( .A1(n6834), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8062) );
  INV_X1 U9355 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8059) );
  XNOR2_X1 U9356 ( .A(n8148), .B(n8059), .ZN(n8230) );
  NAND2_X1 U9357 ( .A1(n5026), .A2(n8230), .ZN(n8061) );
  NAND2_X1 U9358 ( .A1(n8541), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8060) );
  NAND4_X1 U9359 ( .A1(n8063), .A2(n8062), .A3(n8061), .A4(n8060), .ZN(n9803)
         );
  AOI22_X1 U9360 ( .A1(n10993), .A2(n8187), .B1(n9803), .B2(n10990), .ZN(n8064) );
  NAND2_X1 U9361 ( .A1(n8065), .A2(n8064), .ZN(n8066) );
  AOI21_X1 U9362 ( .B1(n11115), .B2(n11062), .A(n8066), .ZN(n11117) );
  INV_X1 U9363 ( .A(n8191), .ZN(n11110) );
  OR2_X1 U9364 ( .A1(n8067), .A2(n11110), .ZN(n8068) );
  NAND2_X1 U9365 ( .A1(n8159), .A2(n8068), .ZN(n11112) );
  AOI22_X1 U9366 ( .A1(n11014), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8185), .B2(
        n11012), .ZN(n8070) );
  NAND2_X1 U9367 ( .A1(n8191), .A2(n9863), .ZN(n8069) );
  OAI211_X1 U9368 ( .C1(n11112), .C2(n9866), .A(n8070), .B(n8069), .ZN(n8071)
         );
  AOI21_X1 U9369 ( .B1(n11115), .B2(n11010), .A(n8071), .ZN(n8072) );
  OAI21_X1 U9370 ( .B1(n11117), .B2(n11014), .A(n8072), .ZN(P1_U3276) );
  INV_X1 U9371 ( .A(n7783), .ZN(n8076) );
  NOR3_X1 U9372 ( .A1(n8074), .A2(n8073), .A3(n10607), .ZN(n8075) );
  AOI21_X1 U9373 ( .B1(n8076), .B2(n10623), .A(n8075), .ZN(n8085) );
  OAI21_X1 U9374 ( .B1(n9314), .B2(n8518), .A(n8077), .ZN(n8078) );
  AOI21_X1 U9375 ( .B1(n10617), .B2(n9326), .A(n8078), .ZN(n8079) );
  OAI21_X1 U9376 ( .B1(n8080), .B2(n9294), .A(n8079), .ZN(n8083) );
  NOR2_X1 U9377 ( .A1(n8081), .A2(n9306), .ZN(n8082) );
  AOI211_X1 U9378 ( .C1(n10611), .C2(n11065), .A(n8083), .B(n8082), .ZN(n8084)
         );
  OAI21_X1 U9379 ( .B1(n8086), .B2(n8085), .A(n8084), .ZN(P2_U3226) );
  INV_X1 U9380 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8087) );
  OAI222_X1 U9381 ( .A1(n8089), .A2(n9691), .B1(n9684), .B2(n8088), .C1(n8087), 
        .C2(n9687), .ZN(P2_U3334) );
  INV_X1 U9382 ( .A(n8945), .ZN(n8091) );
  NAND2_X1 U9383 ( .A1(n8090), .A2(n8091), .ZN(n8093) );
  INV_X1 U9384 ( .A(n8035), .ZN(n8092) );
  AOI21_X1 U9385 ( .B1(n8946), .B2(n8093), .A(n8092), .ZN(n8094) );
  OAI222_X1 U9386 ( .A1(n9548), .A2(n9068), .B1(n9550), .B2(n9081), .C1(n9546), 
        .C2(n8094), .ZN(n11086) );
  INV_X1 U9387 ( .A(n11086), .ZN(n8105) );
  OAI22_X1 U9388 ( .A1(n10933), .A2(n8095), .B1(n9065), .B2(n9554), .ZN(n8098)
         );
  INV_X1 U9389 ( .A(n9067), .ZN(n11084) );
  OAI21_X1 U9390 ( .B1(n8096), .B2(n11084), .A(n8203), .ZN(n11085) );
  NOR2_X1 U9391 ( .A1(n11085), .A2(n9398), .ZN(n8097) );
  AOI211_X1 U9392 ( .C1(n9542), .C2(n9067), .A(n8098), .B(n8097), .ZN(n8104)
         );
  NOR2_X1 U9393 ( .A1(n8099), .A2(n8946), .ZN(n11083) );
  INV_X1 U9394 ( .A(n11083), .ZN(n8102) );
  NAND3_X1 U9395 ( .A1(n8102), .A2(n8101), .A3(n8100), .ZN(n8103) );
  OAI211_X1 U9396 ( .C1(n8105), .C2(n9566), .A(n8104), .B(n8103), .ZN(P2_U3283) );
  NAND2_X1 U9397 ( .A1(n9843), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8107) );
  OAI21_X1 U9398 ( .B1(n9843), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8107), .ZN(
        n8108) );
  AOI211_X1 U9399 ( .C1(n8109), .C2(n8108), .A(n9842), .B(n10808), .ZN(n8118)
         );
  AOI21_X1 U9400 ( .B1(n8145), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8110), .ZN(
        n8112) );
  XNOR2_X1 U9401 ( .A(n9843), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8111) );
  NOR2_X1 U9402 ( .A1(n8112), .A2(n8111), .ZN(n9837) );
  AOI211_X1 U9403 ( .C1(n8112), .C2(n8111), .A(n9837), .B(n10702), .ZN(n8113)
         );
  INV_X1 U9404 ( .A(n8113), .ZN(n8115) );
  NAND2_X1 U9405 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n8114) );
  OAI211_X1 U9406 ( .C1(n10809), .C2(n8116), .A(n8115), .B(n8114), .ZN(n8117)
         );
  AOI211_X1 U9407 ( .C1(n10813), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n8118), .B(
        n8117), .ZN(n8119) );
  INV_X1 U9408 ( .A(n8119), .ZN(P1_U3258) );
  NAND2_X1 U9409 ( .A1(n8121), .A2(n8120), .ZN(n8123) );
  NAND2_X1 U9410 ( .A1(n8123), .A2(n8122), .ZN(n8125) );
  XNOR2_X1 U9411 ( .A(n9349), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8124) );
  NOR2_X1 U9412 ( .A1(n8125), .A2(n8124), .ZN(n9355) );
  AOI21_X1 U9413 ( .B1(n8125), .B2(n8124), .A(n9355), .ZN(n8139) );
  NAND2_X1 U9414 ( .A1(n8127), .A2(n8126), .ZN(n8129) );
  NAND2_X1 U9415 ( .A1(n8129), .A2(n8128), .ZN(n8132) );
  MUX2_X1 U9416 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n6101), .S(n9349), .Z(n8130)
         );
  INV_X1 U9417 ( .A(n8130), .ZN(n8131) );
  NOR2_X1 U9418 ( .A1(n8132), .A2(n8131), .ZN(n9348) );
  AOI211_X1 U9419 ( .C1(n8132), .C2(n8131), .A(n9348), .B(n10788), .ZN(n8133)
         );
  INV_X1 U9420 ( .A(n8133), .ZN(n8137) );
  NOR2_X1 U9421 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10474), .ZN(n8135) );
  NOR2_X1 U9422 ( .A1(n10763), .A2(n9357), .ZN(n8134) );
  AOI211_X1 U9423 ( .C1(n10787), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8135), .B(
        n8134), .ZN(n8136) );
  OAI211_X1 U9424 ( .C1(n8139), .C2(n8138), .A(n8137), .B(n8136), .ZN(P2_U3261) );
  INV_X1 U9425 ( .A(n8763), .ZN(n8140) );
  NAND2_X1 U9426 ( .A1(n8141), .A2(n8140), .ZN(n8143) );
  NAND2_X1 U9427 ( .A1(n8191), .A2(n9804), .ZN(n8142) );
  NAND2_X1 U9428 ( .A1(n8143), .A2(n8142), .ZN(n8308) );
  NAND2_X1 U9429 ( .A1(n8144), .A2(n8546), .ZN(n8147) );
  AOI22_X1 U9430 ( .A1(n8421), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8320), .B2(
        n8145), .ZN(n8146) );
  INV_X1 U9431 ( .A(n9803), .ZN(n10029) );
  NAND2_X1 U9432 ( .A1(n10119), .A2(n10029), .ZN(n8680) );
  XNOR2_X1 U9433 ( .A(n8308), .B(n8683), .ZN(n10121) );
  NAND2_X1 U9434 ( .A1(n8401), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8154) );
  AOI21_X1 U9435 ( .B1(n8148), .B2(P1_REG3_REG_16__SCAN_IN), .A(
        P1_REG3_REG_17__SCAN_IN), .ZN(n8149) );
  OR2_X1 U9436 ( .A1(n8150), .A2(n8149), .ZN(n8256) );
  INV_X1 U9437 ( .A(n8256), .ZN(n10039) );
  NAND2_X1 U9438 ( .A1(n10039), .A2(n5026), .ZN(n8153) );
  NAND2_X1 U9439 ( .A1(n8541), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U9440 ( .A1(n6834), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8151) );
  NAND4_X1 U9441 ( .A1(n8154), .A2(n8153), .A3(n8152), .A4(n8151), .ZN(n9802)
         );
  XNOR2_X1 U9442 ( .A(n8457), .B(n8683), .ZN(n8157) );
  OAI222_X1 U9443 ( .A1(n10030), .A2(n10018), .B1(n8157), .B2(n10867), .C1(
        n10028), .C2(n8156), .ZN(n10117) );
  INV_X1 U9444 ( .A(n10119), .ZN(n8162) );
  INV_X1 U9445 ( .A(n10038), .ZN(n8158) );
  AOI211_X1 U9446 ( .C1(n10119), .C2(n8159), .A(n11111), .B(n8158), .ZN(n10118) );
  NAND2_X1 U9447 ( .A1(n10118), .A2(n10005), .ZN(n8161) );
  AOI22_X1 U9448 ( .A1(n11014), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8230), .B2(
        n11012), .ZN(n8160) );
  OAI211_X1 U9449 ( .C1(n8162), .C2(n11016), .A(n8161), .B(n8160), .ZN(n8163)
         );
  AOI21_X1 U9450 ( .B1(n10117), .B2(n11019), .A(n8163), .ZN(n8164) );
  OAI21_X1 U9451 ( .B1(n10025), .B2(n10121), .A(n8164), .ZN(P1_U3275) );
  NAND2_X1 U9452 ( .A1(n8166), .A2(n8165), .ZN(n8168) );
  NAND2_X1 U9453 ( .A1(n8191), .A2(n9133), .ZN(n8170) );
  NAND2_X1 U9454 ( .A1(n9804), .A2(n9160), .ZN(n8169) );
  NAND2_X1 U9455 ( .A1(n8170), .A2(n8169), .ZN(n8171) );
  XNOR2_X1 U9456 ( .A(n8171), .B(n9152), .ZN(n8175) );
  NAND2_X1 U9457 ( .A1(n8174), .A2(n8175), .ZN(n8178) );
  NAND2_X1 U9458 ( .A1(n8191), .A2(n9160), .ZN(n8173) );
  NAND2_X1 U9459 ( .A1(n9804), .A2(n9159), .ZN(n8172) );
  NAND2_X1 U9460 ( .A1(n8173), .A2(n8172), .ZN(n8182) );
  INV_X1 U9461 ( .A(n8174), .ZN(n8177) );
  INV_X1 U9462 ( .A(n8175), .ZN(n8176) );
  INV_X1 U9463 ( .A(n8227), .ZN(n8184) );
  INV_X1 U9464 ( .A(n8179), .ZN(n8181) );
  NAND2_X1 U9465 ( .A1(n8181), .A2(n8180), .ZN(n8183) );
  AOI22_X1 U9466 ( .A1(n8184), .A2(n8178), .B1(n8183), .B2(n8182), .ZN(n8193)
         );
  NAND2_X1 U9467 ( .A1(n9796), .A2(n8185), .ZN(n8189) );
  AOI21_X1 U9468 ( .B1(n9758), .B2(n8187), .A(n8186), .ZN(n8188) );
  OAI211_X1 U9469 ( .C1(n10029), .C2(n9756), .A(n8189), .B(n8188), .ZN(n8190)
         );
  AOI21_X1 U9470 ( .B1(n8191), .B2(n9773), .A(n8190), .ZN(n8192) );
  OAI21_X1 U9471 ( .B1(n8193), .B2(n9785), .A(n8192), .ZN(P1_U3239) );
  INV_X1 U9472 ( .A(n8385), .ZN(n8197) );
  OAI222_X1 U9473 ( .A1(P2_U3152), .A2(n8195), .B1(n9684), .B2(n8197), .C1(
        n8194), .C2(n9687), .ZN(P2_U3333) );
  OAI222_X1 U9474 ( .A1(n10144), .A2(n8198), .B1(n10147), .B2(n8197), .C1(
        n8196), .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9475 ( .A(n9081), .ZN(n9323) );
  OR2_X1 U9476 ( .A1(n11101), .A2(n9323), .ZN(n8199) );
  OR2_X1 U9477 ( .A1(n9079), .A2(n8511), .ZN(n8960) );
  NAND2_X1 U9478 ( .A1(n9079), .A2(n8511), .ZN(n8961) );
  NAND2_X1 U9479 ( .A1(n8960), .A2(n8961), .ZN(n8270) );
  XNOR2_X1 U9480 ( .A(n8271), .B(n8270), .ZN(n11130) );
  INV_X1 U9481 ( .A(n11130), .ZN(n8210) );
  NAND2_X1 U9482 ( .A1(n8201), .A2(n8956), .ZN(n8277) );
  INV_X1 U9483 ( .A(n8270), .ZN(n8958) );
  XNOR2_X1 U9484 ( .A(n8277), .B(n8958), .ZN(n8202) );
  OAI222_X1 U9485 ( .A1(n9550), .A2(n9074), .B1(n9548), .B2(n9081), .C1(n9546), 
        .C2(n8202), .ZN(n11127) );
  INV_X1 U9486 ( .A(n9079), .ZN(n11124) );
  OAI21_X1 U9487 ( .B1(n8204), .B2(n11124), .A(n8293), .ZN(n11126) );
  OAI22_X1 U9488 ( .A1(n10933), .A2(n8205), .B1(n9077), .B2(n9554), .ZN(n8206)
         );
  AOI21_X1 U9489 ( .B1(n9079), .B2(n9542), .A(n8206), .ZN(n8207) );
  OAI21_X1 U9490 ( .B1(n11126), .B2(n9398), .A(n8207), .ZN(n8208) );
  AOI21_X1 U9491 ( .B1(n11127), .B2(n10933), .A(n8208), .ZN(n8209) );
  OAI21_X1 U9492 ( .B1(n8210), .B2(n9581), .A(n8209), .ZN(P2_U3281) );
  NAND2_X1 U9493 ( .A1(n9573), .A2(n9574), .ZN(n8211) );
  OAI21_X1 U9494 ( .B1(n8511), .B2(n9548), .A(n8211), .ZN(n8300) );
  AOI22_X1 U9495 ( .A1(n8300), .A2(n9251), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8212) );
  OAI21_X1 U9496 ( .B1(n8294), .B2(n9294), .A(n8212), .ZN(n8213) );
  AOI21_X1 U9497 ( .B1(n9658), .B2(n10611), .A(n8213), .ZN(n8220) );
  INV_X1 U9498 ( .A(n8215), .ZN(n8218) );
  OAI22_X1 U9499 ( .A1(n8216), .A2(n9306), .B1(n8511), .B2(n10607), .ZN(n8217)
         );
  NAND3_X1 U9500 ( .A1(n8214), .A2(n8218), .A3(n8217), .ZN(n8219) );
  OAI211_X1 U9501 ( .C1(n8221), .C2(n9306), .A(n8220), .B(n8219), .ZN(P2_U3228) );
  INV_X1 U9502 ( .A(n8398), .ZN(n8239) );
  OAI222_X1 U9503 ( .A1(n10147), .A2(n8239), .B1(n10144), .B2(n5753), .C1(
        n8222), .C2(P1_U3084), .ZN(P1_U3327) );
  NAND2_X1 U9504 ( .A1(n10119), .A2(n9133), .ZN(n8224) );
  NAND2_X1 U9505 ( .A1(n9803), .A2(n9160), .ZN(n8223) );
  NAND2_X1 U9506 ( .A1(n8224), .A2(n8223), .ZN(n8225) );
  XNOR2_X1 U9507 ( .A(n8225), .B(n9152), .ZN(n8244) );
  AND2_X1 U9508 ( .A1(n9803), .A2(n9159), .ZN(n8226) );
  AOI21_X1 U9509 ( .B1(n10119), .B2(n9143), .A(n8226), .ZN(n8243) );
  XNOR2_X1 U9510 ( .A(n8244), .B(n8243), .ZN(n8229) );
  INV_X1 U9511 ( .A(n8246), .ZN(n8228) );
  AOI21_X1 U9512 ( .B1(n8229), .B2(n8227), .A(n8228), .ZN(n8235) );
  NAND2_X1 U9513 ( .A1(n9796), .A2(n8230), .ZN(n8232) );
  AOI22_X1 U9514 ( .A1(n9758), .A2(n9804), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8231) );
  OAI211_X1 U9515 ( .C1(n10018), .C2(n9756), .A(n8232), .B(n8231), .ZN(n8233)
         );
  AOI21_X1 U9516 ( .B1(n10119), .B2(n9773), .A(n8233), .ZN(n8234) );
  OAI21_X1 U9517 ( .B1(n8235), .B2(n9785), .A(n8234), .ZN(P1_U3224) );
  INV_X1 U9518 ( .A(n8412), .ZN(n9689) );
  AOI21_X1 U9519 ( .B1(n10141), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n8236), .ZN(
        n8237) );
  OAI21_X1 U9520 ( .B1(n9689), .B2(n10147), .A(n8237), .ZN(P1_U3326) );
  OAI222_X1 U9521 ( .A1(n8240), .A2(P2_U3152), .B1(n9684), .B2(n8239), .C1(
        n8238), .C2(n9687), .ZN(P2_U3332) );
  INV_X1 U9522 ( .A(n8420), .ZN(n9202) );
  AOI21_X1 U9523 ( .B1(n10141), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n8241), .ZN(
        n8242) );
  OAI21_X1 U9524 ( .B1(n9202), .B2(n10147), .A(n8242), .ZN(P1_U3325) );
  NAND2_X1 U9525 ( .A1(n8244), .A2(n8243), .ZN(n8245) );
  NAND2_X1 U9526 ( .A1(n8247), .A2(n8546), .ZN(n8249) );
  AOI22_X1 U9527 ( .A1(n8421), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8320), .B2(
        n9843), .ZN(n8248) );
  NAND2_X1 U9528 ( .A1(n10112), .A2(n9133), .ZN(n8251) );
  NAND2_X1 U9529 ( .A1(n9802), .A2(n9160), .ZN(n8250) );
  NAND2_X1 U9530 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  XNOR2_X1 U9531 ( .A(n8252), .B(n9157), .ZN(n9089) );
  AND2_X1 U9532 ( .A1(n9802), .A2(n9159), .ZN(n8253) );
  AOI21_X1 U9533 ( .B1(n10112), .B2(n9143), .A(n8253), .ZN(n9090) );
  XNOR2_X1 U9534 ( .A(n9089), .B(n9090), .ZN(n9093) );
  XOR2_X1 U9535 ( .A(n9094), .B(n9093), .Z(n8259) );
  AOI22_X1 U9536 ( .A1(n9791), .A2(n10000), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8255) );
  NAND2_X1 U9537 ( .A1(n9758), .A2(n9803), .ZN(n8254) );
  OAI211_X1 U9538 ( .C1(n9760), .C2(n8256), .A(n8255), .B(n8254), .ZN(n8257)
         );
  AOI21_X1 U9539 ( .B1(n10112), .B2(n9773), .A(n8257), .ZN(n8258) );
  OAI21_X1 U9540 ( .B1(n8259), .B2(n9785), .A(n8258), .ZN(P1_U3226) );
  INV_X1 U9541 ( .A(n8261), .ZN(n8263) );
  NAND2_X1 U9542 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  XNOR2_X1 U9543 ( .A(n8260), .B(n8264), .ZN(n8269) );
  NOR2_X1 U9544 ( .A1(n9294), .A2(n8283), .ZN(n8267) );
  INV_X1 U9545 ( .A(n9074), .ZN(n9321) );
  NAND2_X1 U9546 ( .A1(n10617), .A2(n9321), .ZN(n8265) );
  NAND2_X1 U9547 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n9353) );
  OAI211_X1 U9548 ( .C1(n9547), .C2(n9314), .A(n8265), .B(n9353), .ZN(n8266)
         );
  AOI211_X1 U9549 ( .C1(n9653), .C2(n10611), .A(n8267), .B(n8266), .ZN(n8268)
         );
  OAI21_X1 U9550 ( .B1(n8269), .B2(n9306), .A(n8268), .ZN(P2_U3230) );
  OR2_X1 U9551 ( .A1(n9658), .A2(n9074), .ZN(n8966) );
  NAND2_X1 U9552 ( .A1(n9658), .A2(n9074), .ZN(n8965) );
  NAND2_X1 U9553 ( .A1(n9658), .A2(n9321), .ZN(n8273) );
  NAND2_X1 U9554 ( .A1(n9653), .A2(n9573), .ZN(n8274) );
  OAI21_X1 U9555 ( .B1(n5092), .B2(n8870), .A(n9174), .ZN(n9650) );
  INV_X1 U9556 ( .A(n8275), .ZN(n8282) );
  XOR2_X1 U9557 ( .A(n9653), .B(n9189), .Z(n8276) );
  NAND2_X1 U9558 ( .A1(n8276), .A2(n11067), .ZN(n9651) );
  INV_X1 U9559 ( .A(n8960), .ZN(n8298) );
  OAI211_X1 U9560 ( .C1(n8277), .C2(n8298), .A(n8965), .B(n8961), .ZN(n8278)
         );
  NAND2_X1 U9561 ( .A1(n8278), .A2(n8966), .ZN(n8813) );
  XNOR2_X1 U9562 ( .A(n8813), .B(n8870), .ZN(n8280) );
  OAI22_X1 U9563 ( .A1(n9074), .A2(n9548), .B1(n9547), .B2(n9550), .ZN(n8279)
         );
  AOI21_X1 U9564 ( .B1(n8280), .B2(n9576), .A(n8279), .ZN(n9655) );
  OAI21_X1 U9565 ( .B1(n9555), .B2(n9651), .A(n9655), .ZN(n8281) );
  AOI21_X1 U9566 ( .B1(n9650), .B2(n8282), .A(n8281), .ZN(n8289) );
  OAI22_X1 U9567 ( .A1(n10933), .A2(n8284), .B1(n8283), .B2(n9554), .ZN(n8285)
         );
  AOI21_X1 U9568 ( .B1(n9653), .B2(n9542), .A(n8285), .ZN(n8288) );
  NAND2_X1 U9569 ( .A1(n9650), .A2(n8286), .ZN(n8287) );
  OAI211_X1 U9570 ( .C1(n8289), .C2(n9541), .A(n8288), .B(n8287), .ZN(P2_U3279) );
  OAI21_X1 U9571 ( .B1(n8291), .B2(n8272), .A(n8290), .ZN(n9661) );
  INV_X1 U9572 ( .A(n9189), .ZN(n8292) );
  AOI211_X1 U9573 ( .C1(n9658), .C2(n8293), .A(n11125), .B(n8292), .ZN(n9657)
         );
  INV_X1 U9574 ( .A(n9658), .ZN(n8297) );
  INV_X1 U9575 ( .A(n8294), .ZN(n8295) );
  AOI22_X1 U9576 ( .A1(n9566), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8295), .B2(
        n10927), .ZN(n8296) );
  OAI21_X1 U9577 ( .B1(n8297), .B2(n9568), .A(n8296), .ZN(n8303) );
  AOI21_X1 U9578 ( .B1(n8277), .B2(n8961), .A(n8298), .ZN(n8299) );
  XNOR2_X1 U9579 ( .A(n8299), .B(n8963), .ZN(n8301) );
  AOI21_X1 U9580 ( .B1(n8301), .B2(n9576), .A(n8300), .ZN(n9660) );
  NOR2_X1 U9581 ( .A1(n9660), .A2(n9541), .ZN(n8302) );
  AOI211_X1 U9582 ( .C1(n9657), .C2(n9467), .A(n8303), .B(n8302), .ZN(n8304)
         );
  OAI21_X1 U9583 ( .B1(n9581), .B2(n9661), .A(n8304), .ZN(P2_U3280) );
  OAI222_X1 U9584 ( .A1(n8307), .A2(P2_U3152), .B1(n9684), .B2(n8306), .C1(
        n8305), .C2(n9687), .ZN(P2_U3338) );
  NAND2_X1 U9585 ( .A1(n8308), .A2(n8683), .ZN(n8310) );
  NAND2_X1 U9586 ( .A1(n10119), .A2(n9803), .ZN(n8309) );
  NAND2_X1 U9587 ( .A1(n8310), .A2(n8309), .ZN(n10032) );
  OR2_X1 U9588 ( .A1(n10112), .A2(n9802), .ZN(n8311) );
  NAND2_X1 U9589 ( .A1(n10032), .A2(n8311), .ZN(n8313) );
  NAND2_X1 U9590 ( .A1(n10112), .A2(n9802), .ZN(n8312) );
  NAND2_X1 U9591 ( .A1(n8313), .A2(n8312), .ZN(n10007) );
  NAND2_X1 U9592 ( .A1(n8314), .A2(n8546), .ZN(n8316) );
  AOI22_X1 U9593 ( .A1(n8421), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8320), .B2(
        n9846), .ZN(n8315) );
  INV_X1 U9594 ( .A(n10000), .ZN(n10031) );
  OR2_X1 U9595 ( .A1(n10107), .A2(n10031), .ZN(n8688) );
  NAND2_X1 U9596 ( .A1(n10107), .A2(n10031), .ZN(n8689) );
  NAND2_X1 U9597 ( .A1(n8688), .A2(n8689), .ZN(n10017) );
  NAND2_X1 U9598 ( .A1(n10007), .A2(n10017), .ZN(n8318) );
  NAND2_X1 U9599 ( .A1(n10107), .A2(n10000), .ZN(n8317) );
  NAND2_X1 U9600 ( .A1(n8318), .A2(n8317), .ZN(n9991) );
  NAND2_X1 U9601 ( .A1(n8319), .A2(n8546), .ZN(n8322) );
  AOI22_X1 U9602 ( .A1(n8421), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8320), .B2(
        n9850), .ZN(n8321) );
  NOR2_X1 U9603 ( .A1(n9998), .A2(n10019), .ZN(n8324) );
  NAND2_X1 U9604 ( .A1(n9998), .A2(n10019), .ZN(n8323) );
  OAI21_X1 U9605 ( .B1(n9991), .B2(n8324), .A(n8323), .ZN(n9976) );
  NAND2_X1 U9606 ( .A1(n8325), .A2(n8546), .ZN(n8327) );
  NAND2_X1 U9607 ( .A1(n8421), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8326) );
  INV_X1 U9608 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9755) );
  AND2_X1 U9609 ( .A1(n8328), .A2(n9755), .ZN(n8329) );
  OR2_X1 U9610 ( .A1(n8329), .A2(n8337), .ZN(n9978) );
  INV_X1 U9611 ( .A(n5026), .ZN(n8339) );
  AOI22_X1 U9612 ( .A1(n8401), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n6834), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U9613 ( .A1(n8541), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8330) );
  OAI211_X1 U9614 ( .C1(n9978), .C2(n8339), .A(n8331), .B(n8330), .ZN(n10001)
         );
  INV_X1 U9615 ( .A(n10001), .ZN(n8332) );
  OR2_X1 U9616 ( .A1(n10097), .A2(n8332), .ZN(n8555) );
  NAND2_X1 U9617 ( .A1(n10097), .A2(n8332), .ZN(n8551) );
  INV_X1 U9618 ( .A(n9984), .ZN(n8333) );
  AOI21_X2 U9619 ( .B1(n9976), .B2(n8333), .A(n5046), .ZN(n9960) );
  NAND2_X1 U9620 ( .A1(n8334), .A2(n8546), .ZN(n8336) );
  NAND2_X1 U9621 ( .A1(n8421), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8335) );
  OR2_X1 U9622 ( .A1(n8337), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U9623 ( .A1(n8337), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U9624 ( .A1(n8338), .A2(n8352), .ZN(n9964) );
  OR2_X1 U9625 ( .A1(n9964), .A2(n8339), .ZN(n8345) );
  INV_X1 U9626 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U9627 ( .A1(n8401), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U9628 ( .A1(n6834), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8340) );
  OAI211_X1 U9629 ( .C1(n8342), .C2(n6600), .A(n8341), .B(n8340), .ZN(n8343)
         );
  INV_X1 U9630 ( .A(n8343), .ZN(n8344) );
  NAND2_X1 U9631 ( .A1(n8345), .A2(n8344), .ZN(n9986) );
  INV_X1 U9632 ( .A(n9986), .ZN(n9771) );
  OR2_X1 U9633 ( .A1(n10093), .A2(n9771), .ZN(n8556) );
  NAND2_X1 U9634 ( .A1(n10093), .A2(n9771), .ZN(n8700) );
  NAND2_X1 U9635 ( .A1(n10093), .A2(n9986), .ZN(n8347) );
  NAND2_X1 U9636 ( .A1(n8348), .A2(n8546), .ZN(n8350) );
  NAND2_X1 U9637 ( .A1(n8421), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U9638 ( .A1(n8401), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8357) );
  NAND2_X1 U9639 ( .A1(n8541), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8356) );
  INV_X1 U9640 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8353) );
  INV_X1 U9641 ( .A(n8352), .ZN(n8351) );
  NAND2_X1 U9642 ( .A1(n8351), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8362) );
  AOI21_X1 U9643 ( .B1(n8353), .B2(n8352), .A(n8364), .ZN(n9948) );
  NAND2_X1 U9644 ( .A1(n5026), .A2(n9948), .ZN(n8355) );
  NAND2_X1 U9645 ( .A1(n6834), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8354) );
  NAND4_X1 U9646 ( .A1(n8357), .A2(n8356), .A3(n8355), .A4(n8354), .ZN(n9971)
         );
  OR2_X1 U9647 ( .A1(n10087), .A2(n9971), .ZN(n8358) );
  NAND2_X1 U9648 ( .A1(n8359), .A2(n8546), .ZN(n8361) );
  NAND2_X1 U9649 ( .A1(n8421), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U9650 ( .A1(n8541), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U9651 ( .A1(n8401), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8368) );
  INV_X1 U9652 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U9653 ( .A1(n8363), .A2(n8362), .ZN(n8365) );
  NAND2_X1 U9654 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n8364), .ZN(n8378) );
  AND2_X1 U9655 ( .A1(n8365), .A2(n8378), .ZN(n9936) );
  NAND2_X1 U9656 ( .A1(n5026), .A2(n9936), .ZN(n8367) );
  NAND2_X1 U9657 ( .A1(n6834), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8366) );
  NAND4_X1 U9658 ( .A1(n8369), .A2(n8368), .A3(n8367), .A4(n8366), .ZN(n9954)
         );
  OR2_X1 U9659 ( .A1(n10082), .A2(n9954), .ZN(n8370) );
  NAND2_X1 U9660 ( .A1(n9931), .A2(n8370), .ZN(n8372) );
  NAND2_X1 U9661 ( .A1(n10082), .A2(n9954), .ZN(n8371) );
  NAND2_X1 U9662 ( .A1(n8372), .A2(n8371), .ZN(n9913) );
  NAND2_X1 U9663 ( .A1(n8373), .A2(n8546), .ZN(n8375) );
  NAND2_X1 U9664 ( .A1(n8421), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U9665 ( .A1(n8401), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U9666 ( .A1(n8541), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8382) );
  INV_X1 U9667 ( .A(n8378), .ZN(n8376) );
  NAND2_X1 U9668 ( .A1(n8376), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8390) );
  INV_X1 U9669 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U9670 ( .A1(n8378), .A2(n8377), .ZN(n8379) );
  AND2_X1 U9671 ( .A1(n8390), .A2(n8379), .ZN(n9925) );
  NAND2_X1 U9672 ( .A1(n5026), .A2(n9925), .ZN(n8381) );
  NAND2_X1 U9673 ( .A1(n6834), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8380) );
  NAND4_X1 U9674 ( .A1(n8383), .A2(n8382), .A3(n8381), .A4(n8380), .ZN(n9942)
         );
  OR2_X1 U9675 ( .A1(n10078), .A2(n9942), .ZN(n8384) );
  NAND2_X1 U9676 ( .A1(n8385), .A2(n8546), .ZN(n8387) );
  NAND2_X1 U9677 ( .A1(n8421), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U9678 ( .A1(n8541), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U9679 ( .A1(n8401), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8394) );
  INV_X1 U9680 ( .A(n8390), .ZN(n8388) );
  NAND2_X1 U9681 ( .A1(n8388), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8404) );
  INV_X1 U9682 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U9683 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  AND2_X1 U9684 ( .A1(n8404), .A2(n8391), .ZN(n9902) );
  NAND2_X1 U9685 ( .A1(n5026), .A2(n9902), .ZN(n8393) );
  NAND2_X1 U9686 ( .A1(n6834), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8392) );
  NAND4_X1 U9687 ( .A1(n8395), .A2(n8394), .A3(n8393), .A4(n8392), .ZN(n9920)
         );
  INV_X1 U9688 ( .A(n9920), .ZN(n9794) );
  OR2_X1 U9689 ( .A1(n10072), .A2(n9794), .ZN(n8712) );
  NAND2_X1 U9690 ( .A1(n10072), .A2(n9794), .ZN(n8711) );
  NAND2_X1 U9691 ( .A1(n8712), .A2(n8711), .ZN(n8769) );
  OR2_X1 U9692 ( .A1(n10072), .A2(n9920), .ZN(n8396) );
  NAND2_X1 U9693 ( .A1(n8397), .A2(n8396), .ZN(n9885) );
  NAND2_X1 U9694 ( .A1(n8398), .A2(n8546), .ZN(n8400) );
  NAND2_X1 U9695 ( .A1(n8421), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U9696 ( .A1(n8541), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U9697 ( .A1(n8401), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8408) );
  INV_X1 U9698 ( .A(n8404), .ZN(n8402) );
  INV_X1 U9699 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U9700 ( .A1(n8404), .A2(n8403), .ZN(n8405) );
  NAND2_X1 U9701 ( .A1(n5026), .A2(n9887), .ZN(n8407) );
  NAND2_X1 U9702 ( .A1(n6834), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8406) );
  NAND4_X1 U9703 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n9908)
         );
  NOR2_X1 U9704 ( .A1(n10067), .A2(n9908), .ZN(n8410) );
  NAND2_X1 U9705 ( .A1(n10067), .A2(n9908), .ZN(n8411) );
  NAND2_X1 U9706 ( .A1(n8412), .A2(n8546), .ZN(n8414) );
  NAND2_X1 U9707 ( .A1(n8421), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U9708 ( .A1(n8401), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U9709 ( .A1(n6834), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U9710 ( .A(n8428), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U9711 ( .A1(n5026), .A2(n9878), .ZN(n8416) );
  NAND2_X1 U9712 ( .A1(n8541), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8415) );
  NAND4_X1 U9713 ( .A1(n8418), .A2(n8417), .A3(n8416), .A4(n8415), .ZN(n9893)
         );
  INV_X1 U9714 ( .A(n9893), .ZN(n8419) );
  NAND2_X1 U9715 ( .A1(n10062), .A2(n8419), .ZN(n8720) );
  NAND2_X1 U9716 ( .A1(n8420), .A2(n8546), .ZN(n8423) );
  NAND2_X1 U9717 ( .A1(n8421), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U9718 ( .A1(n8401), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U9719 ( .A1(n6834), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8432) );
  INV_X1 U9720 ( .A(n8428), .ZN(n8425) );
  AND2_X1 U9721 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n8424) );
  NAND2_X1 U9722 ( .A1(n8425), .A2(n8424), .ZN(n8469) );
  INV_X1 U9723 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8427) );
  INV_X1 U9724 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8426) );
  OAI21_X1 U9725 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(n8429) );
  NAND2_X1 U9726 ( .A1(n5026), .A2(n9164), .ZN(n8431) );
  NAND2_X1 U9727 ( .A1(n8541), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8430) );
  NAND4_X1 U9728 ( .A1(n8433), .A2(n8432), .A3(n8431), .A4(n8430), .ZN(n9870)
         );
  INV_X1 U9729 ( .A(n9870), .ZN(n9700) );
  OR2_X1 U9730 ( .A1(n10057), .A2(n9700), .ZN(n8549) );
  NAND2_X1 U9731 ( .A1(n10057), .A2(n9700), .ZN(n8725) );
  NAND2_X1 U9732 ( .A1(n8492), .A2(n8496), .ZN(n8494) );
  INV_X1 U9733 ( .A(n8439), .ZN(n8434) );
  AND2_X1 U9734 ( .A1(n8435), .A2(n8434), .ZN(n8436) );
  INV_X1 U9735 ( .A(n8440), .ZN(n8442) );
  INV_X1 U9736 ( .A(SI_28_), .ZN(n8441) );
  MUX2_X1 U9737 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5752), .Z(n8528) );
  INV_X1 U9738 ( .A(n8443), .ZN(n8445) );
  INV_X1 U9739 ( .A(SI_29_), .ZN(n8444) );
  NAND2_X1 U9740 ( .A1(n8445), .A2(n8444), .ZN(n8446) );
  NAND2_X1 U9741 ( .A1(n8531), .A2(n8446), .ZN(n10146) );
  NAND2_X1 U9742 ( .A1(n8421), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U9743 ( .A1(n8541), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U9744 ( .A1(n8401), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8453) );
  INV_X1 U9745 ( .A(n8469), .ZN(n8450) );
  NAND2_X1 U9746 ( .A1(n5026), .A2(n8450), .ZN(n8452) );
  NAND2_X1 U9747 ( .A1(n6834), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8451) );
  NAND4_X1 U9748 ( .A1(n8454), .A2(n8453), .A3(n8452), .A4(n8451), .ZN(n9801)
         );
  INV_X1 U9749 ( .A(n9801), .ZN(n8455) );
  NOR2_X1 U9750 ( .A1(n10112), .A2(n10018), .ZN(n8685) );
  INV_X1 U9751 ( .A(n8685), .ZN(n8679) );
  NAND2_X1 U9752 ( .A1(n10112), .A2(n10018), .ZN(n10012) );
  INV_X1 U9753 ( .A(n10012), .ZN(n8686) );
  NOR2_X1 U9754 ( .A1(n10017), .A2(n8686), .ZN(n8458) );
  NAND2_X1 U9755 ( .A1(n8689), .A2(n8685), .ZN(n8459) );
  AND2_X1 U9756 ( .A1(n8459), .A2(n8688), .ZN(n8553) );
  NAND2_X1 U9757 ( .A1(n9998), .A2(n9985), .ZN(n8694) );
  NAND2_X1 U9758 ( .A1(n8695), .A2(n8694), .ZN(n9992) );
  NAND2_X1 U9759 ( .A1(n5646), .A2(n8460), .ZN(n9999) );
  NAND2_X1 U9760 ( .A1(n9999), .A2(n8695), .ZN(n9983) );
  NAND2_X1 U9761 ( .A1(n9983), .A2(n9984), .ZN(n9982) );
  NAND2_X1 U9762 ( .A1(n9982), .A2(n8551), .ZN(n9969) );
  NAND2_X1 U9763 ( .A1(n9969), .A2(n9970), .ZN(n9968) );
  NAND2_X1 U9764 ( .A1(n9968), .A2(n8700), .ZN(n9952) );
  INV_X1 U9765 ( .A(n9971), .ZN(n9711) );
  NAND2_X1 U9766 ( .A1(n10087), .A2(n9711), .ZN(n8619) );
  INV_X1 U9767 ( .A(n9954), .ZN(n9122) );
  OR2_X1 U9768 ( .A1(n10082), .A2(n9122), .ZN(n8550) );
  NAND2_X1 U9769 ( .A1(n10082), .A2(n9122), .ZN(n8624) );
  NAND2_X1 U9770 ( .A1(n8550), .A2(n8624), .ZN(n9932) );
  INV_X1 U9771 ( .A(n9932), .ZN(n9941) );
  INV_X1 U9772 ( .A(n9942), .ZN(n9127) );
  OR2_X1 U9773 ( .A1(n10078), .A2(n9127), .ZN(n8706) );
  NAND2_X1 U9774 ( .A1(n10078), .A2(n9127), .ZN(n8707) );
  NAND2_X1 U9775 ( .A1(n8706), .A2(n8707), .ZN(n9915) );
  INV_X1 U9776 ( .A(n9915), .ZN(n9919) );
  INV_X1 U9777 ( .A(n9908), .ZN(n9740) );
  OR2_X1 U9778 ( .A1(n10067), .A2(n9740), .ZN(n8718) );
  XNOR2_X1 U9779 ( .A(n8462), .B(n8461), .ZN(n8468) );
  NAND2_X1 U9780 ( .A1(n9870), .A2(n10993), .ZN(n8466) );
  INV_X1 U9781 ( .A(n10675), .ZN(n9819) );
  NAND2_X1 U9782 ( .A1(n9819), .A2(P1_B_REG_SCAN_IN), .ZN(n8463) );
  AND2_X1 U9783 ( .A1(n10990), .A2(n8463), .ZN(n9854) );
  NAND2_X1 U9784 ( .A1(n9854), .A2(n8464), .ZN(n8465) );
  AOI21_X2 U9785 ( .B1(n8468), .B2(n10998), .A(n8467), .ZN(n10055) );
  OAI21_X1 U9786 ( .B1(n8469), .B2(n10879), .A(n10055), .ZN(n8470) );
  NAND2_X1 U9787 ( .A1(n8470), .A2(n11019), .ZN(n8476) );
  INV_X1 U9788 ( .A(n10072), .ZN(n9904) );
  INV_X1 U9789 ( .A(n10093), .ZN(n9967) );
  INV_X1 U9790 ( .A(n10107), .ZN(n10011) );
  NAND2_X1 U9791 ( .A1(n10008), .A2(n9998), .ZN(n9993) );
  NAND2_X1 U9792 ( .A1(n9904), .A2(n9924), .ZN(n9899) );
  INV_X1 U9793 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8472) );
  OAI22_X1 U9794 ( .A1(n8473), .A2(n11016), .B1(n8472), .B2(n11019), .ZN(n8474) );
  AOI21_X1 U9795 ( .B1(n5042), .B2(n11009), .A(n8474), .ZN(n8475) );
  OAI211_X1 U9796 ( .C1(n10056), .C2(n10025), .A(n8476), .B(n8475), .ZN(
        P1_U3355) );
  NAND2_X1 U9797 ( .A1(n10617), .A2(n10612), .ZN(n8478) );
  OAI211_X1 U9798 ( .C1(n7559), .C2(n9314), .A(n8478), .B(n8477), .ZN(n8481)
         );
  NOR2_X1 U9799 ( .A1(n9294), .A2(n8479), .ZN(n8480) );
  AOI211_X1 U9800 ( .C1(n10611), .C2(n8916), .A(n8481), .B(n8480), .ZN(n8490)
         );
  NAND2_X1 U9801 ( .A1(n8482), .A2(n8483), .ZN(n8484) );
  NAND2_X1 U9802 ( .A1(n8484), .A2(n9057), .ZN(n9061) );
  OAI22_X1 U9803 ( .A1(n9306), .A2(n8487), .B1(n10607), .B2(n8486), .ZN(n8488)
         );
  NAND3_X1 U9804 ( .A1(n9061), .A2(n5908), .A3(n8488), .ZN(n8489) );
  OAI211_X1 U9805 ( .C1(n8491), .C2(n9306), .A(n8490), .B(n8489), .ZN(P2_U3241) );
  INV_X1 U9806 ( .A(n8492), .ZN(n8493) );
  NAND2_X1 U9807 ( .A1(n8493), .A2(n8771), .ZN(n8495) );
  NAND2_X1 U9808 ( .A1(n8497), .A2(n8496), .ZN(n8498) );
  NAND2_X1 U9809 ( .A1(n8499), .A2(n8498), .ZN(n8500) );
  NAND2_X1 U9810 ( .A1(n8500), .A2(n10998), .ZN(n8502) );
  AOI22_X1 U9811 ( .A1(n10993), .A2(n9893), .B1(n9801), .B2(n10990), .ZN(n8501) );
  AOI21_X1 U9812 ( .B1(n10057), .B2(n9877), .A(n8503), .ZN(n10058) );
  AOI22_X1 U9813 ( .A1(n11014), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9164), .B2(
        n11012), .ZN(n8504) );
  OAI21_X1 U9814 ( .B1(n5220), .B2(n11016), .A(n8504), .ZN(n8507) );
  NOR2_X1 U9815 ( .A1(n10061), .A2(n10042), .ZN(n8506) );
  OAI21_X1 U9816 ( .B1(n10060), .B2(n11014), .A(n8508), .ZN(P1_U3263) );
  OAI21_X1 U9817 ( .B1(n9314), .B2(n8511), .A(n8510), .ZN(n8512) );
  AOI21_X1 U9818 ( .B1(n10617), .B2(n9324), .A(n8512), .ZN(n8513) );
  OAI21_X1 U9819 ( .B1(n8514), .B2(n9294), .A(n8513), .ZN(n8515) );
  AOI21_X1 U9820 ( .B1(n11101), .B2(n10611), .A(n8515), .ZN(n8523) );
  INV_X1 U9821 ( .A(n8517), .ZN(n8521) );
  OAI22_X1 U9822 ( .A1(n8519), .A2(n9306), .B1(n8518), .B2(n10607), .ZN(n8520)
         );
  NAND3_X1 U9823 ( .A1(n8516), .A2(n8521), .A3(n8520), .ZN(n8522) );
  OAI211_X1 U9824 ( .C1(n8509), .C2(n9306), .A(n8523), .B(n8522), .ZN(P2_U3217) );
  NOR4_X1 U9825 ( .A1(n10028), .A2(n10151), .A3(n8524), .A4(n10675), .ZN(n8812) );
  INV_X1 U9826 ( .A(n8808), .ZN(n8526) );
  OAI21_X1 U9827 ( .B1(n8525), .B2(n8526), .A(P1_B_REG_SCAN_IN), .ZN(n8811) );
  INV_X1 U9828 ( .A(n8527), .ZN(n8529) );
  NAND2_X1 U9829 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  MUX2_X1 U9830 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5752), .Z(n8532) );
  NAND2_X1 U9831 ( .A1(n8532), .A2(SI_30_), .ZN(n8534) );
  OAI21_X1 U9832 ( .B1(n8532), .B2(SI_30_), .A(n8534), .ZN(n8545) );
  INV_X1 U9833 ( .A(n8545), .ZN(n8533) );
  MUX2_X1 U9834 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5752), .Z(n8536) );
  XNOR2_X1 U9835 ( .A(n8536), .B(SI_31_), .ZN(n8537) );
  NAND2_X1 U9836 ( .A1(n9678), .A2(n8546), .ZN(n8540) );
  NAND2_X1 U9837 ( .A1(n8421), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U9838 ( .A1(n8541), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U9839 ( .A1(n8401), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U9840 ( .A1(n6834), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8542) );
  AND2_X1 U9841 ( .A1(n9852), .A2(n9856), .ZN(n8793) );
  NAND2_X1 U9842 ( .A1(n9171), .A2(n8546), .ZN(n8548) );
  NAND2_X1 U9843 ( .A1(n8421), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8547) );
  NOR2_X1 U9844 ( .A1(n10049), .A2(n8614), .ZN(n8794) );
  NOR2_X1 U9845 ( .A1(n8793), .A2(n8794), .ZN(n8775) );
  INV_X1 U9846 ( .A(n8791), .ZN(n8721) );
  INV_X1 U9847 ( .A(n9868), .ZN(n9880) );
  AND2_X1 U9848 ( .A1(n8718), .A2(n8712), .ZN(n8782) );
  AND2_X1 U9849 ( .A1(n8706), .A2(n8550), .ZN(n8618) );
  NAND2_X1 U9850 ( .A1(n8700), .A2(n8551), .ZN(n8552) );
  NAND2_X1 U9851 ( .A1(n8552), .A2(n8556), .ZN(n8625) );
  NAND3_X1 U9852 ( .A1(n8619), .A2(n8625), .A3(n8695), .ZN(n8603) );
  AND2_X1 U9853 ( .A1(n8553), .A2(n8694), .ZN(n8554) );
  OR2_X1 U9854 ( .A1(n8603), .A2(n8554), .ZN(n8559) );
  NAND2_X1 U9855 ( .A1(n8556), .A2(n8555), .ZN(n8701) );
  NAND3_X1 U9856 ( .A1(n8619), .A2(n8625), .A3(n8701), .ZN(n8557) );
  AND2_X1 U9857 ( .A1(n8557), .A2(n8620), .ZN(n8558) );
  NAND2_X1 U9858 ( .A1(n8559), .A2(n8558), .ZN(n8605) );
  AND2_X1 U9859 ( .A1(n10012), .A2(n8680), .ZN(n8560) );
  NAND2_X1 U9860 ( .A1(n8689), .A2(n8560), .ZN(n8599) );
  NAND2_X1 U9861 ( .A1(n8673), .A2(n8670), .ZN(n8598) );
  AND2_X1 U9862 ( .A1(n8663), .A2(n8563), .ZN(n8660) );
  OAI21_X1 U9863 ( .B1(n8656), .B2(n8561), .A(n8660), .ZN(n8568) );
  AND3_X1 U9864 ( .A1(n8563), .A2(n8646), .A3(n8562), .ZN(n8564) );
  NAND2_X1 U9865 ( .A1(n8663), .A2(n8564), .ZN(n8596) );
  AND2_X1 U9866 ( .A1(n8649), .A2(n8565), .ZN(n8593) );
  AND2_X1 U9867 ( .A1(n8649), .A2(n8643), .ZN(n8566) );
  OR3_X1 U9868 ( .A1(n8596), .A2(n8593), .A3(n8566), .ZN(n8567) );
  AND4_X1 U9869 ( .A1(n8568), .A2(n8661), .A3(n8662), .A4(n8567), .ZN(n8569)
         );
  OAI211_X1 U9870 ( .C1(n8598), .C2(n8569), .A(n8681), .B(n8674), .ZN(n8570)
         );
  INV_X1 U9871 ( .A(n8570), .ZN(n8571) );
  OR2_X1 U9872 ( .A1(n8599), .A2(n8571), .ZN(n8601) );
  NAND2_X1 U9873 ( .A1(n8601), .A2(n8632), .ZN(n8572) );
  NOR2_X1 U9874 ( .A1(n8605), .A2(n8572), .ZN(n8573) );
  NAND2_X1 U9875 ( .A1(n8618), .A2(n8573), .ZN(n8781) );
  NAND2_X1 U9876 ( .A1(n7085), .A2(n10824), .ZN(n8574) );
  NAND3_X1 U9877 ( .A1(n8575), .A2(n6636), .A3(n8574), .ZN(n8576) );
  NAND2_X1 U9878 ( .A1(n8577), .A2(n8576), .ZN(n8580) );
  NAND2_X1 U9879 ( .A1(n10863), .A2(n10842), .ZN(n8578) );
  OAI211_X1 U9880 ( .C1(n8581), .C2(n8580), .A(n8579), .B(n8578), .ZN(n8585)
         );
  INV_X1 U9881 ( .A(n8582), .ZN(n8584) );
  NAND3_X1 U9882 ( .A1(n8585), .A2(n8584), .A3(n8583), .ZN(n8587) );
  NAND2_X1 U9883 ( .A1(n8587), .A2(n8586), .ZN(n8590) );
  NAND3_X1 U9884 ( .A1(n8590), .A2(n8589), .A3(n8588), .ZN(n8592) );
  NAND2_X1 U9885 ( .A1(n8592), .A2(n8591), .ZN(n8608) );
  NAND2_X1 U9886 ( .A1(n8711), .A2(n8707), .ZN(n8784) );
  INV_X1 U9887 ( .A(n8784), .ZN(n8607) );
  INV_X1 U9888 ( .A(n8593), .ZN(n8594) );
  NAND3_X1 U9889 ( .A1(n8594), .A2(n8639), .A3(n10996), .ZN(n8595) );
  OR2_X1 U9890 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  OR3_X1 U9891 ( .A1(n8599), .A2(n8598), .A3(n8597), .ZN(n8600) );
  AND2_X1 U9892 ( .A1(n8601), .A2(n8600), .ZN(n8602) );
  NOR2_X1 U9893 ( .A1(n8603), .A2(n8602), .ZN(n8604) );
  OAI21_X1 U9894 ( .B1(n8605), .B2(n8604), .A(n8624), .ZN(n8606) );
  NAND2_X1 U9895 ( .A1(n8618), .A2(n8606), .ZN(n8779) );
  OAI211_X1 U9896 ( .C1(n8781), .C2(n8608), .A(n8607), .B(n8779), .ZN(n8609)
         );
  NAND2_X1 U9897 ( .A1(n8782), .A2(n8609), .ZN(n8611) );
  NAND2_X1 U9898 ( .A1(n8778), .A2(n8610), .ZN(n8785) );
  OAI21_X1 U9899 ( .B1(n9880), .B2(n8611), .A(n8785), .ZN(n8613) );
  AND2_X1 U9900 ( .A1(n8725), .A2(n8720), .ZN(n8786) );
  INV_X1 U9901 ( .A(n8786), .ZN(n8612) );
  NOR2_X1 U9902 ( .A1(n8613), .A2(n8612), .ZN(n8615) );
  NAND2_X1 U9903 ( .A1(n10049), .A2(n8614), .ZN(n8745) );
  OAI211_X1 U9904 ( .C1(n8721), .C2(n8615), .A(n8745), .B(n8726), .ZN(n8616)
         );
  INV_X1 U9905 ( .A(n9856), .ZN(n9800) );
  AOI21_X1 U9906 ( .B1(n8775), .B2(n8616), .A(n8796), .ZN(n8617) );
  XNOR2_X1 U9907 ( .A(n8617), .B(n9850), .ZN(n8803) );
  INV_X1 U9908 ( .A(n8618), .ZN(n8627) );
  INV_X1 U9909 ( .A(n8619), .ZN(n8622) );
  INV_X1 U9910 ( .A(n8620), .ZN(n8621) );
  MUX2_X1 U9911 ( .A(n8622), .B(n8621), .S(n8735), .Z(n8623) );
  OR2_X1 U9912 ( .A1(n9932), .A2(n8623), .ZN(n8705) );
  OAI211_X1 U9913 ( .C1(n8705), .C2(n8625), .A(n8624), .B(n8707), .ZN(n8626)
         );
  MUX2_X1 U9914 ( .A(n8627), .B(n8626), .S(n8735), .Z(n8710) );
  INV_X1 U9915 ( .A(n8628), .ZN(n8629) );
  INV_X1 U9916 ( .A(n8735), .ZN(n8741) );
  XNOR2_X1 U9917 ( .A(n8629), .B(n8741), .ZN(n8630) );
  NAND2_X1 U9918 ( .A1(n8630), .A2(n8751), .ZN(n8636) );
  NAND2_X1 U9919 ( .A1(n8636), .A2(n9810), .ZN(n8631) );
  AOI21_X1 U9920 ( .B1(n8631), .B2(n8632), .A(n5386), .ZN(n8655) );
  NAND3_X1 U9921 ( .A1(n8632), .A2(n8741), .A3(n10935), .ZN(n8633) );
  OAI21_X1 U9922 ( .B1(n8754), .B2(n8634), .A(n8633), .ZN(n8635) );
  NAND2_X1 U9923 ( .A1(n8636), .A2(n8635), .ZN(n8653) );
  AND2_X1 U9924 ( .A1(n8637), .A2(n8735), .ZN(n8641) );
  NAND4_X1 U9925 ( .A1(n8653), .A2(n8641), .A3(n8649), .A4(n8638), .ZN(n8654)
         );
  AND4_X1 U9926 ( .A1(n8645), .A2(n8741), .A3(n8639), .A4(n10996), .ZN(n8640)
         );
  AND2_X1 U9927 ( .A1(n8646), .A2(n8640), .ZN(n8652) );
  NAND2_X1 U9928 ( .A1(n8649), .A2(n8641), .ZN(n8642) );
  AOI21_X1 U9929 ( .B1(n8645), .B2(n10996), .A(n8642), .ZN(n8651) );
  NAND4_X1 U9930 ( .A1(n8646), .A2(n8741), .A3(n8645), .A4(n8644), .ZN(n8648)
         );
  OR2_X1 U9931 ( .A1(n8646), .A2(n8741), .ZN(n8647) );
  OAI211_X1 U9932 ( .C1(n8649), .C2(n8735), .A(n8648), .B(n8647), .ZN(n8650)
         );
  MUX2_X1 U9933 ( .A(n8657), .B(n8656), .S(n8735), .Z(n8658) );
  NOR2_X1 U9934 ( .A1(n8760), .A2(n8658), .ZN(n8659) );
  NAND2_X1 U9935 ( .A1(n8669), .A2(n8661), .ZN(n8672) );
  INV_X1 U9936 ( .A(n8662), .ZN(n8668) );
  INV_X1 U9937 ( .A(n8663), .ZN(n8664) );
  AOI21_X1 U9938 ( .B1(n8666), .B2(n8665), .A(n8664), .ZN(n8667) );
  MUX2_X1 U9939 ( .A(n8672), .B(n8671), .S(n8741), .Z(n8678) );
  INV_X1 U9940 ( .A(n8673), .ZN(n8676) );
  INV_X1 U9941 ( .A(n8674), .ZN(n8675) );
  MUX2_X1 U9942 ( .A(n8676), .B(n8675), .S(n8735), .Z(n8677) );
  AOI21_X1 U9943 ( .B1(n8678), .B2(n8763), .A(n8677), .ZN(n8684) );
  NAND2_X1 U9944 ( .A1(n8679), .A2(n10012), .ZN(n10033) );
  INV_X1 U9945 ( .A(n10033), .ZN(n10026) );
  MUX2_X1 U9946 ( .A(n8681), .B(n8680), .S(n8741), .Z(n8682) );
  OAI211_X1 U9947 ( .C1(n8684), .C2(n8683), .A(n10026), .B(n8682), .ZN(n8693)
         );
  MUX2_X1 U9948 ( .A(n8686), .B(n8685), .S(n8741), .Z(n8687) );
  NOR2_X1 U9949 ( .A1(n10017), .A2(n8687), .ZN(n8692) );
  MUX2_X1 U9950 ( .A(n8689), .B(n8688), .S(n8735), .Z(n8690) );
  NAND2_X1 U9951 ( .A1(n8460), .A2(n8690), .ZN(n8691) );
  AOI21_X1 U9952 ( .B1(n8693), .B2(n8692), .A(n8691), .ZN(n8699) );
  INV_X1 U9953 ( .A(n8694), .ZN(n8697) );
  INV_X1 U9954 ( .A(n8695), .ZN(n8696) );
  MUX2_X1 U9955 ( .A(n8697), .B(n8696), .S(n8735), .Z(n8698) );
  OAI211_X1 U9956 ( .C1(n8699), .C2(n8698), .A(n9970), .B(n9984), .ZN(n8703)
         );
  NAND3_X1 U9957 ( .A1(n8701), .A2(n8741), .A3(n8700), .ZN(n8702) );
  AND3_X1 U9958 ( .A1(n9953), .A2(n8703), .A3(n8702), .ZN(n8704) );
  NOR2_X1 U9959 ( .A1(n8705), .A2(n8704), .ZN(n8709) );
  MUX2_X1 U9960 ( .A(n8707), .B(n8706), .S(n8735), .Z(n8708) );
  OAI211_X1 U9961 ( .C1(n8710), .C2(n8709), .A(n9907), .B(n8708), .ZN(n8717)
         );
  INV_X1 U9962 ( .A(n8711), .ZN(n8714) );
  INV_X1 U9963 ( .A(n8712), .ZN(n8713) );
  MUX2_X1 U9964 ( .A(n8714), .B(n8713), .S(n8741), .Z(n8715) );
  INV_X1 U9965 ( .A(n8715), .ZN(n8716) );
  MUX2_X1 U9966 ( .A(n9867), .B(n8718), .S(n8735), .Z(n8719) );
  INV_X1 U9967 ( .A(n8720), .ZN(n8722) );
  NAND2_X1 U9968 ( .A1(n8723), .A2(n8726), .ZN(n8730) );
  NAND3_X1 U9969 ( .A1(n8726), .A2(n8725), .A3(n8724), .ZN(n8728) );
  NAND2_X1 U9970 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  NAND2_X1 U9971 ( .A1(n8794), .A2(n9852), .ZN(n8731) );
  INV_X1 U9972 ( .A(n8793), .ZN(n8736) );
  AND2_X1 U9973 ( .A1(n8731), .A2(n8736), .ZN(n8740) );
  NAND2_X1 U9974 ( .A1(n10049), .A2(n9856), .ZN(n8732) );
  NAND2_X1 U9975 ( .A1(n8745), .A2(n8732), .ZN(n8788) );
  NAND2_X1 U9976 ( .A1(n8736), .A2(n8735), .ZN(n8737) );
  NAND2_X1 U9977 ( .A1(n8737), .A2(n8788), .ZN(n8738) );
  INV_X1 U9978 ( .A(n8740), .ZN(n8742) );
  NAND2_X1 U9979 ( .A1(n8742), .A2(n8741), .ZN(n8743) );
  INV_X1 U9980 ( .A(n8796), .ZN(n8804) );
  INV_X1 U9981 ( .A(n8745), .ZN(n8774) );
  NOR4_X1 U9982 ( .A1(n8748), .A2(n10860), .A3(n8747), .A4(n8746), .ZN(n8752)
         );
  NAND4_X1 U9983 ( .A1(n8751), .A2(n8752), .A3(n8750), .A4(n8749), .ZN(n8755)
         );
  NOR4_X1 U9984 ( .A1(n8755), .A2(n10995), .A3(n8754), .A4(n8753), .ZN(n8757)
         );
  NAND2_X1 U9985 ( .A1(n8757), .A2(n8756), .ZN(n8759) );
  NOR4_X1 U9986 ( .A1(n8761), .A2(n8760), .A3(n8759), .A4(n8758), .ZN(n8762)
         );
  NAND4_X1 U9987 ( .A1(n8765), .A2(n8764), .A3(n8763), .A4(n8762), .ZN(n8766)
         );
  NOR4_X1 U9988 ( .A1(n9992), .A2(n10017), .A3(n10033), .A4(n8766), .ZN(n8767)
         );
  NAND4_X1 U9989 ( .A1(n9953), .A2(n9970), .A3(n9984), .A4(n8767), .ZN(n8768)
         );
  NOR4_X1 U9990 ( .A1(n8769), .A2(n9915), .A3(n9932), .A4(n8768), .ZN(n8770)
         );
  NAND4_X1 U9991 ( .A1(n8771), .A2(n9892), .A3(n9868), .A4(n8770), .ZN(n8772)
         );
  AOI21_X1 U9992 ( .B1(n8776), .B2(n8775), .A(n6636), .ZN(n8798) );
  OAI21_X1 U9993 ( .B1(n8781), .B2(n8780), .A(n8779), .ZN(n8783) );
  OAI21_X1 U9994 ( .B1(n8784), .B2(n8783), .A(n8782), .ZN(n8787) );
  OAI211_X1 U9995 ( .C1(n5208), .C2(n8787), .A(n8786), .B(n8785), .ZN(n8790)
         );
  AOI211_X1 U9996 ( .C1(n8791), .C2(n8790), .A(n8789), .B(n8788), .ZN(n8792)
         );
  AOI211_X1 U9997 ( .C1(n8794), .C2(n9800), .A(n8793), .B(n8792), .ZN(n8797)
         );
  NOR3_X1 U9998 ( .A1(n8797), .A2(n8796), .A3(n8795), .ZN(n8799) );
  NOR2_X1 U9999 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  AND4_X1 U10000 ( .A1(n8807), .A2(n8806), .A3(n8805), .A4(n8804), .ZN(n8809)
         );
  INV_X1 U10001 ( .A(n8870), .ZN(n8967) );
  NAND2_X1 U10002 ( .A1(n8813), .A2(n8967), .ZN(n8815) );
  INV_X1 U10003 ( .A(n9573), .ZN(n9291) );
  OR2_X1 U10004 ( .A1(n9653), .A2(n9291), .ZN(n8814) );
  NAND2_X1 U10005 ( .A1(n8815), .A2(n8814), .ZN(n9570) );
  XNOR2_X1 U10006 ( .A(n9645), .B(n9547), .ZN(n9571) );
  INV_X1 U10007 ( .A(n9571), .ZN(n9561) );
  OR2_X1 U10008 ( .A1(n9645), .A2(n9547), .ZN(n8816) );
  NAND2_X1 U10009 ( .A1(n9642), .A2(n9273), .ZN(n8976) );
  NAND2_X1 U10010 ( .A1(n8977), .A2(n8976), .ZN(n9539) );
  INV_X1 U10011 ( .A(n9539), .ZN(n9543) );
  XNOR2_X1 U10012 ( .A(n9635), .B(n9549), .ZN(n9531) );
  INV_X1 U10013 ( .A(n9531), .ZN(n8871) );
  NAND2_X1 U10014 ( .A1(n9532), .A2(n8871), .ZN(n8818) );
  OR2_X1 U10015 ( .A1(n9635), .A2(n9549), .ZN(n8817) );
  NAND2_X1 U10016 ( .A1(n8818), .A2(n8817), .ZN(n9516) );
  NAND2_X1 U10017 ( .A1(n9630), .A2(n9533), .ZN(n8987) );
  NAND2_X1 U10018 ( .A1(n8988), .A2(n8987), .ZN(n9517) );
  NAND2_X1 U10019 ( .A1(n9516), .A2(n9517), .ZN(n8820) );
  INV_X1 U10020 ( .A(n9533), .ZN(n9275) );
  OR2_X1 U10021 ( .A1(n9630), .A2(n9275), .ZN(n8819) );
  NAND2_X1 U10022 ( .A1(n8820), .A2(n8819), .ZN(n9502) );
  NAND2_X1 U10023 ( .A1(n9502), .A2(n9182), .ZN(n8821) );
  INV_X1 U10024 ( .A(n9519), .ZN(n9224) );
  OR2_X1 U10025 ( .A1(n9625), .A2(n9224), .ZN(n8992) );
  OR2_X1 U10026 ( .A1(n9620), .A2(n9284), .ZN(n8996) );
  NAND2_X1 U10027 ( .A1(n9620), .A2(n9284), .ZN(n9474) );
  NAND2_X1 U10028 ( .A1(n9615), .A2(n9261), .ZN(n8998) );
  NAND2_X1 U10029 ( .A1(n8997), .A2(n8998), .ZN(n9476) );
  INV_X1 U10030 ( .A(n9474), .ZN(n8822) );
  NOR2_X1 U10031 ( .A1(n9476), .A2(n8822), .ZN(n8823) );
  NAND2_X1 U10032 ( .A1(n9611), .A2(n9442), .ZN(n9007) );
  NAND2_X1 U10033 ( .A1(n9006), .A2(n9007), .ZN(n9461) );
  INV_X1 U10034 ( .A(n9461), .ZN(n9453) );
  NAND2_X1 U10035 ( .A1(n9462), .A2(n9453), .ZN(n8824) );
  NAND2_X1 U10036 ( .A1(n8824), .A2(n9006), .ZN(n9440) );
  NAND2_X1 U10037 ( .A1(n9607), .A2(n9250), .ZN(n9012) );
  NAND2_X1 U10038 ( .A1(n9440), .A2(n9012), .ZN(n8825) );
  NAND2_X1 U10039 ( .A1(n8825), .A2(n9011), .ZN(n9428) );
  NAND2_X1 U10040 ( .A1(n9600), .A2(n9443), .ZN(n9016) );
  NAND2_X1 U10041 ( .A1(n9428), .A2(n9427), .ZN(n9426) );
  NAND2_X1 U10042 ( .A1(n5934), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U10043 ( .A1(n9589), .A2(n8829), .ZN(n9023) );
  NAND2_X1 U10044 ( .A1(n9191), .A2(n9412), .ZN(n9022) );
  NAND2_X1 U10045 ( .A1(n8830), .A2(n9022), .ZN(n8845) );
  INV_X1 U10046 ( .A(n8845), .ZN(n8847) );
  NAND2_X1 U10047 ( .A1(n9171), .A2(n8848), .ZN(n8833) );
  NAND2_X1 U10048 ( .A1(n8831), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8832) );
  INV_X1 U10049 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U10050 ( .A1(n8834), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U10051 ( .A1(n5921), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8835) );
  OAI211_X1 U10052 ( .C1(n8842), .C2(n8837), .A(n8836), .B(n8835), .ZN(n9320)
         );
  INV_X1 U10053 ( .A(n9320), .ZN(n8850) );
  NOR2_X1 U10054 ( .A1(n9400), .A2(n8850), .ZN(n8855) );
  INV_X1 U10055 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U10056 ( .A1(n5921), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8840) );
  INV_X1 U10057 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8838) );
  OR2_X1 U10058 ( .A1(n5922), .A2(n8838), .ZN(n8839) );
  OAI211_X1 U10059 ( .C1(n8842), .C2(n8841), .A(n8840), .B(n8839), .ZN(n9394)
         );
  OR2_X1 U10060 ( .A1(n9394), .A2(n8843), .ZN(n8844) );
  OAI21_X1 U10061 ( .B1(n8847), .B2(n9400), .A(n8846), .ZN(n8853) );
  NAND2_X1 U10062 ( .A1(n5934), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8849) );
  INV_X1 U10063 ( .A(n9394), .ZN(n9029) );
  NAND2_X1 U10064 ( .A1(n9400), .A2(n8850), .ZN(n9024) );
  AND2_X1 U10065 ( .A1(n8851), .A2(n9029), .ZN(n8854) );
  INV_X1 U10066 ( .A(n8854), .ZN(n8856) );
  INV_X1 U10067 ( .A(n8855), .ZN(n9025) );
  NAND2_X1 U10068 ( .A1(n8856), .A2(n9025), .ZN(n8882) );
  NAND2_X1 U10069 ( .A1(n9022), .A2(n9023), .ZN(n9193) );
  NAND2_X1 U10070 ( .A1(n9011), .A2(n9012), .ZN(n9437) );
  INV_X1 U10071 ( .A(n9437), .ZN(n9439) );
  NOR3_X1 U10072 ( .A1(n8884), .A2(n8885), .A3(n8307), .ZN(n8859) );
  INV_X1 U10073 ( .A(n8857), .ZN(n8906) );
  NAND4_X1 U10074 ( .A1(n8859), .A2(n8906), .A3(n7263), .A4(n8858), .ZN(n8863)
         );
  NOR4_X1 U10075 ( .A1(n8863), .A2(n8862), .A3(n8861), .A4(n8860), .ZN(n8865)
         );
  NAND4_X1 U10076 ( .A1(n8865), .A2(n8923), .A3(n8864), .A4(n7753), .ZN(n8867)
         );
  NOR4_X1 U10077 ( .A1(n8867), .A2(n8946), .A3(n5370), .A4(n8866), .ZN(n8868)
         );
  NAND4_X1 U10078 ( .A1(n8963), .A2(n8953), .A3(n8958), .A4(n8868), .ZN(n8869)
         );
  NOR4_X1 U10079 ( .A1(n9539), .A2(n9571), .A3(n8870), .A4(n8869), .ZN(n8872)
         );
  NAND4_X1 U10080 ( .A1(n9490), .A2(n8872), .A3(n8871), .A4(n9517), .ZN(n8873)
         );
  NOR4_X1 U10081 ( .A1(n9461), .A2(n8873), .A3(n9476), .A4(n9503), .ZN(n8874)
         );
  NAND4_X1 U10082 ( .A1(n5345), .A2(n9439), .A3(n9427), .A4(n8874), .ZN(n8875)
         );
  NOR4_X1 U10083 ( .A1(n8882), .A2(n8883), .A3(n9193), .A4(n8875), .ZN(n8876)
         );
  XNOR2_X1 U10084 ( .A(n8876), .B(n9555), .ZN(n8878) );
  OAI22_X1 U10085 ( .A1(n8878), .A2(n8891), .B1(n8877), .B2(n9033), .ZN(n9037)
         );
  NOR2_X1 U10086 ( .A1(n10922), .A2(n8880), .ZN(n8881) );
  NAND2_X2 U10087 ( .A1(n8881), .A2(n9033), .ZN(n9028) );
  MUX2_X1 U10088 ( .A(n8883), .B(n8882), .S(n9028), .Z(n9032) );
  INV_X1 U10089 ( .A(n8884), .ZN(n8887) );
  INV_X1 U10090 ( .A(n8885), .ZN(n8886) );
  NAND3_X1 U10091 ( .A1(n8887), .A2(n7263), .A3(n8886), .ZN(n8888) );
  NAND2_X1 U10092 ( .A1(n8889), .A2(n8888), .ZN(n8895) );
  NAND3_X1 U10093 ( .A1(n8892), .A2(n8891), .A3(n8890), .ZN(n8893) );
  OAI21_X1 U10094 ( .B1(n8897), .B2(n9028), .A(n8896), .ZN(n8901) );
  MUX2_X1 U10095 ( .A(n7347), .B(n8898), .S(n9028), .Z(n8899) );
  OAI21_X1 U10096 ( .B1(n10886), .B2(n10605), .A(n8899), .ZN(n8900) );
  OAI21_X1 U10097 ( .B1(n8902), .B2(n8901), .A(n8900), .ZN(n8909) );
  NAND2_X1 U10098 ( .A1(n8909), .A2(n5356), .ZN(n8905) );
  MUX2_X1 U10099 ( .A(n10610), .B(n9054), .S(n9028), .Z(n8904) );
  NAND2_X1 U10100 ( .A1(n8905), .A2(n8904), .ZN(n8907) );
  OAI211_X1 U10101 ( .C1(n8909), .C2(n8908), .A(n8907), .B(n8906), .ZN(n8913)
         );
  MUX2_X1 U10102 ( .A(n8911), .B(n8910), .S(n9028), .Z(n8912) );
  NAND2_X1 U10103 ( .A1(n8913), .A2(n8912), .ZN(n8919) );
  MUX2_X1 U10104 ( .A(n9331), .B(n8916), .S(n9028), .Z(n8917) );
  MUX2_X1 U10105 ( .A(n8921), .B(n8920), .S(n9028), .Z(n8922) );
  INV_X1 U10106 ( .A(n9028), .ZN(n9010) );
  MUX2_X1 U10107 ( .A(n8925), .B(n8924), .S(n9010), .Z(n8926) );
  AND2_X1 U10108 ( .A1(n8931), .A2(n8932), .ZN(n8927) );
  MUX2_X1 U10109 ( .A(n8928), .B(n8927), .S(n9028), .Z(n8929) );
  OAI211_X1 U10110 ( .C1(n5090), .C2(n8932), .A(n8931), .B(n8930), .ZN(n8936)
         );
  NAND2_X1 U10111 ( .A1(n8934), .A2(n8933), .ZN(n8935) );
  MUX2_X1 U10112 ( .A(n8936), .B(n8935), .S(n9028), .Z(n8937) );
  INV_X1 U10113 ( .A(n8937), .ZN(n8938) );
  NAND3_X1 U10114 ( .A1(n8940), .A2(n8939), .A3(n8938), .ZN(n8949) );
  INV_X1 U10115 ( .A(n8941), .ZN(n8942) );
  NOR2_X1 U10116 ( .A1(n8943), .A2(n8942), .ZN(n8944) );
  MUX2_X1 U10117 ( .A(n8945), .B(n8944), .S(n9028), .Z(n8947) );
  NOR2_X1 U10118 ( .A1(n8947), .A2(n8946), .ZN(n8948) );
  NAND2_X1 U10119 ( .A1(n8949), .A2(n8948), .ZN(n8954) );
  MUX2_X1 U10120 ( .A(n8951), .B(n8950), .S(n9010), .Z(n8952) );
  NAND3_X1 U10121 ( .A1(n8954), .A2(n8953), .A3(n8952), .ZN(n8959) );
  MUX2_X1 U10122 ( .A(n8956), .B(n8955), .S(n9028), .Z(n8957) );
  NAND3_X1 U10123 ( .A1(n8959), .A2(n8958), .A3(n8957), .ZN(n8964) );
  MUX2_X1 U10124 ( .A(n8961), .B(n8960), .S(n9028), .Z(n8962) );
  MUX2_X1 U10125 ( .A(n8966), .B(n8965), .S(n9028), .Z(n8968) );
  NAND2_X1 U10126 ( .A1(n9573), .A2(n9028), .ZN(n8970) );
  NAND2_X1 U10127 ( .A1(n9291), .A2(n9010), .ZN(n8969) );
  MUX2_X1 U10128 ( .A(n8970), .B(n8969), .S(n9653), .Z(n8971) );
  OR2_X1 U10129 ( .A1(n9547), .A2(n9028), .ZN(n8973) );
  NAND2_X1 U10130 ( .A1(n9547), .A2(n9028), .ZN(n8972) );
  MUX2_X1 U10131 ( .A(n8973), .B(n8972), .S(n9645), .Z(n8974) );
  NAND2_X1 U10132 ( .A1(n8975), .A2(n9543), .ZN(n8979) );
  MUX2_X1 U10133 ( .A(n8977), .B(n8976), .S(n9028), .Z(n8978) );
  NAND2_X1 U10134 ( .A1(n8979), .A2(n8978), .ZN(n8983) );
  INV_X1 U10135 ( .A(n9549), .ZN(n9518) );
  NAND2_X1 U10136 ( .A1(n9635), .A2(n9518), .ZN(n9179) );
  INV_X1 U10137 ( .A(n9179), .ZN(n8980) );
  NAND2_X1 U10138 ( .A1(n8983), .A2(n8980), .ZN(n8982) );
  MUX2_X1 U10139 ( .A(n9635), .B(n9518), .S(n9028), .Z(n8981) );
  NAND2_X1 U10140 ( .A1(n8982), .A2(n8981), .ZN(n8985) );
  OR3_X1 U10141 ( .A1(n8983), .A2(n9635), .A3(n9518), .ZN(n8984) );
  NAND2_X1 U10142 ( .A1(n8985), .A2(n8984), .ZN(n8989) );
  MUX2_X1 U10143 ( .A(n9533), .B(n9630), .S(n9010), .Z(n8986) );
  OAI21_X1 U10144 ( .B1(n8989), .B2(n8987), .A(n8986), .ZN(n8991) );
  INV_X1 U10145 ( .A(n8988), .ZN(n9180) );
  NAND2_X1 U10146 ( .A1(n8989), .A2(n9180), .ZN(n8990) );
  NAND2_X1 U10147 ( .A1(n9490), .A2(n8992), .ZN(n8995) );
  NAND2_X1 U10148 ( .A1(n9474), .A2(n9010), .ZN(n8994) );
  NOR2_X1 U10149 ( .A1(n9519), .A2(n9028), .ZN(n8993) );
  AOI22_X1 U10150 ( .A1(n8995), .A2(n8994), .B1(n8993), .B2(n9625), .ZN(n9002)
         );
  NAND2_X1 U10151 ( .A1(n8997), .A2(n8996), .ZN(n9000) );
  NAND2_X1 U10152 ( .A1(n8998), .A2(n9474), .ZN(n8999) );
  MUX2_X1 U10153 ( .A(n9000), .B(n8999), .S(n9028), .Z(n9001) );
  INV_X1 U10154 ( .A(n9261), .ZN(n9491) );
  MUX2_X1 U10155 ( .A(n9491), .B(n9615), .S(n9010), .Z(n9004) );
  NAND2_X1 U10156 ( .A1(n9615), .A2(n9491), .ZN(n9003) );
  AND2_X1 U10157 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  MUX2_X1 U10158 ( .A(n9007), .B(n9006), .S(n9028), .Z(n9008) );
  NAND3_X1 U10159 ( .A1(n9009), .A2(n9439), .A3(n9008), .ZN(n9014) );
  MUX2_X1 U10160 ( .A(n9012), .B(n9011), .S(n9010), .Z(n9013) );
  NAND3_X1 U10161 ( .A1(n9427), .A2(n9014), .A3(n9013), .ZN(n9018) );
  MUX2_X1 U10162 ( .A(n9016), .B(n9015), .S(n9028), .Z(n9017) );
  NAND2_X1 U10163 ( .A1(n9018), .A2(n9017), .ZN(n9021) );
  NAND3_X1 U10164 ( .A1(n9595), .A2(n9213), .A3(n9028), .ZN(n9020) );
  OR3_X1 U10165 ( .A1(n9595), .A2(n9213), .A3(n9028), .ZN(n9019) );
  MUX2_X1 U10166 ( .A(n9023), .B(n9022), .S(n9028), .Z(n9027) );
  NAND2_X1 U10167 ( .A1(n9025), .A2(n9024), .ZN(n9026) );
  INV_X1 U10168 ( .A(n8851), .ZN(n9395) );
  MUX2_X1 U10169 ( .A(n9029), .B(n9395), .S(n9028), .Z(n9030) );
  OAI21_X1 U10170 ( .B1(n9394), .B2(n8851), .A(n9030), .ZN(n9031) );
  NAND3_X1 U10171 ( .A1(n9036), .A2(n9034), .A3(n9033), .ZN(n9035) );
  NAND2_X1 U10172 ( .A1(n9035), .A2(n8307), .ZN(n9041) );
  INV_X1 U10173 ( .A(n9036), .ZN(n9038) );
  INV_X1 U10174 ( .A(n9690), .ZN(n9042) );
  NAND3_X1 U10175 ( .A1(n9043), .A2(n9042), .A3(n9572), .ZN(n9044) );
  OAI211_X1 U10176 ( .C1(n9045), .C2(n9047), .A(n9044), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9046) );
  INV_X1 U10177 ( .A(n9048), .ZN(n10926) );
  AOI22_X1 U10178 ( .A1(n10617), .A2(n9054), .B1(n10611), .B2(n10925), .ZN(
        n9051) );
  INV_X1 U10179 ( .A(n9049), .ZN(n9050) );
  OAI211_X1 U10180 ( .C1(n9052), .C2(n9314), .A(n9051), .B(n9050), .ZN(n9059)
         );
  INV_X1 U10181 ( .A(n8482), .ZN(n10624) );
  AOI22_X1 U10182 ( .A1(n9055), .A2(n9054), .B1(n10623), .B2(n9053), .ZN(n9056) );
  NOR3_X1 U10183 ( .A1(n10624), .A2(n9057), .A3(n9056), .ZN(n9058) );
  AOI211_X1 U10184 ( .C1(n10616), .C2(n10926), .A(n9059), .B(n9058), .ZN(n9060) );
  OAI21_X1 U10185 ( .B1(n9061), .B2(n9306), .A(n9060), .ZN(P2_U3229) );
  OAI21_X1 U10186 ( .B1(n9314), .B2(n9081), .A(n9062), .ZN(n9063) );
  AOI21_X1 U10187 ( .B1(n10617), .B2(n9325), .A(n9063), .ZN(n9064) );
  OAI21_X1 U10188 ( .B1(n9065), .B2(n9294), .A(n9064), .ZN(n9066) );
  AOI21_X1 U10189 ( .B1(n10611), .B2(n9067), .A(n9066), .ZN(n9072) );
  OAI22_X1 U10190 ( .A1(n9069), .A2(n9306), .B1(n9068), .B2(n10607), .ZN(n9070) );
  NAND3_X1 U10191 ( .A1(n8081), .A2(n5095), .A3(n9070), .ZN(n9071) );
  OAI211_X1 U10192 ( .C1(n8516), .C2(n9306), .A(n9072), .B(n9071), .ZN(
        P2_U3236) );
  OAI21_X1 U10193 ( .B1(n9314), .B2(n9074), .A(n9073), .ZN(n9075) );
  AOI21_X1 U10194 ( .B1(n10617), .B2(n9323), .A(n9075), .ZN(n9076) );
  OAI21_X1 U10195 ( .B1(n9077), .B2(n9294), .A(n9076), .ZN(n9078) );
  AOI21_X1 U10196 ( .B1(n9079), .B2(n10611), .A(n9078), .ZN(n9086) );
  INV_X1 U10197 ( .A(n9080), .ZN(n9084) );
  OAI22_X1 U10198 ( .A1(n9082), .A2(n9306), .B1(n9081), .B2(n10607), .ZN(n9083) );
  NAND3_X1 U10199 ( .A1(n8509), .A2(n9084), .A3(n9083), .ZN(n9085) );
  OAI211_X1 U10200 ( .C1(n8214), .C2(n9306), .A(n9086), .B(n9085), .ZN(
        P2_U3243) );
  INV_X1 U10201 ( .A(n9159), .ZN(n9126) );
  OAI22_X1 U10202 ( .A1(n9998), .A2(n9128), .B1(n10019), .B2(n9126), .ZN(n9100) );
  INV_X1 U10203 ( .A(n9100), .ZN(n9103) );
  OAI22_X1 U10204 ( .A1(n9998), .A2(n9087), .B1(n10019), .B2(n9128), .ZN(n9088) );
  XNOR2_X1 U10205 ( .A(n9088), .B(n9157), .ZN(n9101) );
  INV_X1 U10206 ( .A(n9101), .ZN(n9102) );
  INV_X1 U10207 ( .A(n9089), .ZN(n9091) );
  AND2_X1 U10208 ( .A1(n9091), .A2(n9090), .ZN(n9092) );
  NAND2_X1 U10209 ( .A1(n10107), .A2(n9133), .ZN(n9096) );
  NAND2_X1 U10210 ( .A1(n10000), .A2(n9160), .ZN(n9095) );
  NAND2_X1 U10211 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  XNOR2_X1 U10212 ( .A(n9097), .B(n9157), .ZN(n9098) );
  AOI22_X1 U10213 ( .A1(n10107), .A2(n9160), .B1(n9159), .B2(n10000), .ZN(
        n9779) );
  XNOR2_X1 U10214 ( .A(n9101), .B(n9100), .ZN(n9717) );
  AOI22_X1 U10215 ( .A1(n10097), .A2(n9133), .B1(n9143), .B2(n10001), .ZN(
        n9104) );
  XOR2_X1 U10216 ( .A(n9157), .B(n9104), .Z(n9753) );
  INV_X1 U10217 ( .A(n9753), .ZN(n9105) );
  AOI22_X1 U10218 ( .A1(n10097), .A2(n9160), .B1(n9159), .B2(n10001), .ZN(
        n9752) );
  INV_X1 U10219 ( .A(n9752), .ZN(n9106) );
  NAND2_X1 U10220 ( .A1(n10093), .A2(n9133), .ZN(n9108) );
  NAND2_X1 U10221 ( .A1(n9986), .A2(n9160), .ZN(n9107) );
  NAND2_X1 U10222 ( .A1(n9108), .A2(n9107), .ZN(n9109) );
  XNOR2_X1 U10223 ( .A(n9109), .B(n9152), .ZN(n9114) );
  INV_X1 U10224 ( .A(n9114), .ZN(n9112) );
  AND2_X1 U10225 ( .A1(n9986), .A2(n9159), .ZN(n9110) );
  AOI21_X1 U10226 ( .B1(n10093), .B2(n9160), .A(n9110), .ZN(n9113) );
  INV_X1 U10227 ( .A(n9113), .ZN(n9111) );
  NAND2_X1 U10228 ( .A1(n9112), .A2(n9111), .ZN(n9724) );
  AND2_X1 U10229 ( .A1(n9114), .A2(n9113), .ZN(n9723) );
  NAND2_X1 U10230 ( .A1(n10087), .A2(n9133), .ZN(n9116) );
  NAND2_X1 U10231 ( .A1(n9971), .A2(n9160), .ZN(n9115) );
  NAND2_X1 U10232 ( .A1(n9116), .A2(n9115), .ZN(n9117) );
  XNOR2_X1 U10233 ( .A(n9117), .B(n9152), .ZN(n9120) );
  AND2_X1 U10234 ( .A1(n9971), .A2(n9159), .ZN(n9118) );
  AOI21_X1 U10235 ( .B1(n10087), .B2(n9160), .A(n9118), .ZN(n9119) );
  NOR2_X1 U10236 ( .A1(n9120), .A2(n9119), .ZN(n9766) );
  NAND2_X1 U10237 ( .A1(n9120), .A2(n9119), .ZN(n9764) );
  AOI22_X1 U10238 ( .A1(n10082), .A2(n9133), .B1(n9143), .B2(n9954), .ZN(n9121) );
  XNOR2_X1 U10239 ( .A(n9121), .B(n9157), .ZN(n9123) );
  INV_X1 U10240 ( .A(n10082), .ZN(n9938) );
  OAI22_X1 U10241 ( .A1(n9938), .A2(n9128), .B1(n9122), .B2(n9126), .ZN(n9707)
         );
  AOI22_X1 U10242 ( .A1(n10078), .A2(n9133), .B1(n9143), .B2(n9942), .ZN(n9125) );
  XOR2_X1 U10243 ( .A(n9157), .B(n9125), .Z(n9130) );
  INV_X1 U10244 ( .A(n10078), .ZN(n9916) );
  OAI22_X1 U10245 ( .A1(n9916), .A2(n9128), .B1(n9127), .B2(n9126), .ZN(n9129)
         );
  NOR2_X1 U10246 ( .A1(n9130), .A2(n9129), .ZN(n9131) );
  AOI21_X1 U10247 ( .B1(n9130), .B2(n9129), .A(n9131), .ZN(n9746) );
  INV_X1 U10248 ( .A(n9131), .ZN(n9132) );
  NAND2_X1 U10249 ( .A1(n10072), .A2(n9133), .ZN(n9135) );
  NAND2_X1 U10250 ( .A1(n9920), .A2(n9143), .ZN(n9134) );
  NAND2_X1 U10251 ( .A1(n9135), .A2(n9134), .ZN(n9136) );
  XNOR2_X1 U10252 ( .A(n9136), .B(n9152), .ZN(n9138) );
  AND2_X1 U10253 ( .A1(n9920), .A2(n9159), .ZN(n9137) );
  AOI21_X1 U10254 ( .B1(n10072), .B2(n9160), .A(n9137), .ZN(n9139) );
  AND2_X1 U10255 ( .A1(n9138), .A2(n9139), .ZN(n9733) );
  INV_X1 U10256 ( .A(n9138), .ZN(n9141) );
  INV_X1 U10257 ( .A(n9139), .ZN(n9140) );
  NAND2_X1 U10258 ( .A1(n9141), .A2(n9140), .ZN(n9734) );
  OAI21_X2 U10259 ( .B1(n9737), .B2(n9733), .A(n9734), .ZN(n9790) );
  AND2_X1 U10260 ( .A1(n9908), .A2(n9159), .ZN(n9142) );
  AOI21_X1 U10261 ( .B1(n10067), .B2(n9143), .A(n9142), .ZN(n9146) );
  AOI22_X1 U10262 ( .A1(n10067), .A2(n9133), .B1(n9143), .B2(n9908), .ZN(n9144) );
  XNOR2_X1 U10263 ( .A(n9144), .B(n9157), .ZN(n9145) );
  XOR2_X1 U10264 ( .A(n9146), .B(n9145), .Z(n9789) );
  INV_X1 U10265 ( .A(n9145), .ZN(n9148) );
  NAND2_X1 U10266 ( .A1(n10062), .A2(n9133), .ZN(n9151) );
  NAND2_X1 U10267 ( .A1(n9893), .A2(n9160), .ZN(n9150) );
  NAND2_X1 U10268 ( .A1(n9151), .A2(n9150), .ZN(n9153) );
  XNOR2_X1 U10269 ( .A(n9153), .B(n9152), .ZN(n9156) );
  AND2_X1 U10270 ( .A1(n9893), .A2(n9159), .ZN(n9154) );
  AOI21_X1 U10271 ( .B1(n10062), .B2(n9160), .A(n9154), .ZN(n9155) );
  NOR2_X1 U10272 ( .A1(n9156), .A2(n9155), .ZN(n9695) );
  NAND2_X1 U10273 ( .A1(n9156), .A2(n9155), .ZN(n9693) );
  AOI22_X1 U10274 ( .A1(n10057), .A2(n9133), .B1(n9160), .B2(n9870), .ZN(n9158) );
  XNOR2_X1 U10275 ( .A(n9158), .B(n9157), .ZN(n9162) );
  AOI22_X1 U10276 ( .A1(n10057), .A2(n9160), .B1(n9159), .B2(n9870), .ZN(n9161) );
  XNOR2_X1 U10277 ( .A(n9162), .B(n9161), .ZN(n9163) );
  INV_X1 U10278 ( .A(n9164), .ZN(n9167) );
  AOI22_X1 U10279 ( .A1(n9758), .A2(n9893), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n9166) );
  NAND2_X1 U10280 ( .A1(n9791), .A2(n9801), .ZN(n9165) );
  OAI211_X1 U10281 ( .C1(n9760), .C2(n9167), .A(n9166), .B(n9165), .ZN(n9168)
         );
  AOI21_X1 U10282 ( .B1(n10057), .B2(n9773), .A(n9168), .ZN(n9169) );
  OAI21_X1 U10283 ( .B1(n9170), .B2(n9785), .A(n9169), .ZN(P1_U3218) );
  INV_X1 U10284 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10505) );
  INV_X1 U10285 ( .A(n9171), .ZN(n9204) );
  OAI222_X1 U10286 ( .A1(n10144), .A2(n10505), .B1(n10147), .B2(n9204), .C1(
        P1_U3084), .C2(n9172), .ZN(P1_U3323) );
  INV_X1 U10287 ( .A(n9645), .ZN(n9569) );
  INV_X1 U10288 ( .A(n9547), .ZN(n9175) );
  NAND2_X1 U10289 ( .A1(n9540), .A2(n9539), .ZN(n9538) );
  NAND2_X1 U10290 ( .A1(n9538), .A2(n9178), .ZN(n9526) );
  OR2_X1 U10291 ( .A1(n9625), .A2(n9519), .ZN(n9181) );
  INV_X1 U10292 ( .A(n9284), .ZN(n9504) );
  NAND2_X1 U10293 ( .A1(n9469), .A2(n9476), .ZN(n9470) );
  INV_X1 U10294 ( .A(n9611), .ZN(n9460) );
  INV_X1 U10295 ( .A(n9443), .ZN(n9413) );
  INV_X1 U10296 ( .A(n9630), .ZN(n9514) );
  INV_X1 U10297 ( .A(n9625), .ZN(n9501) );
  NAND2_X1 U10298 ( .A1(n9456), .A2(n9450), .ZN(n9444) );
  AOI21_X1 U10299 ( .B1(n9589), .B2(n9406), .A(n9399), .ZN(n9590) );
  INV_X1 U10300 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9190) );
  OAI22_X1 U10301 ( .A1(n9191), .A2(n9568), .B1(n9190), .B2(n10933), .ZN(n9192) );
  AOI21_X1 U10302 ( .B1(n9590), .B2(n9579), .A(n9192), .ZN(n9200) );
  XNOR2_X1 U10303 ( .A(n9194), .B(n9193), .ZN(n9196) );
  NOR2_X1 U10304 ( .A1(n9690), .A2(n10500), .ZN(n9195) );
  NOR2_X1 U10305 ( .A1(n9550), .A2(n9195), .ZN(n9393) );
  AOI222_X1 U10306 ( .A1(n9576), .A2(n9196), .B1(n9430), .B2(n9572), .C1(n9320), .C2(n9393), .ZN(n9591) );
  OAI21_X1 U10307 ( .B1(n9197), .B2(n9554), .A(n9591), .ZN(n9198) );
  NAND2_X1 U10308 ( .A1(n9198), .A2(n10933), .ZN(n9199) );
  OAI211_X1 U10309 ( .C1(n9594), .C2(n9581), .A(n9200), .B(n9199), .ZN(
        P2_U3267) );
  INV_X1 U10310 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9201) );
  OAI222_X1 U10311 ( .A1(n6355), .A2(n9691), .B1(n9684), .B2(n9202), .C1(n9201), .C2(n9687), .ZN(P2_U3330) );
  OAI222_X1 U10312 ( .A1(n5819), .A2(n9691), .B1(n9684), .B2(n9204), .C1(n9687), .C2(n9203), .ZN(P2_U3328) );
  INV_X1 U10313 ( .A(n9600), .ZN(n9425) );
  INV_X1 U10314 ( .A(n9206), .ZN(n9207) );
  AOI21_X1 U10315 ( .B1(n9205), .B2(n9207), .A(n9306), .ZN(n9211) );
  NOR3_X1 U10316 ( .A1(n9208), .A2(n9250), .A3(n10607), .ZN(n9210) );
  OAI21_X1 U10317 ( .B1(n9211), .B2(n9210), .A(n9209), .ZN(n9217) );
  OAI22_X1 U10318 ( .A1(n9250), .A2(n9313), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9212), .ZN(n9215) );
  NOR2_X1 U10319 ( .A1(n9213), .A2(n9314), .ZN(n9214) );
  AOI211_X1 U10320 ( .C1(n10616), .C2(n9423), .A(n9215), .B(n9214), .ZN(n9216)
         );
  OAI211_X1 U10321 ( .C1(n9425), .C2(n9319), .A(n9217), .B(n9216), .ZN(
        P2_U3216) );
  INV_X1 U10322 ( .A(n9620), .ZN(n9488) );
  INV_X1 U10323 ( .A(n9221), .ZN(n9218) );
  OAI22_X1 U10324 ( .A1(n9218), .A2(n9306), .B1(n9284), .B2(n10607), .ZN(n9222) );
  INV_X1 U10325 ( .A(n9219), .ZN(n9220) );
  NAND2_X1 U10326 ( .A1(n9221), .A2(n9220), .ZN(n9258) );
  NAND2_X1 U10327 ( .A1(n9222), .A2(n9258), .ZN(n9228) );
  INV_X1 U10328 ( .A(n9223), .ZN(n9486) );
  OAI22_X1 U10329 ( .A1(n9313), .A2(n9224), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10452), .ZN(n9226) );
  NOR2_X1 U10330 ( .A1(n9261), .A2(n9314), .ZN(n9225) );
  AOI211_X1 U10331 ( .C1(n10616), .C2(n9486), .A(n9226), .B(n9225), .ZN(n9227)
         );
  OAI211_X1 U10332 ( .C1(n9488), .C2(n9319), .A(n9228), .B(n9227), .ZN(
        P2_U3218) );
  XNOR2_X1 U10333 ( .A(n9230), .B(n9229), .ZN(n9231) );
  XNOR2_X1 U10334 ( .A(n9232), .B(n9231), .ZN(n9237) );
  NAND2_X1 U10335 ( .A1(n9691), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9388) );
  OAI21_X1 U10336 ( .B1(n9313), .B2(n9547), .A(n9388), .ZN(n9233) );
  AOI21_X1 U10337 ( .B1(n10613), .B2(n9518), .A(n9233), .ZN(n9234) );
  OAI21_X1 U10338 ( .B1(n9553), .B2(n9294), .A(n9234), .ZN(n9235) );
  AOI21_X1 U10339 ( .B1(n9642), .B2(n10611), .A(n9235), .ZN(n9236) );
  OAI21_X1 U10340 ( .B1(n9237), .B2(n9306), .A(n9236), .ZN(P2_U3221) );
  AOI21_X1 U10341 ( .B1(n9238), .B2(n5586), .A(n9306), .ZN(n9243) );
  NOR3_X1 U10342 ( .A1(n9240), .A2(n9549), .A3(n10607), .ZN(n9242) );
  OAI21_X1 U10343 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9247) );
  OAI22_X1 U10344 ( .A1(n9313), .A2(n9549), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10471), .ZN(n9245) );
  NOR2_X1 U10345 ( .A1(n9294), .A2(n9521), .ZN(n9244) );
  AOI211_X1 U10346 ( .C1(n10613), .C2(n9519), .A(n9245), .B(n9244), .ZN(n9246)
         );
  OAI211_X1 U10347 ( .C1(n9514), .C2(n9319), .A(n9247), .B(n9246), .ZN(
        P2_U3225) );
  OAI211_X1 U10348 ( .C1(n9249), .C2(n9248), .A(n9308), .B(n10623), .ZN(n9256)
         );
  OAI22_X1 U10349 ( .A1(n9250), .A2(n9550), .B1(n9261), .B2(n9548), .ZN(n9463)
         );
  AOI22_X1 U10350 ( .A1(n9463), .A2(n9251), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n9255) );
  NAND2_X1 U10351 ( .A1(n9611), .A2(n10611), .ZN(n9254) );
  INV_X1 U10352 ( .A(n9252), .ZN(n9458) );
  NAND2_X1 U10353 ( .A1(n10616), .A2(n9458), .ZN(n9253) );
  NAND4_X1 U10354 ( .A1(n9256), .A2(n9255), .A3(n9254), .A4(n9253), .ZN(
        P2_U3227) );
  NAND2_X1 U10355 ( .A1(n9258), .A2(n9257), .ZN(n9260) );
  XNOR2_X1 U10356 ( .A(n9260), .B(n9259), .ZN(n9264) );
  OAI22_X1 U10357 ( .A1(n9264), .A2(n9306), .B1(n9261), .B2(n10607), .ZN(n9262) );
  OAI21_X1 U10358 ( .B1(n9264), .B2(n9263), .A(n9262), .ZN(n9268) );
  OAI22_X1 U10359 ( .A1(n9313), .A2(n9284), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10480), .ZN(n9266) );
  NOR2_X1 U10360 ( .A1(n9442), .A2(n9314), .ZN(n9265) );
  AOI211_X1 U10361 ( .C1(n10616), .C2(n9472), .A(n9266), .B(n9265), .ZN(n9267)
         );
  OAI211_X1 U10362 ( .C1(n9184), .C2(n9319), .A(n9268), .B(n9267), .ZN(
        P2_U3231) );
  INV_X1 U10363 ( .A(n9635), .ZN(n9530) );
  AOI21_X1 U10364 ( .B1(n9270), .B2(n9269), .A(n9306), .ZN(n9271) );
  NAND2_X1 U10365 ( .A1(n9271), .A2(n9238), .ZN(n9278) );
  INV_X1 U10366 ( .A(n9272), .ZN(n9528) );
  AOI22_X1 U10367 ( .A1(n10617), .A2(n9177), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3152), .ZN(n9274) );
  OAI21_X1 U10368 ( .B1(n9275), .B2(n9314), .A(n9274), .ZN(n9276) );
  AOI21_X1 U10369 ( .B1(n9528), .B2(n10616), .A(n9276), .ZN(n9277) );
  OAI211_X1 U10370 ( .C1(n9530), .C2(n9319), .A(n9278), .B(n9277), .ZN(
        P2_U3235) );
  OAI21_X1 U10371 ( .B1(n9281), .B2(n9241), .A(n9279), .ZN(n9289) );
  NOR3_X1 U10372 ( .A1(n9281), .A2(n9280), .A3(n10607), .ZN(n9282) );
  OAI21_X1 U10373 ( .B1(n9282), .B2(n10617), .A(n9533), .ZN(n9287) );
  INV_X1 U10374 ( .A(n9283), .ZN(n9499) );
  OAI22_X1 U10375 ( .A1(n9314), .A2(n9284), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10490), .ZN(n9285) );
  AOI21_X1 U10376 ( .B1(n9499), .B2(n10616), .A(n9285), .ZN(n9286) );
  OAI211_X1 U10377 ( .C1(n9501), .C2(n9319), .A(n9287), .B(n9286), .ZN(n9288)
         );
  AOI21_X1 U10378 ( .B1(n9289), .B2(n10623), .A(n9288), .ZN(n9290) );
  INV_X1 U10379 ( .A(n9290), .ZN(P2_U3237) );
  NAND2_X1 U10380 ( .A1(n9691), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9364) );
  OAI21_X1 U10381 ( .B1(n9313), .B2(n9291), .A(n9364), .ZN(n9292) );
  AOI21_X1 U10382 ( .B1(n10613), .B2(n9177), .A(n9292), .ZN(n9293) );
  OAI21_X1 U10383 ( .B1(n9564), .B2(n9294), .A(n9293), .ZN(n9303) );
  INV_X1 U10384 ( .A(n9295), .ZN(n9301) );
  INV_X1 U10385 ( .A(n9296), .ZN(n9298) );
  NAND2_X1 U10386 ( .A1(n9298), .A2(n9297), .ZN(n9300) );
  NOR2_X1 U10387 ( .A1(n9301), .A2(n9300), .ZN(n9299) );
  AOI211_X1 U10388 ( .C1(n9301), .C2(n9300), .A(n9306), .B(n9299), .ZN(n9302)
         );
  AOI211_X1 U10389 ( .C1(n10611), .C2(n9645), .A(n9303), .B(n9302), .ZN(n9304)
         );
  INV_X1 U10390 ( .A(n9304), .ZN(P2_U3240) );
  INV_X1 U10391 ( .A(n9305), .ZN(n9307) );
  AOI21_X1 U10392 ( .B1(n9308), .B2(n9307), .A(n9306), .ZN(n9311) );
  NOR3_X1 U10393 ( .A1(n9309), .A2(n9442), .A3(n10607), .ZN(n9310) );
  OAI21_X1 U10394 ( .B1(n9311), .B2(n9310), .A(n9205), .ZN(n9318) );
  INV_X1 U10395 ( .A(n9312), .ZN(n9447) );
  OAI22_X1 U10396 ( .A1(n9442), .A2(n9313), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10284), .ZN(n9316) );
  NOR2_X1 U10397 ( .A1(n9443), .A2(n9314), .ZN(n9315) );
  AOI211_X1 U10398 ( .C1(n10616), .C2(n9447), .A(n9316), .B(n9315), .ZN(n9317)
         );
  OAI211_X1 U10399 ( .C1(n9450), .C2(n9319), .A(n9318), .B(n9317), .ZN(
        P2_U3242) );
  MUX2_X1 U10400 ( .A(n9394), .B(P2_DATAO_REG_31__SCAN_IN), .S(n9333), .Z(
        P2_U3583) );
  MUX2_X1 U10401 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9320), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10402 ( .A(n9412), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9333), .Z(
        P2_U3581) );
  MUX2_X1 U10403 ( .A(n9430), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9333), .Z(
        P2_U3580) );
  MUX2_X1 U10404 ( .A(n9413), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9333), .Z(
        P2_U3579) );
  INV_X1 U10405 ( .A(n9442), .ZN(n9477) );
  MUX2_X1 U10406 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9477), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10407 ( .A(n9491), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9333), .Z(
        P2_U3576) );
  MUX2_X1 U10408 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9504), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10409 ( .A(n9519), .B(P2_DATAO_REG_22__SCAN_IN), .S(n9333), .Z(
        P2_U3574) );
  MUX2_X1 U10410 ( .A(n9533), .B(P2_DATAO_REG_21__SCAN_IN), .S(n9333), .Z(
        P2_U3573) );
  MUX2_X1 U10411 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9518), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10412 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9177), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10413 ( .A(n9573), .B(P2_DATAO_REG_17__SCAN_IN), .S(n9333), .Z(
        P2_U3569) );
  MUX2_X1 U10414 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9321), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10415 ( .A(n9322), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9333), .Z(
        P2_U3567) );
  MUX2_X1 U10416 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9323), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10417 ( .A(n9324), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9333), .Z(
        P2_U3565) );
  MUX2_X1 U10418 ( .A(n9325), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9333), .Z(
        P2_U3564) );
  MUX2_X1 U10419 ( .A(n9326), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9333), .Z(
        P2_U3563) );
  MUX2_X1 U10420 ( .A(n9327), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9333), .Z(
        P2_U3562) );
  MUX2_X1 U10421 ( .A(n9328), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9333), .Z(
        P2_U3561) );
  MUX2_X1 U10422 ( .A(n9329), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9333), .Z(
        P2_U3560) );
  MUX2_X1 U10423 ( .A(n9330), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9333), .Z(
        P2_U3559) );
  MUX2_X1 U10424 ( .A(n9331), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9333), .Z(
        P2_U3558) );
  MUX2_X1 U10425 ( .A(n10612), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9333), .Z(
        P2_U3557) );
  MUX2_X1 U10426 ( .A(n7347), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9333), .Z(
        P2_U3555) );
  MUX2_X1 U10427 ( .A(n5338), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9333), .Z(
        P2_U3554) );
  MUX2_X1 U10428 ( .A(n7229), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9333), .Z(
        P2_U3553) );
  OAI21_X1 U10429 ( .B1(n9336), .B2(n9335), .A(n9334), .ZN(n9337) );
  NAND2_X1 U10430 ( .A1(n10761), .A2(n9337), .ZN(n9347) );
  NAND2_X1 U10431 ( .A1(n10794), .A2(n9338), .ZN(n9346) );
  NOR2_X1 U10432 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9339), .ZN(n9340) );
  AOI21_X1 U10433 ( .B1(n10787), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9340), .ZN(
        n9345) );
  OAI211_X1 U10434 ( .C1(n9343), .C2(n9342), .A(n10796), .B(n9341), .ZN(n9344)
         );
  NAND4_X1 U10435 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(
        P2_U3256) );
  NAND2_X1 U10436 ( .A1(n9368), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9350) );
  OAI21_X1 U10437 ( .B1(n9368), .B2(P2_REG2_REG_17__SCAN_IN), .A(n9350), .ZN(
        n9351) );
  NOR2_X1 U10438 ( .A1(n9352), .A2(n9351), .ZN(n9367) );
  AOI211_X1 U10439 ( .C1(n9352), .C2(n9351), .A(n9367), .B(n10788), .ZN(n9363)
         );
  INV_X1 U10440 ( .A(n9353), .ZN(n9354) );
  AOI21_X1 U10441 ( .B1(n10787), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9354), .ZN(
        n9361) );
  XNOR2_X1 U10442 ( .A(n9373), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9359) );
  AOI21_X1 U10443 ( .B1(n9357), .B2(n9356), .A(n9355), .ZN(n9358) );
  NAND2_X1 U10444 ( .A1(n9359), .A2(n9358), .ZN(n9372) );
  OAI211_X1 U10445 ( .C1(n9359), .C2(n9358), .A(n10796), .B(n9372), .ZN(n9360)
         );
  OAI211_X1 U10446 ( .C1(n10763), .C2(n9373), .A(n9361), .B(n9360), .ZN(n9362)
         );
  OR2_X1 U10447 ( .A1(n9363), .A2(n9362), .ZN(P2_U3262) );
  INV_X1 U10448 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9365) );
  OAI21_X1 U10449 ( .B1(n10772), .B2(n9365), .A(n9364), .ZN(n9366) );
  AOI21_X1 U10450 ( .B1(n9382), .B2(n10794), .A(n9366), .ZN(n9378) );
  MUX2_X1 U10451 ( .A(n6141), .B(P2_REG2_REG_18__SCAN_IN), .S(n9382), .Z(n9369) );
  INV_X1 U10452 ( .A(n9369), .ZN(n9370) );
  NAND2_X1 U10453 ( .A1(n9370), .A2(n9371), .ZN(n9379) );
  OAI21_X1 U10454 ( .B1(n9371), .B2(n9370), .A(n9379), .ZN(n9376) );
  XNOR2_X1 U10455 ( .A(n9382), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9384) );
  OAI21_X1 U10456 ( .B1(n9374), .B2(n9373), .A(n9372), .ZN(n9383) );
  XNOR2_X1 U10457 ( .A(n9384), .B(n9383), .ZN(n9375) );
  AOI22_X1 U10458 ( .A1(n10761), .A2(n9376), .B1(n10796), .B2(n9375), .ZN(
        n9377) );
  NAND2_X1 U10459 ( .A1(n9378), .A2(n9377), .ZN(P2_U3263) );
  MUX2_X1 U10460 ( .A(n6156), .B(P2_REG2_REG_19__SCAN_IN), .S(n10922), .Z(
        n9381) );
  OAI21_X1 U10461 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n9382), .A(n9379), .ZN(
        n9380) );
  XOR2_X1 U10462 ( .A(n9381), .B(n9380), .Z(n9392) );
  OAI22_X1 U10463 ( .A1(n9384), .A2(n9383), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n9382), .ZN(n9386) );
  XNOR2_X1 U10464 ( .A(n10922), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9385) );
  XNOR2_X1 U10465 ( .A(n9386), .B(n9385), .ZN(n9390) );
  NAND2_X1 U10466 ( .A1(n10787), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9387) );
  OAI211_X1 U10467 ( .C1(n10763), .C2(n10922), .A(n9388), .B(n9387), .ZN(n9389) );
  AOI21_X1 U10468 ( .B1(n10796), .B2(n9390), .A(n9389), .ZN(n9391) );
  OAI21_X1 U10469 ( .B1(n10788), .B2(n9392), .A(n9391), .ZN(P2_U3264) );
  XNOR2_X1 U10470 ( .A(n9585), .B(n8851), .ZN(n9583) );
  NAND2_X1 U10471 ( .A1(n9394), .A2(n9393), .ZN(n9586) );
  NOR2_X1 U10472 ( .A1(n9566), .A2(n9586), .ZN(n9402) );
  NOR2_X1 U10473 ( .A1(n9395), .A2(n9568), .ZN(n9396) );
  AOI211_X1 U10474 ( .C1(n9566), .C2(P2_REG2_REG_31__SCAN_IN), .A(n9402), .B(
        n9396), .ZN(n9397) );
  OAI21_X1 U10475 ( .B1(n9583), .B2(n9398), .A(n9397), .ZN(P2_U3265) );
  INV_X1 U10476 ( .A(n9399), .ZN(n9401) );
  NAND2_X1 U10477 ( .A1(n9401), .A2(n9400), .ZN(n9584) );
  NAND3_X1 U10478 ( .A1(n9585), .A2(n9579), .A3(n9584), .ZN(n9404) );
  AOI21_X1 U10479 ( .B1(n9541), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9402), .ZN(
        n9403) );
  OAI211_X1 U10480 ( .C1(n9588), .C2(n9568), .A(n9404), .B(n9403), .ZN(
        P2_U3266) );
  XNOR2_X1 U10481 ( .A(n9405), .B(n5345), .ZN(n9599) );
  INV_X1 U10482 ( .A(n9406), .ZN(n9407) );
  AOI21_X1 U10483 ( .B1(n9595), .B2(n9422), .A(n9407), .ZN(n9596) );
  AOI22_X1 U10484 ( .A1(n9408), .A2(n10927), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n9541), .ZN(n9409) );
  OAI21_X1 U10485 ( .B1(n5324), .B2(n9568), .A(n9409), .ZN(n9417) );
  OAI211_X1 U10486 ( .C1(n9411), .C2(n5345), .A(n9410), .B(n9576), .ZN(n9415)
         );
  AOI22_X1 U10487 ( .A1(n9413), .A2(n9572), .B1(n9574), .B2(n9412), .ZN(n9414)
         );
  NOR2_X1 U10488 ( .A1(n9598), .A2(n9541), .ZN(n9416) );
  AOI211_X1 U10489 ( .C1(n9579), .C2(n9596), .A(n9417), .B(n9416), .ZN(n9418)
         );
  OAI21_X1 U10490 ( .B1(n9599), .B2(n9581), .A(n9418), .ZN(P2_U3268) );
  INV_X1 U10491 ( .A(n9419), .ZN(n9420) );
  AOI21_X1 U10492 ( .B1(n9427), .B2(n9421), .A(n9420), .ZN(n9604) );
  AOI21_X1 U10493 ( .B1(n9600), .B2(n9444), .A(n5325), .ZN(n9601) );
  AOI22_X1 U10494 ( .A1(n9423), .A2(n10927), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n9541), .ZN(n9424) );
  OAI21_X1 U10495 ( .B1(n9425), .B2(n9568), .A(n9424), .ZN(n9434) );
  OAI211_X1 U10496 ( .C1(n9428), .C2(n9427), .A(n9426), .B(n9576), .ZN(n9432)
         );
  AOI22_X1 U10497 ( .A1(n9430), .A2(n9574), .B1(n9572), .B2(n9429), .ZN(n9431)
         );
  NOR2_X1 U10498 ( .A1(n9603), .A2(n9541), .ZN(n9433) );
  AOI211_X1 U10499 ( .C1(n9601), .C2(n9579), .A(n9434), .B(n9433), .ZN(n9435)
         );
  OAI21_X1 U10500 ( .B1(n9604), .B2(n9581), .A(n9435), .ZN(P2_U3269) );
  OAI21_X1 U10501 ( .B1(n9438), .B2(n9437), .A(n9436), .ZN(n9609) );
  XNOR2_X1 U10502 ( .A(n9440), .B(n9439), .ZN(n9441) );
  OAI222_X1 U10503 ( .A1(n9550), .A2(n9443), .B1(n9548), .B2(n9442), .C1(n9546), .C2(n9441), .ZN(n9605) );
  INV_X1 U10504 ( .A(n9456), .ZN(n9446) );
  INV_X1 U10505 ( .A(n9444), .ZN(n9445) );
  AOI211_X1 U10506 ( .C1(n9607), .C2(n9446), .A(n11125), .B(n9445), .ZN(n9606)
         );
  NAND2_X1 U10507 ( .A1(n9606), .A2(n9467), .ZN(n9449) );
  AOI22_X1 U10508 ( .A1(n9447), .A2(n10927), .B1(n9566), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9448) );
  OAI211_X1 U10509 ( .C1(n9450), .C2(n9568), .A(n9449), .B(n9448), .ZN(n9451)
         );
  AOI21_X1 U10510 ( .B1(n9605), .B2(n10933), .A(n9451), .ZN(n9452) );
  OAI21_X1 U10511 ( .B1(n9609), .B2(n9581), .A(n9452), .ZN(P2_U3270) );
  XNOR2_X1 U10512 ( .A(n9454), .B(n9453), .ZN(n9614) );
  INV_X1 U10513 ( .A(n9455), .ZN(n9457) );
  AOI211_X1 U10514 ( .C1(n9611), .C2(n9457), .A(n11125), .B(n9456), .ZN(n9610)
         );
  AOI22_X1 U10515 ( .A1(n9566), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9458), .B2(
        n10927), .ZN(n9459) );
  OAI21_X1 U10516 ( .B1(n9460), .B2(n9568), .A(n9459), .ZN(n9466) );
  XNOR2_X1 U10517 ( .A(n9462), .B(n9461), .ZN(n9464) );
  AOI21_X1 U10518 ( .B1(n9464), .B2(n9576), .A(n9463), .ZN(n9613) );
  NOR2_X1 U10519 ( .A1(n9613), .A2(n9541), .ZN(n9465) );
  AOI211_X1 U10520 ( .C1(n9610), .C2(n9467), .A(n9466), .B(n9465), .ZN(n9468)
         );
  OAI21_X1 U10521 ( .B1(n9614), .B2(n9581), .A(n9468), .ZN(P2_U3271) );
  OAI21_X1 U10522 ( .B1(n9469), .B2(n9476), .A(n9470), .ZN(n9471) );
  INV_X1 U10523 ( .A(n9471), .ZN(n9619) );
  XOR2_X1 U10524 ( .A(n9615), .B(n9485), .Z(n9616) );
  AOI22_X1 U10525 ( .A1(n9566), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9472), .B2(
        n10927), .ZN(n9473) );
  OAI21_X1 U10526 ( .B1(n9184), .B2(n9568), .A(n9473), .ZN(n9480) );
  NAND2_X1 U10527 ( .A1(n9489), .A2(n9474), .ZN(n9475) );
  XOR2_X1 U10528 ( .A(n9476), .B(n9475), .Z(n9478) );
  AOI222_X1 U10529 ( .A1(n9576), .A2(n9478), .B1(n9477), .B2(n9574), .C1(n9504), .C2(n9572), .ZN(n9618) );
  NOR2_X1 U10530 ( .A1(n9618), .A2(n9541), .ZN(n9479) );
  AOI211_X1 U10531 ( .C1(n9616), .C2(n9579), .A(n9480), .B(n9479), .ZN(n9481)
         );
  OAI21_X1 U10532 ( .B1(n9619), .B2(n9581), .A(n9481), .ZN(P2_U3272) );
  AOI21_X1 U10533 ( .B1(n9490), .B2(n9482), .A(n9483), .ZN(n9484) );
  INV_X1 U10534 ( .A(n9484), .ZN(n9624) );
  AOI21_X1 U10535 ( .B1(n9620), .B2(n9497), .A(n5326), .ZN(n9621) );
  AOI22_X1 U10536 ( .A1(n9566), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9486), .B2(
        n10927), .ZN(n9487) );
  OAI21_X1 U10537 ( .B1(n9488), .B2(n9568), .A(n9487), .ZN(n9494) );
  OAI21_X1 U10538 ( .B1(n5645), .B2(n9490), .A(n9489), .ZN(n9492) );
  AOI222_X1 U10539 ( .A1(n9576), .A2(n9492), .B1(n9519), .B2(n9572), .C1(n9491), .C2(n9574), .ZN(n9623) );
  NOR2_X1 U10540 ( .A1(n9623), .A2(n9566), .ZN(n9493) );
  AOI211_X1 U10541 ( .C1(n9621), .C2(n9579), .A(n9494), .B(n9493), .ZN(n9495)
         );
  OAI21_X1 U10542 ( .B1(n9624), .B2(n9581), .A(n9495), .ZN(P2_U3273) );
  XNOR2_X1 U10543 ( .A(n9496), .B(n9503), .ZN(n9629) );
  INV_X1 U10544 ( .A(n9511), .ZN(n9498) );
  AOI21_X1 U10545 ( .B1(n9625), .B2(n9498), .A(n5327), .ZN(n9626) );
  AOI22_X1 U10546 ( .A1(n9566), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9499), .B2(
        n10927), .ZN(n9500) );
  OAI21_X1 U10547 ( .B1(n9501), .B2(n9568), .A(n9500), .ZN(n9507) );
  XNOR2_X1 U10548 ( .A(n9502), .B(n9503), .ZN(n9505) );
  AOI222_X1 U10549 ( .A1(n9576), .A2(n9505), .B1(n9533), .B2(n9572), .C1(n9504), .C2(n9574), .ZN(n9628) );
  NOR2_X1 U10550 ( .A1(n9628), .A2(n9566), .ZN(n9506) );
  AOI211_X1 U10551 ( .C1(n9626), .C2(n9579), .A(n9507), .B(n9506), .ZN(n9508)
         );
  OAI21_X1 U10552 ( .B1(n9629), .B2(n9581), .A(n9508), .ZN(P2_U3274) );
  AOI21_X1 U10553 ( .B1(n9517), .B2(n9510), .A(n9509), .ZN(n9634) );
  INV_X1 U10554 ( .A(n9527), .ZN(n9512) );
  AOI21_X1 U10555 ( .B1(n9630), .B2(n9512), .A(n9511), .ZN(n9631) );
  INV_X1 U10556 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9513) );
  OAI22_X1 U10557 ( .A1(n9514), .A2(n9568), .B1(n10933), .B2(n9513), .ZN(n9515) );
  AOI21_X1 U10558 ( .B1(n9631), .B2(n9579), .A(n9515), .ZN(n9524) );
  XOR2_X1 U10559 ( .A(n9516), .B(n9517), .Z(n9520) );
  AOI222_X1 U10560 ( .A1(n9576), .A2(n9520), .B1(n9519), .B2(n9574), .C1(n9518), .C2(n9572), .ZN(n9633) );
  OAI21_X1 U10561 ( .B1(n9521), .B2(n9554), .A(n9633), .ZN(n9522) );
  NAND2_X1 U10562 ( .A1(n9522), .A2(n10933), .ZN(n9523) );
  OAI211_X1 U10563 ( .C1(n9634), .C2(n9581), .A(n9524), .B(n9523), .ZN(
        P2_U3275) );
  OAI21_X1 U10564 ( .B1(n9526), .B2(n9531), .A(n9525), .ZN(n9639) );
  AOI21_X1 U10565 ( .B1(n9635), .B2(n9551), .A(n9527), .ZN(n9636) );
  AOI22_X1 U10566 ( .A1(n9566), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9528), .B2(
        n10927), .ZN(n9529) );
  OAI21_X1 U10567 ( .B1(n9530), .B2(n9568), .A(n9529), .ZN(n9536) );
  XNOR2_X1 U10568 ( .A(n9532), .B(n9531), .ZN(n9534) );
  AOI222_X1 U10569 ( .A1(n9576), .A2(n9534), .B1(n9177), .B2(n9572), .C1(n9533), .C2(n9574), .ZN(n9638) );
  NOR2_X1 U10570 ( .A1(n9638), .A2(n9566), .ZN(n9535) );
  AOI211_X1 U10571 ( .C1(n9636), .C2(n9579), .A(n9536), .B(n9535), .ZN(n9537)
         );
  OAI21_X1 U10572 ( .B1(n9581), .B2(n9639), .A(n9537), .ZN(P2_U3276) );
  OAI21_X1 U10573 ( .B1(n9540), .B2(n9539), .A(n9538), .ZN(n9644) );
  AOI22_X1 U10574 ( .A1(n9642), .A2(n9542), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n9541), .ZN(n9559) );
  XNOR2_X1 U10575 ( .A(n9544), .B(n9543), .ZN(n9545) );
  OAI222_X1 U10576 ( .A1(n9550), .A2(n9549), .B1(n9548), .B2(n9547), .C1(n9546), .C2(n9545), .ZN(n9640) );
  INV_X1 U10577 ( .A(n9551), .ZN(n9552) );
  AOI211_X1 U10578 ( .C1(n9642), .C2(n9562), .A(n11125), .B(n9552), .ZN(n9641)
         );
  INV_X1 U10579 ( .A(n9641), .ZN(n9556) );
  OAI22_X1 U10580 ( .A1(n9556), .A2(n9555), .B1(n9554), .B2(n9553), .ZN(n9557)
         );
  OAI21_X1 U10581 ( .B1(n9640), .B2(n9557), .A(n10933), .ZN(n9558) );
  OAI211_X1 U10582 ( .C1(n9644), .C2(n9581), .A(n9559), .B(n9558), .ZN(
        P2_U3277) );
  XNOR2_X1 U10583 ( .A(n9560), .B(n9561), .ZN(n9649) );
  INV_X1 U10584 ( .A(n9562), .ZN(n9563) );
  AOI21_X1 U10585 ( .B1(n9645), .B2(n5088), .A(n9563), .ZN(n9646) );
  INV_X1 U10586 ( .A(n9564), .ZN(n9565) );
  AOI22_X1 U10587 ( .A1(n9566), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9565), .B2(
        n10927), .ZN(n9567) );
  OAI21_X1 U10588 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9578) );
  XNOR2_X1 U10589 ( .A(n9570), .B(n9571), .ZN(n9575) );
  AOI222_X1 U10590 ( .A1(n9576), .A2(n9575), .B1(n9177), .B2(n9574), .C1(n9573), .C2(n9572), .ZN(n9648) );
  NOR2_X1 U10591 ( .A1(n9648), .A2(n9566), .ZN(n9577) );
  AOI211_X1 U10592 ( .C1(n9646), .C2(n9579), .A(n9578), .B(n9577), .ZN(n9580)
         );
  OAI21_X1 U10593 ( .B1(n9581), .B2(n9649), .A(n9580), .ZN(P2_U3278) );
  NAND2_X1 U10594 ( .A1(n8851), .A2(n11066), .ZN(n9582) );
  OAI211_X1 U10595 ( .C1(n9583), .C2(n11125), .A(n9582), .B(n9586), .ZN(n9662)
         );
  MUX2_X1 U10596 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9662), .S(n11132), .Z(
        P2_U3551) );
  NAND3_X1 U10597 ( .A1(n9585), .A2(n11067), .A3(n9584), .ZN(n9587) );
  OAI211_X1 U10598 ( .C1(n9588), .C2(n11123), .A(n9587), .B(n9586), .ZN(n9663)
         );
  MUX2_X1 U10599 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9663), .S(n11132), .Z(
        P2_U3550) );
  AOI22_X1 U10600 ( .A1(n9590), .A2(n11067), .B1(n11066), .B2(n9589), .ZN(
        n9592) );
  AND2_X1 U10601 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  MUX2_X1 U10602 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9664), .S(n11132), .Z(
        P2_U3549) );
  AOI22_X1 U10603 ( .A1(n9596), .A2(n11067), .B1(n11066), .B2(n9595), .ZN(
        n9597) );
  OAI211_X1 U10604 ( .C1(n9599), .C2(n11082), .A(n9598), .B(n9597), .ZN(n9665)
         );
  MUX2_X1 U10605 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9665), .S(n11132), .Z(
        P2_U3548) );
  AOI22_X1 U10606 ( .A1(n9601), .A2(n11067), .B1(n11066), .B2(n9600), .ZN(
        n9602) );
  OAI211_X1 U10607 ( .C1(n9604), .C2(n11082), .A(n9603), .B(n9602), .ZN(n9666)
         );
  MUX2_X1 U10608 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9666), .S(n11132), .Z(
        P2_U3547) );
  AOI211_X1 U10609 ( .C1(n11066), .C2(n9607), .A(n9606), .B(n9605), .ZN(n9608)
         );
  OAI21_X1 U10610 ( .B1(n9609), .B2(n11082), .A(n9608), .ZN(n9667) );
  MUX2_X1 U10611 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9667), .S(n11132), .Z(
        P2_U3546) );
  AOI21_X1 U10612 ( .B1(n11066), .B2(n9611), .A(n9610), .ZN(n9612) );
  OAI211_X1 U10613 ( .C1(n9614), .C2(n11082), .A(n9613), .B(n9612), .ZN(n9668)
         );
  MUX2_X1 U10614 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9668), .S(n11132), .Z(
        P2_U3545) );
  AOI22_X1 U10615 ( .A1(n9616), .A2(n11067), .B1(n11066), .B2(n9615), .ZN(
        n9617) );
  OAI211_X1 U10616 ( .C1(n9619), .C2(n11082), .A(n9618), .B(n9617), .ZN(n9669)
         );
  MUX2_X1 U10617 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9669), .S(n11132), .Z(
        P2_U3544) );
  AOI22_X1 U10618 ( .A1(n9621), .A2(n11067), .B1(n11066), .B2(n9620), .ZN(
        n9622) );
  OAI211_X1 U10619 ( .C1(n9624), .C2(n11082), .A(n9623), .B(n9622), .ZN(n9670)
         );
  MUX2_X1 U10620 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9670), .S(n11132), .Z(
        P2_U3543) );
  AOI22_X1 U10621 ( .A1(n9626), .A2(n11067), .B1(n11066), .B2(n9625), .ZN(
        n9627) );
  OAI211_X1 U10622 ( .C1(n9629), .C2(n11082), .A(n9628), .B(n9627), .ZN(n9671)
         );
  MUX2_X1 U10623 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9671), .S(n11132), .Z(
        P2_U3542) );
  AOI22_X1 U10624 ( .A1(n9631), .A2(n11067), .B1(n11066), .B2(n9630), .ZN(
        n9632) );
  OAI211_X1 U10625 ( .C1(n9634), .C2(n11082), .A(n9633), .B(n9632), .ZN(n9672)
         );
  MUX2_X1 U10626 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9672), .S(n11132), .Z(
        P2_U3541) );
  AOI22_X1 U10627 ( .A1(n9636), .A2(n11067), .B1(n11066), .B2(n9635), .ZN(
        n9637) );
  OAI211_X1 U10628 ( .C1(n9639), .C2(n11082), .A(n9638), .B(n9637), .ZN(n9673)
         );
  MUX2_X1 U10629 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9673), .S(n11132), .Z(
        P2_U3540) );
  AOI211_X1 U10630 ( .C1(n11066), .C2(n9642), .A(n9641), .B(n9640), .ZN(n9643)
         );
  OAI21_X1 U10631 ( .B1(n9644), .B2(n11082), .A(n9643), .ZN(n9674) );
  MUX2_X1 U10632 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9674), .S(n11132), .Z(
        P2_U3539) );
  AOI22_X1 U10633 ( .A1(n9646), .A2(n11067), .B1(n11066), .B2(n9645), .ZN(
        n9647) );
  OAI211_X1 U10634 ( .C1(n9649), .C2(n11082), .A(n9648), .B(n9647), .ZN(n9675)
         );
  MUX2_X1 U10635 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9675), .S(n11132), .Z(
        P2_U3538) );
  INV_X1 U10636 ( .A(n9650), .ZN(n9656) );
  INV_X1 U10637 ( .A(n9651), .ZN(n9652) );
  AOI21_X1 U10638 ( .B1(n11066), .B2(n9653), .A(n9652), .ZN(n9654) );
  OAI211_X1 U10639 ( .C1(n9656), .C2(n11082), .A(n9655), .B(n9654), .ZN(n9676)
         );
  MUX2_X1 U10640 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9676), .S(n11132), .Z(
        P2_U3537) );
  AOI21_X1 U10641 ( .B1(n11066), .B2(n9658), .A(n9657), .ZN(n9659) );
  OAI211_X1 U10642 ( .C1(n9661), .C2(n11082), .A(n9660), .B(n9659), .ZN(n9677)
         );
  MUX2_X1 U10643 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9677), .S(n11132), .Z(
        P2_U3536) );
  MUX2_X1 U10644 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9662), .S(n11135), .Z(
        P2_U3519) );
  MUX2_X1 U10645 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9663), .S(n11135), .Z(
        P2_U3518) );
  MUX2_X1 U10646 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9665), .S(n11135), .Z(
        P2_U3516) );
  MUX2_X1 U10647 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9666), .S(n11135), .Z(
        P2_U3515) );
  MUX2_X1 U10648 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9667), .S(n11135), .Z(
        P2_U3514) );
  MUX2_X1 U10649 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9668), .S(n11135), .Z(
        P2_U3513) );
  MUX2_X1 U10650 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9669), .S(n11135), .Z(
        P2_U3512) );
  MUX2_X1 U10651 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9670), .S(n11135), .Z(
        P2_U3511) );
  MUX2_X1 U10652 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9671), .S(n11135), .Z(
        P2_U3510) );
  MUX2_X1 U10653 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9672), .S(n11135), .Z(
        P2_U3509) );
  MUX2_X1 U10654 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9673), .S(n11135), .Z(
        P2_U3508) );
  MUX2_X1 U10655 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9674), .S(n11135), .Z(
        P2_U3507) );
  MUX2_X1 U10656 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9675), .S(n11135), .Z(
        P2_U3505) );
  MUX2_X1 U10657 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9676), .S(n11135), .Z(
        P2_U3502) );
  MUX2_X1 U10658 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9677), .S(n11135), .Z(
        P2_U3499) );
  INV_X1 U10659 ( .A(n9678), .ZN(n10143) );
  NOR4_X1 U10660 ( .A1(n9680), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n9679), .ZN(n9681) );
  AOI21_X1 U10661 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9682), .A(n9681), .ZN(
        n9683) );
  OAI21_X1 U10662 ( .B1(n10143), .B2(n9684), .A(n9683), .ZN(P2_U3327) );
  INV_X1 U10663 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9685) );
  OAI222_X1 U10664 ( .A1(n9691), .A2(n9686), .B1(n9684), .B2(n10146), .C1(
        n9685), .C2(n9687), .ZN(P2_U3329) );
  INV_X1 U10665 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9688) );
  OAI222_X1 U10666 ( .A1(n9691), .A2(n9690), .B1(n9684), .B2(n9689), .C1(n9688), .C2(n9687), .ZN(P2_U3331) );
  MUX2_X1 U10667 ( .A(n9692), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10668 ( .A(n9693), .ZN(n9694) );
  NOR2_X1 U10669 ( .A1(n9695), .A2(n9694), .ZN(n9696) );
  XNOR2_X1 U10670 ( .A(n9697), .B(n9696), .ZN(n9703) );
  NAND2_X1 U10671 ( .A1(n9796), .A2(n9878), .ZN(n9699) );
  AOI22_X1 U10672 ( .A1(n9758), .A2(n9908), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9698) );
  OAI211_X1 U10673 ( .C1(n9700), .C2(n9756), .A(n9699), .B(n9698), .ZN(n9701)
         );
  AOI21_X1 U10674 ( .B1(n10062), .B2(n9773), .A(n9701), .ZN(n9702) );
  OAI21_X1 U10675 ( .B1(n9703), .B2(n9785), .A(n9702), .ZN(P1_U3212) );
  INV_X1 U10676 ( .A(n9704), .ZN(n9705) );
  NOR2_X1 U10677 ( .A1(n9706), .A2(n9705), .ZN(n9708) );
  XNOR2_X1 U10678 ( .A(n9708), .B(n9707), .ZN(n9714) );
  NAND2_X1 U10679 ( .A1(n9796), .A2(n9936), .ZN(n9710) );
  AOI22_X1 U10680 ( .A1(n9791), .A2(n9942), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9709) );
  OAI211_X1 U10681 ( .C1(n9711), .C2(n9793), .A(n9710), .B(n9709), .ZN(n9712)
         );
  AOI21_X1 U10682 ( .B1(n10082), .B2(n9773), .A(n9712), .ZN(n9713) );
  OAI21_X1 U10683 ( .B1(n9714), .B2(n9785), .A(n9713), .ZN(P1_U3214) );
  AOI21_X1 U10684 ( .B1(n9717), .B2(n9715), .A(n9716), .ZN(n9722) );
  NAND2_X1 U10685 ( .A1(n10001), .A2(n9791), .ZN(n9718) );
  NAND2_X1 U10686 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9841) );
  OAI211_X1 U10687 ( .C1(n10031), .C2(n9793), .A(n9718), .B(n9841), .ZN(n9720)
         );
  NOR2_X1 U10688 ( .A1(n9998), .A2(n9799), .ZN(n9719) );
  AOI211_X1 U10689 ( .C1(n9996), .C2(n9796), .A(n9720), .B(n9719), .ZN(n9721)
         );
  OAI21_X1 U10690 ( .B1(n9722), .B2(n9785), .A(n9721), .ZN(P1_U3217) );
  INV_X1 U10691 ( .A(n9723), .ZN(n9725) );
  NAND2_X1 U10692 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  XNOR2_X1 U10693 ( .A(n9727), .B(n9726), .ZN(n9732) );
  AOI22_X1 U10694 ( .A1(n9791), .A2(n9971), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9729) );
  NAND2_X1 U10695 ( .A1(n10001), .A2(n9758), .ZN(n9728) );
  OAI211_X1 U10696 ( .C1(n9760), .C2(n9964), .A(n9729), .B(n9728), .ZN(n9730)
         );
  AOI21_X1 U10697 ( .B1(n10093), .B2(n9773), .A(n9730), .ZN(n9731) );
  OAI21_X1 U10698 ( .B1(n9732), .B2(n9785), .A(n9731), .ZN(P1_U3221) );
  INV_X1 U10699 ( .A(n9733), .ZN(n9735) );
  NAND2_X1 U10700 ( .A1(n9735), .A2(n9734), .ZN(n9736) );
  XNOR2_X1 U10701 ( .A(n9737), .B(n9736), .ZN(n9743) );
  NAND2_X1 U10702 ( .A1(n9796), .A2(n9902), .ZN(n9739) );
  AOI22_X1 U10703 ( .A1(n9758), .A2(n9942), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9738) );
  OAI211_X1 U10704 ( .C1(n9740), .C2(n9756), .A(n9739), .B(n9738), .ZN(n9741)
         );
  AOI21_X1 U10705 ( .B1(n10072), .B2(n9773), .A(n9741), .ZN(n9742) );
  OAI21_X1 U10706 ( .B1(n9743), .B2(n9785), .A(n9742), .ZN(P1_U3223) );
  OAI21_X1 U10707 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(n9747) );
  NAND2_X1 U10708 ( .A1(n9747), .A2(n9787), .ZN(n9751) );
  AOI22_X1 U10709 ( .A1(n9758), .A2(n9954), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9748) );
  OAI21_X1 U10710 ( .B1(n9794), .B2(n9756), .A(n9748), .ZN(n9749) );
  AOI21_X1 U10711 ( .B1(n9796), .B2(n9925), .A(n9749), .ZN(n9750) );
  OAI211_X1 U10712 ( .C1(n9916), .C2(n9799), .A(n9751), .B(n9750), .ZN(
        P1_U3227) );
  XNOR2_X1 U10713 ( .A(n9753), .B(n9752), .ZN(n9754) );
  XNOR2_X1 U10714 ( .A(n5050), .B(n9754), .ZN(n9763) );
  OAI22_X1 U10715 ( .A1(n9771), .A2(n9756), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9755), .ZN(n9757) );
  AOI21_X1 U10716 ( .B1(n9758), .B2(n9985), .A(n9757), .ZN(n9759) );
  OAI21_X1 U10717 ( .B1(n9760), .B2(n9978), .A(n9759), .ZN(n9761) );
  AOI21_X1 U10718 ( .B1(n10097), .B2(n9773), .A(n9761), .ZN(n9762) );
  OAI21_X1 U10719 ( .B1(n9763), .B2(n9785), .A(n9762), .ZN(P1_U3231) );
  INV_X1 U10720 ( .A(n9764), .ZN(n9765) );
  NOR2_X1 U10721 ( .A1(n9766), .A2(n9765), .ZN(n9767) );
  XNOR2_X1 U10722 ( .A(n9768), .B(n9767), .ZN(n9775) );
  NAND2_X1 U10723 ( .A1(n9796), .A2(n9948), .ZN(n9770) );
  AOI22_X1 U10724 ( .A1(n9791), .A2(n9954), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9769) );
  OAI211_X1 U10725 ( .C1(n9771), .C2(n9793), .A(n9770), .B(n9769), .ZN(n9772)
         );
  AOI21_X1 U10726 ( .B1(n10087), .B2(n9773), .A(n9772), .ZN(n9774) );
  OAI21_X1 U10727 ( .B1(n9775), .B2(n9785), .A(n9774), .ZN(P1_U3233) );
  INV_X1 U10728 ( .A(n9776), .ZN(n9778) );
  NAND2_X1 U10729 ( .A1(n9778), .A2(n9777), .ZN(n9780) );
  XNOR2_X1 U10730 ( .A(n9780), .B(n9779), .ZN(n9786) );
  NAND2_X1 U10731 ( .A1(n9985), .A2(n9791), .ZN(n9781) );
  NAND2_X1 U10732 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10725)
         );
  OAI211_X1 U10733 ( .C1(n9793), .C2(n10018), .A(n9781), .B(n10725), .ZN(n9783) );
  NOR2_X1 U10734 ( .A1(n10011), .A2(n9799), .ZN(n9782) );
  AOI211_X1 U10735 ( .C1(n10009), .C2(n9796), .A(n9783), .B(n9782), .ZN(n9784)
         );
  OAI21_X1 U10736 ( .B1(n9786), .B2(n9785), .A(n9784), .ZN(P1_U3236) );
  INV_X1 U10737 ( .A(n10067), .ZN(n9889) );
  OAI211_X1 U10738 ( .C1(n9790), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9798)
         );
  AOI22_X1 U10739 ( .A1(n9791), .A2(n9893), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9792) );
  OAI21_X1 U10740 ( .B1(n9794), .B2(n9793), .A(n9792), .ZN(n9795) );
  AOI21_X1 U10741 ( .B1(n9796), .B2(n9887), .A(n9795), .ZN(n9797) );
  OAI211_X1 U10742 ( .C1(n9889), .C2(n9799), .A(n9798), .B(n9797), .ZN(
        P1_U3238) );
  MUX2_X1 U10743 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9800), .S(P1_U4006), .Z(
        P1_U3586) );
  INV_X2 U10744 ( .A(P1_U4006), .ZN(n9822) );
  MUX2_X1 U10745 ( .A(n9801), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9822), .Z(
        P1_U3584) );
  MUX2_X1 U10746 ( .A(n9870), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9822), .Z(
        P1_U3583) );
  MUX2_X1 U10747 ( .A(n9893), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9822), .Z(
        P1_U3582) );
  MUX2_X1 U10748 ( .A(n9908), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9822), .Z(
        P1_U3581) );
  MUX2_X1 U10749 ( .A(n9920), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9822), .Z(
        P1_U3580) );
  MUX2_X1 U10750 ( .A(n9942), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9822), .Z(
        P1_U3579) );
  MUX2_X1 U10751 ( .A(n9954), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9822), .Z(
        P1_U3578) );
  MUX2_X1 U10752 ( .A(n9971), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9822), .Z(
        P1_U3577) );
  MUX2_X1 U10753 ( .A(n9986), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9822), .Z(
        P1_U3576) );
  MUX2_X1 U10754 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10001), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10755 ( .A(n9802), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9822), .Z(
        P1_U3572) );
  MUX2_X1 U10756 ( .A(n9803), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9822), .Z(
        P1_U3571) );
  MUX2_X1 U10757 ( .A(n9804), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9822), .Z(
        P1_U3570) );
  MUX2_X1 U10758 ( .A(n9805), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9822), .Z(
        P1_U3568) );
  MUX2_X1 U10759 ( .A(n9806), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9822), .Z(
        P1_U3567) );
  MUX2_X1 U10760 ( .A(n9807), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9822), .Z(
        P1_U3566) );
  MUX2_X1 U10761 ( .A(n10991), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9822), .Z(
        P1_U3565) );
  MUX2_X1 U10762 ( .A(n9808), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9822), .Z(
        P1_U3564) );
  MUX2_X1 U10763 ( .A(n10992), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9822), .Z(
        P1_U3563) );
  MUX2_X1 U10764 ( .A(n9809), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9822), .Z(
        P1_U3562) );
  MUX2_X1 U10765 ( .A(n9810), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9822), .Z(
        P1_U3561) );
  MUX2_X1 U10766 ( .A(n9811), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9822), .Z(
        P1_U3560) );
  MUX2_X1 U10767 ( .A(n10862), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9822), .Z(
        P1_U3559) );
  MUX2_X1 U10768 ( .A(n5603), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9822), .Z(
        P1_U3558) );
  MUX2_X1 U10769 ( .A(n10863), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9822), .Z(
        P1_U3557) );
  MUX2_X1 U10770 ( .A(n7085), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9822), .Z(
        P1_U3556) );
  MUX2_X1 U10771 ( .A(n9812), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9822), .Z(
        P1_U3555) );
  INV_X1 U10772 ( .A(n9813), .ZN(n9815) );
  MUX2_X1 U10773 ( .A(n9815), .B(n9814), .S(n10675), .Z(n9817) );
  NOR2_X1 U10774 ( .A1(n9817), .A2(n9816), .ZN(n9823) );
  NAND2_X1 U10775 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  NAND2_X1 U10776 ( .A1(n9821), .A2(n9820), .ZN(n10670) );
  AND2_X1 U10777 ( .A1(n10670), .A2(n10674), .ZN(n10681) );
  NOR3_X1 U10778 ( .A1(n9823), .A2(n10681), .A3(n9822), .ZN(n10811) );
  INV_X1 U10779 ( .A(n10811), .ZN(n9836) );
  OAI21_X1 U10780 ( .B1(n9825), .B2(n5041), .A(n9824), .ZN(n9832) );
  AOI21_X1 U10781 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9830) );
  OAI21_X1 U10782 ( .B1(n10702), .B2(n9830), .A(n9829), .ZN(n9831) );
  AOI21_X1 U10783 ( .B1(n10746), .B2(n9832), .A(n9831), .ZN(n9835) );
  AOI22_X1 U10784 ( .A1(n10813), .A2(P1_ADDR_REG_4__SCAN_IN), .B1(n10744), 
        .B2(n9833), .ZN(n9834) );
  NAND3_X1 U10785 ( .A1(n9836), .A2(n9835), .A3(n9834), .ZN(P1_U3245) );
  AOI21_X1 U10786 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9843), .A(n9837), .ZN(
        n10719) );
  INV_X1 U10787 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9838) );
  AOI22_X1 U10788 ( .A1(n9846), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9838), .B2(
        n10727), .ZN(n10718) );
  NAND2_X1 U10789 ( .A1(n10719), .A2(n10718), .ZN(n10717) );
  OAI21_X1 U10790 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9846), .A(n10717), .ZN(
        n9840) );
  XNOR2_X1 U10791 ( .A(n9850), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9839) );
  XNOR2_X1 U10792 ( .A(n9840), .B(n9839), .ZN(n9851) );
  OR2_X1 U10793 ( .A1(n9846), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U10794 ( .A1(n9846), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U10795 ( .A1(n9845), .A2(n9844), .ZN(n10723) );
  AOI21_X1 U10796 ( .B1(n9846), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10721), .ZN(
        n9848) );
  XNOR2_X1 U10797 ( .A(n9850), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9847) );
  NOR2_X1 U10798 ( .A1(n9859), .A2(n10049), .ZN(n9853) );
  XNOR2_X1 U10799 ( .A(n9853), .B(n9852), .ZN(n10046) );
  NAND2_X1 U10800 ( .A1(n10046), .A2(n11009), .ZN(n9858) );
  INV_X1 U10801 ( .A(n9854), .ZN(n9855) );
  OR2_X1 U10802 ( .A1(n9856), .A2(n9855), .ZN(n10051) );
  NOR2_X1 U10803 ( .A1(n11014), .A2(n10051), .ZN(n9862) );
  AOI21_X1 U10804 ( .B1(n11014), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9862), .ZN(
        n9857) );
  OAI211_X1 U10805 ( .C1(n10048), .C2(n11016), .A(n9858), .B(n9857), .ZN(
        P1_U3261) );
  XNOR2_X1 U10806 ( .A(n10049), .B(n9859), .ZN(n10052) );
  INV_X1 U10807 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U10808 ( .A1(n11019), .A2(n9860), .ZN(n9861) );
  NOR2_X1 U10809 ( .A1(n9862), .A2(n9861), .ZN(n9865) );
  NAND2_X1 U10810 ( .A1(n10049), .A2(n9863), .ZN(n9864) );
  OAI211_X1 U10811 ( .C1(n10052), .C2(n9866), .A(n9865), .B(n9864), .ZN(
        P1_U3262) );
  NAND2_X1 U10812 ( .A1(n9890), .A2(n9867), .ZN(n9869) );
  XNOR2_X1 U10813 ( .A(n9869), .B(n9868), .ZN(n9874) );
  NAND2_X1 U10814 ( .A1(n9870), .A2(n10990), .ZN(n9872) );
  NAND2_X1 U10815 ( .A1(n9908), .A2(n10993), .ZN(n9871) );
  NAND2_X1 U10816 ( .A1(n10062), .A2(n9886), .ZN(n9876) );
  AND2_X1 U10817 ( .A1(n9877), .A2(n9876), .ZN(n10063) );
  AOI22_X1 U10818 ( .A1(n11014), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9878), 
        .B2(n11012), .ZN(n9879) );
  OAI21_X1 U10819 ( .B1(n8471), .B2(n11016), .A(n9879), .ZN(n9883) );
  XNOR2_X1 U10820 ( .A(n9881), .B(n9880), .ZN(n10066) );
  NOR2_X1 U10821 ( .A1(n10066), .A2(n10025), .ZN(n9882) );
  AOI211_X1 U10822 ( .C1(n10063), .C2(n11009), .A(n9883), .B(n9882), .ZN(n9884) );
  OAI21_X1 U10823 ( .B1(n10065), .B2(n11014), .A(n9884), .ZN(P1_U3264) );
  XNOR2_X1 U10824 ( .A(n9885), .B(n9892), .ZN(n10071) );
  AOI21_X1 U10825 ( .B1(n10067), .B2(n9899), .A(n9875), .ZN(n10068) );
  AOI22_X1 U10826 ( .A1(n11014), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9887), 
        .B2(n11012), .ZN(n9888) );
  OAI21_X1 U10827 ( .B1(n9889), .B2(n11016), .A(n9888), .ZN(n9896) );
  OAI21_X1 U10828 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9894) );
  NOR2_X1 U10829 ( .A1(n10070), .A2(n11014), .ZN(n9895) );
  AOI211_X1 U10830 ( .C1(n10068), .C2(n11009), .A(n9896), .B(n9895), .ZN(n9897) );
  OAI21_X1 U10831 ( .B1(n10071), .B2(n10025), .A(n9897), .ZN(P1_U3265) );
  XNOR2_X1 U10832 ( .A(n9898), .B(n9907), .ZN(n10076) );
  INV_X1 U10833 ( .A(n9924), .ZN(n9901) );
  INV_X1 U10834 ( .A(n9899), .ZN(n9900) );
  AOI21_X1 U10835 ( .B1(n10072), .B2(n9901), .A(n9900), .ZN(n10073) );
  AOI22_X1 U10836 ( .A1(n11014), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9902), 
        .B2(n11012), .ZN(n9903) );
  OAI21_X1 U10837 ( .B1(n9904), .B2(n11016), .A(n9903), .ZN(n9911) );
  OAI21_X1 U10838 ( .B1(n9907), .B2(n9906), .A(n9905), .ZN(n9909) );
  AOI222_X1 U10839 ( .A1(n10998), .A2(n9909), .B1(n9908), .B2(n10990), .C1(
        n9942), .C2(n10993), .ZN(n10075) );
  NOR2_X1 U10840 ( .A1(n10075), .A2(n11014), .ZN(n9910) );
  AOI211_X1 U10841 ( .C1(n10073), .C2(n11009), .A(n9911), .B(n9910), .ZN(n9912) );
  OAI21_X1 U10842 ( .B1(n10076), .B2(n10025), .A(n9912), .ZN(P1_U3266) );
  XNOR2_X1 U10843 ( .A(n9914), .B(n9915), .ZN(n10081) );
  NOR2_X1 U10844 ( .A1(n9916), .A2(n11016), .ZN(n9929) );
  OAI21_X1 U10845 ( .B1(n9919), .B2(n9918), .A(n9917), .ZN(n9921) );
  NAND2_X1 U10846 ( .A1(n10078), .A2(n9934), .ZN(n9922) );
  NAND2_X1 U10847 ( .A1(n9922), .A2(n10968), .ZN(n9923) );
  NOR2_X1 U10848 ( .A1(n9924), .A2(n9923), .ZN(n10077) );
  AOI22_X1 U10849 ( .A1(n10077), .A2(n9926), .B1(n11012), .B2(n9925), .ZN(
        n9927) );
  AOI21_X1 U10850 ( .B1(n10080), .B2(n9927), .A(n11014), .ZN(n9928) );
  AOI211_X1 U10851 ( .C1(n11014), .C2(P1_REG2_REG_24__SCAN_IN), .A(n9929), .B(
        n9928), .ZN(n9930) );
  OAI21_X1 U10852 ( .B1(n10025), .B2(n10081), .A(n9930), .ZN(P1_U3267) );
  XNOR2_X1 U10853 ( .A(n9931), .B(n9932), .ZN(n10086) );
  INV_X1 U10854 ( .A(n9934), .ZN(n9935) );
  AOI21_X1 U10855 ( .B1(n10082), .B2(n5232), .A(n9935), .ZN(n10083) );
  AOI22_X1 U10856 ( .A1(n11014), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9936), 
        .B2(n11012), .ZN(n9937) );
  OAI21_X1 U10857 ( .B1(n9938), .B2(n11016), .A(n9937), .ZN(n9945) );
  OAI21_X1 U10858 ( .B1(n9941), .B2(n9940), .A(n5109), .ZN(n9943) );
  AOI222_X1 U10859 ( .A1(n10998), .A2(n9943), .B1(n9942), .B2(n10990), .C1(
        n9971), .C2(n10993), .ZN(n10085) );
  NOR2_X1 U10860 ( .A1(n10085), .A2(n11014), .ZN(n9944) );
  AOI211_X1 U10861 ( .C1(n10083), .C2(n11009), .A(n9945), .B(n9944), .ZN(n9946) );
  OAI21_X1 U10862 ( .B1(n10025), .B2(n10086), .A(n9946), .ZN(P1_U3268) );
  XOR2_X1 U10863 ( .A(n9947), .B(n9953), .Z(n10091) );
  AOI21_X1 U10864 ( .B1(n10087), .B2(n9961), .A(n9933), .ZN(n10088) );
  INV_X1 U10865 ( .A(n10087), .ZN(n9950) );
  AOI22_X1 U10866 ( .A1(n11014), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9948), 
        .B2(n11012), .ZN(n9949) );
  OAI21_X1 U10867 ( .B1(n9950), .B2(n11016), .A(n9949), .ZN(n9957) );
  OAI21_X1 U10868 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9955) );
  AOI222_X1 U10869 ( .A1(n10998), .A2(n9955), .B1(n9954), .B2(n10990), .C1(
        n9986), .C2(n10993), .ZN(n10090) );
  NOR2_X1 U10870 ( .A1(n10090), .A2(n11014), .ZN(n9956) );
  AOI211_X1 U10871 ( .C1(n10088), .C2(n11009), .A(n9957), .B(n9956), .ZN(n9958) );
  OAI21_X1 U10872 ( .B1(n10025), .B2(n10091), .A(n9958), .ZN(P1_U3269) );
  OAI21_X1 U10873 ( .B1(n9960), .B2(n8346), .A(n9959), .ZN(n10096) );
  INV_X1 U10874 ( .A(n9977), .ZN(n9963) );
  INV_X1 U10875 ( .A(n9961), .ZN(n9962) );
  AOI211_X1 U10876 ( .C1(n10093), .C2(n9963), .A(n11111), .B(n9962), .ZN(
        n10092) );
  INV_X1 U10877 ( .A(n9964), .ZN(n9965) );
  AOI22_X1 U10878 ( .A1(n9965), .A2(n11012), .B1(n11014), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9966) );
  OAI21_X1 U10879 ( .B1(n9967), .B2(n11016), .A(n9966), .ZN(n9974) );
  OAI21_X1 U10880 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9972) );
  AOI222_X1 U10881 ( .A1(n10998), .A2(n9972), .B1(n9971), .B2(n10990), .C1(
        n10001), .C2(n10993), .ZN(n10095) );
  NOR2_X1 U10882 ( .A1(n10095), .A2(n11014), .ZN(n9973) );
  AOI211_X1 U10883 ( .C1(n10092), .C2(n10005), .A(n9974), .B(n9973), .ZN(n9975) );
  OAI21_X1 U10884 ( .B1(n10025), .B2(n10096), .A(n9975), .ZN(P1_U3270) );
  XNOR2_X1 U10885 ( .A(n9976), .B(n9984), .ZN(n10101) );
  AOI21_X1 U10886 ( .B1(n10097), .B2(n9993), .A(n9977), .ZN(n10098) );
  INV_X1 U10887 ( .A(n10097), .ZN(n9981) );
  INV_X1 U10888 ( .A(n9978), .ZN(n9979) );
  AOI22_X1 U10889 ( .A1(n9979), .A2(n11012), .B1(n11014), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9980) );
  OAI21_X1 U10890 ( .B1(n9981), .B2(n11016), .A(n9980), .ZN(n9989) );
  OAI21_X1 U10891 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(n9987) );
  AOI222_X1 U10892 ( .A1(n10998), .A2(n9987), .B1(n9986), .B2(n10990), .C1(
        n9985), .C2(n10993), .ZN(n10100) );
  NOR2_X1 U10893 ( .A1(n10100), .A2(n11014), .ZN(n9988) );
  AOI211_X1 U10894 ( .C1(n10098), .C2(n11009), .A(n9989), .B(n9988), .ZN(n9990) );
  OAI21_X1 U10895 ( .B1(n10101), .B2(n10025), .A(n9990), .ZN(P1_U3271) );
  XNOR2_X1 U10896 ( .A(n9991), .B(n9992), .ZN(n10106) );
  INV_X1 U10897 ( .A(n9998), .ZN(n10103) );
  INV_X1 U10898 ( .A(n10008), .ZN(n9995) );
  INV_X1 U10899 ( .A(n9993), .ZN(n9994) );
  AOI211_X1 U10900 ( .C1(n10103), .C2(n9995), .A(n11111), .B(n9994), .ZN(
        n10102) );
  AOI22_X1 U10901 ( .A1(n11014), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9996), 
        .B2(n11012), .ZN(n9997) );
  OAI21_X1 U10902 ( .B1(n9998), .B2(n11016), .A(n9997), .ZN(n10004) );
  OAI21_X1 U10903 ( .B1(n5646), .B2(n8460), .A(n9999), .ZN(n10002) );
  AOI222_X1 U10904 ( .A1(n10998), .A2(n10002), .B1(n10001), .B2(n10990), .C1(
        n10000), .C2(n10993), .ZN(n10105) );
  NOR2_X1 U10905 ( .A1(n10105), .A2(n11014), .ZN(n10003) );
  AOI211_X1 U10906 ( .C1(n10005), .C2(n10102), .A(n10004), .B(n10003), .ZN(
        n10006) );
  OAI21_X1 U10907 ( .B1(n10025), .B2(n10106), .A(n10006), .ZN(P1_U3272) );
  XNOR2_X1 U10908 ( .A(n10007), .B(n10017), .ZN(n10111) );
  AOI21_X1 U10909 ( .B1(n10107), .B2(n5236), .A(n10008), .ZN(n10108) );
  AOI22_X1 U10910 ( .A1(n11014), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10009), 
        .B2(n11012), .ZN(n10010) );
  OAI21_X1 U10911 ( .B1(n10011), .B2(n11016), .A(n10010), .ZN(n10023) );
  NAND2_X1 U10912 ( .A1(n10013), .A2(n10012), .ZN(n10016) );
  INV_X1 U10913 ( .A(n10014), .ZN(n10015) );
  AOI211_X1 U10914 ( .C1(n10017), .C2(n10016), .A(n10867), .B(n10015), .ZN(
        n10021) );
  OAI22_X1 U10915 ( .A1(n10019), .A2(n10030), .B1(n10018), .B2(n10028), .ZN(
        n10020) );
  NOR2_X1 U10916 ( .A1(n10021), .A2(n10020), .ZN(n10110) );
  NOR2_X1 U10917 ( .A1(n10110), .A2(n11014), .ZN(n10022) );
  AOI211_X1 U10918 ( .C1(n10108), .C2(n11009), .A(n10023), .B(n10022), .ZN(
        n10024) );
  OAI21_X1 U10919 ( .B1(n10025), .B2(n10111), .A(n10024), .ZN(P1_U3273) );
  XNOR2_X1 U10920 ( .A(n10027), .B(n10026), .ZN(n10036) );
  OAI22_X1 U10921 ( .A1(n10031), .A2(n10030), .B1(n10029), .B2(n10028), .ZN(
        n10035) );
  XNOR2_X1 U10922 ( .A(n10032), .B(n10033), .ZN(n10116) );
  NOR2_X1 U10923 ( .A1(n10116), .A2(n7103), .ZN(n10034) );
  AOI211_X1 U10924 ( .C1(n10036), .C2(n10998), .A(n10035), .B(n10034), .ZN(
        n10115) );
  AOI21_X1 U10925 ( .B1(n10112), .B2(n10038), .A(n10037), .ZN(n10113) );
  INV_X1 U10926 ( .A(n10112), .ZN(n10041) );
  AOI22_X1 U10927 ( .A1(n11014), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10039), 
        .B2(n11012), .ZN(n10040) );
  OAI21_X1 U10928 ( .B1(n10041), .B2(n11016), .A(n10040), .ZN(n10044) );
  NOR2_X1 U10929 ( .A1(n10116), .A2(n10042), .ZN(n10043) );
  AOI211_X1 U10930 ( .C1(n10113), .C2(n11009), .A(n10044), .B(n10043), .ZN(
        n10045) );
  OAI21_X1 U10931 ( .B1(n10115), .B2(n11014), .A(n10045), .ZN(P1_U3274) );
  NAND2_X1 U10932 ( .A1(n10046), .A2(n10968), .ZN(n10047) );
  OAI211_X1 U10933 ( .C1(n10048), .C2(n11109), .A(n10047), .B(n10051), .ZN(
        n10122) );
  MUX2_X1 U10934 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10122), .S(n10847), .Z(
        P1_U3554) );
  NAND2_X1 U10935 ( .A1(n10049), .A2(n11053), .ZN(n10050) );
  OAI211_X1 U10936 ( .C1(n10052), .C2(n11111), .A(n10051), .B(n10050), .ZN(
        n10123) );
  MUX2_X1 U10937 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10123), .S(n10847), .Z(
        P1_U3553) );
  AOI22_X1 U10938 ( .A1(n5042), .A2(n10968), .B1(n11053), .B2(n10053), .ZN(
        n10054) );
  OAI211_X1 U10939 ( .C1(n10911), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        n10124) );
  MUX2_X1 U10940 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10124), .S(n10847), .Z(
        P1_U3552) );
  AOI22_X1 U10941 ( .A1(n10058), .A2(n10968), .B1(n11053), .B2(n10057), .ZN(
        n10059) );
  AOI22_X1 U10942 ( .A1(n10063), .A2(n10968), .B1(n11053), .B2(n10062), .ZN(
        n10064) );
  OAI211_X1 U10943 ( .C1(n10911), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        n10126) );
  MUX2_X1 U10944 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10126), .S(n10900), .Z(
        P1_U3550) );
  AOI22_X1 U10945 ( .A1(n10068), .A2(n10968), .B1(n11053), .B2(n10067), .ZN(
        n10069) );
  OAI211_X1 U10946 ( .C1(n10911), .C2(n10071), .A(n10070), .B(n10069), .ZN(
        n10127) );
  MUX2_X1 U10947 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10127), .S(n10900), .Z(
        P1_U3549) );
  AOI22_X1 U10948 ( .A1(n10073), .A2(n10968), .B1(n11053), .B2(n10072), .ZN(
        n10074) );
  OAI211_X1 U10949 ( .C1(n10911), .C2(n10076), .A(n10075), .B(n10074), .ZN(
        n10128) );
  MUX2_X1 U10950 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10128), .S(n10847), .Z(
        P1_U3548) );
  AOI21_X1 U10951 ( .B1(n11053), .B2(n10078), .A(n10077), .ZN(n10079) );
  OAI211_X1 U10952 ( .C1(n10911), .C2(n10081), .A(n10080), .B(n10079), .ZN(
        n10129) );
  MUX2_X1 U10953 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10129), .S(n10847), .Z(
        P1_U3547) );
  AOI22_X1 U10954 ( .A1(n10083), .A2(n10968), .B1(n11053), .B2(n10082), .ZN(
        n10084) );
  OAI211_X1 U10955 ( .C1(n10911), .C2(n10086), .A(n10085), .B(n10084), .ZN(
        n10130) );
  MUX2_X1 U10956 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10130), .S(n10847), .Z(
        P1_U3546) );
  AOI22_X1 U10957 ( .A1(n10088), .A2(n10968), .B1(n11053), .B2(n10087), .ZN(
        n10089) );
  OAI211_X1 U10958 ( .C1(n10091), .C2(n10911), .A(n10090), .B(n10089), .ZN(
        n10131) );
  MUX2_X1 U10959 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10131), .S(n10847), .Z(
        P1_U3545) );
  AOI21_X1 U10960 ( .B1(n11053), .B2(n10093), .A(n10092), .ZN(n10094) );
  OAI211_X1 U10961 ( .C1(n10911), .C2(n10096), .A(n10095), .B(n10094), .ZN(
        n10132) );
  MUX2_X1 U10962 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10132), .S(n10847), .Z(
        P1_U3544) );
  AOI22_X1 U10963 ( .A1(n10098), .A2(n10968), .B1(n11053), .B2(n10097), .ZN(
        n10099) );
  OAI211_X1 U10964 ( .C1(n10911), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10133) );
  MUX2_X1 U10965 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10133), .S(n10847), .Z(
        P1_U3543) );
  AOI21_X1 U10966 ( .B1(n11053), .B2(n10103), .A(n10102), .ZN(n10104) );
  OAI211_X1 U10967 ( .C1(n10911), .C2(n10106), .A(n10105), .B(n10104), .ZN(
        n10134) );
  MUX2_X1 U10968 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10134), .S(n10847), .Z(
        P1_U3542) );
  AOI22_X1 U10969 ( .A1(n10108), .A2(n10968), .B1(n11053), .B2(n10107), .ZN(
        n10109) );
  OAI211_X1 U10970 ( .C1(n10911), .C2(n10111), .A(n10110), .B(n10109), .ZN(
        n10135) );
  MUX2_X1 U10971 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10135), .S(n10847), .Z(
        P1_U3541) );
  AOI22_X1 U10972 ( .A1(n10113), .A2(n10968), .B1(n11053), .B2(n10112), .ZN(
        n10114) );
  OAI211_X1 U10973 ( .C1(n11057), .C2(n10116), .A(n10115), .B(n10114), .ZN(
        n10136) );
  MUX2_X1 U10974 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10136), .S(n10847), .Z(
        P1_U3540) );
  AOI211_X1 U10975 ( .C1(n11053), .C2(n10119), .A(n10118), .B(n10117), .ZN(
        n10120) );
  OAI21_X1 U10976 ( .B1(n10911), .B2(n10121), .A(n10120), .ZN(n10138) );
  MUX2_X1 U10977 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10138), .S(n10847), .Z(
        P1_U3539) );
  MUX2_X1 U10978 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10122), .S(n10137), .Z(
        P1_U3522) );
  MUX2_X1 U10979 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10123), .S(n10137), .Z(
        P1_U3521) );
  MUX2_X1 U10980 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10124), .S(n10137), .Z(
        P1_U3520) );
  MUX2_X1 U10981 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10125), .S(n10137), .Z(
        P1_U3519) );
  MUX2_X1 U10982 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10126), .S(n10137), .Z(
        P1_U3518) );
  MUX2_X1 U10983 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10127), .S(n10137), .Z(
        P1_U3517) );
  MUX2_X1 U10984 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10128), .S(n10137), .Z(
        P1_U3516) );
  MUX2_X1 U10985 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10129), .S(n10137), .Z(
        P1_U3515) );
  MUX2_X1 U10986 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10130), .S(n10137), .Z(
        P1_U3514) );
  MUX2_X1 U10987 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10131), .S(n10137), .Z(
        P1_U3513) );
  MUX2_X1 U10988 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10132), .S(n10137), .Z(
        P1_U3512) );
  MUX2_X1 U10989 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10133), .S(n10137), .Z(
        P1_U3511) );
  MUX2_X1 U10990 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10134), .S(n10137), .Z(
        P1_U3510) );
  MUX2_X1 U10991 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10135), .S(n10137), .Z(
        P1_U3508) );
  MUX2_X1 U10992 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10136), .S(n10137), .Z(
        P1_U3505) );
  MUX2_X1 U10993 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10138), .S(n10137), .Z(
        P1_U3502) );
  NOR4_X1 U10994 ( .A1(n6470), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n10139), .ZN(n10140) );
  AOI21_X1 U10995 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10141), .A(n10140), 
        .ZN(n10142) );
  OAI21_X1 U10996 ( .B1(n10143), .B2(n10147), .A(n10142), .ZN(P1_U3322) );
  INV_X1 U10997 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10381) );
  OAI222_X1 U10998 ( .A1(n10147), .A2(n10146), .B1(n10145), .B2(P1_U3084), 
        .C1(n10381), .C2(n10144), .ZN(P1_U3324) );
  INV_X1 U10999 ( .A(n10148), .ZN(n10149) );
  MUX2_X1 U11000 ( .A(n10149), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11001 ( .A1(n10151), .A2(n10150), .ZN(n10181) );
  INV_X1 U11002 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10372) );
  NOR2_X1 U11003 ( .A1(n10169), .A2(n10372), .ZN(P1_U3321) );
  INV_X1 U11004 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10188) );
  NOR2_X1 U11005 ( .A1(n10169), .A2(n10188), .ZN(P1_U3320) );
  INV_X1 U11006 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10152) );
  NOR2_X1 U11007 ( .A1(n10169), .A2(n10152), .ZN(P1_U3319) );
  INV_X1 U11008 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10153) );
  NOR2_X1 U11009 ( .A1(n10169), .A2(n10153), .ZN(P1_U3318) );
  INV_X1 U11010 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10154) );
  NOR2_X1 U11011 ( .A1(n10169), .A2(n10154), .ZN(P1_U3317) );
  INV_X1 U11012 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10155) );
  NOR2_X1 U11013 ( .A1(n10169), .A2(n10155), .ZN(P1_U3316) );
  INV_X1 U11014 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10156) );
  NOR2_X1 U11015 ( .A1(n10169), .A2(n10156), .ZN(P1_U3315) );
  INV_X1 U11016 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10157) );
  NOR2_X1 U11017 ( .A1(n10169), .A2(n10157), .ZN(P1_U3314) );
  INV_X1 U11018 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10158) );
  NOR2_X1 U11019 ( .A1(n10169), .A2(n10158), .ZN(P1_U3313) );
  INV_X1 U11020 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10159) );
  NOR2_X1 U11021 ( .A1(n10169), .A2(n10159), .ZN(P1_U3312) );
  INV_X1 U11022 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10160) );
  NOR2_X1 U11023 ( .A1(n10169), .A2(n10160), .ZN(P1_U3311) );
  INV_X1 U11024 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10161) );
  NOR2_X1 U11025 ( .A1(n10169), .A2(n10161), .ZN(P1_U3310) );
  INV_X1 U11026 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10162) );
  NOR2_X1 U11027 ( .A1(n10169), .A2(n10162), .ZN(P1_U3309) );
  INV_X1 U11028 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10163) );
  NOR2_X1 U11029 ( .A1(n10169), .A2(n10163), .ZN(P1_U3308) );
  INV_X1 U11030 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10164) );
  NOR2_X1 U11031 ( .A1(n10169), .A2(n10164), .ZN(P1_U3307) );
  INV_X1 U11032 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10165) );
  NOR2_X1 U11033 ( .A1(n10169), .A2(n10165), .ZN(P1_U3306) );
  INV_X1 U11034 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10166) );
  NOR2_X1 U11035 ( .A1(n10169), .A2(n10166), .ZN(P1_U3305) );
  INV_X1 U11036 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10167) );
  NOR2_X1 U11037 ( .A1(n10169), .A2(n10167), .ZN(P1_U3304) );
  INV_X1 U11038 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10168) );
  NOR2_X1 U11039 ( .A1(n10169), .A2(n10168), .ZN(P1_U3303) );
  INV_X1 U11040 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10170) );
  NOR2_X1 U11041 ( .A1(n10181), .A2(n10170), .ZN(P1_U3302) );
  INV_X1 U11042 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10171) );
  NOR2_X1 U11043 ( .A1(n10181), .A2(n10171), .ZN(P1_U3301) );
  INV_X1 U11044 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10172) );
  NOR2_X1 U11045 ( .A1(n10181), .A2(n10172), .ZN(P1_U3300) );
  INV_X1 U11046 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10173) );
  NOR2_X1 U11047 ( .A1(n10181), .A2(n10173), .ZN(P1_U3299) );
  INV_X1 U11048 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10174) );
  NOR2_X1 U11049 ( .A1(n10181), .A2(n10174), .ZN(P1_U3298) );
  INV_X1 U11050 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10175) );
  NOR2_X1 U11051 ( .A1(n10181), .A2(n10175), .ZN(P1_U3297) );
  INV_X1 U11052 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10176) );
  NOR2_X1 U11053 ( .A1(n10181), .A2(n10176), .ZN(P1_U3296) );
  INV_X1 U11054 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10177) );
  NOR2_X1 U11055 ( .A1(n10181), .A2(n10177), .ZN(P1_U3295) );
  INV_X1 U11056 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10178) );
  NOR2_X1 U11057 ( .A1(n10181), .A2(n10178), .ZN(P1_U3294) );
  INV_X1 U11058 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10179) );
  NOR2_X1 U11059 ( .A1(n10181), .A2(n10179), .ZN(P1_U3293) );
  INV_X1 U11060 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10180) );
  NOR2_X1 U11061 ( .A1(n10181), .A2(n10180), .ZN(P1_U3292) );
  INV_X1 U11062 ( .A(n10182), .ZN(n10187) );
  INV_X1 U11063 ( .A(n10183), .ZN(n10184) );
  AOI22_X1 U11064 ( .A1(n10760), .A2(n10187), .B1(n10186), .B2(n10757), .ZN(
        P2_U3438) );
  AND2_X1 U11065 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10757), .ZN(P2_U3326) );
  AND2_X1 U11066 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10757), .ZN(P2_U3325) );
  AND2_X1 U11067 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10757), .ZN(P2_U3324) );
  AND2_X1 U11068 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10757), .ZN(P2_U3323) );
  AND2_X1 U11069 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10757), .ZN(P2_U3322) );
  AND2_X1 U11070 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10757), .ZN(P2_U3321) );
  AND2_X1 U11071 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10757), .ZN(P2_U3320) );
  AND2_X1 U11072 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10757), .ZN(P2_U3319) );
  AND2_X1 U11073 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10757), .ZN(P2_U3318) );
  AND2_X1 U11074 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10757), .ZN(P2_U3317) );
  AND2_X1 U11075 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10757), .ZN(P2_U3316) );
  AND2_X1 U11076 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10757), .ZN(P2_U3315) );
  AND2_X1 U11077 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10757), .ZN(P2_U3314) );
  AND2_X1 U11078 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10757), .ZN(P2_U3313) );
  AND2_X1 U11079 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10757), .ZN(P2_U3312) );
  AND2_X1 U11080 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10757), .ZN(P2_U3311) );
  AND2_X1 U11081 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10757), .ZN(P2_U3310) );
  AND2_X1 U11082 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10757), .ZN(P2_U3309) );
  AND2_X1 U11083 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10757), .ZN(P2_U3308) );
  AND2_X1 U11084 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10757), .ZN(P2_U3307) );
  AND2_X1 U11085 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10757), .ZN(P2_U3306) );
  AND2_X1 U11086 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10757), .ZN(P2_U3305) );
  AND2_X1 U11087 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10757), .ZN(P2_U3304) );
  AND2_X1 U11088 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10757), .ZN(P2_U3303) );
  AND2_X1 U11089 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10757), .ZN(P2_U3302) );
  AND2_X1 U11090 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10757), .ZN(P2_U3301) );
  AND2_X1 U11091 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10757), .ZN(P2_U3300) );
  AND2_X1 U11092 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10757), .ZN(P2_U3299) );
  AND2_X1 U11093 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10757), .ZN(P2_U3298) );
  AND2_X1 U11094 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10757), .ZN(P2_U3297) );
  XNOR2_X1 U11095 ( .A(keyinput_126), .B(n10188), .ZN(n10604) );
  INV_X1 U11096 ( .A(keyinput_107), .ZN(n10346) );
  OAI22_X1 U11097 ( .A1(n10190), .A2(keyinput_105), .B1(keyinput_106), .B2(
        P1_IR_REG_15__SCAN_IN), .ZN(n10189) );
  AOI221_X1 U11098 ( .B1(n10190), .B2(keyinput_105), .C1(P1_IR_REG_15__SCAN_IN), .C2(keyinput_106), .A(n10189), .ZN(n10345) );
  INV_X1 U11099 ( .A(keyinput_87), .ZN(n10319) );
  INV_X1 U11100 ( .A(keyinput_86), .ZN(n10318) );
  INV_X1 U11101 ( .A(keyinput_85), .ZN(n10317) );
  OAI22_X1 U11102 ( .A1(n10525), .A2(keyinput_84), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_83), .ZN(n10191) );
  AOI221_X1 U11103 ( .B1(n10525), .B2(keyinput_84), .C1(keyinput_83), .C2(
        P2_DATAO_REG_13__SCAN_IN), .A(n10191), .ZN(n10315) );
  INV_X1 U11104 ( .A(keyinput_66), .ZN(n10294) );
  INV_X1 U11105 ( .A(keyinput_64), .ZN(n10290) );
  OAI22_X1 U11106 ( .A1(n10490), .A2(keyinput_57), .B1(keyinput_56), .B2(
        P2_REG3_REG_13__SCAN_IN), .ZN(n10192) );
  AOI221_X1 U11107 ( .B1(n10490), .B2(keyinput_57), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_56), .A(n10192), .ZN(n10282) );
  INV_X1 U11108 ( .A(keyinput_52), .ZN(n10273) );
  INV_X1 U11109 ( .A(keyinput_51), .ZN(n10272) );
  XNOR2_X1 U11110 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n10270)
         );
  INV_X1 U11111 ( .A(keyinput_45), .ZN(n10264) );
  INV_X1 U11112 ( .A(keyinput_41), .ZN(n10256) );
  INV_X1 U11113 ( .A(keyinput_40), .ZN(n10254) );
  INV_X1 U11114 ( .A(keyinput_38), .ZN(n10248) );
  AOI22_X1 U11115 ( .A1(n9212), .A2(keyinput_36), .B1(n10445), .B2(keyinput_35), .ZN(n10193) );
  OAI221_X1 U11116 ( .B1(n9212), .B2(keyinput_36), .C1(n10445), .C2(
        keyinput_35), .A(n10193), .ZN(n10246) );
  INV_X1 U11117 ( .A(SI_0_), .ZN(n10438) );
  AOI22_X1 U11118 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_33), .B1(n10438), 
        .B2(keyinput_32), .ZN(n10194) );
  OAI221_X1 U11119 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_33), .C1(n10438), 
        .C2(keyinput_32), .A(n10194), .ZN(n10243) );
  INV_X1 U11120 ( .A(SI_1_), .ZN(n10436) );
  INV_X1 U11121 ( .A(keyinput_31), .ZN(n10242) );
  INV_X1 U11122 ( .A(SI_6_), .ZN(n10427) );
  OAI22_X1 U11123 ( .A1(n10427), .A2(keyinput_26), .B1(SI_5_), .B2(keyinput_27), .ZN(n10195) );
  AOI221_X1 U11124 ( .B1(n10427), .B2(keyinput_26), .C1(keyinput_27), .C2(
        SI_5_), .A(n10195), .ZN(n10241) );
  AOI22_X1 U11125 ( .A1(SI_27_), .A2(keyinput_5), .B1(n10395), .B2(keyinput_7), 
        .ZN(n10196) );
  OAI221_X1 U11126 ( .B1(SI_27_), .B2(keyinput_5), .C1(n10395), .C2(keyinput_7), .A(n10196), .ZN(n10197) );
  INV_X1 U11127 ( .A(n10197), .ZN(n10204) );
  AOI22_X1 U11128 ( .A1(SI_29_), .A2(keyinput_3), .B1(SI_24_), .B2(keyinput_8), 
        .ZN(n10198) );
  OAI221_X1 U11129 ( .B1(SI_29_), .B2(keyinput_3), .C1(SI_24_), .C2(keyinput_8), .A(n10198), .ZN(n10199) );
  INV_X1 U11130 ( .A(n10199), .ZN(n10203) );
  AOI22_X1 U11131 ( .A1(SI_28_), .A2(keyinput_4), .B1(SI_23_), .B2(keyinput_9), 
        .ZN(n10200) );
  OAI221_X1 U11132 ( .B1(SI_28_), .B2(keyinput_4), .C1(SI_23_), .C2(keyinput_9), .A(n10200), .ZN(n10201) );
  INV_X1 U11133 ( .A(n10201), .ZN(n10202) );
  AND4_X1 U11134 ( .A1(n5633), .A2(n10204), .A3(n10203), .A4(n10202), .ZN(
        n10213) );
  INV_X1 U11135 ( .A(keyinput_2), .ZN(n10206) );
  INV_X1 U11136 ( .A(SI_30_), .ZN(n10401) );
  OAI221_X1 U11137 ( .B1(SI_30_), .B2(n10206), .C1(n10401), .C2(keyinput_2), 
        .A(n10205), .ZN(n10212) );
  AOI22_X1 U11138 ( .A1(SI_22_), .A2(keyinput_10), .B1(n10208), .B2(
        keyinput_13), .ZN(n10207) );
  OAI221_X1 U11139 ( .B1(SI_22_), .B2(keyinput_10), .C1(n10208), .C2(
        keyinput_13), .A(n10207), .ZN(n10211) );
  AOI22_X1 U11140 ( .A1(SI_20_), .A2(keyinput_12), .B1(SI_21_), .B2(
        keyinput_11), .ZN(n10209) );
  OAI221_X1 U11141 ( .B1(SI_20_), .B2(keyinput_12), .C1(SI_21_), .C2(
        keyinput_11), .A(n10209), .ZN(n10210) );
  AOI211_X1 U11142 ( .C1(n10213), .C2(n10212), .A(n10211), .B(n10210), .ZN(
        n10214) );
  INV_X1 U11143 ( .A(SI_18_), .ZN(n10414) );
  AOI22_X1 U11144 ( .A1(SI_17_), .A2(keyinput_15), .B1(n10414), .B2(
        keyinput_14), .ZN(n10215) );
  OAI221_X1 U11145 ( .B1(SI_17_), .B2(keyinput_15), .C1(n10414), .C2(
        keyinput_14), .A(n10215), .ZN(n10216) );
  INV_X1 U11146 ( .A(n10216), .ZN(n10219) );
  AOI21_X1 U11147 ( .B1(n10220), .B2(n10219), .A(n10218), .ZN(n10226) );
  AOI22_X1 U11148 ( .A1(SI_15_), .A2(keyinput_17), .B1(n10222), .B2(
        keyinput_18), .ZN(n10221) );
  OAI221_X1 U11149 ( .B1(SI_15_), .B2(keyinput_17), .C1(n10222), .C2(
        keyinput_18), .A(n10221), .ZN(n10225) );
  AOI22_X1 U11150 ( .A1(SI_12_), .A2(keyinput_20), .B1(SI_13_), .B2(
        keyinput_19), .ZN(n10223) );
  OAI221_X1 U11151 ( .B1(SI_12_), .B2(keyinput_20), .C1(SI_13_), .C2(
        keyinput_19), .A(n10223), .ZN(n10224) );
  NOR3_X1 U11152 ( .A1(n10226), .A2(n10225), .A3(n10224), .ZN(n10232) );
  AOI22_X1 U11153 ( .A1(SI_11_), .A2(keyinput_21), .B1(n10228), .B2(
        keyinput_22), .ZN(n10227) );
  OAI221_X1 U11154 ( .B1(SI_11_), .B2(keyinput_21), .C1(n10228), .C2(
        keyinput_22), .A(n10227), .ZN(n10231) );
  OAI22_X1 U11155 ( .A1(n10234), .A2(keyinput_24), .B1(SI_7_), .B2(keyinput_25), .ZN(n10233) );
  AOI221_X1 U11156 ( .B1(n10234), .B2(keyinput_24), .C1(keyinput_25), .C2(
        SI_7_), .A(n10233), .ZN(n10235) );
  XOR2_X1 U11157 ( .A(SI_2_), .B(keyinput_30), .Z(n10239) );
  INV_X1 U11158 ( .A(SI_4_), .ZN(n10429) );
  AOI22_X1 U11159 ( .A1(SI_3_), .A2(keyinput_29), .B1(n10429), .B2(keyinput_28), .ZN(n10237) );
  OAI221_X1 U11160 ( .B1(SI_3_), .B2(keyinput_29), .C1(n10429), .C2(
        keyinput_28), .A(n10237), .ZN(n10238) );
  NAND2_X1 U11161 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .ZN(n10244) );
  OAI221_X1 U11162 ( .B1(n10246), .B2(n10245), .C1(P2_REG3_REG_14__SCAN_IN), 
        .C2(keyinput_37), .A(n10244), .ZN(n10247) );
  OAI221_X1 U11163 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        n10452), .C2(n10248), .A(n10247), .ZN(n10252) );
  INV_X1 U11164 ( .A(keyinput_39), .ZN(n10249) );
  OAI22_X1 U11165 ( .A1(n10455), .A2(n10249), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(keyinput_39), .ZN(n10250) );
  INV_X1 U11166 ( .A(n10250), .ZN(n10251) );
  NAND2_X1 U11167 ( .A1(n10252), .A2(n10251), .ZN(n10253) );
  OAI221_X1 U11168 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10254), .C1(n10458), 
        .C2(keyinput_40), .A(n10253), .ZN(n10255) );
  OAI221_X1 U11169 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n10256), .C1(n6158), 
        .C2(keyinput_41), .A(n10255), .ZN(n10261) );
  OAI22_X1 U11170 ( .A1(n10258), .A2(keyinput_43), .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_42), .ZN(n10257) );
  AOI221_X1 U11171 ( .B1(n10258), .B2(keyinput_43), .C1(keyinput_42), .C2(
        P2_REG3_REG_28__SCAN_IN), .A(n10257), .ZN(n10260) );
  XNOR2_X1 U11172 ( .A(keyinput_44), .B(P2_REG3_REG_1__SCAN_IN), .ZN(n10259)
         );
  INV_X1 U11173 ( .A(n10262), .ZN(n10263) );
  OAI221_X1 U11174 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(n10264), .C1(n10471), 
        .C2(keyinput_45), .A(n10263), .ZN(n10269) );
  AOI22_X1 U11175 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_49), .B1(n10474), 
        .B2(keyinput_48), .ZN(n10265) );
  OAI221_X1 U11176 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(n10474), .C2(keyinput_48), .A(n10265), .ZN(n10268) );
  AOI22_X1 U11177 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_47), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .ZN(n10266) );
  OAI221_X1 U11178 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_50), .A(n10266), .ZN(n10267) );
  AOI211_X1 U11179 ( .C1(n10270), .C2(n10269), .A(n10268), .B(n10267), .ZN(
        n10271) );
  AOI22_X1 U11180 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_55), .B1(n5992), 
        .B2(keyinput_53), .ZN(n10274) );
  OAI221_X1 U11181 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(n5992), .C2(keyinput_53), .A(n10274), .ZN(n10276) );
  XOR2_X1 U11182 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .Z(n10280) );
  AOI22_X1 U11183 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .ZN(n10278) );
  OAI221_X1 U11184 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_58), .A(n10278), .ZN(n10279) );
  AOI211_X1 U11185 ( .C1(n10282), .C2(n10281), .A(n10280), .B(n10279), .ZN(
        n10289) );
  AOI22_X1 U11186 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_63), .B1(n10284), .B2(keyinput_62), .ZN(n10283) );
  OAI221_X1 U11187 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_63), .C1(
        n10284), .C2(keyinput_62), .A(n10283), .ZN(n10285) );
  INV_X1 U11188 ( .A(n10285), .ZN(n10287) );
  INV_X1 U11189 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10502) );
  INV_X1 U11190 ( .A(keyinput_65), .ZN(n10291) );
  OAI22_X1 U11191 ( .A1(n10502), .A2(keyinput_65), .B1(n10291), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n10292) );
  INV_X1 U11192 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U11193 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_73), .B1(
        n10379), .B2(keyinput_68), .ZN(n10295) );
  OAI221_X1 U11194 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_73), .C1(
        n10379), .C2(keyinput_68), .A(n10295), .ZN(n10302) );
  AOI22_X1 U11195 ( .A1(n5753), .A2(keyinput_70), .B1(keyinput_72), .B2(n10382), .ZN(n10296) );
  OAI221_X1 U11196 ( .B1(n5753), .B2(keyinput_70), .C1(n10382), .C2(
        keyinput_72), .A(n10296), .ZN(n10301) );
  AOI22_X1 U11197 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_67), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_74), .ZN(n10297) );
  OAI221_X1 U11198 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_67), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput_74), .A(n10297), .ZN(n10300)
         );
  AOI22_X1 U11199 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput_71), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_69), .ZN(n10298) );
  OAI221_X1 U11200 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_71), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_69), .A(n10298), .ZN(n10299)
         );
  NOR4_X1 U11201 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10304) );
  XNOR2_X1 U11202 ( .A(n10510), .B(keyinput_75), .ZN(n10303) );
  AOI22_X1 U11203 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput_77), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_76), .ZN(n10307) );
  OAI221_X1 U11204 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_77), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_76), .A(n10307), .ZN(n10309)
         );
  NAND2_X1 U11205 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_78), .ZN(
        n10308) );
  OAI22_X1 U11206 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_79), .B1(
        keyinput_80), .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n10310) );
  AOI221_X1 U11207 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_79), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_80), .A(n10310), .ZN(n10312)
         );
  OAI211_X1 U11208 ( .C1(n10522), .C2(keyinput_82), .A(n10315), .B(n10314), 
        .ZN(n10316) );
  AOI22_X1 U11209 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_89), .B1(n10321), .B2(keyinput_88), .ZN(n10320) );
  OAI221_X1 U11210 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_89), .C1(
        n10321), .C2(keyinput_88), .A(n10320), .ZN(n10329) );
  OAI22_X1 U11211 ( .A1(n10674), .A2(keyinput_91), .B1(n10540), .B2(
        keyinput_93), .ZN(n10322) );
  AOI221_X1 U11212 ( .B1(n10674), .B2(keyinput_91), .C1(keyinput_93), .C2(
        n10540), .A(n10322), .ZN(n10328) );
  XNOR2_X1 U11213 ( .A(n10543), .B(keyinput_90), .ZN(n10326) );
  XNOR2_X1 U11214 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n10325) );
  XNOR2_X1 U11215 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .ZN(n10324) );
  XNOR2_X1 U11216 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .ZN(n10323) );
  AND4_X1 U11217 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10327) );
  OAI211_X1 U11218 ( .C1(n10330), .C2(n10329), .A(n10328), .B(n10327), .ZN(
        n10339) );
  OAI22_X1 U11219 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_97), .B1(
        keyinput_99), .B2(P1_IR_REG_8__SCAN_IN), .ZN(n10331) );
  AOI221_X1 U11220 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_97), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_99), .A(n10331), .ZN(n10338) );
  AOI22_X1 U11221 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_101), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput_100), .ZN(n10332) );
  OAI221_X1 U11222 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_101), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_100), .A(n10332), .ZN(n10336) );
  XNOR2_X1 U11223 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .ZN(n10334) );
  XNOR2_X1 U11224 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_98), .ZN(n10333) );
  NAND3_X1 U11225 ( .A1(n10339), .A2(n10338), .A3(n10337), .ZN(n10343) );
  INV_X1 U11226 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10341) );
  OAI22_X1 U11227 ( .A1(n10341), .A2(keyinput_102), .B1(keyinput_103), .B2(
        P1_IR_REG_12__SCAN_IN), .ZN(n10340) );
  AOI221_X1 U11228 ( .B1(n10341), .B2(keyinput_102), .C1(P1_IR_REG_12__SCAN_IN), .C2(keyinput_103), .A(n10340), .ZN(n10342) );
  NAND2_X1 U11229 ( .A1(n10343), .A2(n10342), .ZN(n10344) );
  AOI22_X1 U11230 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_109), .B1(n10572), 
        .B2(keyinput_108), .ZN(n10347) );
  OAI221_X1 U11231 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_109), .C1(n10572), .C2(keyinput_108), .A(n10347), .ZN(n10349) );
  OAI22_X1 U11232 ( .A1(n10353), .A2(keyinput_111), .B1(keyinput_112), .B2(
        P1_IR_REG_21__SCAN_IN), .ZN(n10352) );
  AOI221_X1 U11233 ( .B1(n10353), .B2(keyinput_111), .C1(P1_IR_REG_21__SCAN_IN), .C2(keyinput_112), .A(n10352), .ZN(n10358) );
  XOR2_X1 U11234 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_113), .Z(n10357) );
  XNOR2_X1 U11235 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_115), .ZN(n10355)
         );
  XNOR2_X1 U11236 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_114), .ZN(n10354)
         );
  NAND2_X1 U11237 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  AOI211_X1 U11238 ( .C1(n10359), .C2(n10358), .A(n10357), .B(n10356), .ZN(
        n10362) );
  XOR2_X1 U11239 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .Z(n10361) );
  XOR2_X1 U11240 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_117), .Z(n10360) );
  OAI22_X1 U11241 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_120), .B1(
        keyinput_121), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n10363) );
  AOI221_X1 U11242 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_120), .C1(
        P1_IR_REG_30__SCAN_IN), .C2(keyinput_121), .A(n10363), .ZN(n10370) );
  INV_X1 U11243 ( .A(keyinput_118), .ZN(n10364) );
  XNOR2_X1 U11244 ( .A(n10364), .B(P1_IR_REG_27__SCAN_IN), .ZN(n10366) );
  XNOR2_X1 U11245 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_119), .ZN(n10365)
         );
  AND2_X1 U11246 ( .A1(n10366), .A2(n10365), .ZN(n10369) );
  XNOR2_X1 U11247 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_123), .ZN(n10368) );
  XNOR2_X1 U11248 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .ZN(n10367)
         );
  NAND4_X1 U11249 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n10374) );
  OAI22_X1 U11250 ( .A1(n10372), .A2(keyinput_125), .B1(P1_D_REG_1__SCAN_IN), 
        .B2(keyinput_124), .ZN(n10371) );
  AOI221_X1 U11251 ( .B1(n10372), .B2(keyinput_125), .C1(keyinput_124), .C2(
        P1_D_REG_1__SCAN_IN), .A(n10371), .ZN(n10373) );
  OAI21_X1 U11252 ( .B1(n10375), .B2(n10374), .A(n10373), .ZN(n10603) );
  AOI22_X1 U11253 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_253), .B1(n6430), 
        .B2(keyinput_252), .ZN(n10376) );
  OAI221_X1 U11254 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_253), .C1(n6430), 
        .C2(keyinput_252), .A(n10376), .ZN(n10595) );
  AOI22_X1 U11255 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_240), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_239), .ZN(n10377) );
  OAI221_X1 U11256 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_240), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_239), .A(n10377), .ZN(n10580) );
  INV_X1 U11257 ( .A(keyinput_215), .ZN(n10534) );
  INV_X1 U11258 ( .A(keyinput_213), .ZN(n10526) );
  OAI22_X1 U11259 ( .A1(n5753), .A2(keyinput_198), .B1(n10379), .B2(
        keyinput_196), .ZN(n10378) );
  AOI221_X1 U11260 ( .B1(n5753), .B2(keyinput_198), .C1(keyinput_196), .C2(
        n10379), .A(n10378), .ZN(n10388) );
  OAI22_X1 U11261 ( .A1(n10382), .A2(keyinput_200), .B1(n10381), .B2(
        keyinput_195), .ZN(n10380) );
  AOI221_X1 U11262 ( .B1(n10382), .B2(keyinput_200), .C1(keyinput_195), .C2(
        n10381), .A(n10380), .ZN(n10387) );
  OAI22_X1 U11263 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_201), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_202), .ZN(n10383) );
  AOI221_X1 U11264 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_201), .C1(
        keyinput_202), .C2(P2_DATAO_REG_22__SCAN_IN), .A(n10383), .ZN(n10386)
         );
  OAI22_X1 U11265 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_197), .B1(
        keyinput_199), .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10384) );
  AOI221_X1 U11266 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_197), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_199), .A(n10384), .ZN(n10385)
         );
  NAND4_X1 U11267 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10508) );
  INV_X1 U11268 ( .A(keyinput_194), .ZN(n10504) );
  INV_X1 U11269 ( .A(keyinput_193), .ZN(n10503) );
  INV_X1 U11270 ( .A(keyinput_192), .ZN(n10501) );
  INV_X1 U11271 ( .A(keyinput_180), .ZN(n10482) );
  INV_X1 U11272 ( .A(keyinput_179), .ZN(n10481) );
  XNOR2_X1 U11273 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n10479)
         );
  INV_X1 U11274 ( .A(keyinput_173), .ZN(n10470) );
  INV_X1 U11275 ( .A(keyinput_168), .ZN(n10457) );
  INV_X1 U11276 ( .A(keyinput_166), .ZN(n10453) );
  INV_X1 U11277 ( .A(keyinput_159), .ZN(n10435) );
  OAI22_X1 U11278 ( .A1(SI_11_), .A2(keyinput_149), .B1(keyinput_150), .B2(
        SI_10_), .ZN(n10389) );
  AOI221_X1 U11279 ( .B1(SI_11_), .B2(keyinput_149), .C1(SI_10_), .C2(
        keyinput_150), .A(n10389), .ZN(n10422) );
  OAI22_X1 U11280 ( .A1(n10391), .A2(keyinput_148), .B1(keyinput_145), .B2(
        SI_15_), .ZN(n10390) );
  AOI221_X1 U11281 ( .B1(n10391), .B2(keyinput_148), .C1(SI_15_), .C2(
        keyinput_145), .A(n10390), .ZN(n10421) );
  OAI22_X1 U11282 ( .A1(SI_14_), .A2(keyinput_146), .B1(keyinput_147), .B2(
        SI_13_), .ZN(n10392) );
  AOI221_X1 U11283 ( .B1(SI_14_), .B2(keyinput_146), .C1(SI_13_), .C2(
        keyinput_147), .A(n10392), .ZN(n10420) );
  AOI22_X1 U11284 ( .A1(n10395), .A2(keyinput_135), .B1(n10394), .B2(
        keyinput_134), .ZN(n10393) );
  OAI221_X1 U11285 ( .B1(n10395), .B2(keyinput_135), .C1(n10394), .C2(
        keyinput_134), .A(n10393), .ZN(n10412) );
  OAI22_X1 U11286 ( .A1(SI_24_), .A2(keyinput_136), .B1(SI_28_), .B2(
        keyinput_132), .ZN(n10396) );
  AOI221_X1 U11287 ( .B1(SI_24_), .B2(keyinput_136), .C1(keyinput_132), .C2(
        SI_28_), .A(n10396), .ZN(n10405) );
  OAI22_X1 U11288 ( .A1(SI_27_), .A2(keyinput_133), .B1(SI_29_), .B2(
        keyinput_131), .ZN(n10397) );
  INV_X1 U11289 ( .A(keyinput_130), .ZN(n10400) );
  OAI22_X1 U11290 ( .A1(SI_31_), .A2(keyinput_129), .B1(keyinput_128), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n10398) );
  AOI221_X1 U11291 ( .B1(SI_31_), .B2(keyinput_129), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_128), .A(n10398), .ZN(n10399) );
  OAI221_X1 U11292 ( .B1(SI_30_), .B2(keyinput_130), .C1(n10401), .C2(n10400), 
        .A(n10399), .ZN(n10403) );
  XNOR2_X1 U11293 ( .A(SI_23_), .B(keyinput_137), .ZN(n10402) );
  NAND4_X1 U11294 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10411) );
  OAI22_X1 U11295 ( .A1(n10407), .A2(keyinput_139), .B1(keyinput_138), .B2(
        SI_22_), .ZN(n10406) );
  AOI221_X1 U11296 ( .B1(n10407), .B2(keyinput_139), .C1(SI_22_), .C2(
        keyinput_138), .A(n10406), .ZN(n10410) );
  OAI22_X1 U11297 ( .A1(SI_20_), .A2(keyinput_140), .B1(SI_19_), .B2(
        keyinput_141), .ZN(n10408) );
  AOI221_X1 U11298 ( .B1(SI_20_), .B2(keyinput_140), .C1(keyinput_141), .C2(
        SI_19_), .A(n10408), .ZN(n10409) );
  OAI211_X1 U11299 ( .C1(n10412), .C2(n10411), .A(n10410), .B(n10409), .ZN(
        n10416) );
  OAI22_X1 U11300 ( .A1(n10414), .A2(keyinput_142), .B1(keyinput_143), .B2(
        SI_17_), .ZN(n10413) );
  AOI221_X1 U11301 ( .B1(n10414), .B2(keyinput_142), .C1(SI_17_), .C2(
        keyinput_143), .A(n10413), .ZN(n10415) );
  NAND2_X1 U11302 ( .A1(n10416), .A2(n10415), .ZN(n10419) );
  AOI22_X1 U11303 ( .A1(SI_7_), .A2(keyinput_153), .B1(SI_8_), .B2(
        keyinput_152), .ZN(n10423) );
  OAI221_X1 U11304 ( .B1(SI_7_), .B2(keyinput_153), .C1(SI_8_), .C2(
        keyinput_152), .A(n10423), .ZN(n10424) );
  AOI22_X1 U11305 ( .A1(SI_5_), .A2(keyinput_155), .B1(n10427), .B2(
        keyinput_154), .ZN(n10426) );
  OAI221_X1 U11306 ( .B1(SI_5_), .B2(keyinput_155), .C1(n10427), .C2(
        keyinput_154), .A(n10426), .ZN(n10432) );
  OAI22_X1 U11307 ( .A1(n10429), .A2(keyinput_156), .B1(SI_3_), .B2(
        keyinput_157), .ZN(n10428) );
  AOI221_X1 U11308 ( .B1(n10429), .B2(keyinput_156), .C1(keyinput_157), .C2(
        SI_3_), .A(n10428), .ZN(n10431) );
  XNOR2_X1 U11309 ( .A(SI_2_), .B(keyinput_158), .ZN(n10430) );
  OAI211_X1 U11310 ( .C1(n10433), .C2(n10432), .A(n10431), .B(n10430), .ZN(
        n10434) );
  OAI221_X1 U11311 ( .B1(SI_1_), .B2(keyinput_159), .C1(n10436), .C2(n10435), 
        .A(n10434), .ZN(n10440) );
  OAI22_X1 U11312 ( .A1(n10438), .A2(keyinput_160), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_161), .ZN(n10437) );
  AOI221_X1 U11313 ( .B1(n10438), .B2(keyinput_160), .C1(keyinput_161), .C2(
        P2_RD_REG_SCAN_IN), .A(n10437), .ZN(n10439) );
  OAI22_X1 U11314 ( .A1(n10445), .A2(keyinput_163), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_164), .ZN(n10444) );
  AOI221_X1 U11315 ( .B1(n10445), .B2(keyinput_163), .C1(keyinput_164), .C2(
        P2_REG3_REG_27__SCAN_IN), .A(n10444), .ZN(n10446) );
  NAND2_X1 U11316 ( .A1(n10447), .A2(n10446), .ZN(n10451) );
  INV_X1 U11317 ( .A(keyinput_167), .ZN(n10454) );
  INV_X1 U11318 ( .A(keyinput_169), .ZN(n10459) );
  NAND2_X1 U11319 ( .A1(n10462), .A2(n10461), .ZN(n10465) );
  OAI22_X1 U11320 ( .A1(n6366), .A2(keyinput_170), .B1(keyinput_171), .B2(
        P2_REG3_REG_8__SCAN_IN), .ZN(n10463) );
  AOI221_X1 U11321 ( .B1(n6366), .B2(keyinput_170), .C1(P2_REG3_REG_8__SCAN_IN), .C2(keyinput_171), .A(n10463), .ZN(n10464) );
  NAND2_X1 U11322 ( .A1(n10468), .A2(n10467), .ZN(n10469) );
  OAI221_X1 U11323 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_173), .C1(
        n10471), .C2(n10470), .A(n10469), .ZN(n10478) );
  AOI22_X1 U11324 ( .A1(n10474), .A2(keyinput_176), .B1(n10473), .B2(
        keyinput_177), .ZN(n10472) );
  OAI221_X1 U11325 ( .B1(n10474), .B2(keyinput_176), .C1(n10473), .C2(
        keyinput_177), .A(n10472), .ZN(n10477) );
  AOI22_X1 U11326 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_175), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_178), .ZN(n10475) );
  OAI221_X1 U11327 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_175), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_178), .A(n10475), .ZN(n10476)
         );
  OAI22_X1 U11328 ( .A1(n10485), .A2(keyinput_182), .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_181), .ZN(n10484) );
  AOI221_X1 U11329 ( .B1(n10485), .B2(keyinput_182), .C1(keyinput_181), .C2(
        P2_REG3_REG_9__SCAN_IN), .A(n10484), .ZN(n10486) );
  OAI21_X1 U11330 ( .B1(keyinput_183), .B2(n10488), .A(n10486), .ZN(n10487) );
  AOI22_X1 U11331 ( .A1(n10490), .A2(keyinput_185), .B1(n6045), .B2(
        keyinput_184), .ZN(n10489) );
  OAI221_X1 U11332 ( .B1(n10490), .B2(keyinput_185), .C1(n6045), .C2(
        keyinput_184), .A(n10489), .ZN(n10494) );
  OAI22_X1 U11333 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_186), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput_187), .ZN(n10491) );
  AOI221_X1 U11334 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_186), .C1(
        keyinput_187), .C2(P2_REG3_REG_2__SCAN_IN), .A(n10491), .ZN(n10493) );
  XNOR2_X1 U11335 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n10492)
         );
  OAI211_X1 U11336 ( .C1(n5091), .C2(n10494), .A(n10493), .B(n10492), .ZN(
        n10499) );
  OAI22_X1 U11337 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_191), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_190), .ZN(n10495) );
  AOI221_X1 U11338 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_191), .C1(
        keyinput_190), .C2(P2_REG3_REG_26__SCAN_IN), .A(n10495), .ZN(n10498)
         );
  NAND2_X1 U11339 ( .A1(keyinput_205), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(
        n10506) );
  OAI221_X1 U11340 ( .B1(n10508), .B2(n10507), .C1(keyinput_205), .C2(
        P2_DATAO_REG_19__SCAN_IN), .A(n10506), .ZN(n10514) );
  AOI22_X1 U11341 ( .A1(n10511), .A2(keyinput_204), .B1(n10510), .B2(
        keyinput_203), .ZN(n10509) );
  OAI221_X1 U11342 ( .B1(n10511), .B2(keyinput_204), .C1(n10510), .C2(
        keyinput_203), .A(n10509), .ZN(n10513) );
  NAND2_X1 U11343 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_206), .ZN(
        n10512) );
  OAI221_X1 U11344 ( .B1(n10514), .B2(n10513), .C1(P2_DATAO_REG_18__SCAN_IN), 
        .C2(keyinput_206), .A(n10512), .ZN(n10520) );
  OAI22_X1 U11345 ( .A1(n10517), .A2(keyinput_207), .B1(n10516), .B2(
        keyinput_208), .ZN(n10515) );
  AOI221_X1 U11346 ( .B1(n10517), .B2(keyinput_207), .C1(keyinput_208), .C2(
        n10516), .A(n10515), .ZN(n10519) );
  NOR2_X1 U11347 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_209), .ZN(
        n10518) );
  AOI22_X1 U11348 ( .A1(n10523), .A2(keyinput_211), .B1(n10522), .B2(
        keyinput_210), .ZN(n10521) );
  OAI221_X1 U11349 ( .B1(n10523), .B2(keyinput_211), .C1(n10522), .C2(
        keyinput_210), .A(n10521), .ZN(n10524) );
  INV_X1 U11350 ( .A(keyinput_214), .ZN(n10529) );
  NAND2_X1 U11351 ( .A1(n10532), .A2(n10531), .ZN(n10533) );
  OAI221_X1 U11352 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_215), .C1(
        n10535), .C2(n10534), .A(n10533), .ZN(n10538) );
  OAI22_X1 U11353 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_216), .B1(
        keyinput_217), .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n10536) );
  AOI221_X1 U11354 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_216), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_217), .A(n10536), .ZN(n10537)
         );
  NAND2_X1 U11355 ( .A1(n10538), .A2(n10537), .ZN(n10550) );
  OAI22_X1 U11356 ( .A1(n10540), .A2(keyinput_221), .B1(keyinput_220), .B2(
        P1_IR_REG_1__SCAN_IN), .ZN(n10539) );
  AOI221_X1 U11357 ( .B1(n10540), .B2(keyinput_221), .C1(P1_IR_REG_1__SCAN_IN), 
        .C2(keyinput_220), .A(n10539), .ZN(n10541) );
  INV_X1 U11358 ( .A(n10541), .ZN(n10548) );
  XOR2_X1 U11359 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_222), .Z(n10547) );
  AOI22_X1 U11360 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_219), .B1(n10543), 
        .B2(keyinput_218), .ZN(n10542) );
  OAI221_X1 U11361 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_219), .C1(n10543), 
        .C2(keyinput_218), .A(n10542), .ZN(n10546) );
  XNOR2_X1 U11362 ( .A(n10544), .B(keyinput_223), .ZN(n10545) );
  NOR4_X1 U11363 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n10549) );
  INV_X1 U11364 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U11365 ( .A1(n10553), .A2(keyinput_226), .B1(keyinput_229), .B2(
        n10552), .ZN(n10551) );
  OAI221_X1 U11366 ( .B1(n10553), .B2(keyinput_226), .C1(n10552), .C2(
        keyinput_229), .A(n10551), .ZN(n10559) );
  XNOR2_X1 U11367 ( .A(n6457), .B(keyinput_225), .ZN(n10557) );
  XNOR2_X1 U11368 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_228), .ZN(n10556) );
  XNOR2_X1 U11369 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_227), .ZN(n10555) );
  XNOR2_X1 U11370 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_224), .ZN(n10554) );
  NAND4_X1 U11371 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n10558) );
  NOR2_X1 U11372 ( .A1(n10559), .A2(n10558), .ZN(n10562) );
  XOR2_X1 U11373 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_230), .Z(n10561) );
  XNOR2_X1 U11374 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_231), .ZN(n10560)
         );
  AOI22_X1 U11375 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_233), .B1(n6874), 
        .B2(keyinput_232), .ZN(n10563) );
  OAI221_X1 U11376 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_233), .C1(n6874), 
        .C2(keyinput_232), .A(n10563), .ZN(n10564) );
  INV_X1 U11377 ( .A(keyinput_235), .ZN(n10566) );
  INV_X1 U11378 ( .A(n10567), .ZN(n10577) );
  INV_X1 U11379 ( .A(keyinput_236), .ZN(n10570) );
  XNOR2_X1 U11380 ( .A(n10568), .B(keyinput_238), .ZN(n10569) );
  AOI21_X1 U11381 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(n10570), .A(n10569), .ZN(
        n10575) );
  XNOR2_X1 U11382 ( .A(n10571), .B(keyinput_237), .ZN(n10574) );
  NAND3_X1 U11383 ( .A1(n10575), .A2(n10574), .A3(n10573), .ZN(n10576) );
  OAI22_X1 U11384 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_241), .B1(
        keyinput_242), .B2(P1_IR_REG_23__SCAN_IN), .ZN(n10581) );
  AOI221_X1 U11385 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_241), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_242), .A(n10581), .ZN(n10582) );
  XOR2_X1 U11386 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_244), .Z(n10584) );
  XOR2_X1 U11387 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_245), .Z(n10583) );
  NOR2_X1 U11388 ( .A1(n10584), .A2(n10583), .ZN(n10592) );
  AOI22_X1 U11389 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_249), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput_248), .ZN(n10585) );
  OAI221_X1 U11390 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_249), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput_248), .A(n10585), .ZN(n10591) );
  XNOR2_X1 U11391 ( .A(n10668), .B(keyinput_251), .ZN(n10589) );
  XNOR2_X1 U11392 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n10588)
         );
  XNOR2_X1 U11393 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_246), .ZN(n10587)
         );
  XNOR2_X1 U11394 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_250), .ZN(n10586)
         );
  NAND4_X1 U11395 ( .A1(n10589), .A2(n10588), .A3(n10587), .A4(n10586), .ZN(
        n10590) );
  NAND2_X1 U11396 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_254), .ZN(n10593)
         );
  OAI221_X1 U11397 ( .B1(n10595), .B2(n10594), .C1(P1_D_REG_3__SCAN_IN), .C2(
        keyinput_254), .A(n10593), .ZN(n10597) );
  AOI21_X1 U11398 ( .B1(n10597), .B2(keyinput_255), .A(keyinput_127), .ZN(
        n10601) );
  INV_X1 U11399 ( .A(keyinput_255), .ZN(n10596) );
  NAND2_X1 U11400 ( .A1(n10597), .A2(n10596), .ZN(n10600) );
  INV_X1 U11401 ( .A(keyinput_127), .ZN(n10598) );
  AOI22_X1 U11402 ( .A1(n10601), .A2(P1_D_REG_4__SCAN_IN), .B1(n10600), .B2(
        n10599), .ZN(n10602) );
  AOI21_X1 U11403 ( .B1(n10604), .B2(n10603), .A(n10602), .ZN(n10629) );
  INV_X1 U11404 ( .A(n7021), .ZN(n10609) );
  NOR3_X1 U11405 ( .A1(n10607), .A2(n10606), .A3(n10605), .ZN(n10608) );
  AOI21_X1 U11406 ( .B1(n10609), .B2(n10623), .A(n10608), .ZN(n10627) );
  AOI22_X1 U11407 ( .A1(n10613), .A2(n10612), .B1(n10611), .B2(n10610), .ZN(
        n10621) );
  INV_X1 U11408 ( .A(n10614), .ZN(n10615) );
  NAND2_X1 U11409 ( .A1(n10616), .A2(n10615), .ZN(n10620) );
  NAND2_X1 U11410 ( .A1(n9691), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10619) );
  NAND2_X1 U11411 ( .A1(n10617), .A2(n7347), .ZN(n10618) );
  NAND4_X1 U11412 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10622) );
  AOI21_X1 U11413 ( .B1(n10624), .B2(n10623), .A(n10622), .ZN(n10625) );
  OAI21_X1 U11414 ( .B1(n10627), .B2(n10626), .A(n10625), .ZN(n10628) );
  XOR2_X1 U11415 ( .A(n10629), .B(n10628), .Z(P2_U3232) );
  XOR2_X1 U11416 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11417 ( .A(n10630), .ZN(n10631) );
  NAND2_X1 U11418 ( .A1(n10632), .A2(n10631), .ZN(n10633) );
  XOR2_X1 U11419 ( .A(n10771), .B(n10633), .Z(ADD_1071_U5) );
  XOR2_X1 U11420 ( .A(n10635), .B(n10634), .Z(ADD_1071_U54) );
  XOR2_X1 U11421 ( .A(n10637), .B(n10636), .Z(ADD_1071_U53) );
  XNOR2_X1 U11422 ( .A(n10639), .B(n10638), .ZN(ADD_1071_U52) );
  NOR2_X1 U11423 ( .A1(n10641), .A2(n10640), .ZN(n10642) );
  XOR2_X1 U11424 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10642), .Z(ADD_1071_U51) );
  XOR2_X1 U11425 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10643), .Z(ADD_1071_U50) );
  XOR2_X1 U11426 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10644), .Z(ADD_1071_U49) );
  XOR2_X1 U11427 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10645), .Z(ADD_1071_U48) );
  XOR2_X1 U11428 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10646), .Z(ADD_1071_U47) );
  XOR2_X1 U11429 ( .A(n10648), .B(n10647), .Z(ADD_1071_U63) );
  XOR2_X1 U11430 ( .A(n10650), .B(n10649), .Z(ADD_1071_U62) );
  XNOR2_X1 U11431 ( .A(n10652), .B(n10651), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11432 ( .A(n10654), .B(n10653), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11433 ( .A(n10656), .B(n10655), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11434 ( .A(n10658), .B(n10657), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11435 ( .A(n10660), .B(n10659), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11436 ( .A(n10662), .B(n10661), .ZN(ADD_1071_U56) );
  NOR2_X1 U11437 ( .A1(n10664), .A2(n10663), .ZN(n10665) );
  XOR2_X1 U11438 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10665), .Z(ADD_1071_U55)
         );
  NAND2_X1 U11439 ( .A1(n10666), .A2(n10669), .ZN(n10667) );
  OAI21_X1 U11440 ( .B1(n10669), .B2(n10668), .A(n10667), .ZN(P1_U3440) );
  OAI211_X1 U11441 ( .C1(n10670), .C2(n10674), .A(P1_STATE_REG_SCAN_IN), .B(
        n6681), .ZN(n10672) );
  OAI22_X1 U11442 ( .A1(n10702), .A2(P1_REG1_REG_0__SCAN_IN), .B1(n10672), 
        .B2(n10671), .ZN(n10677) );
  NAND3_X1 U11443 ( .A1(n10675), .A2(n10674), .A3(n10673), .ZN(n10676) );
  NAND2_X1 U11444 ( .A1(n10677), .A2(n10676), .ZN(n10680) );
  AOI22_X1 U11445 ( .A1(n10813), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10679) );
  OAI21_X1 U11446 ( .B1(n10681), .B2(n10680), .A(n10679), .ZN(P1_U3241) );
  AOI22_X1 U11447 ( .A1(n10813), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10744), 
        .B2(n10682), .ZN(n10692) );
  OAI211_X1 U11448 ( .C1(n10685), .C2(n10684), .A(n10683), .B(n10746), .ZN(
        n10690) );
  OAI211_X1 U11449 ( .C1(n10688), .C2(n10687), .A(n10686), .B(n10815), .ZN(
        n10689) );
  NAND4_X1 U11450 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        P1_U3247) );
  NOR2_X1 U11451 ( .A1(n10693), .A2(n10710), .ZN(n10699) );
  INV_X1 U11452 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10696) );
  INV_X1 U11453 ( .A(n10694), .ZN(n10695) );
  OAI21_X1 U11454 ( .B1(n10697), .B2(n10696), .A(n10695), .ZN(n10698) );
  AOI21_X1 U11455 ( .B1(n10700), .B2(n10699), .A(n10698), .ZN(n10716) );
  INV_X1 U11456 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10701) );
  NOR3_X1 U11457 ( .A1(n10702), .A2(n10701), .A3(n10709), .ZN(n10704) );
  OAI21_X1 U11458 ( .B1(n10704), .B2(n10744), .A(n10703), .ZN(n10715) );
  INV_X1 U11459 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U11460 ( .A1(n10710), .A2(n10705), .ZN(n10707) );
  OAI211_X1 U11461 ( .C1(n10708), .C2(n10707), .A(n10706), .B(n10746), .ZN(
        n10714) );
  NAND3_X1 U11462 ( .A1(n10710), .A2(n10701), .A3(n10709), .ZN(n10711) );
  NAND3_X1 U11463 ( .A1(n10815), .A2(n10712), .A3(n10711), .ZN(n10713) );
  NAND4_X1 U11464 ( .A1(n10716), .A2(n10715), .A3(n10714), .A4(n10713), .ZN(
        P1_U3252) );
  OAI21_X1 U11465 ( .B1(n10719), .B2(n10718), .A(n10717), .ZN(n10720) );
  AOI22_X1 U11466 ( .A1(n10720), .A2(n10815), .B1(n10813), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n10730) );
  AOI21_X1 U11467 ( .B1(n10723), .B2(n10722), .A(n10721), .ZN(n10724) );
  NAND2_X1 U11468 ( .A1(n10746), .A2(n10724), .ZN(n10726) );
  OAI211_X1 U11469 ( .C1(n10727), .C2(n10809), .A(n10726), .B(n10725), .ZN(
        n10728) );
  INV_X1 U11470 ( .A(n10728), .ZN(n10729) );
  NAND2_X1 U11471 ( .A1(n10730), .A2(n10729), .ZN(P1_U3259) );
  AOI22_X1 U11472 ( .A1(n10813), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n10744), 
        .B2(n10731), .ZN(n10742) );
  AOI21_X1 U11473 ( .B1(n10734), .B2(n10733), .A(n10732), .ZN(n10735) );
  OR2_X1 U11474 ( .A1(n10735), .A2(n10808), .ZN(n10740) );
  OAI211_X1 U11475 ( .C1(n10738), .C2(n10737), .A(n10736), .B(n10815), .ZN(
        n10739) );
  NAND4_X1 U11476 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        P1_U3246) );
  AOI22_X1 U11477 ( .A1(n10813), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(n10744), 
        .B2(n10743), .ZN(n10755) );
  OAI211_X1 U11478 ( .C1(n10748), .C2(n10747), .A(n10746), .B(n10745), .ZN(
        n10753) );
  OAI211_X1 U11479 ( .C1(n10751), .C2(n10750), .A(n10815), .B(n10749), .ZN(
        n10752) );
  NAND4_X1 U11480 ( .A1(n10755), .A2(n10754), .A3(n10753), .A4(n10752), .ZN(
        P1_U3244) );
  INV_X1 U11481 ( .A(n10756), .ZN(n10759) );
  AOI22_X1 U11482 ( .A1(n10760), .A2(n10759), .B1(n10758), .B2(n10757), .ZN(
        P2_U3437) );
  AOI22_X1 U11483 ( .A1(n10761), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10796), .ZN(n10769) );
  NAND2_X1 U11484 ( .A1(n10796), .A2(n10762), .ZN(n10764) );
  OAI211_X1 U11485 ( .C1(n10788), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10764), .B(
        n10763), .ZN(n10765) );
  INV_X1 U11486 ( .A(n10765), .ZN(n10768) );
  AOI21_X1 U11487 ( .B1(n10787), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n10766), .ZN(
        n10767) );
  OAI221_X1 U11488 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10769), .C1(n10779), .C2(
        n10768), .A(n10767), .ZN(P2_U3245) );
  OAI22_X1 U11489 ( .A1(n10772), .A2(n10771), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10770), .ZN(n10777) );
  NAND2_X1 U11490 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10775) );
  AOI211_X1 U11491 ( .C1(n10775), .C2(n10774), .A(n10773), .B(n10788), .ZN(
        n10776) );
  AOI211_X1 U11492 ( .C1(n10794), .C2(n10778), .A(n10777), .B(n10776), .ZN(
        n10784) );
  NOR2_X1 U11493 ( .A1(n10779), .A2(n10762), .ZN(n10782) );
  OAI211_X1 U11494 ( .C1(n10782), .C2(n10781), .A(n10796), .B(n10780), .ZN(
        n10783) );
  NAND2_X1 U11495 ( .A1(n10784), .A2(n10783), .ZN(P2_U3246) );
  INV_X1 U11496 ( .A(n10785), .ZN(n10786) );
  AOI21_X1 U11497 ( .B1(n10787), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n10786), .ZN(
        n10801) );
  AOI211_X1 U11498 ( .C1(n10791), .C2(n10790), .A(n10789), .B(n10788), .ZN(
        n10792) );
  AOI21_X1 U11499 ( .B1(n10794), .B2(n10793), .A(n10792), .ZN(n10800) );
  OAI211_X1 U11500 ( .C1(n10798), .C2(n10797), .A(n10796), .B(n10795), .ZN(
        n10799) );
  NAND3_X1 U11501 ( .A1(n10801), .A2(n10800), .A3(n10799), .ZN(P2_U3247) );
  XNOR2_X1 U11502 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U11503 ( .A(n6533), .B(P1_REG2_REG_2__SCAN_IN), .S(n10802), .Z(
        n10803) );
  NAND2_X1 U11504 ( .A1(n10804), .A2(n10803), .ZN(n10806) );
  NAND2_X1 U11505 ( .A1(n10806), .A2(n10805), .ZN(n10807) );
  OAI22_X1 U11506 ( .A1(n10810), .A2(n10809), .B1(n10808), .B2(n10807), .ZN(
        n10812) );
  AOI211_X1 U11507 ( .C1(n10813), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n10812), .B(
        n10811), .ZN(n10819) );
  OAI211_X1 U11508 ( .C1(n10817), .C2(n10816), .A(n10815), .B(n10814), .ZN(
        n10818) );
  OAI211_X1 U11509 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n10820), .A(n10819), .B(
        n10818), .ZN(P1_U3243) );
  INV_X1 U11510 ( .A(n10821), .ZN(n10827) );
  NOR2_X1 U11511 ( .A1(n10821), .A2(n11057), .ZN(n10826) );
  OAI211_X1 U11512 ( .C1(n10824), .C2(n11109), .A(n10823), .B(n10822), .ZN(
        n10825) );
  AOI211_X1 U11513 ( .C1(n10827), .C2(n11062), .A(n10826), .B(n10825), .ZN(
        n10829) );
  AOI22_X1 U11514 ( .A1(n10900), .A2(n10829), .B1(n6554), .B2(n11118), .ZN(
        P1_U3524) );
  INV_X1 U11515 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U11516 ( .A1(n10137), .A2(n10829), .B1(n10828), .B2(n11120), .ZN(
        P1_U3457) );
  INV_X1 U11517 ( .A(n10830), .ZN(n10838) );
  INV_X1 U11518 ( .A(n10831), .ZN(n10833) );
  NAND3_X1 U11519 ( .A1(n10833), .A2(n11067), .A3(n10832), .ZN(n10834) );
  OAI211_X1 U11520 ( .C1(n10836), .C2(n11123), .A(n10835), .B(n10834), .ZN(
        n10837) );
  AOI21_X1 U11521 ( .B1(n11129), .B2(n10838), .A(n10837), .ZN(n10840) );
  AOI22_X1 U11522 ( .A1(n11132), .A2(n10840), .B1(n6738), .B2(n11131), .ZN(
        P2_U3521) );
  INV_X1 U11523 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U11524 ( .A1(n11135), .A2(n10840), .B1(n10839), .B2(n5340), .ZN(
        P2_U3454) );
  INV_X1 U11525 ( .A(n11057), .ZN(n11114) );
  INV_X1 U11526 ( .A(n10841), .ZN(n10846) );
  OAI22_X1 U11527 ( .A1(n10843), .A2(n11111), .B1(n10842), .B2(n11109), .ZN(
        n10845) );
  AOI211_X1 U11528 ( .C1(n11114), .C2(n10846), .A(n10845), .B(n10844), .ZN(
        n10849) );
  AOI22_X1 U11529 ( .A1(n10847), .A2(n10849), .B1(n6555), .B2(n11118), .ZN(
        P1_U3525) );
  INV_X1 U11530 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U11531 ( .A1(n10137), .A2(n10849), .B1(n10848), .B2(n11120), .ZN(
        P1_U3460) );
  INV_X1 U11532 ( .A(n10850), .ZN(n11036) );
  INV_X1 U11533 ( .A(n10851), .ZN(n10856) );
  OAI22_X1 U11534 ( .A1(n10853), .A2(n11125), .B1(n10852), .B2(n11123), .ZN(
        n10855) );
  AOI211_X1 U11535 ( .C1(n11036), .C2(n10856), .A(n10855), .B(n10854), .ZN(
        n10858) );
  AOI22_X1 U11536 ( .A1(n11132), .A2(n10858), .B1(n6737), .B2(n11131), .ZN(
        P2_U3522) );
  INV_X1 U11537 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U11538 ( .A1(n11135), .A2(n10858), .B1(n10857), .B2(n5340), .ZN(
        P2_U3457) );
  XNOR2_X1 U11539 ( .A(n10860), .B(n10859), .ZN(n10866) );
  XNOR2_X1 U11540 ( .A(n10861), .B(n10860), .ZN(n10877) );
  NAND2_X1 U11541 ( .A1(n10877), .A2(n11062), .ZN(n10865) );
  AOI22_X1 U11542 ( .A1(n10993), .A2(n10863), .B1(n10862), .B2(n10990), .ZN(
        n10864) );
  OAI211_X1 U11543 ( .C1(n10867), .C2(n10866), .A(n10865), .B(n10864), .ZN(
        n10878) );
  AND2_X1 U11544 ( .A1(n10877), .A2(n11114), .ZN(n10872) );
  OR2_X1 U11545 ( .A1(n10868), .A2(n10880), .ZN(n10869) );
  NAND2_X1 U11546 ( .A1(n10870), .A2(n10869), .ZN(n10875) );
  OAI22_X1 U11547 ( .A1(n10875), .A2(n11111), .B1(n10880), .B2(n11109), .ZN(
        n10871) );
  NOR3_X1 U11548 ( .A1(n10878), .A2(n10872), .A3(n10871), .ZN(n10874) );
  AOI22_X1 U11549 ( .A1(n10900), .A2(n10874), .B1(n6551), .B2(n11118), .ZN(
        P1_U3526) );
  INV_X1 U11550 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U11551 ( .A1(n10137), .A2(n10874), .B1(n10873), .B2(n11120), .ZN(
        P1_U3463) );
  INV_X1 U11552 ( .A(n10875), .ZN(n10876) );
  AOI22_X1 U11553 ( .A1(n10877), .A2(n11010), .B1(n11009), .B2(n10876), .ZN(
        n10884) );
  MUX2_X1 U11554 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10878), .S(n11019), .Z(
        n10882) );
  OAI22_X1 U11555 ( .A1(n11016), .A2(n10880), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n10879), .ZN(n10881) );
  NOR2_X1 U11556 ( .A1(n10882), .A2(n10881), .ZN(n10883) );
  NAND2_X1 U11557 ( .A1(n10884), .A2(n10883), .ZN(P1_U3288) );
  INV_X1 U11558 ( .A(n10885), .ZN(n10890) );
  OAI22_X1 U11559 ( .A1(n10887), .A2(n11125), .B1(n10886), .B2(n11123), .ZN(
        n10889) );
  AOI211_X1 U11560 ( .C1(n11036), .C2(n10890), .A(n10889), .B(n10888), .ZN(
        n10892) );
  AOI22_X1 U11561 ( .A1(n11132), .A2(n10892), .B1(n6736), .B2(n11131), .ZN(
        P2_U3523) );
  INV_X1 U11562 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U11563 ( .A1(n11135), .A2(n10892), .B1(n10891), .B2(n5340), .ZN(
        P2_U3460) );
  AND2_X1 U11564 ( .A1(n10893), .A2(n11114), .ZN(n10897) );
  OAI22_X1 U11565 ( .A1(n10895), .A2(n11111), .B1(n10894), .B2(n11109), .ZN(
        n10896) );
  NOR3_X1 U11566 ( .A1(n10898), .A2(n10897), .A3(n10896), .ZN(n10902) );
  AOI22_X1 U11567 ( .A1(n10900), .A2(n10902), .B1(n10899), .B2(n11118), .ZN(
        P1_U3527) );
  INV_X1 U11568 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U11569 ( .A1(n10137), .A2(n10902), .B1(n10901), .B2(n11120), .ZN(
        P1_U3466) );
  NOR2_X1 U11570 ( .A1(n10903), .A2(n11082), .ZN(n10908) );
  OAI22_X1 U11571 ( .A1(n10905), .A2(n11125), .B1(n10904), .B2(n11123), .ZN(
        n10907) );
  AOI211_X1 U11572 ( .C1(n10908), .C2(n7469), .A(n10907), .B(n10906), .ZN(
        n10910) );
  AOI22_X1 U11573 ( .A1(n11132), .A2(n10910), .B1(n6734), .B2(n11131), .ZN(
        P2_U3524) );
  INV_X1 U11574 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U11575 ( .A1(n11135), .A2(n10910), .B1(n10909), .B2(n5340), .ZN(
        P2_U3463) );
  INV_X1 U11576 ( .A(n10911), .ZN(n11091) );
  OAI21_X1 U11577 ( .B1(n10913), .B2(n11109), .A(n10912), .ZN(n10915) );
  AOI211_X1 U11578 ( .C1(n10916), .C2(n11091), .A(n10915), .B(n10914), .ZN(
        n10918) );
  AOI22_X1 U11579 ( .A1(n10900), .A2(n10918), .B1(n6560), .B2(n11118), .ZN(
        P1_U3528) );
  INV_X1 U11580 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U11581 ( .A1(n10137), .A2(n10918), .B1(n10917), .B2(n11120), .ZN(
        P1_U3469) );
  INV_X1 U11582 ( .A(n10919), .ZN(n10920) );
  NOR2_X1 U11583 ( .A1(n10921), .A2(n10920), .ZN(n10932) );
  NAND2_X1 U11584 ( .A1(n10923), .A2(n10922), .ZN(n10929) );
  AOI22_X1 U11585 ( .A1(n10927), .A2(n10926), .B1(n10925), .B2(n10924), .ZN(
        n10928) );
  NAND2_X1 U11586 ( .A1(n10929), .A2(n10928), .ZN(n10930) );
  NOR3_X1 U11587 ( .A1(n10932), .A2(n10931), .A3(n10930), .ZN(n10934) );
  AOI22_X1 U11588 ( .A1(n9566), .A2(n6719), .B1(n10934), .B2(n10933), .ZN(
        P2_U3291) );
  AOI22_X1 U11589 ( .A1(n10936), .A2(n10968), .B1(n11053), .B2(n10935), .ZN(
        n10937) );
  OAI211_X1 U11590 ( .C1(n10939), .C2(n11057), .A(n10938), .B(n10937), .ZN(
        n10940) );
  INV_X1 U11591 ( .A(n10940), .ZN(n10942) );
  AOI22_X1 U11592 ( .A1(n10900), .A2(n10942), .B1(n6550), .B2(n11118), .ZN(
        P1_U3529) );
  INV_X1 U11593 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U11594 ( .A1(n10137), .A2(n10942), .B1(n10941), .B2(n11120), .ZN(
        P1_U3472) );
  OAI22_X1 U11595 ( .A1(n10944), .A2(n11125), .B1(n10943), .B2(n11123), .ZN(
        n10946) );
  AOI211_X1 U11596 ( .C1(n11129), .C2(n10947), .A(n10946), .B(n10945), .ZN(
        n10949) );
  AOI22_X1 U11597 ( .A1(n11132), .A2(n10949), .B1(n6742), .B2(n11131), .ZN(
        P2_U3526) );
  INV_X1 U11598 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U11599 ( .A1(n11135), .A2(n10949), .B1(n10948), .B2(n5340), .ZN(
        P2_U3469) );
  OAI211_X1 U11600 ( .C1(n10952), .C2(n11109), .A(n10951), .B(n10950), .ZN(
        n10955) );
  AOI21_X1 U11601 ( .B1(n7103), .B2(n11057), .A(n10953), .ZN(n10954) );
  NOR2_X1 U11602 ( .A1(n10955), .A2(n10954), .ZN(n10958) );
  AOI22_X1 U11603 ( .A1(n10847), .A2(n10958), .B1(n10956), .B2(n11118), .ZN(
        P1_U3530) );
  INV_X1 U11604 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U11605 ( .A1(n10137), .A2(n10958), .B1(n10957), .B2(n11120), .ZN(
        P1_U3475) );
  AOI22_X1 U11606 ( .A1(n10960), .A2(n11067), .B1(n11066), .B2(n10959), .ZN(
        n10961) );
  OAI211_X1 U11607 ( .C1(n11082), .C2(n10963), .A(n10962), .B(n10961), .ZN(
        n10964) );
  INV_X1 U11608 ( .A(n10964), .ZN(n10966) );
  AOI22_X1 U11609 ( .A1(n11132), .A2(n10966), .B1(n6796), .B2(n11131), .ZN(
        P2_U3527) );
  INV_X1 U11610 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U11611 ( .A1(n11135), .A2(n10966), .B1(n10965), .B2(n5340), .ZN(
        P2_U3472) );
  AOI22_X1 U11612 ( .A1(n10969), .A2(n10968), .B1(n11053), .B2(n10967), .ZN(
        n10970) );
  OAI21_X1 U11613 ( .B1(n10971), .B2(n11057), .A(n10970), .ZN(n10972) );
  NOR2_X1 U11614 ( .A1(n10973), .A2(n10972), .ZN(n10976) );
  AOI22_X1 U11615 ( .A1(n10847), .A2(n10976), .B1(n10974), .B2(n11118), .ZN(
        P1_U3531) );
  INV_X1 U11616 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U11617 ( .A1(n10137), .A2(n10976), .B1(n10975), .B2(n11120), .ZN(
        P1_U3478) );
  NAND3_X1 U11618 ( .A1(n10978), .A2(n11129), .A3(n10977), .ZN(n10980) );
  OAI211_X1 U11619 ( .C1(n10981), .C2(n11123), .A(n10980), .B(n10979), .ZN(
        n10982) );
  INV_X1 U11620 ( .A(n10982), .ZN(n10984) );
  AOI22_X1 U11621 ( .A1(n11132), .A2(n10985), .B1(n6812), .B2(n11131), .ZN(
        P2_U3528) );
  AOI22_X1 U11622 ( .A1(n11135), .A2(n10985), .B1(n5946), .B2(n5340), .ZN(
        P2_U3475) );
  XNOR2_X1 U11623 ( .A(n10986), .B(n10995), .ZN(n11003) );
  INV_X1 U11624 ( .A(n11003), .ZN(n11011) );
  INV_X1 U11625 ( .A(n10987), .ZN(n11017) );
  INV_X1 U11626 ( .A(n10988), .ZN(n10989) );
  OAI21_X1 U11627 ( .B1(n11017), .B2(n10989), .A(n5094), .ZN(n11007) );
  OAI22_X1 U11628 ( .A1(n11007), .A2(n11111), .B1(n11017), .B2(n11109), .ZN(
        n11004) );
  AOI22_X1 U11629 ( .A1(n10993), .A2(n10992), .B1(n10991), .B2(n10990), .ZN(
        n11002) );
  INV_X1 U11630 ( .A(n10994), .ZN(n11000) );
  AND3_X1 U11631 ( .A1(n10997), .A2(n10996), .A3(n10995), .ZN(n10999) );
  OAI21_X1 U11632 ( .B1(n11000), .B2(n10999), .A(n10998), .ZN(n11001) );
  OAI211_X1 U11633 ( .C1(n11003), .C2(n7103), .A(n11002), .B(n11001), .ZN(
        n11020) );
  AOI211_X1 U11634 ( .C1(n11114), .C2(n11011), .A(n11004), .B(n11020), .ZN(
        n11006) );
  AOI22_X1 U11635 ( .A1(n10847), .A2(n11006), .B1(n6668), .B2(n11118), .ZN(
        P1_U3532) );
  INV_X1 U11636 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U11637 ( .A1(n10137), .A2(n11006), .B1(n11005), .B2(n11120), .ZN(
        P1_U3481) );
  INV_X1 U11638 ( .A(n11007), .ZN(n11008) );
  AOI22_X1 U11639 ( .A1(n11011), .A2(n11010), .B1(n11009), .B2(n11008), .ZN(
        n11022) );
  AOI22_X1 U11640 ( .A1(n11014), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11013), 
        .B2(n11012), .ZN(n11015) );
  OAI21_X1 U11641 ( .B1(n11017), .B2(n11016), .A(n11015), .ZN(n11018) );
  AOI21_X1 U11642 ( .B1(n11020), .B2(n11019), .A(n11018), .ZN(n11021) );
  NAND2_X1 U11643 ( .A1(n11022), .A2(n11021), .ZN(P1_U3282) );
  INV_X1 U11644 ( .A(n11023), .ZN(n11028) );
  OAI22_X1 U11645 ( .A1(n11025), .A2(n11125), .B1(n11024), .B2(n11123), .ZN(
        n11027) );
  AOI211_X1 U11646 ( .C1(n11036), .C2(n11028), .A(n11027), .B(n11026), .ZN(
        n11029) );
  AOI22_X1 U11647 ( .A1(n11132), .A2(n11029), .B1(n6866), .B2(n11131), .ZN(
        P2_U3529) );
  AOI22_X1 U11648 ( .A1(n11135), .A2(n11029), .B1(n5971), .B2(n5340), .ZN(
        P2_U3478) );
  INV_X1 U11649 ( .A(n11030), .ZN(n11035) );
  OAI22_X1 U11650 ( .A1(n11032), .A2(n11125), .B1(n11031), .B2(n11123), .ZN(
        n11034) );
  AOI211_X1 U11651 ( .C1(n11036), .C2(n11035), .A(n11034), .B(n11033), .ZN(
        n11037) );
  AOI22_X1 U11652 ( .A1(n11132), .A2(n11037), .B1(n6970), .B2(n11131), .ZN(
        P2_U3530) );
  AOI22_X1 U11653 ( .A1(n11135), .A2(n11037), .B1(n5991), .B2(n5340), .ZN(
        P2_U3481) );
  OAI22_X1 U11654 ( .A1(n11039), .A2(n11111), .B1(n11038), .B2(n11109), .ZN(
        n11041) );
  AOI211_X1 U11655 ( .C1(n11091), .C2(n11042), .A(n11041), .B(n11040), .ZN(
        n11044) );
  AOI22_X1 U11656 ( .A1(n10847), .A2(n11044), .B1(n10701), .B2(n11118), .ZN(
        P1_U3534) );
  INV_X1 U11657 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U11658 ( .A1(n10137), .A2(n11044), .B1(n11043), .B2(n11120), .ZN(
        P1_U3487) );
  NAND2_X1 U11659 ( .A1(n11045), .A2(n11066), .ZN(n11046) );
  AND2_X1 U11660 ( .A1(n11047), .A2(n11046), .ZN(n11050) );
  OR2_X1 U11661 ( .A1(n11048), .A2(n11082), .ZN(n11049) );
  AOI22_X1 U11662 ( .A1(n11132), .A2(n11052), .B1(n7391), .B2(n11131), .ZN(
        P2_U3531) );
  AOI22_X1 U11663 ( .A1(n11135), .A2(n11052), .B1(n6012), .B2(n5340), .ZN(
        P2_U3484) );
  INV_X1 U11664 ( .A(n11058), .ZN(n11061) );
  NAND2_X1 U11665 ( .A1(n11054), .A2(n11053), .ZN(n11055) );
  OAI211_X1 U11666 ( .C1(n11058), .C2(n11057), .A(n11056), .B(n11055), .ZN(
        n11059) );
  AOI211_X1 U11667 ( .C1(n11062), .C2(n11061), .A(n11060), .B(n11059), .ZN(
        n11064) );
  AOI22_X1 U11668 ( .A1(n10847), .A2(n11064), .B1(n6992), .B2(n11118), .ZN(
        P1_U3535) );
  INV_X1 U11669 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U11670 ( .A1(n10137), .A2(n11064), .B1(n11063), .B2(n11120), .ZN(
        P1_U3490) );
  AOI22_X1 U11671 ( .A1(n11068), .A2(n11067), .B1(n11066), .B2(n11065), .ZN(
        n11069) );
  OAI211_X1 U11672 ( .C1(n11071), .C2(n11082), .A(n11070), .B(n11069), .ZN(
        n11072) );
  INV_X1 U11673 ( .A(n11072), .ZN(n11074) );
  AOI22_X1 U11674 ( .A1(n11132), .A2(n11074), .B1(n7395), .B2(n11131), .ZN(
        P2_U3532) );
  INV_X1 U11675 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U11676 ( .A1(n11135), .A2(n11074), .B1(n11073), .B2(n5340), .ZN(
        P2_U3487) );
  OAI22_X1 U11677 ( .A1(n11076), .A2(n11111), .B1(n11075), .B2(n11109), .ZN(
        n11078) );
  AOI211_X1 U11678 ( .C1(n11114), .C2(n11079), .A(n11078), .B(n11077), .ZN(
        n11081) );
  AOI22_X1 U11679 ( .A1(n10847), .A2(n11081), .B1(n7131), .B2(n11118), .ZN(
        P1_U3536) );
  INV_X1 U11680 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U11681 ( .A1(n10137), .A2(n11081), .B1(n11080), .B2(n11120), .ZN(
        P1_U3493) );
  NOR2_X1 U11682 ( .A1(n11083), .A2(n11082), .ZN(n11088) );
  OAI22_X1 U11683 ( .A1(n11085), .A2(n11125), .B1(n11084), .B2(n11123), .ZN(
        n11087) );
  AOI211_X1 U11684 ( .C1(n11088), .C2(n8100), .A(n11087), .B(n11086), .ZN(
        n11090) );
  AOI22_X1 U11685 ( .A1(n11132), .A2(n11090), .B1(n6049), .B2(n11131), .ZN(
        P2_U3533) );
  INV_X1 U11686 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U11687 ( .A1(n11135), .A2(n11090), .B1(n11089), .B2(n5340), .ZN(
        P2_U3490) );
  NAND2_X1 U11688 ( .A1(n11092), .A2(n11091), .ZN(n11098) );
  OAI21_X1 U11689 ( .B1(n11094), .B2(n11109), .A(n11093), .ZN(n11095) );
  NOR2_X1 U11690 ( .A1(n11096), .A2(n11095), .ZN(n11097) );
  AOI22_X1 U11691 ( .A1(n10847), .A2(n11100), .B1(n7319), .B2(n11118), .ZN(
        P1_U3537) );
  INV_X1 U11692 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U11693 ( .A1(n10137), .A2(n11100), .B1(n11099), .B2(n11120), .ZN(
        P1_U3496) );
  INV_X1 U11694 ( .A(n11101), .ZN(n11102) );
  OAI22_X1 U11695 ( .A1(n11103), .A2(n11125), .B1(n11102), .B2(n11123), .ZN(
        n11104) );
  AOI211_X1 U11696 ( .C1(n11106), .C2(n11129), .A(n11105), .B(n11104), .ZN(
        n11108) );
  AOI22_X1 U11697 ( .A1(n11132), .A2(n11108), .B1(n6064), .B2(n11131), .ZN(
        P2_U3534) );
  INV_X1 U11698 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U11699 ( .A1(n11135), .A2(n11108), .B1(n11107), .B2(n5340), .ZN(
        P2_U3493) );
  OAI22_X1 U11700 ( .A1(n11112), .A2(n11111), .B1(n11110), .B2(n11109), .ZN(
        n11113) );
  AOI21_X1 U11701 ( .B1(n11115), .B2(n11114), .A(n11113), .ZN(n11116) );
  AND2_X1 U11702 ( .A1(n11117), .A2(n11116), .ZN(n11122) );
  AOI22_X1 U11703 ( .A1(n10847), .A2(n11122), .B1(n11119), .B2(n11118), .ZN(
        P1_U3538) );
  INV_X1 U11704 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11121) );
  AOI22_X1 U11705 ( .A1(n10137), .A2(n11122), .B1(n11121), .B2(n11120), .ZN(
        P1_U3499) );
  OAI22_X1 U11706 ( .A1(n11126), .A2(n11125), .B1(n11124), .B2(n11123), .ZN(
        n11128) );
  AOI211_X1 U11707 ( .C1(n11130), .C2(n11129), .A(n11128), .B(n11127), .ZN(
        n11134) );
  AOI22_X1 U11708 ( .A1(n11132), .A2(n11134), .B1(n6087), .B2(n11131), .ZN(
        P2_U3535) );
  INV_X1 U11709 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U11710 ( .A1(n11135), .A2(n11134), .B1(n11133), .B2(n5340), .ZN(
        P2_U3496) );
  XNOR2_X1 U11711 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NOR2_X1 U5111 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5773) );
  CLKBUF_X1 U5249 ( .A(n9939), .Z(n5109) );
  CLKBUF_X1 U5549 ( .A(n5024), .Z(n8541) );
endmodule

