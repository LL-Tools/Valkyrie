

module b17_C_SARLock_k_64_2 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9586, n9587, n9588, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963;

  CLKBUF_X2 U11031 ( .A(n14555), .Z(n14591) );
  OAI21_X2 U11032 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18756), .A(n16440), 
        .ZN(n17759) );
  OAI21_X1 U11033 ( .B1(n14617), .B2(n9822), .A(n9820), .ZN(n14610) );
  NAND2_X1 U11034 ( .A1(n17255), .A2(n17139), .ZN(n17230) );
  INV_X2 U11035 ( .A(n9624), .ZN(n10791) );
  XNOR2_X1 U11036 ( .A(n10146), .B(n10144), .ZN(n13520) );
  OR2_X1 U11037 ( .A1(n11985), .A2(n11996), .ZN(n12190) );
  OR2_X1 U11038 ( .A1(n11998), .A2(n11996), .ZN(n12191) );
  NOR2_X1 U11039 ( .A1(n11300), .A2(n14814), .ZN(n9881) );
  BUF_X2 U11040 ( .A(n16903), .Z(n17082) );
  CLKBUF_X2 U11041 ( .A(n12134), .Z(n9593) );
  BUF_X1 U11042 ( .A(n12012), .Z(n12275) );
  AND2_X1 U11043 ( .A1(n12845), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10192) );
  AND2_X1 U11044 ( .A1(n10401), .A2(n16220), .ZN(n12249) );
  AND2_X1 U11045 ( .A1(n10401), .A2(n10172), .ZN(n12251) );
  AND2_X1 U11046 ( .A1(n12845), .A2(n10529), .ZN(n10276) );
  CLKBUF_X2 U11047 ( .A(n11053), .Z(n11672) );
  CLKBUF_X2 U11048 ( .A(n11205), .Z(n11786) );
  INV_X4 U11049 ( .A(n10692), .ZN(n17030) );
  INV_X1 U11050 ( .A(n11892), .ZN(n11878) );
  NAND2_X1 U11051 ( .A1(n9963), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12260) );
  NAND2_X1 U11052 ( .A1(n10183), .A2(n10529), .ZN(n12268) );
  NAND2_X1 U11053 ( .A1(n12790), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12008) );
  CLKBUF_X2 U11054 ( .A(n10002), .Z(n16235) );
  NAND2_X1 U11055 ( .A1(n10663), .A2(n16781), .ZN(n15507) );
  NAND2_X2 U11056 ( .A1(n9648), .A2(n9632), .ZN(n11129) );
  NAND2_X1 U11057 ( .A1(n11120), .A2(n9594), .ZN(n11130) );
  INV_X1 U11058 ( .A(n13012), .ZN(n9996) );
  NAND4_X1 U11059 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11112) );
  AND4_X1 U11060 ( .A1(n11083), .A2(n11082), .A3(n11081), .A4(n11080), .ZN(
        n11099) );
  INV_X1 U11061 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10529) );
  AND2_X1 U11062 ( .A1(n11006), .A2(n13824), .ZN(n11205) );
  AND2_X1 U11063 ( .A1(n11004), .A2(n13813), .ZN(n11241) );
  AND2_X1 U11064 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16220) );
  OR2_X1 U11065 ( .A1(n11387), .A2(n11384), .ZN(n11290) );
  AND2_X1 U11066 ( .A1(n11005), .A2(n13813), .ZN(n11354) );
  INV_X1 U11067 ( .A(n11122), .ZN(n9594) );
  NAND2_X1 U11069 ( .A1(n9963), .A2(n10529), .ZN(n12017) );
  AND2_X1 U11070 ( .A1(n12877), .A2(n20926), .ZN(n12901) );
  INV_X1 U11071 ( .A(n10061), .ZN(n10047) );
  AND4_X1 U11072 ( .A1(n11091), .A2(n11090), .A3(n11089), .A4(n11088), .ZN(
        n11097) );
  INV_X1 U11073 ( .A(n10621), .ZN(n13207) );
  AOI21_X1 U11074 ( .B1(n14878), .B2(n14879), .A(n9846), .ZN(n12788) );
  AND2_X1 U11075 ( .A1(n16006), .A2(n16008), .ZN(n14856) );
  AND2_X1 U11076 ( .A1(n12875), .A2(n12874), .ZN(n12956) );
  INV_X1 U11077 ( .A(n17011), .ZN(n16903) );
  INV_X2 U11078 ( .A(n15507), .ZN(n10721) );
  INV_X2 U11079 ( .A(n17061), .ZN(n17027) );
  NOR2_X1 U11080 ( .A1(n11136), .A2(n19999), .ZN(n13875) );
  CLKBUF_X2 U11081 ( .A(n11100), .Z(n13810) );
  NAND2_X1 U11082 ( .A1(n13469), .A2(n19076), .ZN(n12857) );
  NAND2_X1 U11083 ( .A1(n15089), .A2(n12397), .ZN(n15229) );
  INV_X2 U11084 ( .A(n16821), .ZN(n17091) );
  NOR2_X1 U11086 ( .A1(n14125), .A2(n14114), .ZN(n15682) );
  CLKBUF_X3 U11087 ( .A(n11112), .Z(n19999) );
  XNOR2_X1 U11088 ( .A(n9847), .B(n10500), .ZN(n14878) );
  NAND2_X1 U11089 ( .A1(n9707), .A2(n12179), .ZN(n14084) );
  INV_X1 U11090 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19780) );
  NAND2_X1 U11091 ( .A1(n17141), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17286) );
  NOR2_X1 U11092 ( .A1(n17763), .A2(n15517), .ZN(n17627) );
  INV_X1 U11093 ( .A(n17744), .ZN(n17472) );
  AND2_X1 U11094 ( .A1(n12681), .A2(n11928), .ZN(n13440) );
  XNOR2_X1 U11095 ( .A(n12692), .B(n12691), .ZN(n14429) );
  INV_X1 U11096 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20926) );
  OR3_X1 U11097 ( .A1(n10651), .A2(n18711), .A3(n10658), .ZN(n9586) );
  OR3_X1 U11098 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n10667), .ZN(n9587) );
  NAND2_X1 U11099 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18711), .ZN(
        n10666) );
  NOR2_X2 U11100 ( .A1(n14907), .A2(n14901), .ZN(n13276) );
  OAI21_X2 U11101 ( .B1(n14320), .B2(n14322), .A(n14321), .ZN(n14577) );
  AND2_X1 U11102 ( .A1(n12602), .A2(n12623), .ZN(n9588) );
  INV_X2 U11103 ( .A(n13798), .ZN(n10219) );
  NAND2_X1 U11104 ( .A1(n13785), .A2(n13799), .ZN(n13798) );
  NAND2_X2 U11105 ( .A1(n15331), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16032) );
  AND2_X4 U11106 ( .A1(n15144), .A2(n15293), .ZN(n15331) );
  NAND2_X2 U11107 ( .A1(n19043), .A2(n19059), .ZN(n19042) );
  NOR2_X2 U11108 ( .A1(n17658), .A2(n10983), .ZN(n16606) );
  CLKBUF_X1 U11110 ( .A(n10701), .Z(n9592) );
  INV_X1 U11111 ( .A(n9591), .ZN(n17087) );
  NAND2_X2 U11112 ( .A1(n15061), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12511) );
  NOR2_X4 U11113 ( .A1(n15094), .A2(n9843), .ZN(n15061) );
  NOR2_X2 U11114 ( .A1(n15272), .A2(n16082), .ZN(n15355) );
  INV_X1 U11115 ( .A(n10692), .ZN(n9590) );
  NAND2_X2 U11116 ( .A1(n10124), .A2(n10123), .ZN(n10146) );
  OAI21_X2 U11117 ( .B1(n12320), .B2(n9899), .A(n9898), .ZN(n15146) );
  BUF_X1 U11118 ( .A(n10701), .Z(n9591) );
  NOR2_X1 U11119 ( .A1(n9915), .A2(n10666), .ZN(n10701) );
  NAND2_X2 U11120 ( .A1(n14642), .A2(n14146), .ZN(n14617) );
  NAND2_X2 U11121 ( .A1(n9825), .A2(n9823), .ZN(n14642) );
  NOR2_X2 U11122 ( .A1(n15123), .A2(n15122), .ZN(n15289) );
  NOR2_X2 U11123 ( .A1(n16046), .A2(n15093), .ZN(n15123) );
  INV_X2 U11124 ( .A(n16730), .ZN(n10901) );
  AOI211_X4 U11125 ( .C1(n9599), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n10854), .B(n10853), .ZN(n16730) );
  XNOR2_X1 U11126 ( .A(n13159), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14271) );
  AND2_X1 U11127 ( .A1(n9891), .A2(n12538), .ZN(n12539) );
  NAND2_X2 U11128 ( .A1(n15144), .A2(n13193), .ZN(n15094) );
  NAND2_X1 U11129 ( .A1(n12505), .A2(n12504), .ZN(n15156) );
  NOR2_X1 U11130 ( .A1(n13203), .A2(n13202), .ZN(n9749) );
  XNOR2_X1 U11131 ( .A(n10481), .B(n10477), .ZN(n14887) );
  OR2_X1 U11132 ( .A1(n15961), .A2(n18939), .ZN(n9710) );
  XNOR2_X1 U11133 ( .A(n12284), .B(n14193), .ZN(n14187) );
  CLKBUF_X1 U11134 ( .A(n12495), .Z(n12496) );
  NAND2_X1 U11135 ( .A1(n13731), .A2(n13733), .ZN(n13732) );
  NAND2_X1 U11136 ( .A1(n12108), .A2(n12107), .ZN(n9841) );
  NOR2_X2 U11137 ( .A1(n14836), .A2(n18939), .ZN(n15532) );
  XNOR2_X1 U11138 ( .A(n12602), .B(n11390), .ZN(n12617) );
  INV_X1 U11139 ( .A(n19508), .ZN(n12027) );
  BUF_X1 U11140 ( .A(n12195), .Z(n19191) );
  OR2_X1 U11141 ( .A1(n11985), .A2(n11992), .ZN(n19431) );
  INV_X1 U11142 ( .A(n11973), .ZN(n14023) );
  INV_X1 U11143 ( .A(n13050), .ZN(n9620) );
  NOR2_X1 U11144 ( .A1(n10139), .A2(n13573), .ZN(n19507) );
  AND2_X1 U11145 ( .A1(n10078), .A2(n10077), .ZN(n10079) );
  NOR2_X1 U11146 ( .A1(n12141), .A2(n12149), .ZN(n12140) );
  AND4_X1 U11147 ( .A1(n9647), .A2(n11155), .A3(n11154), .A4(n12703), .ZN(
        n11157) );
  INV_X2 U11148 ( .A(n12874), .ZN(n13571) );
  INV_X2 U11149 ( .A(n11878), .ZN(n11928) );
  NAND2_X1 U11150 ( .A1(n11864), .A2(n13882), .ZN(n11134) );
  INV_X2 U11151 ( .A(n12134), .ZN(n9692) );
  NAND2_X1 U11152 ( .A1(n11013), .A2(n11012), .ZN(n11116) );
  BUF_X2 U11153 ( .A(n12046), .Z(n12170) );
  INV_X1 U11154 ( .A(n12258), .ZN(n12049) );
  AND4_X1 U11155 ( .A1(n11095), .A2(n11094), .A3(n11093), .A4(n11092), .ZN(
        n11096) );
  BUF_X2 U11156 ( .A(n11241), .Z(n11739) );
  CLKBUF_X2 U11158 ( .A(n11219), .Z(n11220) );
  BUF_X2 U11159 ( .A(n11036), .Z(n11712) );
  CLKBUF_X2 U11161 ( .A(n9939), .Z(n12845) );
  BUF_X2 U11162 ( .A(n11354), .Z(n11787) );
  BUF_X2 U11163 ( .A(n11227), .Z(n11785) );
  BUF_X2 U11164 ( .A(n11106), .Z(n11620) );
  INV_X4 U11165 ( .A(n9644), .ZN(n9595) );
  INV_X4 U11166 ( .A(n17065), .ZN(n9596) );
  AND2_X2 U11167 ( .A1(n16220), .A2(n9883), .ZN(n10185) );
  INV_X1 U11169 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10922) );
  NOR2_X4 U11170 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13824) );
  AND3_X1 U11171 ( .A1(n9751), .A2(n9685), .A3(n9637), .ZN(n14272) );
  OAI21_X1 U11172 ( .B1(n14239), .B2(n14240), .A(n13134), .ZN(n13141) );
  AOI21_X1 U11173 ( .B1(n12539), .B2(n9894), .A(n9661), .ZN(n12543) );
  AND2_X1 U11174 ( .A1(n14560), .A2(n14559), .ZN(n14574) );
  CLKBUF_X1 U11175 ( .A(n13131), .Z(n9603) );
  OR2_X1 U11176 ( .A1(n14562), .A2(n14558), .ZN(n14560) );
  AOI21_X1 U11177 ( .B1(n15102), .B2(n13222), .A(n13221), .ZN(n13226) );
  OAI21_X1 U11178 ( .B1(n15132), .B2(n15131), .A(n12521), .ZN(n15102) );
  NAND2_X1 U11179 ( .A1(n15316), .A2(n12519), .ZN(n15132) );
  CLKBUF_X1 U11180 ( .A(n15229), .Z(n9612) );
  AND2_X1 U11181 ( .A1(n14725), .A2(n15579), .ZN(n14726) );
  AOI211_X1 U11182 ( .C1(n18958), .C2(n18961), .A(n14280), .B(n14279), .ZN(
        n14281) );
  NAND2_X1 U11183 ( .A1(n15144), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16082) );
  AOI211_X1 U11184 ( .C1(n15781), .C2(n14580), .A(n14579), .B(n14578), .ZN(
        n14581) );
  AOI21_X1 U11185 ( .B1(n14247), .B2(n16199), .A(n15049), .ZN(n14248) );
  XNOR2_X1 U11186 ( .A(n13169), .B(n13168), .ZN(n18961) );
  NAND2_X1 U11187 ( .A1(n12516), .A2(n15147), .ZN(n16051) );
  NOR2_X1 U11188 ( .A1(n17400), .A2(n12755), .ZN(n12767) );
  NAND3_X1 U11189 ( .A1(n9842), .A2(n15156), .A3(n16093), .ZN(n16092) );
  NAND2_X1 U11190 ( .A1(n14885), .A2(n10482), .ZN(n9847) );
  XNOR2_X1 U11191 ( .A(n9749), .B(n13208), .ZN(n14865) );
  NAND2_X1 U11192 ( .A1(n12506), .A2(n12304), .ZN(n9842) );
  NOR2_X1 U11193 ( .A1(n17401), .A2(n17402), .ZN(n17400) );
  NAND2_X1 U11194 ( .A1(n9633), .A2(n9733), .ZN(n15198) );
  NAND2_X1 U11195 ( .A1(n14887), .A2(n14886), .ZN(n14885) );
  XNOR2_X1 U11196 ( .A(n13203), .B(n13202), .ZN(n15052) );
  NAND2_X1 U11197 ( .A1(n12500), .A2(n12499), .ZN(n15158) );
  NOR2_X1 U11198 ( .A1(n16308), .A2(n15514), .ZN(n16288) );
  NOR2_X1 U11199 ( .A1(n17420), .A2(n10791), .ZN(n17419) );
  OR2_X1 U11200 ( .A1(n10481), .A2(n10480), .ZN(n10482) );
  AOI21_X1 U11201 ( .B1(n12724), .B2(n19967), .A(n12723), .ZN(n12725) );
  CLKBUF_X1 U11202 ( .A(n14960), .Z(n14970) );
  CLKBUF_X1 U11203 ( .A(n12469), .Z(n10643) );
  XNOR2_X1 U11204 ( .A(n9718), .B(n9717), .ZN(n14287) );
  MUX2_X1 U11205 ( .A(n12690), .B(n11928), .S(n14301), .Z(n12692) );
  CLKBUF_X1 U11206 ( .A(n13279), .Z(n14995) );
  NAND2_X1 U11207 ( .A1(n14309), .A2(n14302), .ZN(n14301) );
  NAND2_X1 U11208 ( .A1(n12283), .A2(n14012), .ZN(n12284) );
  NOR2_X1 U11209 ( .A1(n10805), .A2(n10791), .ZN(n17451) );
  AND2_X2 U11210 ( .A1(n14328), .A2(n14307), .ZN(n14309) );
  OR2_X1 U11211 ( .A1(n12494), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14086) );
  NAND2_X1 U11212 ( .A1(n10617), .A2(n10616), .ZN(n14853) );
  NAND2_X1 U11213 ( .A1(n14856), .A2(n9734), .ZN(n15004) );
  OR2_X1 U11214 ( .A1(n15964), .A2(n12419), .ZN(n12540) );
  NOR2_X1 U11215 ( .A1(n9667), .A2(n12912), .ZN(n12486) );
  NAND2_X1 U11216 ( .A1(n12139), .A2(n13924), .ZN(n16118) );
  NAND2_X1 U11217 ( .A1(n14362), .A2(n9687), .ZN(n15625) );
  NOR2_X1 U11218 ( .A1(n13732), .A2(n13781), .ZN(n13796) );
  NAND2_X1 U11219 ( .A1(n9803), .A2(n10791), .ZN(n17474) );
  NOR2_X1 U11220 ( .A1(n15531), .A2(n18939), .ZN(n15996) );
  AND2_X1 U11221 ( .A1(n10797), .A2(n9654), .ZN(n9631) );
  AND2_X1 U11222 ( .A1(n14031), .A2(n14037), .ZN(n14107) );
  OR2_X1 U11223 ( .A1(n11298), .A2(n11297), .ZN(n13795) );
  NAND2_X1 U11224 ( .A1(n10170), .A2(n10169), .ZN(n13606) );
  NOR2_X1 U11225 ( .A1(n12592), .A2(n11481), .ZN(n11298) );
  OAI21_X1 U11226 ( .B1(n12577), .B2(n11481), .A(n11338), .ZN(n13733) );
  AND2_X1 U11227 ( .A1(n9712), .A2(n9711), .ZN(n14836) );
  NAND2_X1 U11228 ( .A1(n13949), .A2(n13043), .ZN(n9712) );
  NAND2_X1 U11229 ( .A1(n11329), .A2(n11340), .ZN(n12577) );
  AND3_X1 U11230 ( .A1(n9881), .A2(n9880), .A3(n11339), .ZN(n11387) );
  OAI22_X1 U11231 ( .A1(n12009), .A2(n19463), .B1(n19431), .B2(n11984), .ZN(
        n11989) );
  OR2_X1 U11232 ( .A1(n11299), .A2(n11300), .ZN(n11328) );
  OR2_X1 U11233 ( .A1(n11985), .A2(n11997), .ZN(n12186) );
  NAND2_X1 U11234 ( .A1(n11312), .A2(n11311), .ZN(n13840) );
  NAND2_X1 U11235 ( .A1(n11978), .A2(n9694), .ZN(n19463) );
  CLKBUF_X1 U11236 ( .A(n13256), .Z(n14527) );
  XNOR2_X1 U11237 ( .A(n13018), .B(n13017), .ZN(n14267) );
  NAND2_X1 U11238 ( .A1(n9696), .A2(n9694), .ZN(n19082) );
  AND2_X1 U11239 ( .A1(n15682), .A2(n15681), .ZN(n15684) );
  OR2_X1 U11240 ( .A1(n11983), .A2(n11996), .ZN(n19543) );
  OR2_X1 U11241 ( .A1(n11983), .A2(n11992), .ZN(n12198) );
  NAND2_X1 U11242 ( .A1(n10164), .A2(n10163), .ZN(n10168) );
  XNOR2_X1 U11243 ( .A(n11185), .B(n11184), .ZN(n11300) );
  NAND2_X1 U11244 ( .A1(n11311), .A2(n11265), .ZN(n11299) );
  AND2_X1 U11245 ( .A1(n11201), .A2(n11200), .ZN(n14814) );
  NOR2_X2 U11246 ( .A1(n12544), .A2(n12462), .ZN(n13054) );
  OR2_X1 U11247 ( .A1(n11974), .A2(n11973), .ZN(n11998) );
  OAI22_X1 U11248 ( .A1(n13582), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12578), 
        .B2(n11260), .ZN(n11185) );
  NOR2_X1 U11249 ( .A1(n18127), .A2(n17287), .ZN(n17209) );
  NAND2_X2 U11250 ( .A1(n14539), .A2(n13672), .ZN(n14543) );
  NOR2_X2 U11251 ( .A1(n17332), .A2(n16440), .ZN(n17752) );
  OR2_X1 U11252 ( .A1(n11264), .A2(n11263), .ZN(n11265) );
  NAND2_X1 U11253 ( .A1(n9621), .A2(n9620), .ZN(n12544) );
  NAND2_X2 U11254 ( .A1(n13746), .A2(n13532), .ZN(n13694) );
  NAND2_X2 U11255 ( .A1(n10119), .A2(n10118), .ZN(n11973) );
  NAND2_X1 U11256 ( .A1(n10117), .A2(n10116), .ZN(n10118) );
  OAI21_X1 U11257 ( .B1(n18539), .B2(n15487), .A(n9903), .ZN(n18593) );
  OR2_X1 U11258 ( .A1(n15393), .A2(n15402), .ZN(n11997) );
  NAND2_X1 U11259 ( .A1(n13048), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13050) );
  NOR2_X2 U11260 ( .A1(n12328), .A2(n12327), .ZN(n12331) );
  NAND2_X1 U11261 ( .A1(n10136), .A2(n10133), .ZN(n15393) );
  AND2_X1 U11262 ( .A1(n10113), .A2(n10149), .ZN(n10115) );
  NAND2_X1 U11263 ( .A1(n10131), .A2(n10130), .ZN(n10139) );
  NAND2_X1 U11264 ( .A1(n12322), .A2(n12321), .ZN(n12328) );
  CLKBUF_X1 U11265 ( .A(n10132), .Z(n10133) );
  NOR2_X1 U11266 ( .A1(n10968), .A2(n17702), .ZN(n10970) );
  NAND2_X1 U11267 ( .A1(n18571), .A2(n18546), .ZN(n17768) );
  NOR2_X1 U11268 ( .A1(n13044), .A2(n15095), .ZN(n13045) );
  NOR2_X1 U11269 ( .A1(n19037), .A2(n19003), .ZN(n19036) );
  NAND2_X1 U11270 ( .A1(n15914), .A2(n11896), .ZN(n15906) );
  NAND2_X1 U11271 ( .A1(n11203), .A2(n11202), .ZN(n11256) );
  NOR2_X1 U11272 ( .A1(n10966), .A2(n17714), .ZN(n17704) );
  XNOR2_X1 U11273 ( .A(n10562), .B(n10564), .ZN(n10560) );
  CLKBUF_X1 U11274 ( .A(n11164), .Z(n11165) );
  NOR2_X1 U11275 ( .A1(n9785), .A2(n17715), .ZN(n17714) );
  INV_X1 U11276 ( .A(n13020), .ZN(n9616) );
  NAND2_X1 U11277 ( .A1(n10080), .A2(n10079), .ZN(n10082) );
  NAND2_X1 U11278 ( .A1(n11882), .A2(n11881), .ZN(n13939) );
  NAND2_X1 U11279 ( .A1(n13022), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13020) );
  NOR2_X2 U11280 ( .A1(n9769), .A2(n12226), .ZN(n12292) );
  NOR2_X1 U11281 ( .A1(n10902), .A2(n12738), .ZN(n16439) );
  OR2_X2 U11282 ( .A1(n17330), .A2(n18597), .ZN(n17398) );
  NAND2_X1 U11283 ( .A1(n9887), .A2(n10089), .ZN(n10153) );
  NAND2_X1 U11284 ( .A1(n12140), .A2(n12138), .ZN(n12226) );
  AND2_X1 U11285 ( .A1(n11873), .A2(n9724), .ZN(n13934) );
  NAND2_X1 U11286 ( .A1(n9650), .A2(n12887), .ZN(n13310) );
  XNOR2_X1 U11287 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n10728), .ZN(
        n17726) );
  OR2_X1 U11288 ( .A1(n11128), .A2(n11125), .ZN(n11156) );
  XNOR2_X1 U11289 ( .A(n10730), .B(n10952), .ZN(n10728) );
  AND2_X1 U11290 ( .A1(n10064), .A2(n12857), .ZN(n9635) );
  AND2_X2 U11291 ( .A1(n13145), .A2(n10076), .ZN(n10098) );
  INV_X1 U11292 ( .A(n9845), .ZN(n13145) );
  NAND2_X1 U11293 ( .A1(n12889), .A2(n12888), .ZN(n9727) );
  AND2_X1 U11294 ( .A1(n13175), .A2(n13468), .ZN(n12872) );
  INV_X2 U11295 ( .A(n10949), .ZN(n17291) );
  AND2_X1 U11296 ( .A1(n10074), .A2(n13173), .ZN(n10092) );
  NOR2_X1 U11297 ( .A1(n13027), .A2(n15151), .ZN(n13028) );
  OR2_X1 U11298 ( .A1(n10727), .A2(n10726), .ZN(n10952) );
  AND2_X1 U11299 ( .A1(n12874), .A2(n10056), .ZN(n13173) );
  AND2_X1 U11300 ( .A1(n11862), .A2(n11129), .ZN(n11152) );
  AOI211_X2 U11301 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n10771), .B(n10770), .ZN(n17264) );
  NOR2_X1 U11302 ( .A1(n11130), .A2(n14210), .ZN(n11132) );
  CLKBUF_X2 U11303 ( .A(n11888), .Z(n9625) );
  INV_X1 U11304 ( .A(n12775), .ZN(n11818) );
  NAND4_X1 U11305 ( .A1(n10670), .A2(n9924), .A3(n10669), .A4(n10668), .ZN(
        n17758) );
  AND4_X1 U11306 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n17280) );
  CLKBUF_X2 U11307 ( .A(n12900), .Z(n13164) );
  NAND2_X1 U11308 ( .A1(n11291), .A2(n11135), .ZN(n11121) );
  NAND2_X2 U11309 ( .A1(n11151), .A2(n19999), .ZN(n20800) );
  CLKBUF_X1 U11310 ( .A(n11151), .Z(n13532) );
  CLKBUF_X1 U11311 ( .A(n12901), .Z(n13163) );
  INV_X1 U11312 ( .A(n13029), .ZN(n9614) );
  NAND2_X1 U11313 ( .A1(n9692), .A2(n13012), .ZN(n10053) );
  AND2_X1 U11314 ( .A1(n9983), .A2(n10062), .ZN(n9613) );
  NAND2_X1 U11315 ( .A1(n10062), .A2(n9983), .ZN(n10074) );
  INV_X1 U11316 ( .A(n11046), .ZN(n11131) );
  NAND2_X1 U11317 ( .A1(n9622), .A2(n9714), .ZN(n13029) );
  INV_X1 U11318 ( .A(n11116), .ZN(n11291) );
  NOR2_X2 U11319 ( .A1(n11122), .A2(n11120), .ZN(n11864) );
  INV_X1 U11320 ( .A(n11129), .ZN(n14210) );
  CLKBUF_X1 U11321 ( .A(n11122), .Z(n11123) );
  OR2_X2 U11322 ( .A1(n16389), .A2(n16337), .ZN(n16391) );
  NAND2_X1 U11323 ( .A1(n10022), .A2(n10021), .ZN(n13182) );
  NAND2_X1 U11324 ( .A1(n11129), .A2(n11116), .ZN(n13258) );
  NOR2_X1 U11325 ( .A1(n17507), .A2(n17506), .ZN(n17487) );
  NAND2_X1 U11326 ( .A1(n11033), .A2(n11032), .ZN(n11046) );
  NAND2_X1 U11327 ( .A1(n9649), .A2(n9931), .ZN(n11122) );
  NAND2_X2 U11328 ( .A1(n11023), .A2(n11022), .ZN(n11135) );
  AOI211_X1 U11329 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n10696), .B(n10695), .ZN(n10708) );
  INV_X2 U11330 ( .A(U212), .ZN(n16388) );
  AND2_X1 U11331 ( .A1(n13034), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9622) );
  NAND2_X1 U11332 ( .A1(n10036), .A2(n9914), .ZN(n10037) );
  MUX2_X1 U11333 ( .A(n9969), .B(n9968), .S(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10048) );
  NAND2_X1 U11334 ( .A1(n10184), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12046) );
  NOR2_X1 U11335 ( .A1(n13033), .A2(n15164), .ZN(n13034) );
  AND4_X1 U11336 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n11078) );
  AND4_X1 U11337 ( .A1(n11063), .A2(n11062), .A3(n11061), .A4(n11060), .ZN(
        n11079) );
  AND4_X1 U11338 ( .A1(n11021), .A2(n11020), .A3(n11019), .A4(n11018), .ZN(
        n11022) );
  AND4_X1 U11339 ( .A1(n11017), .A2(n11016), .A3(n11015), .A4(n11014), .ZN(
        n11023) );
  AND4_X1 U11340 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11013) );
  AND4_X1 U11341 ( .A1(n11087), .A2(n11086), .A3(n11085), .A4(n11084), .ZN(
        n11098) );
  INV_X2 U11342 ( .A(U214), .ZN(n16389) );
  AND4_X1 U11343 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11033) );
  AND4_X1 U11344 ( .A1(n11031), .A2(n11030), .A3(n11029), .A4(n11028), .ZN(
        n11032) );
  AND4_X1 U11345 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n11012) );
  NAND2_X2 U11346 ( .A1(n18745), .A2(n18629), .ZN(n18689) );
  AND4_X1 U11347 ( .A1(n11075), .A2(n11074), .A3(n11073), .A4(n11072), .ZN(
        n11076) );
  AND4_X1 U11348 ( .A1(n11071), .A2(n11070), .A3(n11069), .A4(n11068), .ZN(
        n11077) );
  AOI21_X1 U11349 ( .B1(n11172), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10998), .ZN(n11001) );
  BUF_X2 U11350 ( .A(n11035), .Z(n11784) );
  AND2_X1 U11351 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  AND2_X1 U11352 ( .A1(n10032), .A2(n10031), .ZN(n10036) );
  OR2_X2 U11353 ( .A1(n12810), .A2(n10529), .ZN(n12266) );
  AND4_X1 U11354 ( .A1(n9962), .A2(n9961), .A3(n9960), .A4(n9959), .ZN(n9969)
         );
  AND4_X1 U11355 ( .A1(n9967), .A2(n9966), .A3(n9965), .A4(n9964), .ZN(n9968)
         );
  BUF_X2 U11356 ( .A(n11226), .Z(n11211) );
  INV_X2 U11357 ( .A(n18628), .ZN(n18685) );
  INV_X2 U11358 ( .A(n16425), .ZN(U215) );
  NAND3_X2 U11359 ( .A1(n18556), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17011) );
  CLKBUF_X2 U11360 ( .A(n10699), .Z(n9598) );
  INV_X4 U11361 ( .A(n10714), .ZN(n9599) );
  NAND2_X2 U11362 ( .A1(n16235), .A2(n10529), .ZN(n12258) );
  BUF_X2 U11363 ( .A(n11172), .Z(n11756) );
  AND2_X2 U11364 ( .A1(n11007), .A2(n10996), .ZN(n11226) );
  INV_X1 U11365 ( .A(n13035), .ZN(n9618) );
  AND2_X1 U11366 ( .A1(n11212), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10998) );
  AND2_X2 U11367 ( .A1(n18774), .A2(n19780), .ZN(n19040) );
  INV_X2 U11368 ( .A(n16428), .ZN(n16430) );
  NOR2_X2 U11370 ( .A1(n10656), .A2(n10658), .ZN(n17066) );
  NAND2_X1 U11371 ( .A1(n13038), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13035) );
  INV_X2 U11372 ( .A(n18763), .ZN(n18745) );
  INV_X1 U11373 ( .A(n9915), .ZN(n18556) );
  NAND2_X2 U11374 ( .A1(n10185), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12272) );
  INV_X2 U11375 ( .A(n20792), .ZN(n20794) );
  AND2_X1 U11376 ( .A1(n11007), .A2(n13824), .ZN(n11036) );
  AND2_X2 U11377 ( .A1(n10996), .A2(n9861), .ZN(n11107) );
  AND2_X2 U11378 ( .A1(n11006), .A2(n10996), .ZN(n11210) );
  INV_X2 U11379 ( .A(n13104), .ZN(n9600) );
  AND2_X1 U11380 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11048) );
  NOR2_X1 U11381 ( .A1(n18894), .A2(n9715), .ZN(n9714) );
  NOR2_X2 U11382 ( .A1(n13037), .A2(n16125), .ZN(n13038) );
  AND2_X1 U11383 ( .A1(n16733), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17701) );
  AND2_X1 U11384 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10994), .ZN(
        n11006) );
  OR3_X2 U11385 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18711), .A3(
        n18562), .ZN(n10732) );
  AND3_X1 U11386 ( .A1(n18727), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10665) );
  AND2_X1 U11387 ( .A1(n13652), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11004) );
  NOR2_X1 U11388 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10997), .ZN(
        n10999) );
  CLKBUF_X1 U11389 ( .A(n10922), .Z(n18733) );
  AND2_X1 U11390 ( .A1(n9933), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14075) );
  AND2_X1 U11391 ( .A1(n10172), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9939) );
  BUF_X2 U11392 ( .A(n10001), .Z(n9601) );
  INV_X2 U11393 ( .A(n11800), .ZN(n9602) );
  INV_X2 U11394 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18711) );
  NAND2_X2 U11395 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18562) );
  NAND2_X2 U11396 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13037) );
  INV_X1 U11397 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16125) );
  NOR2_X2 U11398 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13811) );
  AND2_X1 U11399 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13581) );
  NOR2_X1 U11400 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10172) );
  AND2_X1 U11401 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9861) );
  NOR2_X2 U11402 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16236) );
  NOR2_X1 U11403 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11005) );
  AND2_X1 U11404 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13813) );
  OR2_X2 U11405 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10658) );
  INV_X1 U11406 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18727) );
  NOR2_X4 U11408 ( .A1(n17230), .A2(n17399), .ZN(n17222) );
  AOI211_X4 U11409 ( .C1(n17090), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n10878), .B(n10877), .ZN(n18122) );
  NAND2_X1 U11410 ( .A1(n12433), .A2(n12432), .ZN(n13131) );
  NAND2_X1 U11411 ( .A1(n12228), .A2(n18923), .ZN(n12229) );
  NAND2_X1 U11412 ( .A1(n17627), .A2(n17969), .ZN(n9604) );
  NAND2_X1 U11413 ( .A1(n12757), .A2(n17749), .ZN(n9605) );
  AND2_X1 U11414 ( .A1(n9604), .A2(n9605), .ZN(n17657) );
  NOR2_X2 U11415 ( .A1(n18749), .A2(n16440), .ZN(n17749) );
  NOR2_X2 U11416 ( .A1(n17657), .A2(n17876), .ZN(n17549) );
  INV_X1 U11417 ( .A(n12810), .ZN(n9606) );
  NAND2_X1 U11418 ( .A1(n13617), .A2(n11973), .ZN(n9607) );
  NAND2_X1 U11419 ( .A1(n13617), .A2(n11973), .ZN(n11991) );
  NAND2_X1 U11420 ( .A1(n10150), .A2(n10149), .ZN(n10561) );
  BUF_X1 U11421 ( .A(n10150), .Z(n10119) );
  NAND2_X1 U11422 ( .A1(n10115), .A2(n10114), .ZN(n10150) );
  NAND2_X2 U11423 ( .A1(n9635), .A2(n10066), .ZN(n13210) );
  NOR2_X2 U11424 ( .A1(n12401), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12422) );
  CLKBUF_X1 U11425 ( .A(n19044), .Z(n9608) );
  INV_X1 U11426 ( .A(n19076), .ZN(n9609) );
  INV_X1 U11427 ( .A(n10179), .ZN(n9610) );
  NAND2_X1 U11428 ( .A1(n10096), .A2(n10060), .ZN(n9611) );
  XOR2_X1 U11429 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n13089), .Z(
        n16717) );
  NOR2_X1 U11430 ( .A1(n16467), .A2(n16468), .ZN(n16466) );
  INV_X1 U11431 ( .A(n16717), .ZN(n16297) );
  NOR2_X2 U11432 ( .A1(n15004), .A2(n15005), .ZN(n14994) );
  AND2_X1 U11433 ( .A1(n12874), .A2(n12134), .ZN(n12883) );
  NAND2_X1 U11434 ( .A1(n15610), .A2(n15609), .ZN(n15611) );
  INV_X1 U11435 ( .A(n12877), .ZN(n12874) );
  NAND2_X1 U11436 ( .A1(n9706), .A2(n12230), .ZN(n14188) );
  NOR2_X2 U11437 ( .A1(n14142), .A2(n14207), .ZN(n14386) );
  NOR2_X2 U11438 ( .A1(n9868), .A2(n13794), .ZN(n13860) );
  NOR2_X2 U11439 ( .A1(n14373), .A2(n14374), .ZN(n14455) );
  NOR2_X2 U11440 ( .A1(n15906), .A2(n14404), .ZN(n9726) );
  NOR2_X4 U11441 ( .A1(n14440), .A2(n14361), .ZN(n14362) );
  OR2_X2 U11442 ( .A1(n14449), .A2(n14438), .ZN(n14440) );
  NAND2_X2 U11443 ( .A1(n13901), .A2(n11878), .ZN(n11874) );
  INV_X4 U11444 ( .A(n11888), .ZN(n13901) );
  AND2_X1 U11445 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n9615) );
  AND2_X1 U11446 ( .A1(n9614), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13030) );
  AND2_X1 U11447 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9617) );
  AND2_X1 U11448 ( .A1(n9616), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13021) );
  AND2_X1 U11449 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9619) );
  AND2_X1 U11450 ( .A1(n9618), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13036) );
  AND2_X1 U11451 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n9621) );
  AND2_X1 U11452 ( .A1(n9620), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9713) );
  NAND2_X2 U11453 ( .A1(n14104), .A2(n10399), .ZN(n10439) );
  OAI21_X2 U11454 ( .B1(n12817), .B2(n14873), .A(n14875), .ZN(n14868) );
  NOR2_X2 U11455 ( .A1(n10524), .A2(n10523), .ZN(n12817) );
  NOR2_X4 U11456 ( .A1(n14039), .A2(n12952), .ZN(n14104) );
  NAND2_X2 U11457 ( .A1(n10219), .A2(n9856), .ZN(n14039) );
  NAND2_X2 U11458 ( .A1(n9897), .A2(n9896), .ZN(n16061) );
  NOR2_X2 U11459 ( .A1(n13763), .A2(n13764), .ZN(n13762) );
  NAND2_X1 U11460 ( .A1(n11974), .A2(n14023), .ZN(n11985) );
  NAND2_X1 U11461 ( .A1(n12494), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14085) );
  XNOR2_X2 U11462 ( .A(n10785), .B(n10786), .ZN(n17684) );
  OAI21_X2 U11463 ( .B1(n17582), .B2(n17911), .A(n10791), .ZN(n10797) );
  NOR2_X2 U11464 ( .A1(n17738), .A2(n10710), .ZN(n17727) );
  INV_X1 U11465 ( .A(n9622), .ZN(n13031) );
  NOR2_X1 U11466 ( .A1(n10656), .A2(n10658), .ZN(n9623) );
  NOR2_X2 U11467 ( .A1(n13771), .A2(n12930), .ZN(n13785) );
  NOR2_X1 U11468 ( .A1(n17261), .A2(n12727), .ZN(n17670) );
  AND2_X2 U11469 ( .A1(n12778), .A2(n11776), .ZN(n13121) );
  NOR3_X2 U11470 ( .A1(n14347), .A2(n9878), .A3(n14311), .ZN(n12778) );
  OAI21_X2 U11471 ( .B1(n12516), .B2(n12382), .A(n12381), .ZN(n15086) );
  NAND2_X1 U11472 ( .A1(n19999), .A2(n11136), .ZN(n11888) );
  XNOR2_X2 U11473 ( .A(n12487), .B(n12231), .ZN(n12494) );
  NAND3_X2 U11474 ( .A1(n12109), .A2(n9708), .A3(n12912), .ZN(n12487) );
  AND2_X1 U11475 ( .A1(n16220), .A2(n9883), .ZN(n9626) );
  AND2_X2 U11476 ( .A1(n16220), .A2(n9883), .ZN(n9627) );
  INV_X1 U11477 ( .A(n9626), .ZN(n9628) );
  OAI21_X2 U11478 ( .B1(n15229), .B2(n15231), .A(n15230), .ZN(n15066) );
  NOR2_X2 U11479 ( .A1(n13024), .A2(n15139), .ZN(n12528) );
  NOR2_X2 U11480 ( .A1(n13025), .A2(n18830), .ZN(n13026) );
  NOR2_X2 U11481 ( .A1(n13023), .A2(n20810), .ZN(n13022) );
  NAND2_X1 U11482 ( .A1(n18556), .A2(n10663), .ZN(n10699) );
  NAND2_X1 U11483 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10651), .ZN(
        n10656) );
  NOR2_X1 U11484 ( .A1(n11997), .A2(n11999), .ZN(n9695) );
  NAND2_X1 U11485 ( .A1(n10074), .A2(n10067), .ZN(n10058) );
  OR2_X1 U11486 ( .A1(n19999), .A2(n19998), .ZN(n11189) );
  AND2_X1 U11487 ( .A1(n14892), .A2(n14899), .ZN(n9850) );
  INV_X1 U11488 ( .A(n12487), .ZN(n9902) );
  NAND2_X1 U11489 ( .A1(n9888), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9887) );
  NAND3_X1 U11490 ( .A1(n9884), .A2(n9885), .A3(n10107), .ZN(n10149) );
  AND2_X1 U11491 ( .A1(n12134), .A2(n13012), .ZN(n10062) );
  NAND2_X1 U11492 ( .A1(n12134), .A2(n9996), .ZN(n10054) );
  NAND2_X1 U11493 ( .A1(n13664), .A2(n12576), .ZN(n12581) );
  AND2_X1 U11494 ( .A1(n11135), .A2(n11136), .ZN(n12621) );
  NAND2_X1 U11495 ( .A1(n12686), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11260) );
  AND3_X1 U11496 ( .A1(n11046), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n19999), 
        .ZN(n11853) );
  XNOR2_X1 U11497 ( .A(n13825), .B(n20157), .ZN(n13808) );
  NAND2_X1 U11498 ( .A1(n11260), .A2(n11189), .ZN(n11840) );
  CLKBUF_X1 U11499 ( .A(n12673), .Z(n12674) );
  AND2_X1 U11500 ( .A1(n14921), .A2(n12335), .ZN(n9773) );
  INV_X1 U11501 ( .A(n13790), .ZN(n9738) );
  NAND2_X1 U11502 ( .A1(n14188), .A2(n14187), .ZN(n9897) );
  AND2_X1 U11503 ( .A1(n10075), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10076) );
  AND2_X1 U11504 ( .A1(n10089), .A2(n10088), .ZN(n10090) );
  NAND2_X1 U11505 ( .A1(n10126), .A2(n10127), .ZN(n10134) );
  NAND2_X1 U11506 ( .A1(n9696), .A2(n11993), .ZN(n12195) );
  NOR2_X1 U11507 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10663) );
  INV_X1 U11508 ( .A(n10713), .ZN(n10720) );
  INV_X1 U11509 ( .A(n10683), .ZN(n17065) );
  NOR2_X1 U11510 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n9797), .ZN(
        n9796) );
  INV_X1 U11511 ( .A(n9918), .ZN(n9797) );
  AND2_X1 U11512 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n10728), .ZN(
        n10729) );
  XNOR2_X1 U11513 ( .A(n17280), .B(n17291), .ZN(n10709) );
  NOR2_X1 U11514 ( .A1(n18134), .A2(n10901), .ZN(n10908) );
  NAND2_X1 U11515 ( .A1(n13623), .A2(n13901), .ZN(n9724) );
  NAND2_X1 U11516 ( .A1(n11346), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11345) );
  NAND2_X1 U11517 ( .A1(n9916), .A2(n9832), .ZN(n9831) );
  INV_X1 U11518 ( .A(n14679), .ZN(n9832) );
  AND2_X1 U11519 ( .A1(n14589), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12643) );
  NOR2_X2 U11520 ( .A1(n12511), .A2(n14244), .ZN(n14243) );
  OR2_X1 U11521 ( .A1(n9900), .A2(n9683), .ZN(n9898) );
  AND2_X1 U11522 ( .A1(n9900), .A2(n12325), .ZN(n9899) );
  OR2_X1 U11523 ( .A1(n13473), .A2(n13472), .ZN(n13475) );
  OR2_X1 U11524 ( .A1(n19730), .A2(n19336), .ZN(n19368) );
  NOR2_X1 U11525 ( .A1(n9764), .A2(n9763), .ZN(n16467) );
  NOR2_X1 U11526 ( .A1(n17587), .A2(n17586), .ZN(n13090) );
  NAND2_X1 U11527 ( .A1(n16606), .A2(n17600), .ZN(n17587) );
  NAND2_X1 U11528 ( .A1(n9696), .A2(n9636), .ZN(n9697) );
  CLKBUF_X1 U11529 ( .A(n11712), .Z(n11738) );
  NAND2_X1 U11530 ( .A1(n12660), .A2(n13649), .ZN(n11150) );
  NAND2_X1 U11531 ( .A1(n11120), .A2(n11121), .ZN(n11126) );
  NOR2_X1 U11532 ( .A1(n9772), .A2(n12353), .ZN(n9771) );
  INV_X1 U11533 ( .A(n9904), .ZN(n9772) );
  NOR2_X1 U11534 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10401) );
  AND3_X1 U11535 ( .A1(n12176), .A2(n12175), .A3(n12174), .ZN(n12180) );
  INV_X1 U11536 ( .A(n15068), .ZN(n12412) );
  AND2_X1 U11537 ( .A1(n12224), .A2(n12223), .ZN(n12231) );
  NAND2_X1 U11538 ( .A1(n9611), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10152) );
  NAND2_X1 U11539 ( .A1(n10552), .A2(n9634), .ZN(n10089) );
  NAND2_X1 U11540 ( .A1(n10132), .A2(n10106), .ZN(n10114) );
  NAND2_X1 U11541 ( .A1(n9988), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9995) );
  NAND2_X1 U11542 ( .A1(n9993), .A2(n10529), .ZN(n9994) );
  NAND2_X1 U11543 ( .A1(n17267), .A2(n10760), .ZN(n10783) );
  OR2_X1 U11544 ( .A1(n17291), .A2(n17280), .ZN(n10730) );
  NAND2_X1 U11545 ( .A1(n11133), .A2(n19999), .ZN(n13235) );
  AND3_X1 U11546 ( .A1(n11291), .A2(n11826), .A3(n11131), .ZN(n13446) );
  INV_X1 U11547 ( .A(n11136), .ZN(n11151) );
  NAND2_X1 U11548 ( .A1(n9879), .A2(n14322), .ZN(n9878) );
  NOR2_X1 U11549 ( .A1(n14334), .A2(n14491), .ZN(n9879) );
  AOI21_X1 U11550 ( .B1(n9866), .B2(n11481), .A(n14403), .ZN(n9865) );
  NAND2_X1 U11551 ( .A1(n9863), .A2(n9866), .ZN(n9862) );
  NOR2_X1 U11552 ( .A1(n11129), .A2(n20689), .ZN(n11322) );
  NOR2_X1 U11553 ( .A1(n14610), .A2(n12638), .ZN(n14723) );
  INV_X1 U11554 ( .A(n9816), .ZN(n14608) );
  AOI21_X1 U11555 ( .B1(n14617), .B2(n9820), .A(n9817), .ZN(n9816) );
  INV_X1 U11556 ( .A(n9818), .ZN(n9817) );
  AOI21_X1 U11557 ( .B1(n9822), .B2(n9820), .A(n9819), .ZN(n9818) );
  OAI21_X1 U11558 ( .B1(n15805), .B2(n9814), .A(n12610), .ZN(n9813) );
  INV_X1 U11559 ( .A(n9813), .ZN(n9812) );
  NAND2_X1 U11560 ( .A1(n11361), .A2(n11383), .ZN(n12603) );
  INV_X1 U11561 ( .A(n11853), .ZN(n11845) );
  CLKBUF_X1 U11562 ( .A(n12661), .Z(n12662) );
  NAND2_X1 U11563 ( .A1(n11188), .A2(n11187), .ZN(n20157) );
  NAND2_X1 U11564 ( .A1(n12386), .A2(n12420), .ZN(n12383) );
  NAND2_X1 U11565 ( .A1(n12333), .A2(n12332), .ZN(n12343) );
  INV_X1 U11566 ( .A(n12348), .ZN(n12333) );
  NAND2_X1 U11567 ( .A1(n12306), .A2(n9774), .ZN(n12323) );
  AND2_X1 U11568 ( .A1(n18883), .A2(n13997), .ZN(n9774) );
  NAND2_X1 U11569 ( .A1(n10125), .A2(n13571), .ZN(n10517) );
  INV_X1 U11570 ( .A(n12180), .ZN(n12912) );
  NAND2_X1 U11571 ( .A1(n9615), .A2(n9614), .ZN(n13027) );
  INV_X1 U11572 ( .A(n14939), .ZN(n9746) );
  INV_X1 U11573 ( .A(n16165), .ZN(n9728) );
  NOR2_X1 U11574 ( .A1(n13800), .A2(n9740), .ZN(n9739) );
  INV_X1 U11575 ( .A(n13856), .ZN(n9740) );
  AND2_X1 U11576 ( .A1(n12507), .A2(n13138), .ZN(n12508) );
  AND3_X1 U11577 ( .A1(n12280), .A2(n12279), .A3(n12278), .ZN(n12920) );
  INV_X1 U11578 ( .A(n18941), .ZN(n9730) );
  INV_X1 U11579 ( .A(n18942), .ZN(n9729) );
  AND2_X1 U11580 ( .A1(n12496), .A2(n14085), .ZN(n9837) );
  INV_X1 U11581 ( .A(n13612), .ZN(n10570) );
  NAND2_X1 U11582 ( .A1(n12907), .A2(n13146), .ZN(n12024) );
  NAND2_X1 U11583 ( .A1(n10106), .A2(n10083), .ZN(n11967) );
  OAI21_X1 U11584 ( .B1(n12449), .B2(n10042), .A(n9845), .ZN(n10553) );
  OR2_X1 U11585 ( .A1(n12874), .A2(n10047), .ZN(n10042) );
  NAND2_X2 U11586 ( .A1(n16265), .A2(n12877), .ZN(n12144) );
  NAND2_X1 U11587 ( .A1(n9885), .A2(n10107), .ZN(n10112) );
  NAND2_X1 U11588 ( .A1(n13145), .A2(n16265), .ZN(n10066) );
  OR2_X1 U11589 ( .A1(n10517), .A2(n12098), .ZN(n10144) );
  NAND2_X1 U11590 ( .A1(n10013), .A2(n10529), .ZN(n10022) );
  NAND2_X1 U11591 ( .A1(n10020), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10021) );
  NAND2_X1 U11592 ( .A1(n9938), .A2(n10529), .ZN(n9946) );
  NAND3_X1 U11593 ( .A1(n18127), .A2(n18111), .A3(n18119), .ZN(n10906) );
  NOR2_X1 U11594 ( .A1(n17683), .A2(n10787), .ZN(n10789) );
  NOR2_X1 U11595 ( .A1(n10783), .A2(n17264), .ZN(n10784) );
  NOR2_X1 U11596 ( .A1(n18134), .A2(n18115), .ZN(n10937) );
  NAND2_X1 U11597 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17680), .ZN(
        n10978) );
  NOR2_X1 U11598 ( .A1(n10972), .A2(n17695), .ZN(n10975) );
  XOR2_X1 U11599 ( .A(n10783), .B(n17264), .Z(n10772) );
  AND2_X1 U11600 ( .A1(n10747), .A2(n10963), .ZN(n10760) );
  NOR2_X1 U11601 ( .A1(n17726), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9779) );
  INV_X1 U11602 ( .A(n10729), .ZN(n9784) );
  NOR2_X1 U11603 ( .A1(n17277), .A2(n10730), .ZN(n10747) );
  CLKBUF_X1 U11604 ( .A(n13235), .Z(n13236) );
  NOR2_X1 U11605 ( .A1(n11752), .A2(n14568), .ZN(n11753) );
  NAND2_X1 U11606 ( .A1(n11727), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11752) );
  AND2_X1 U11607 ( .A1(n9675), .A2(n11619), .ZN(n9874) );
  AND2_X1 U11608 ( .A1(n11563), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11564) );
  AND2_X1 U11609 ( .A1(n9671), .A2(n14143), .ZN(n9870) );
  AOI21_X1 U11610 ( .B1(n12583), .B2(n11495), .A(n11349), .ZN(n13781) );
  NOR2_X2 U11611 ( .A1(n15625), .A2(n14335), .ZN(n14336) );
  BUF_X1 U11612 ( .A(n14554), .Z(n15740) );
  NAND2_X1 U11613 ( .A1(n14651), .A2(n12629), .ZN(n9825) );
  NAND2_X1 U11614 ( .A1(n9726), .A2(n9725), .ZN(n13976) );
  INV_X1 U11615 ( .A(n13905), .ZN(n9725) );
  AND2_X1 U11616 ( .A1(n13940), .A2(n13850), .ZN(n15914) );
  NOR2_X2 U11617 ( .A1(n13939), .A2(n13938), .ZN(n13940) );
  NAND2_X1 U11618 ( .A1(n12555), .A2(n12621), .ZN(n12559) );
  MUX2_X1 U11619 ( .A(n11874), .B(n11867), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n11870) );
  NAND2_X1 U11620 ( .A1(n11861), .A2(n11860), .ZN(n13601) );
  NOR2_X1 U11621 ( .A1(n9670), .A2(n12226), .ZN(n12291) );
  NOR2_X1 U11622 ( .A1(n13912), .A2(n9859), .ZN(n9858) );
  INV_X1 U11623 ( .A(n9917), .ZN(n9859) );
  OR2_X1 U11624 ( .A1(n14929), .A2(n14923), .ZN(n14925) );
  INV_X1 U11625 ( .A(n14032), .ZN(n9741) );
  OAI21_X1 U11626 ( .B1(n16118), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n16116), .ZN(n12152) );
  AOI21_X1 U11627 ( .B1(n12431), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12537), .ZN(n12432) );
  INV_X1 U11628 ( .A(n12540), .ZN(n9895) );
  OR2_X1 U11629 ( .A1(n9844), .A2(n15069), .ZN(n9843) );
  INV_X1 U11630 ( .A(n13217), .ZN(n10616) );
  INV_X1 U11631 ( .A(n12524), .ZN(n10617) );
  NAND2_X1 U11632 ( .A1(n16061), .A2(n12313), .ZN(n12320) );
  NAND2_X1 U11633 ( .A1(n9736), .A2(n9679), .ZN(n13763) );
  INV_X1 U11634 ( .A(n13675), .ZN(n9736) );
  INV_X1 U11635 ( .A(n13676), .ZN(n9735) );
  XNOR2_X1 U11636 ( .A(n12302), .B(n12508), .ZN(n16093) );
  INV_X1 U11637 ( .A(n15159), .ZN(n12504) );
  AND2_X2 U11638 ( .A1(n10128), .A2(n10134), .ZN(n15402) );
  NAND2_X1 U11639 ( .A1(n13142), .A2(n10551), .ZN(n16263) );
  OAI21_X1 U11640 ( .B1(n19078), .B2(n19725), .A(n19724), .ZN(n19086) );
  NOR2_X1 U11641 ( .A1(n19077), .A2(n19119), .ZN(n19078) );
  INV_X1 U11642 ( .A(n19631), .ZN(n19077) );
  NOR2_X1 U11643 ( .A1(n9763), .A2(n17421), .ZN(n9765) );
  NOR2_X1 U11644 ( .A1(n16487), .A2(n16488), .ZN(n16486) );
  CLKBUF_X1 U11645 ( .A(n16717), .Z(n9763) );
  NOR2_X1 U11646 ( .A1(n10863), .A2(n10862), .ZN(n10864) );
  NOR2_X1 U11647 ( .A1(n17087), .A2(n16979), .ZN(n10863) );
  NOR3_X1 U11648 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n10922), .ZN(n10650) );
  OAI21_X1 U11649 ( .B1(n9598), .B2(n20883), .A(n10700), .ZN(n10704) );
  OR2_X1 U11650 ( .A1(n10689), .A2(n10688), .ZN(n10949) );
  NAND2_X1 U11651 ( .A1(n10982), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10983) );
  NAND2_X1 U11652 ( .A1(n10789), .A2(n17997), .ZN(n10790) );
  OR2_X1 U11653 ( .A1(n12728), .A2(n9907), .ZN(n15514) );
  NAND2_X1 U11654 ( .A1(n10809), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12728) );
  AND2_X1 U11655 ( .A1(n9791), .A2(n9800), .ZN(n10809) );
  NOR2_X1 U11656 ( .A1(n17451), .A2(n10808), .ZN(n9791) );
  INV_X1 U11657 ( .A(n10784), .ZN(n12727) );
  NAND2_X1 U11658 ( .A1(n10808), .A2(n9795), .ZN(n9792) );
  NAND2_X1 U11659 ( .A1(n17451), .A2(n9795), .ZN(n9794) );
  NAND2_X1 U11660 ( .A1(n9653), .A2(n9798), .ZN(n9800) );
  NAND2_X1 U11661 ( .A1(n9799), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9798) );
  INV_X1 U11662 ( .A(n10805), .ZN(n9799) );
  NAND2_X1 U11663 ( .A1(n10801), .A2(n10800), .ZN(n17455) );
  INV_X1 U11664 ( .A(n17457), .ZN(n10801) );
  NAND3_X1 U11665 ( .A1(n10797), .A2(n10796), .A3(n9801), .ZN(n9803) );
  NOR2_X1 U11666 ( .A1(n9802), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9801) );
  INV_X1 U11667 ( .A(n10795), .ZN(n9802) );
  NOR2_X1 U11668 ( .A1(n17640), .A2(n10793), .ZN(n17628) );
  XNOR2_X1 U11669 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n10772), .ZN(
        n17691) );
  NAND2_X1 U11670 ( .A1(n17705), .A2(n9790), .ZN(n9787) );
  INV_X1 U11671 ( .A(n17691), .ZN(n9790) );
  NAND2_X1 U11672 ( .A1(n10759), .A2(n9788), .ZN(n9786) );
  NOR2_X1 U11673 ( .A1(n17691), .A2(n9789), .ZN(n9788) );
  NAND2_X1 U11674 ( .A1(n17718), .A2(n10746), .ZN(n17707) );
  XNOR2_X1 U11675 ( .A(n10760), .B(n17267), .ZN(n17706) );
  NAND2_X1 U11676 ( .A1(n17720), .A2(n17719), .ZN(n17718) );
  INV_X1 U11677 ( .A(n10658), .ZN(n16781) );
  NAND2_X1 U11678 ( .A1(n18533), .A2(n10904), .ZN(n18564) );
  AND2_X1 U11679 ( .A1(n14417), .A2(n13874), .ZN(n19847) );
  INV_X1 U11680 ( .A(n12690), .ZN(n9717) );
  NAND2_X1 U11681 ( .A1(n9720), .A2(n9719), .ZN(n9718) );
  INV_X1 U11682 ( .A(n14464), .ZN(n14468) );
  INV_X1 U11683 ( .A(n14539), .ZN(n14532) );
  INV_X1 U11684 ( .A(n14287), .ZN(n14661) );
  XNOR2_X1 U11685 ( .A(n9831), .B(n14550), .ZN(n9830) );
  OR2_X1 U11686 ( .A1(n12709), .A2(n12694), .ZN(n19983) );
  OR2_X1 U11687 ( .A1(n13608), .A2(n19116), .ZN(n14942) );
  OR2_X1 U11688 ( .A1(n18995), .A2(n12996), .ZN(n16003) );
  NAND2_X1 U11689 ( .A1(n14243), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13159) );
  OR2_X1 U11690 ( .A1(n14865), .A2(n15384), .ZN(n13214) );
  INV_X1 U11691 ( .A(n16207), .ZN(n19063) );
  INV_X1 U11692 ( .A(n19507), .ZN(n19752) );
  AND2_X1 U11693 ( .A1(n13475), .A2(n13474), .ZN(n19744) );
  NAND2_X1 U11694 ( .A1(n16581), .A2(n9651), .ZN(n13287) );
  AND2_X1 U11695 ( .A1(n17426), .A2(n10981), .ZN(n10991) );
  OR2_X1 U11696 ( .A1(n17413), .A2(n17412), .ZN(n17414) );
  NAND2_X1 U11697 ( .A1(n17404), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17410) );
  NOR2_X1 U11698 ( .A1(n17483), .A2(n17418), .ZN(n9806) );
  NOR2_X1 U11699 ( .A1(n18714), .A2(n17689), .ZN(n17615) );
  INV_X1 U11700 ( .A(n17622), .ZN(n17671) );
  INV_X1 U11701 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10995) );
  NAND2_X1 U11702 ( .A1(n9701), .A2(n10065), .ZN(n10081) );
  AOI22_X1 U11703 ( .A1(n13210), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n10099), .ZN(n10065) );
  NAND2_X1 U11704 ( .A1(n10084), .A2(n9702), .ZN(n9701) );
  NOR2_X1 U11705 ( .A1(n9854), .A2(n19780), .ZN(n9702) );
  NOR2_X1 U11706 ( .A1(n12877), .A2(n19076), .ZN(n9889) );
  INV_X1 U11707 ( .A(n14609), .ZN(n9819) );
  INV_X1 U11708 ( .A(n11189), .ZN(n11252) );
  INV_X1 U11709 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10997) );
  NOR2_X1 U11710 ( .A1(n11182), .A2(n11181), .ZN(n12578) );
  AOI22_X1 U11711 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U11712 ( .A1(n11205), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U11713 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11002) );
  XNOR2_X1 U11714 ( .A(n11147), .B(n11159), .ZN(n20124) );
  INV_X1 U11715 ( .A(n12227), .ZN(n9770) );
  CLKBUF_X1 U11716 ( .A(n12845), .Z(n12827) );
  NAND2_X1 U11717 ( .A1(n14994), .A2(n14996), .ZN(n13279) );
  NAND2_X1 U11718 ( .A1(n12331), .A2(n9680), .ZN(n12348) );
  XNOR2_X1 U11719 ( .A(n12501), .B(n12502), .ZN(n12495) );
  OAI21_X1 U11720 ( .B1(n12181), .B2(n12033), .A(n9697), .ZN(n12034) );
  NAND2_X1 U11721 ( .A1(n9696), .A2(n9695), .ZN(n9693) );
  AND3_X1 U11722 ( .A1(n12081), .A2(n12080), .A3(n12079), .ZN(n12479) );
  NAND2_X1 U11723 ( .A1(n12860), .A2(n10057), .ZN(n13180) );
  NAND2_X1 U11724 ( .A1(n9886), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9885) );
  INV_X1 U11725 ( .A(n11990), .ZN(n11977) );
  AOI22_X1 U11726 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n9943) );
  INV_X1 U11727 ( .A(n9698), .ZN(n9934) );
  OAI22_X1 U11728 ( .A1(n15507), .A2(n10674), .B1(n17061), .B2(n10673), .ZN(
        n10675) );
  INV_X1 U11729 ( .A(n14444), .ZN(n9875) );
  NOR2_X1 U11730 ( .A1(n11467), .A2(n9873), .ZN(n9872) );
  NOR2_X1 U11731 ( .A1(n14139), .A2(n14117), .ZN(n9873) );
  NAND2_X1 U11732 ( .A1(n13972), .A2(n14117), .ZN(n14119) );
  NOR2_X1 U11733 ( .A1(n9662), .A2(n15785), .ZN(n9822) );
  AND2_X1 U11734 ( .A1(n14750), .A2(n9821), .ZN(n9820) );
  NAND2_X1 U11735 ( .A1(n15785), .A2(n9690), .ZN(n9821) );
  NAND2_X1 U11737 ( .A1(n13528), .A2(n12574), .ZN(n12575) );
  NAND2_X1 U11738 ( .A1(n11132), .A2(n13446), .ZN(n12673) );
  NAND2_X1 U11739 ( .A1(n11138), .A2(n11302), .ZN(n12684) );
  OR2_X1 U11740 ( .A1(n11233), .A2(n11232), .ZN(n12565) );
  OAI211_X1 U11741 ( .C1(n11150), .C2(n13532), .A(n11157), .B(n12699), .ZN(
        n11202) );
  NAND2_X1 U11742 ( .A1(n11239), .A2(n11238), .ZN(n11264) );
  INV_X1 U11743 ( .A(n11299), .ZN(n9880) );
  AOI22_X1 U11744 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U11745 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_8__3__SCAN_IN), .B2(n11205), .ZN(n11051) );
  OAI21_X1 U11746 ( .B1(n20801), .B2(n13835), .A(n14819), .ZN(n19997) );
  AOI22_X1 U11747 ( .A1(n12826), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n9997) );
  AOI22_X1 U11748 ( .A1(n12826), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U11749 ( .A1(n12416), .A2(n12420), .ZN(n12414) );
  INV_X1 U11750 ( .A(n12331), .ZN(n12358) );
  NAND2_X1 U11751 ( .A1(n12323), .A2(n12420), .ZN(n12322) );
  AND2_X1 U11752 ( .A1(n12307), .A2(n13806), .ZN(n12306) );
  OR2_X1 U11753 ( .A1(n12286), .A2(n9770), .ZN(n9768) );
  MUX2_X1 U11754 ( .A(n12452), .B(P2_EBX_REG_2__SCAN_IN), .S(n9593), .Z(n12141) );
  INV_X1 U11755 ( .A(n9848), .ZN(n10481) );
  INV_X1 U11756 ( .A(n14892), .ZN(n9851) );
  NAND2_X1 U11757 ( .A1(n9753), .A2(n14881), .ZN(n9752) );
  INV_X1 U11758 ( .A(n14888), .ZN(n9753) );
  NAND2_X1 U11759 ( .A1(n9617), .A2(n9616), .ZN(n13044) );
  NAND2_X1 U11760 ( .A1(n13026), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13024) );
  NAND2_X1 U11761 ( .A1(n13028), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13025) );
  INV_X1 U11762 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U11763 ( .A1(n9619), .A2(n9618), .ZN(n13033) );
  INV_X1 U11764 ( .A(n9733), .ZN(n14944) );
  NAND2_X1 U11765 ( .A1(n9666), .A2(n12412), .ZN(n9703) );
  NAND2_X1 U11766 ( .A1(n14960), .A2(n9732), .ZN(n9733) );
  AND2_X1 U11767 ( .A1(n14961), .A2(n14829), .ZN(n9732) );
  INV_X1 U11768 ( .A(n15066), .ZN(n12413) );
  AND2_X1 U11769 ( .A1(n12412), .A2(n9893), .ZN(n9892) );
  AND2_X1 U11770 ( .A1(n15982), .A2(n13138), .ZN(n12429) );
  NAND2_X1 U11771 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n9844) );
  NOR2_X1 U11772 ( .A1(n13274), .A2(n12419), .ZN(n12403) );
  NAND2_X1 U11773 ( .A1(n13848), .A2(n9678), .ZN(n13958) );
  INV_X1 U11774 ( .A(n9901), .ZN(n9900) );
  INV_X1 U11775 ( .A(n12956), .ZN(n12944) );
  NOR2_X1 U11776 ( .A1(n12501), .A2(n12503), .ZN(n12507) );
  NOR2_X1 U11777 ( .A1(n10157), .A2(n9704), .ZN(n10562) );
  NOR2_X1 U11778 ( .A1(n10154), .A2(n9705), .ZN(n9704) );
  OAI22_X1 U11779 ( .A1(n10152), .A2(n10529), .B1(n10151), .B2(n19734), .ZN(
        n10564) );
  NAND2_X1 U11780 ( .A1(n9921), .A2(n9910), .ZN(n12876) );
  OR2_X1 U11781 ( .A1(n13167), .A2(n19659), .ZN(n12889) );
  OR2_X1 U11782 ( .A1(n12023), .A2(n12022), .ZN(n12907) );
  NAND2_X1 U11783 ( .A1(n12868), .A2(n10071), .ZN(n10072) );
  AND2_X1 U11784 ( .A1(n13143), .A2(n13011), .ZN(n10071) );
  OR2_X1 U11785 ( .A1(n10517), .A2(n11999), .ZN(n10165) );
  NAND2_X1 U11786 ( .A1(n12874), .A2(n9882), .ZN(n10541) );
  INV_X1 U11787 ( .A(n16265), .ZN(n9882) );
  INV_X1 U11788 ( .A(n11967), .ZN(n11969) );
  NAND2_X1 U11789 ( .A1(n9956), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9957) );
  NAND2_X1 U11790 ( .A1(n10040), .A2(n10041), .ZN(n9845) );
  INV_X1 U11791 ( .A(n10054), .ZN(n10040) );
  NOR2_X1 U11792 ( .A1(n10667), .A2(n10656), .ZN(n10676) );
  NAND2_X1 U11793 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n10922), .ZN(
        n10667) );
  NOR2_X1 U11794 ( .A1(n10667), .A2(n10666), .ZN(n10693) );
  NOR4_X1 U11795 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n10922), .ZN(n10683) );
  NOR2_X1 U11796 ( .A1(n17011), .A2(n17130), .ZN(n10672) );
  NAND2_X1 U11797 ( .A1(n17404), .A2(n9642), .ZN(n13098) );
  NOR2_X1 U11798 ( .A1(n9631), .A2(n17538), .ZN(n17500) );
  INV_X1 U11799 ( .A(n18115), .ZN(n10907) );
  OAI21_X1 U11800 ( .B1(n18115), .B2(n10914), .A(n12736), .ZN(n10917) );
  NOR2_X1 U11801 ( .A1(n15612), .A2(n10919), .ZN(n12734) );
  OAI211_X1 U11802 ( .C1(n9598), .C2(n15417), .A(n10831), .B(n10830), .ZN(
        n12731) );
  AND2_X1 U11803 ( .A1(n14459), .A2(n14458), .ZN(n14461) );
  NAND2_X1 U11804 ( .A1(n13409), .A2(n13601), .ZN(n13534) );
  AOI21_X1 U11805 ( .B1(n11804), .B2(n11803), .A(n11802), .ZN(n13120) );
  AND2_X1 U11806 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n11726), .ZN(
        n11727) );
  AND2_X1 U11807 ( .A1(n11731), .A2(n11730), .ZN(n14322) );
  INV_X1 U11808 ( .A(n9879), .ZN(n9877) );
  NOR2_X1 U11809 ( .A1(n11669), .A2(n11668), .ZN(n11670) );
  NOR2_X1 U11810 ( .A1(n11645), .A2(n15630), .ZN(n11646) );
  NOR2_X1 U11811 ( .A1(n11598), .A2(n11597), .ZN(n11599) );
  NAND2_X1 U11812 ( .A1(n11599), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11645) );
  AND2_X1 U11813 ( .A1(n14454), .A2(n14456), .ZN(n9876) );
  NOR2_X1 U11814 ( .A1(n11531), .A2(n11530), .ZN(n11563) );
  OR2_X1 U11815 ( .A1(n11514), .A2(n11499), .ZN(n11531) );
  INV_X1 U11816 ( .A(n14389), .ZN(n11529) );
  NOR2_X1 U11817 ( .A1(n11478), .A2(n14129), .ZN(n11483) );
  AND2_X1 U11818 ( .A1(n14617), .A2(n14620), .ZN(n14765) );
  OR2_X1 U11819 ( .A1(n11463), .A2(n15702), .ZN(n11478) );
  AND2_X1 U11820 ( .A1(n11424), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11425) );
  NOR2_X1 U11821 ( .A1(n11420), .A2(n11419), .ZN(n11424) );
  AND2_X1 U11822 ( .A1(n9865), .A2(n13862), .ZN(n9864) );
  NAND2_X1 U11823 ( .A1(n9869), .A2(n11366), .ZN(n9867) );
  AND2_X1 U11824 ( .A1(n9862), .A2(n9865), .ZN(n9869) );
  AND2_X1 U11825 ( .A1(n11391), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11395) );
  AND2_X1 U11826 ( .A1(n11362), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11391) );
  NOR2_X1 U11827 ( .A1(n11345), .A2(n19856), .ZN(n11362) );
  AND2_X1 U11828 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11292), .ZN(
        n11346) );
  XNOR2_X1 U11829 ( .A(n12581), .B(n19955), .ZN(n13777) );
  XNOR2_X1 U11830 ( .A(n12651), .B(n14550), .ZN(n9828) );
  NOR2_X1 U11831 ( .A1(n12770), .A2(n14679), .ZN(n12771) );
  INV_X1 U11832 ( .A(n14346), .ZN(n9723) );
  NAND2_X1 U11833 ( .A1(n14362), .A2(n14346), .ZN(n15623) );
  NAND2_X1 U11834 ( .A1(n14461), .A2(n14451), .ZN(n14446) );
  NAND2_X1 U11835 ( .A1(n9722), .A2(n9721), .ZN(n14449) );
  INV_X1 U11836 ( .A(n14447), .ZN(n9721) );
  INV_X1 U11837 ( .A(n14446), .ZN(n9722) );
  NOR2_X2 U11839 ( .A1(n9643), .A2(n14380), .ZN(n14459) );
  NAND2_X1 U11840 ( .A1(n15684), .A2(n14208), .ZN(n14391) );
  AND2_X1 U11841 ( .A1(n15785), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15771) );
  OR2_X1 U11842 ( .A1(n14123), .A2(n11912), .ZN(n14125) );
  NOR2_X1 U11843 ( .A1(n9826), .A2(n9824), .ZN(n9823) );
  INV_X1 U11844 ( .A(n9681), .ZN(n9826) );
  INV_X1 U11845 ( .A(n12631), .ZN(n9824) );
  NOR2_X2 U11846 ( .A1(n13976), .A2(n13975), .ZN(n15709) );
  NAND2_X1 U11847 ( .A1(n15772), .A2(n12632), .ZN(n14146) );
  NOR2_X1 U11848 ( .A1(n15785), .A2(n12627), .ZN(n14652) );
  INV_X1 U11849 ( .A(n9726), .ZN(n14406) );
  INV_X1 U11850 ( .A(n9810), .ZN(n9809) );
  OAI21_X1 U11851 ( .B1(n9813), .B2(n12601), .A(n9665), .ZN(n9810) );
  AND2_X1 U11852 ( .A1(n15903), .A2(n15915), .ZN(n11896) );
  AND2_X1 U11853 ( .A1(n12609), .A2(n12608), .ZN(n15800) );
  NAND2_X1 U11854 ( .A1(n15806), .A2(n15805), .ZN(n15804) );
  INV_X1 U11855 ( .A(n13879), .ZN(n11882) );
  XNOR2_X1 U11856 ( .A(n12575), .B(n19990), .ZN(n13663) );
  AND2_X1 U11857 ( .A1(n13630), .A2(n12707), .ZN(n14772) );
  CLKBUF_X1 U11858 ( .A(n12684), .Z(n12685) );
  OR2_X1 U11859 ( .A1(n12709), .A2(n15544), .ZN(n13630) );
  NAND2_X1 U11860 ( .A1(n11204), .A2(n11256), .ZN(n11321) );
  OR2_X1 U11861 ( .A1(n11203), .A2(n11202), .ZN(n11204) );
  XNOR2_X1 U11862 ( .A(n11264), .B(n11262), .ZN(n11308) );
  NAND2_X1 U11863 ( .A1(n11328), .A2(n11301), .ZN(n13841) );
  INV_X1 U11864 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13652) );
  CLKBUF_X1 U11865 ( .A(n13581), .Z(n15541) );
  CLKBUF_X1 U11866 ( .A(n13232), .Z(n13233) );
  OR2_X1 U11867 ( .A1(n13840), .A2(n20528), .ZN(n20476) );
  NAND2_X1 U11868 ( .A1(n19998), .A2(n19997), .ZN(n20165) );
  AND2_X1 U11869 ( .A1(n13840), .A2(n20528), .ZN(n20445) );
  INV_X1 U11870 ( .A(n20165), .ZN(n20051) );
  AND3_X1 U11871 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n19998), .A3(n19997), 
        .ZN(n20039) );
  INV_X1 U11872 ( .A(n20519), .ZN(n20624) );
  INV_X1 U11873 ( .A(n14826), .ZN(n9709) );
  NOR2_X1 U11874 ( .A1(n12425), .A2(n12426), .ZN(n13073) );
  NAND2_X1 U11875 ( .A1(n12414), .A2(n12415), .ZN(n12425) );
  OR2_X1 U11876 ( .A1(n12399), .A2(n12398), .ZN(n12401) );
  NAND2_X1 U11877 ( .A1(n12383), .A2(n12384), .ZN(n12399) );
  NOR2_X1 U11878 ( .A1(n15532), .A2(n15533), .ZN(n15531) );
  NAND2_X1 U11879 ( .A1(n12339), .A2(n14921), .ZN(n12336) );
  CLKBUF_X1 U11880 ( .A(n15027), .Z(n15036) );
  NAND2_X1 U11881 ( .A1(n12331), .A2(n9904), .ZN(n12349) );
  NAND2_X1 U11882 ( .A1(n9767), .A2(n9766), .ZN(n9769) );
  NOR2_X1 U11883 ( .A1(n9768), .A2(n12290), .ZN(n9766) );
  INV_X1 U11884 ( .A(n12225), .ZN(n9767) );
  AND2_X1 U11885 ( .A1(n12292), .A2(n12288), .ZN(n12307) );
  AND2_X1 U11886 ( .A1(n13605), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U11887 ( .A1(n12788), .A2(n12789), .ZN(n14873) );
  NAND2_X1 U11888 ( .A1(n14900), .A2(n14899), .ZN(n14898) );
  AND2_X1 U11889 ( .A1(n14855), .A2(n14844), .ZN(n9734) );
  AND2_X1 U11890 ( .A1(n14218), .A2(n14217), .ZN(n14938) );
  NOR2_X1 U11891 ( .A1(n15359), .A2(n15360), .ZN(n13848) );
  AND3_X1 U11892 ( .A1(n12915), .A2(n12914), .A3(n12913), .ZN(n18942) );
  NOR2_X1 U11893 ( .A1(n18941), .A2(n18942), .ZN(n18943) );
  CLKBUF_X1 U11894 ( .A(n13380), .Z(n19071) );
  NAND2_X1 U11895 ( .A1(n13054), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13018) );
  CLKBUF_X1 U11896 ( .A(n13050), .Z(n13053) );
  CLKBUF_X1 U11897 ( .A(n13048), .Z(n13049) );
  OR2_X1 U11898 ( .A1(n12393), .A2(n15256), .ZN(n15088) );
  CLKBUF_X1 U11899 ( .A(n13045), .Z(n13047) );
  NAND2_X1 U11900 ( .A1(n9748), .A2(n14841), .ZN(n9747) );
  INV_X1 U11901 ( .A(n14852), .ZN(n9748) );
  CLKBUF_X1 U11902 ( .A(n13020), .Z(n13042) );
  CLKBUF_X1 U11903 ( .A(n13024), .Z(n13041) );
  CLKBUF_X1 U11904 ( .A(n13025), .Z(n13040) );
  CLKBUF_X1 U11905 ( .A(n13029), .Z(n13039) );
  NAND2_X1 U11906 ( .A1(n12429), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15082) );
  NAND2_X1 U11907 ( .A1(n14839), .A2(n14906), .ZN(n14907) );
  AND2_X1 U11908 ( .A1(n9674), .A2(n12526), .ZN(n9745) );
  NAND2_X1 U11909 ( .A1(n16031), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15133) );
  AOI21_X1 U11910 ( .B1(n15328), .B2(n12518), .A(n12517), .ZN(n15318) );
  NAND2_X1 U11911 ( .A1(n16051), .A2(n16049), .ZN(n15328) );
  CLKBUF_X1 U11912 ( .A(n13958), .Z(n14156) );
  NAND2_X1 U11913 ( .A1(n14107), .A2(n14108), .ZN(n14171) );
  NAND2_X1 U11914 ( .A1(n13762), .A2(n13784), .ZN(n15359) );
  INV_X1 U11915 ( .A(n13909), .ZN(n9737) );
  AND2_X1 U11916 ( .A1(n12285), .A2(n9676), .ZN(n9896) );
  NOR2_X1 U11917 ( .A1(n16193), .A2(n16195), .ZN(n16172) );
  AND3_X1 U11918 ( .A1(n12933), .A2(n12932), .A3(n12931), .ZN(n13676) );
  NAND2_X1 U11919 ( .A1(n13684), .A2(n13685), .ZN(n13675) );
  NOR2_X1 U11920 ( .A1(n13675), .A2(n13676), .ZN(n13679) );
  NAND2_X1 U11921 ( .A1(n9730), .A2(n9655), .ZN(n9731) );
  INV_X1 U11922 ( .A(n13739), .ZN(n9743) );
  NAND3_X1 U11923 ( .A1(n9838), .A2(n12497), .A3(n19042), .ZN(n9834) );
  INV_X1 U11924 ( .A(n13611), .ZN(n9744) );
  NAND2_X1 U11925 ( .A1(n16120), .A2(n12419), .ZN(n12139) );
  INV_X1 U11926 ( .A(n12876), .ZN(n13315) );
  OR2_X1 U11927 ( .A1(n19738), .A2(n19744), .ZN(n19279) );
  CLKBUF_X1 U11928 ( .A(n13949), .Z(n14070) );
  OAI21_X1 U11929 ( .B1(n10136), .B2(n15603), .A(n9852), .ZN(n13473) );
  INV_X1 U11930 ( .A(n9853), .ZN(n9852) );
  OAI21_X1 U11931 ( .B1(n10133), .B2(n15603), .A(n10138), .ZN(n9853) );
  INV_X1 U11932 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U11933 ( .A1(n10148), .A2(n10147), .ZN(n13616) );
  CLKBUF_X1 U11934 ( .A(n12444), .Z(n12445) );
  INV_X1 U11935 ( .A(n10541), .ZN(n13468) );
  OR2_X1 U11936 ( .A1(n19153), .A2(n19746), .ZN(n19132) );
  OR2_X1 U11937 ( .A1(n19132), .A2(n19752), .ZN(n19154) );
  OR2_X1 U11938 ( .A1(n19153), .A2(n19744), .ZN(n19186) );
  INV_X1 U11939 ( .A(n19112), .ZN(n19114) );
  AND2_X1 U11940 ( .A1(n19428), .A2(n19746), .ZN(n19465) );
  NOR3_X2 U11941 ( .A1(n19070), .A2(n19158), .A3(n19747), .ZN(n19112) );
  INV_X1 U11942 ( .A(n19506), .ZN(n19511) );
  CLKBUF_X1 U11943 ( .A(n12874), .Z(n13146) );
  NOR2_X1 U11944 ( .A1(n19730), .A2(n19279), .ZN(n19580) );
  NOR2_X1 U11945 ( .A1(n16507), .A2(n16508), .ZN(n16506) );
  NOR2_X1 U11946 ( .A1(n9652), .A2(n17473), .ZN(n16527) );
  INV_X1 U11947 ( .A(n17499), .ZN(n9761) );
  NOR2_X1 U11948 ( .A1(n16918), .A2(n16944), .ZN(n16899) );
  NAND2_X1 U11949 ( .A1(n18556), .A2(n10652), .ZN(n17074) );
  INV_X1 U11950 ( .A(n10656), .ZN(n10652) );
  NAND2_X1 U11951 ( .A1(n10720), .A2(n10719), .ZN(n10727) );
  OAI221_X1 U11952 ( .B1(n18563), .B2(n10902), .C1(n18563), .C2(n18749), .A(
        n14230), .ZN(n15610) );
  AOI21_X1 U11953 ( .B1(n14228), .B2(n18597), .A(n18619), .ZN(n17292) );
  NOR2_X1 U11954 ( .A1(n17403), .A2(n9757), .ZN(n9756) );
  NOR2_X1 U11955 ( .A1(n17470), .A2(n17469), .ZN(n17458) );
  NAND2_X1 U11956 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17558) );
  NAND2_X1 U11957 ( .A1(n17701), .A2(n9663), .ZN(n17658) );
  AND2_X1 U11958 ( .A1(n17701), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17688) );
  NAND2_X1 U11959 ( .A1(n17721), .A2(n17759), .ZN(n17689) );
  NOR2_X1 U11960 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15515), .ZN(
        n16287) );
  NOR2_X1 U11961 ( .A1(n17416), .A2(n15587), .ZN(n16307) );
  INV_X1 U11962 ( .A(n12756), .ZN(n12726) );
  NAND2_X1 U11963 ( .A1(n17669), .A2(n10790), .ZN(n17605) );
  INV_X1 U11964 ( .A(n17926), .ZN(n9776) );
  NOR2_X1 U11965 ( .A1(n12731), .A2(n10907), .ZN(n18549) );
  INV_X1 U11966 ( .A(n10790), .ZN(n10792) );
  AOI21_X1 U11967 ( .B1(n10979), .B2(n10978), .A(n10977), .ZN(n17668) );
  NOR2_X1 U11968 ( .A1(n18026), .A2(n17696), .ZN(n17695) );
  NAND2_X1 U11969 ( .A1(n9784), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9783) );
  NOR2_X1 U11970 ( .A1(n17750), .A2(n10691), .ZN(n17740) );
  NOR2_X1 U11971 ( .A1(n17740), .A2(n17739), .ZN(n17738) );
  XNOR2_X1 U11972 ( .A(n10949), .B(n10690), .ZN(n17751) );
  INV_X1 U11973 ( .A(n18541), .ZN(n15487) );
  INV_X1 U11974 ( .A(n12731), .ZN(n18111) );
  AOI211_X2 U11975 ( .C1(n10657), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n10899), .B(n10898), .ZN(n18119) );
  INV_X1 U11976 ( .A(n10921), .ZN(n18127) );
  NOR2_X1 U11977 ( .A1(n14130), .A2(n19857), .ZN(n15701) );
  NAND2_X1 U11978 ( .A1(n15642), .A2(n14254), .ZN(n19857) );
  AND2_X1 U11979 ( .A1(n14417), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19884) );
  INV_X1 U11980 ( .A(n19833), .ZN(n19879) );
  INV_X1 U11981 ( .A(n14472), .ZN(n19899) );
  OAI21_X1 U11982 ( .B1(n13600), .B2(n11866), .A(n11865), .ZN(n14464) );
  CLKBUF_X1 U11983 ( .A(n14211), .Z(n14528) );
  INV_X1 U11984 ( .A(n14518), .ZN(n14526) );
  NOR2_X1 U11985 ( .A1(n14532), .A2(n13672), .ZN(n14534) );
  NAND2_X1 U11986 ( .A1(n13244), .A2(n13243), .ZN(n14539) );
  INV_X1 U11987 ( .A(n14534), .ZN(n14542) );
  AND3_X1 U11988 ( .A1(n13479), .A2(n13478), .A3(n13601), .ZN(n19908) );
  NOR2_X1 U11989 ( .A1(n19908), .A2(n19936), .ZN(n19920) );
  BUF_X1 U11990 ( .A(n19920), .Z(n19935) );
  INV_X1 U11991 ( .A(n13746), .ZN(n13728) );
  OR2_X1 U11992 ( .A1(n13115), .A2(n14545), .ZN(n13116) );
  XNOR2_X1 U11993 ( .A(n13121), .B(n13120), .ZN(n14553) );
  AND2_X2 U11994 ( .A1(n12780), .A2(n20625), .ZN(n19947) );
  AND2_X1 U11995 ( .A1(n14636), .A2(n12784), .ZN(n15781) );
  INV_X1 U11996 ( .A(n19948), .ZN(n19803) );
  INV_X1 U11997 ( .A(n19947), .ZN(n19995) );
  XNOR2_X1 U11998 ( .A(n12655), .B(n12654), .ZN(n13129) );
  NAND2_X1 U11999 ( .A1(n12653), .A2(n12652), .ZN(n12655) );
  OAI21_X1 U12000 ( .B1(n14562), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14561), .ZN(n14563) );
  CLKBUF_X1 U12001 ( .A(n14599), .Z(n14600) );
  XNOR2_X1 U12002 ( .A(n11873), .B(n13623), .ZN(n13902) );
  INV_X1 U12003 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20521) );
  CLKBUF_X1 U12004 ( .A(n11321), .Z(n13963) );
  CLKBUF_X1 U12005 ( .A(n14423), .Z(n20315) );
  INV_X1 U12006 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20394) );
  CLKBUF_X1 U12007 ( .A(n13841), .Z(n13842) );
  AND2_X1 U12008 ( .A1(n14812), .A2(n20625), .ZN(n20621) );
  CLKBUF_X1 U12009 ( .A(n13582), .Z(n13583) );
  NAND2_X1 U12011 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13601), .ZN(n14819) );
  INV_X1 U12012 ( .A(n20231), .ZN(n20214) );
  INV_X1 U12013 ( .A(n20383), .ZN(n20387) );
  INV_X1 U12014 ( .A(n20534), .ZN(n20562) );
  INV_X1 U12015 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20689) );
  INV_X1 U12016 ( .A(n9712), .ZN(n14850) );
  INV_X1 U12017 ( .A(n18922), .ZN(n18947) );
  AND2_X1 U12018 ( .A1(n13076), .A2(n13077), .ZN(n18932) );
  INV_X1 U12019 ( .A(n18912), .ZN(n18922) );
  CLKBUF_X1 U12020 ( .A(n13055), .Z(n18933) );
  INV_X1 U12021 ( .A(n15072), .ZN(n15977) );
  NOR2_X1 U12022 ( .A1(n14174), .A2(n14173), .ZN(n14218) );
  INV_X1 U12023 ( .A(n14104), .ZN(n14174) );
  AND2_X1 U12024 ( .A1(n9672), .A2(n14040), .ZN(n9856) );
  CLKBUF_X1 U12025 ( .A(n13735), .Z(n13736) );
  AND2_X1 U12026 ( .A1(n14925), .A2(n14924), .ZN(n16009) );
  NAND2_X1 U12027 ( .A1(n12873), .A2(n19633), .ZN(n18995) );
  AND2_X1 U12028 ( .A1(n18973), .A2(n19116), .ZN(n18996) );
  CLKBUF_X1 U12030 ( .A(n13356), .Z(n13404) );
  INV_X1 U12031 ( .A(n14269), .ZN(n9750) );
  NAND2_X1 U12032 ( .A1(n14271), .A2(n19048), .ZN(n9751) );
  AND2_X1 U12033 ( .A1(n16124), .A2(n19743), .ZN(n19047) );
  XNOR2_X1 U12034 ( .A(n9603), .B(n9909), .ZN(n15194) );
  NAND2_X1 U12035 ( .A1(n9895), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9894) );
  INV_X1 U12036 ( .A(n15061), .ZN(n15063) );
  AND2_X1 U12037 ( .A1(n15156), .A2(n9842), .ZN(n16094) );
  CLKBUF_X1 U12038 ( .A(n14188), .Z(n14189) );
  INV_X1 U12039 ( .A(n16191), .ZN(n19064) );
  INV_X1 U12040 ( .A(n15384), .ZN(n19053) );
  INV_X1 U12041 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19751) );
  INV_X1 U12042 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19734) );
  NAND2_X1 U12043 ( .A1(n15402), .A2(n10158), .ZN(n10131) );
  OAI21_X1 U12044 ( .B1(n19080), .B2(n19118), .A(n19576), .ZN(n19122) );
  INV_X1 U12045 ( .A(n19152), .ZN(n19119) );
  INV_X1 U12046 ( .A(n19154), .ZN(n19181) );
  INV_X1 U12047 ( .A(n19216), .ZN(n19202) );
  OAI211_X1 U12048 ( .C1(n19228), .C2(n19224), .A(n19576), .B(n19223), .ZN(
        n19245) );
  OAI21_X1 U12049 ( .B1(n19228), .B2(n19227), .A(n19226), .ZN(n19244) );
  OR2_X1 U12050 ( .A1(n19368), .A2(n19337), .ZN(n19386) );
  OAI21_X1 U12051 ( .B1(n19407), .B2(n19422), .A(n19576), .ZN(n19424) );
  NOR2_X2 U12052 ( .A1(n19435), .A2(n19507), .ZN(n19455) );
  INV_X1 U12053 ( .A(n19535), .ZN(n19563) );
  INV_X1 U12054 ( .A(n19568), .ZN(n19627) );
  NOR2_X1 U12055 ( .A1(n16486), .A2(n9763), .ZN(n16479) );
  OAI21_X1 U12056 ( .B1(n16539), .B2(n9760), .A(n9759), .ZN(n13300) );
  NAND2_X1 U12057 ( .A1(n9762), .A2(n9761), .ZN(n9760) );
  NAND2_X1 U12058 ( .A1(n9763), .A2(n9762), .ZN(n9759) );
  INV_X1 U12059 ( .A(n17488), .ZN(n9762) );
  NOR2_X1 U12060 ( .A1(n16538), .A2(n9763), .ZN(n13301) );
  NOR2_X1 U12061 ( .A1(n16539), .A2(n17499), .ZN(n16538) );
  NOR2_X1 U12062 ( .A1(n13287), .A2(n17509), .ZN(n13286) );
  NAND2_X1 U12063 ( .A1(n16297), .A2(n9925), .ZN(n16581) );
  AND2_X1 U12064 ( .A1(n10867), .A2(n9911), .ZN(n18134) );
  INV_X1 U12065 ( .A(n16899), .ZN(n16931) );
  NOR2_X1 U12066 ( .A1(n16572), .A2(n16973), .ZN(n16961) );
  INV_X1 U12067 ( .A(n17114), .ZN(n17129) );
  NOR2_X2 U12068 ( .A1(n17360), .A2(n17155), .ZN(n17149) );
  NOR2_X1 U12069 ( .A1(n17165), .A2(n17356), .ZN(n17159) );
  NOR2_X1 U12070 ( .A1(n17352), .A2(n17175), .ZN(n17169) );
  NAND2_X1 U12071 ( .A1(n17169), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17165) );
  NOR3_X1 U12072 ( .A1(n17259), .A2(n17218), .A3(n17336), .ZN(n17210) );
  AOI211_X1 U12073 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n10756), .B(n10755), .ZN(n10757) );
  OR2_X1 U12074 ( .A1(n10743), .A2(n10742), .ZN(n10744) );
  AOI21_X1 U12075 ( .B1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n9599), .A(
        n10698), .ZN(n10707) );
  NOR2_X1 U12076 ( .A1(n10704), .A2(n10703), .ZN(n10705) );
  AOI21_X1 U12077 ( .B1(n9596), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(n10664), .ZN(n10669) );
  INV_X1 U12078 ( .A(n17290), .ZN(n17268) );
  INV_X1 U12079 ( .A(n17283), .ZN(n17285) );
  CLKBUF_X1 U12080 ( .A(n17318), .Z(n17326) );
  CLKBUF_X1 U12081 ( .A(n18760), .Z(n17327) );
  CLKBUF_X1 U12082 ( .A(n17395), .Z(n17387) );
  NOR2_X1 U12083 ( .A1(n17332), .A2(n17387), .ZN(n17388) );
  NAND2_X1 U12085 ( .A1(n17458), .A2(n9919), .ZN(n17433) );
  NAND2_X1 U12086 ( .A1(n13090), .A2(n9755), .ZN(n17507) );
  AND2_X1 U12087 ( .A1(n9638), .A2(n9923), .ZN(n9755) );
  NAND2_X1 U12088 ( .A1(n13090), .A2(n10984), .ZN(n17544) );
  NOR2_X1 U12089 ( .A1(n17965), .A2(n17876), .ZN(n17827) );
  AND2_X1 U12090 ( .A1(n17749), .A2(n17965), .ZN(n9777) );
  INV_X1 U12091 ( .A(n17627), .ZN(n17674) );
  INV_X1 U12092 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17731) );
  INV_X1 U12093 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17747) );
  INV_X1 U12094 ( .A(n17749), .ZN(n17764) );
  XNOR2_X1 U12095 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n15516), .ZN(
        n16322) );
  NAND2_X1 U12096 ( .A1(n9624), .A2(n12758), .ZN(n12754) );
  AND2_X1 U12097 ( .A1(n12767), .A2(n12730), .ZN(n12753) );
  OR2_X1 U12098 ( .A1(n12728), .A2(n12727), .ZN(n12729) );
  NOR2_X1 U12099 ( .A1(n12762), .A2(n12761), .ZN(n12763) );
  NAND2_X1 U12100 ( .A1(n9798), .A2(n9656), .ZN(n17430) );
  INV_X1 U12101 ( .A(n9803), .ZN(n17541) );
  NOR2_X2 U12102 ( .A1(n13099), .A2(n18564), .ZN(n18546) );
  INV_X1 U12103 ( .A(n17675), .ZN(n17999) );
  NOR2_X1 U12104 ( .A1(n9689), .A2(n17705), .ZN(n17692) );
  NAND2_X1 U12105 ( .A1(n9787), .A2(n9786), .ZN(n17690) );
  NOR2_X1 U12106 ( .A1(n17892), .A2(n18074), .ZN(n18052) );
  AND2_X1 U12107 ( .A1(n13255), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19996)
         );
  CLKBUF_X1 U12108 ( .A(n16420), .Z(n16425) );
  NAND2_X1 U12109 ( .A1(n14659), .A2(n19970), .ZN(n9716) );
  OAI211_X1 U12110 ( .C1(n14273), .C2(n16191), .A(n13216), .B(n9840), .ZN(
        P2_U3015) );
  NAND2_X1 U12111 ( .A1(n14271), .A2(n19063), .ZN(n9840) );
  AND3_X1 U12112 ( .A1(n13215), .A2(n9906), .A3(n13214), .ZN(n13216) );
  AOI21_X1 U12113 ( .B1(n15054), .B2(n19063), .A(n14250), .ZN(n14251) );
  NAND2_X1 U12114 ( .A1(n16779), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9754) );
  AOI21_X1 U12115 ( .B1(n13113), .B2(n16743), .A(n13112), .ZN(n13114) );
  AOI211_X1 U12116 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16794), .A(n16472), .B(
        n16471), .ZN(n16476) );
  NOR2_X1 U12117 ( .A1(n10991), .A2(n10990), .ZN(n10992) );
  NAND2_X1 U12118 ( .A1(n10989), .A2(n10988), .ZN(n10990) );
  NAND2_X1 U12119 ( .A1(n9807), .A2(n9804), .ZN(P3_U2802) );
  NOR3_X1 U12120 ( .A1(n17414), .A2(n9806), .A3(n9805), .ZN(n9804) );
  INV_X1 U12121 ( .A(n17417), .ZN(n9805) );
  INV_X2 U12122 ( .A(n9587), .ZN(n17077) );
  INV_X1 U12123 ( .A(n17066), .ZN(n10811) );
  INV_X1 U12124 ( .A(n10811), .ZN(n15471) );
  INV_X2 U12125 ( .A(n10844), .ZN(n10657) );
  AND2_X1 U12127 ( .A1(n9739), .A2(n9737), .ZN(n9629) );
  INV_X1 U12128 ( .A(n9855), .ZN(n14030) );
  INV_X2 U12129 ( .A(n9586), .ZN(n17090) );
  INV_X1 U12130 ( .A(n9778), .ZN(n17969) );
  NOR2_X1 U12131 ( .A1(n14347), .A2(n14491), .ZN(n14332) );
  OR2_X1 U12132 ( .A1(n15094), .A2(n9844), .ZN(n9630) );
  AOI211_X1 U12133 ( .C1(n16487), .C2(n16297), .A(n9765), .B(n17411), .ZN(
        n9764) );
  AND4_X1 U12134 ( .A1(n11044), .A2(n11043), .A3(n11042), .A4(n11041), .ZN(
        n9632) );
  INV_X1 U12135 ( .A(n11997), .ZN(n9694) );
  INV_X2 U12136 ( .A(n15785), .ZN(n15772) );
  OR2_X1 U12137 ( .A1(n14828), .A2(n14829), .ZN(n9633) );
  INV_X1 U12138 ( .A(n16265), .ZN(n19076) );
  OR2_X1 U12139 ( .A1(n12226), .A2(n9684), .ZN(n12287) );
  AND2_X2 U12140 ( .A1(n9946), .A2(n9945), .ZN(n12134) );
  OR2_X1 U12141 ( .A1(n14347), .A2(n9878), .ZN(n14321) );
  AND2_X1 U12142 ( .A1(n13175), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9634) );
  AND2_X1 U12143 ( .A1(n9694), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n9636)
         );
  INV_X1 U12144 ( .A(n12601), .ZN(n9814) );
  OR2_X1 U12145 ( .A1(n14865), .A2(n16034), .ZN(n9637) );
  AND2_X1 U12146 ( .A1(n10984), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9638) );
  NAND2_X1 U12147 ( .A1(n14455), .A2(n9675), .ZN(n9639) );
  OR2_X1 U12148 ( .A1(n14085), .A2(n12502), .ZN(n9640) );
  AND3_X2 U12149 ( .A1(n12133), .A2(n12132), .A3(n12131), .ZN(n12419) );
  NAND2_X1 U12150 ( .A1(n10219), .A2(n9917), .ZN(n13854) );
  NAND2_X1 U12151 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16795), .ZN(n16724) );
  INV_X1 U12152 ( .A(n16724), .ZN(n16779) );
  NAND2_X1 U12153 ( .A1(n9738), .A2(n9739), .ZN(n13855) );
  AND2_X1 U12154 ( .A1(n13972), .A2(n9671), .ZN(n9641) );
  AOI21_X1 U12155 ( .B1(n12617), .B2(n11495), .A(n11394), .ZN(n14402) );
  AND2_X1 U12156 ( .A1(n14160), .A2(n9674), .ZN(n12525) );
  AND2_X1 U12157 ( .A1(n13848), .A2(n9673), .ZN(n13956) );
  INV_X1 U12158 ( .A(n9871), .ZN(n14065) );
  AND2_X1 U12159 ( .A1(n9756), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9642) );
  NAND2_X1 U12160 ( .A1(n10219), .A2(n9858), .ZN(n9857) );
  NAND2_X1 U12161 ( .A1(n10219), .A2(n9672), .ZN(n9855) );
  AOI21_X1 U12162 ( .B1(n12603), .B2(n11495), .A(n11365), .ZN(n13865) );
  NAND2_X1 U12163 ( .A1(n13738), .A2(n13749), .ZN(n13748) );
  OR2_X1 U12164 ( .A1(n14391), .A2(n14390), .ZN(n9643) );
  OR2_X1 U12166 ( .A1(n17515), .A2(n17500), .ZN(n9645) );
  NAND2_X1 U12167 ( .A1(n10788), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9778) );
  NAND2_X2 U12168 ( .A1(n9995), .A2(n9994), .ZN(n12877) );
  AND2_X1 U12169 ( .A1(n14455), .A2(n14456), .ZN(n14453) );
  NAND2_X1 U12170 ( .A1(n9897), .A2(n12285), .ZN(n15161) );
  NOR3_X1 U12171 ( .A1(n13132), .A2(n12419), .A3(n13190), .ZN(n9646) );
  NOR2_X1 U12172 ( .A1(n13031), .A2(n18894), .ZN(n13032) );
  NOR2_X1 U12173 ( .A1(n15094), .A2(n13196), .ZN(n15077) );
  AND2_X1 U12174 ( .A1(n13576), .A2(n11114), .ZN(n9647) );
  NOR2_X1 U12175 ( .A1(n14358), .A2(n14359), .ZN(n14348) );
  NAND2_X1 U12176 ( .A1(n11974), .A2(n11973), .ZN(n11983) );
  INV_X1 U12177 ( .A(n11112), .ZN(n13882) );
  AND4_X1 U12178 ( .A1(n11040), .A2(n11039), .A3(n11038), .A4(n11037), .ZN(
        n9648) );
  AND4_X1 U12179 ( .A1(n11104), .A2(n11103), .A3(n11102), .A4(n11101), .ZN(
        n9649) );
  OR2_X1 U12180 ( .A1(n13167), .A2(n18789), .ZN(n9650) );
  INV_X1 U12181 ( .A(n13182), .ZN(n10067) );
  OR2_X1 U12182 ( .A1(n16717), .A2(n13091), .ZN(n9651) );
  NAND2_X1 U12183 ( .A1(n11387), .A2(n11386), .ZN(n12602) );
  NOR2_X1 U12184 ( .A1(n13300), .A2(n9763), .ZN(n9652) );
  NOR2_X1 U12185 ( .A1(n13275), .A2(n14888), .ZN(n14880) );
  BUF_X1 U12186 ( .A(n11131), .Z(n12686) );
  AND2_X1 U12187 ( .A1(n10804), .A2(n9796), .ZN(n9653) );
  XNOR2_X1 U12188 ( .A(n10168), .B(n10165), .ZN(n13615) );
  NOR2_X1 U12189 ( .A1(n14825), .A2(n18939), .ZN(n15950) );
  NAND2_X1 U12190 ( .A1(n16120), .A2(n16119), .ZN(n12490) );
  OR2_X1 U12192 ( .A1(n17605), .A2(n17876), .ZN(n9654) );
  AND2_X1 U12193 ( .A1(n9729), .A2(n14097), .ZN(n9655) );
  AND2_X1 U12194 ( .A1(n10804), .A2(n9918), .ZN(n9656) );
  AND2_X1 U12195 ( .A1(n14960), .A2(n14961), .ZN(n14828) );
  OR2_X1 U12196 ( .A1(n12673), .A2(n11888), .ZN(n9657) );
  NOR2_X1 U12197 ( .A1(n17725), .A2(n10729), .ZN(n9658) );
  OR2_X1 U12198 ( .A1(n13313), .A2(n9727), .ZN(n9659) );
  NOR2_X1 U12199 ( .A1(n12429), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15081) );
  INV_X1 U12200 ( .A(n15081), .ZN(n9893) );
  OR2_X1 U12201 ( .A1(n13275), .A2(n9752), .ZN(n9660) );
  AND2_X1 U12202 ( .A1(n12540), .A2(n15062), .ZN(n9661) );
  AND2_X1 U12203 ( .A1(n12637), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9662) );
  AND2_X1 U12204 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9663) );
  INV_X1 U12205 ( .A(n12496), .ZN(n12497) );
  NAND2_X1 U12206 ( .A1(n10570), .A2(n9743), .ZN(n9664) );
  NAND2_X1 U12207 ( .A1(n12611), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9665) );
  AND2_X1 U12208 ( .A1(n12423), .A2(n9893), .ZN(n9666) );
  NAND2_X1 U12209 ( .A1(n9829), .A2(n9827), .ZN(n14659) );
  NAND2_X1 U12210 ( .A1(n9902), .A2(n12231), .ZN(n12501) );
  NAND2_X1 U12211 ( .A1(n12320), .A2(n12319), .ZN(n15362) );
  AND2_X1 U12212 ( .A1(n12109), .A2(n9708), .ZN(n9667) );
  NAND2_X1 U12213 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10772), .ZN(
        n9668) );
  AND2_X1 U12214 ( .A1(n12331), .A2(n9771), .ZN(n9669) );
  INV_X1 U12215 ( .A(n9839), .ZN(n9838) );
  NAND2_X1 U12216 ( .A1(n14086), .A2(n12493), .ZN(n9839) );
  INV_X1 U12217 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9854) );
  INV_X1 U12218 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U12219 ( .A1(n13972), .A2(n9870), .ZN(n14142) );
  AND2_X1 U12220 ( .A1(n14856), .A2(n14855), .ZN(n14843) );
  NAND2_X1 U12221 ( .A1(n13848), .A2(n13849), .ZN(n13847) );
  NAND2_X1 U12222 ( .A1(n10792), .A2(n10791), .ZN(n17640) );
  OR2_X1 U12223 ( .A1(n12225), .A2(n9768), .ZN(n9670) );
  NOR2_X1 U12224 ( .A1(n9742), .A2(n9741), .ZN(n14031) );
  AND2_X1 U12225 ( .A1(n13860), .A2(n13971), .ZN(n13972) );
  OR2_X1 U12226 ( .A1(n13794), .A2(n13865), .ZN(n14401) );
  NAND2_X1 U12227 ( .A1(n14160), .A2(n9745), .ZN(n12524) );
  AND2_X1 U12228 ( .A1(n9872), .A2(n14066), .ZN(n9671) );
  AND2_X1 U12229 ( .A1(n9858), .A2(n9913), .ZN(n9672) );
  XNOR2_X1 U12230 ( .A(n12229), .B(n14093), .ZN(n14083) );
  AND2_X1 U12231 ( .A1(n9728), .A2(n13849), .ZN(n9673) );
  NAND2_X1 U12232 ( .A1(n9811), .A2(n9809), .ZN(n15793) );
  NAND2_X1 U12233 ( .A1(n9825), .A2(n12631), .ZN(n14145) );
  NAND2_X1 U12234 ( .A1(n15804), .A2(n12601), .ZN(n15799) );
  AND2_X1 U12235 ( .A1(n14162), .A2(n9746), .ZN(n9674) );
  NAND2_X1 U12236 ( .A1(n14160), .A2(n14162), .ZN(n14161) );
  NOR2_X1 U12237 ( .A1(n13958), .A2(n14157), .ZN(n14155) );
  NAND2_X1 U12238 ( .A1(n13777), .A2(n13776), .ZN(n13775) );
  AND2_X1 U12239 ( .A1(n11135), .A2(n9594), .ZN(n12567) );
  AND2_X1 U12240 ( .A1(n9876), .A2(n9875), .ZN(n9675) );
  NOR2_X1 U12241 ( .A1(n16098), .A2(n16095), .ZN(n9676) );
  NAND2_X1 U12242 ( .A1(n14455), .A2(n9876), .ZN(n14443) );
  NOR2_X1 U12243 ( .A1(n12226), .A2(n12225), .ZN(n9677) );
  AND2_X1 U12244 ( .A1(n9673), .A2(n13957), .ZN(n9678) );
  AND2_X1 U12245 ( .A1(n9735), .A2(n13680), .ZN(n9679) );
  NAND2_X1 U12246 ( .A1(n13972), .A2(n9872), .ZN(n9871) );
  NOR2_X1 U12247 ( .A1(n14853), .A2(n14852), .ZN(n14840) );
  AND2_X1 U12248 ( .A1(n12346), .A2(n9771), .ZN(n9680) );
  NAND2_X1 U12249 ( .A1(n10541), .A2(n12144), .ZN(n12868) );
  NAND2_X1 U12250 ( .A1(n15785), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9681) );
  INV_X1 U12251 ( .A(n9857), .ZN(n13913) );
  NAND2_X1 U12252 ( .A1(n19042), .A2(n12493), .ZN(n9682) );
  AND2_X1 U12253 ( .A1(n12319), .A2(n12325), .ZN(n9683) );
  NAND2_X1 U12254 ( .A1(n14898), .A2(n10441), .ZN(n14894) );
  NOR2_X1 U12255 ( .A1(n14853), .A2(n9747), .ZN(n14839) );
  OR2_X1 U12256 ( .A1(n12225), .A2(n9770), .ZN(n9684) );
  NOR2_X1 U12257 ( .A1(n14270), .A2(n9750), .ZN(n9685) );
  NOR2_X1 U12258 ( .A1(n9867), .A2(n13794), .ZN(n13861) );
  INV_X2 U12259 ( .A(n12795), .ZN(n10184) );
  INV_X1 U12260 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9785) );
  INV_X1 U12261 ( .A(n19977), .ZN(n19970) );
  INV_X1 U12262 ( .A(n11394), .ZN(n9866) );
  NAND2_X1 U12263 ( .A1(n13606), .A2(n13605), .ZN(n13604) );
  NOR2_X1 U12264 ( .A1(n13790), .A2(n13800), .ZN(n13801) );
  NOR2_X1 U12265 ( .A1(n13611), .A2(n9664), .ZN(n13738) );
  NAND2_X1 U12266 ( .A1(n13767), .A2(n13789), .ZN(n13790) );
  NOR2_X1 U12267 ( .A1(n13748), .A2(n13766), .ZN(n13767) );
  NAND2_X1 U12268 ( .A1(n9744), .A2(n10570), .ZN(n13609) );
  NAND2_X1 U12269 ( .A1(n10552), .A2(n13175), .ZN(n13209) );
  NOR2_X1 U12270 ( .A1(n13500), .A2(n12906), .ZN(n13921) );
  NAND2_X1 U12271 ( .A1(n12926), .A2(n12925), .ZN(n13684) );
  NAND2_X1 U12272 ( .A1(n9731), .A2(n12922), .ZN(n13682) );
  OR3_X1 U12273 ( .A1(n10460), .A2(n10459), .A3(n10458), .ZN(n9686) );
  NAND2_X1 U12274 ( .A1(n11978), .A2(n11977), .ZN(n19508) );
  OAI21_X1 U12275 ( .B1(n13841), .B2(n11481), .A(n11307), .ZN(n13656) );
  NOR2_X1 U12276 ( .A1(n15622), .A2(n9723), .ZN(n9687) );
  INV_X1 U12277 ( .A(n9713), .ZN(n13052) );
  OR2_X1 U12278 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n9688) );
  NAND2_X1 U12279 ( .A1(n9738), .A2(n9629), .ZN(n9742) );
  INV_X1 U12280 ( .A(n9598), .ZN(n17089) );
  INV_X1 U12281 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9705) );
  INV_X1 U12282 ( .A(n10676), .ZN(n10714) );
  AND2_X1 U12283 ( .A1(n13090), .A2(n9638), .ZN(n16548) );
  INV_X1 U12284 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9789) );
  NOR2_X1 U12285 ( .A1(n13098), .A2(n16469), .ZN(n13088) );
  NAND2_X1 U12286 ( .A1(n13934), .A2(n13933), .ZN(n13879) );
  NOR2_X1 U12287 ( .A1(n17433), .A2(n17432), .ZN(n17404) );
  AND2_X1 U12288 ( .A1(n10759), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9689) );
  NAND2_X1 U12289 ( .A1(n14618), .A2(n12554), .ZN(n9690) );
  NAND2_X1 U12290 ( .A1(n17404), .A2(n9756), .ZN(n9758) );
  AND2_X1 U12291 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16733) );
  INV_X1 U12292 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n9757) );
  INV_X1 U12293 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9795) );
  OAI21_X1 U12294 ( .B1(n17446), .B2(n17755), .A(n18201), .ZN(n17612) );
  OAI22_X2 U12295 ( .A1(n14517), .A2(n19115), .B1(n19097), .B2(n19114), .ZN(
        n19482) );
  OAI22_X2 U12296 ( .A1(n19101), .A2(n19115), .B1(n15022), .B2(n19114), .ZN(
        n19486) );
  OAI22_X2 U12297 ( .A1(n14998), .A2(n19115), .B1(n14999), .B2(n19114), .ZN(
        n19500) );
  AOI22_X2 U12298 ( .A1(DATAI_23_), .A2(n20037), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20036), .ZN(n20686) );
  AOI22_X2 U12299 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20036), .B1(DATAI_27_), 
        .B2(n20037), .ZN(n20651) );
  AOI22_X2 U12300 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20036), .B1(DATAI_24_), 
        .B2(n20037), .ZN(n20630) );
  OAI22_X2 U12301 ( .A1(n15015), .A2(n19115), .B1(n15016), .B2(n19114), .ZN(
        n19490) );
  INV_X1 U12302 ( .A(n19113), .ZN(n19115) );
  CLKBUF_X1 U12303 ( .A(n18946), .Z(n9691) );
  NOR4_X1 U12304 ( .A1(n19040), .A2(n18933), .A3(n19786), .A4(n16218), .ZN(
        n18946) );
  NOR2_X1 U12305 ( .A1(n18760), .A2(n17293), .ZN(n17318) );
  AOI22_X2 U12306 ( .A1(DATAI_20_), .A2(n20037), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20036), .ZN(n20657) );
  NOR2_X1 U12307 ( .A1(n12134), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12875) );
  NAND2_X1 U12308 ( .A1(n9593), .A2(n9688), .ZN(n9904) );
  AND2_X1 U12309 ( .A1(n9593), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12353) );
  AND2_X1 U12310 ( .A1(n9593), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12327) );
  AND2_X1 U12311 ( .A1(n9593), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12344) );
  AND2_X1 U12312 ( .A1(n9593), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12341) );
  AND2_X1 U12313 ( .A1(n9593), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12398) );
  AND2_X1 U12314 ( .A1(n9593), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12426) );
  NAND2_X2 U12315 ( .A1(n9996), .A2(n9692), .ZN(n10056) );
  MUX2_X1 U12316 ( .A(n12916), .B(n13743), .S(n9593), .Z(n12227) );
  MUX2_X1 U12317 ( .A(n12479), .B(n12135), .S(n9593), .Z(n12149) );
  MUX2_X1 U12318 ( .A(n12920), .B(P2_EBX_REG_6__SCAN_IN), .S(n9593), .Z(n12286) );
  MUX2_X1 U12319 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n12419), .S(n9692), .Z(n12290) );
  MUX2_X1 U12320 ( .A(n12450), .B(P2_EBX_REG_4__SCAN_IN), .S(n9593), .Z(n12225) );
  NAND2_X1 U12321 ( .A1(n12292), .A2(n9692), .ZN(n12420) );
  NOR2_X1 U12322 ( .A1(n12293), .A2(n9692), .ZN(n12294) );
  OAI21_X1 U12323 ( .B1(n12191), .B2(n12000), .A(n9693), .ZN(n12001) );
  INV_X2 U12324 ( .A(n11998), .ZN(n9696) );
  INV_X2 U12325 ( .A(n12802), .ZN(n10002) );
  NAND3_X2 U12326 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12802) );
  OAI21_X1 U12327 ( .B1(n12802), .B2(n9699), .A(n9700), .ZN(n9698) );
  NAND3_X1 U12328 ( .A1(n12444), .A2(n10085), .A3(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n9700) );
  INV_X2 U12329 ( .A(n12841), .ZN(n12826) );
  NAND2_X2 U12330 ( .A1(n12444), .A2(n10085), .ZN(n12841) );
  AND2_X2 U12331 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12444) );
  INV_X2 U12332 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10085) );
  NOR2_X2 U12333 ( .A1(n15066), .A2(n9703), .ZN(n12431) );
  INV_X2 U12334 ( .A(n10154), .ZN(n13204) );
  XNOR2_X2 U12335 ( .A(n10561), .B(n10560), .ZN(n11974) );
  NAND2_X1 U12336 ( .A1(n14084), .A2(n14083), .ZN(n9706) );
  NAND2_X1 U12337 ( .A1(n19044), .A2(n19045), .ZN(n9707) );
  NAND2_X1 U12338 ( .A1(n15146), .A2(n15148), .ZN(n12516) );
  NAND2_X2 U12339 ( .A1(n12025), .A2(n12024), .ZN(n9708) );
  XNOR2_X2 U12340 ( .A(n9708), .B(n9841), .ZN(n16120) );
  INV_X1 U12341 ( .A(n9710), .ZN(n14824) );
  AND2_X2 U12342 ( .A1(n9710), .A2(n9709), .ZN(n14825) );
  NOR2_X1 U12343 ( .A1(n15960), .A2(n15962), .ZN(n15961) );
  INV_X1 U12344 ( .A(n15113), .ZN(n9711) );
  NAND2_X1 U12345 ( .A1(n12528), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13023) );
  NAND2_X1 U12346 ( .A1(n13045), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13046) );
  NAND3_X1 U12347 ( .A1(n14665), .A2(n14664), .A3(n9716), .ZN(P1_U3001) );
  NAND2_X1 U12348 ( .A1(n14309), .A2(n11962), .ZN(n9719) );
  NAND2_X1 U12349 ( .A1(n14301), .A2(n11878), .ZN(n9720) );
  INV_X1 U12350 ( .A(n9727), .ZN(n12890) );
  INV_X2 U12351 ( .A(n12841), .ZN(n9963) );
  NAND2_X1 U12352 ( .A1(n13682), .A2(n13683), .ZN(n12926) );
  NOR2_X1 U12353 ( .A1(n15198), .A2(n19058), .ZN(n15199) );
  INV_X1 U12354 ( .A(n9742), .ZN(n13910) );
  NOR3_X2 U12355 ( .A1(n13275), .A2(n9752), .A3(n10644), .ZN(n12469) );
  NAND2_X1 U12356 ( .A1(n12469), .A2(n12468), .ZN(n12473) );
  NAND3_X1 U12357 ( .A1(n16463), .A2(n16464), .A3(n9754), .ZN(P3_U2640) );
  INV_X1 U12358 ( .A(n9758), .ZN(n16310) );
  NAND2_X1 U12359 ( .A1(n12339), .A2(n9773), .ZN(n12386) );
  OAI21_X1 U12360 ( .B1(n12422), .B2(n9775), .A(n12420), .ZN(n12421) );
  NAND2_X1 U12361 ( .A1(n9593), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U12362 ( .A1(n9778), .A2(n10790), .ZN(n17675) );
  AND2_X1 U12363 ( .A1(n17969), .A2(n9624), .ZN(n17629) );
  AND2_X1 U12364 ( .A1(n17969), .A2(n9776), .ZN(n17944) );
  AOI21_X1 U12365 ( .B1(n17627), .B2(n9778), .A(n9777), .ZN(n17656) );
  NAND2_X2 U12366 ( .A1(n10665), .A2(n18711), .ZN(n10692) );
  INV_X1 U12367 ( .A(n17727), .ZN(n9780) );
  NOR2_X2 U12368 ( .A1(n17727), .A2(n17726), .ZN(n17725) );
  NAND2_X1 U12369 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  OAI211_X2 U12370 ( .C1(n17725), .C2(n9783), .A(n9782), .B(n9781), .ZN(n17720) );
  NAND2_X1 U12371 ( .A1(n10729), .A2(n9785), .ZN(n9782) );
  AND3_X2 U12372 ( .A1(n9787), .A2(n9786), .A3(n9668), .ZN(n10785) );
  NAND3_X1 U12373 ( .A1(n9794), .A2(n9793), .A3(n9792), .ZN(n12756) );
  NAND3_X1 U12374 ( .A1(n9653), .A2(n9798), .A3(n9795), .ZN(n9793) );
  INV_X1 U12375 ( .A(n9800), .ZN(n17429) );
  INV_X1 U12376 ( .A(n17474), .ZN(n17515) );
  NAND3_X1 U12377 ( .A1(n10796), .A2(n10797), .A3(n10795), .ZN(n17542) );
  NAND2_X1 U12378 ( .A1(n9808), .A2(n17415), .ZN(n9807) );
  NOR2_X1 U12379 ( .A1(n17400), .A2(n17622), .ZN(n9808) );
  NAND2_X1 U12380 ( .A1(n15806), .A2(n9812), .ZN(n9811) );
  OAI21_X2 U12381 ( .B1(n12563), .B2(n12591), .A(n12562), .ZN(n13494) );
  XNOR2_X2 U12382 ( .A(n11319), .B(n11318), .ZN(n12563) );
  OAI21_X2 U12383 ( .B1(n11321), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9815), 
        .ZN(n11319) );
  INV_X1 U12384 ( .A(n11234), .ZN(n9815) );
  NAND2_X1 U12385 ( .A1(n12770), .A2(n12651), .ZN(n14548) );
  OR2_X1 U12386 ( .A1(n12770), .A2(n9831), .ZN(n14549) );
  NAND2_X1 U12387 ( .A1(n12770), .A2(n9828), .ZN(n9827) );
  OR2_X1 U12388 ( .A1(n12770), .A2(n9830), .ZN(n9829) );
  NAND2_X1 U12389 ( .A1(n9837), .A2(n9833), .ZN(n9835) );
  INV_X1 U12390 ( .A(n19042), .ZN(n9833) );
  NAND2_X1 U12391 ( .A1(n14090), .A2(n14085), .ZN(n12498) );
  NAND2_X1 U12392 ( .A1(n9838), .A2(n19042), .ZN(n14090) );
  NAND4_X1 U12393 ( .A1(n9836), .A2(n9640), .A3(n9835), .A4(n9834), .ZN(n14186) );
  NAND2_X1 U12394 ( .A1(n9839), .A2(n9837), .ZN(n9836) );
  INV_X1 U12395 ( .A(n9841), .ZN(n12109) );
  NAND2_X2 U12396 ( .A1(n16092), .A2(n12509), .ZN(n15144) );
  AND2_X1 U12397 ( .A1(n9847), .A2(n10501), .ZN(n9846) );
  OAI211_X1 U12398 ( .C1(n9851), .C2(n10441), .A(n9849), .B(n9686), .ZN(n9848)
         );
  NAND2_X1 U12399 ( .A1(n14900), .A2(n9850), .ZN(n9849) );
  XNOR2_X2 U12400 ( .A(n10439), .B(n10437), .ZN(n14900) );
  AND2_X2 U12401 ( .A1(n9854), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14074) );
  NAND2_X1 U12402 ( .A1(n13606), .A2(n9860), .ZN(n13735) );
  INV_X1 U12403 ( .A(n13735), .ZN(n10171) );
  NAND2_X1 U12404 ( .A1(n10081), .A2(n10082), .ZN(n10083) );
  OR2_X2 U12405 ( .A1(n10081), .A2(n10082), .ZN(n10106) );
  AND2_X2 U12406 ( .A1(n13581), .A2(n9861), .ZN(n11053) );
  AND2_X2 U12407 ( .A1(n13824), .A2(n9861), .ZN(n11105) );
  NOR2_X1 U12408 ( .A1(n13812), .A2(n9861), .ZN(n13816) );
  INV_X1 U12409 ( .A(n11135), .ZN(n11826) );
  INV_X1 U12410 ( .A(n12617), .ZN(n9863) );
  NAND3_X1 U12411 ( .A1(n11366), .A2(n9864), .A3(n9862), .ZN(n9868) );
  NAND2_X1 U12412 ( .A1(n14455), .A2(n9874), .ZN(n14358) );
  NOR2_X1 U12413 ( .A1(n14347), .A2(n9877), .ZN(n14320) );
  NAND2_X1 U12414 ( .A1(n9881), .A2(n9880), .ZN(n11340) );
  AND3_X2 U12415 ( .A1(n9883), .A2(n9854), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10001) );
  INV_X2 U12416 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9883) );
  INV_X1 U12417 ( .A(n10111), .ZN(n9884) );
  INV_X1 U12418 ( .A(n10152), .ZN(n9886) );
  NAND3_X1 U12419 ( .A1(n10106), .A2(n10083), .A3(n10134), .ZN(n10132) );
  NAND3_X1 U12420 ( .A1(n9890), .A2(n10064), .A3(n12857), .ZN(n9888) );
  NAND2_X1 U12421 ( .A1(n13145), .A2(n9889), .ZN(n9890) );
  NAND2_X1 U12422 ( .A1(n12413), .A2(n9892), .ZN(n9891) );
  XNOR2_X1 U12423 ( .A(n12539), .B(n12540), .ZN(n15057) );
  OAI21_X1 U12424 ( .B1(n12319), .B2(n12325), .A(n15363), .ZN(n9901) );
  NAND2_X2 U12425 ( .A1(n12649), .A2(n12648), .ZN(n12770) );
  CLKBUF_X1 U12426 ( .A(n13808), .Z(n20314) );
  XNOR2_X1 U12427 ( .A(n14242), .B(n14241), .ZN(n15056) );
  NAND2_X1 U12428 ( .A1(n11328), .A2(n14814), .ZN(n11329) );
  CLKBUF_X1 U12429 ( .A(n12656), .Z(n12697) );
  INV_X1 U12430 ( .A(n12656), .ZN(n11047) );
  AOI22_X1 U12431 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11053), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U12432 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11712), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11050) );
  AND2_X1 U12433 ( .A1(n13840), .A2(n12563), .ZN(n20572) );
  XNOR2_X1 U12434 ( .A(n13519), .B(n13520), .ZN(n19738) );
  NAND2_X1 U12435 ( .A1(n11170), .A2(n11169), .ZN(n13825) );
  OR2_X1 U12436 ( .A1(n11170), .A2(n11169), .ZN(n11171) );
  NAND2_X1 U12437 ( .A1(n11258), .A2(n20522), .ZN(n14423) );
  NAND2_X1 U12438 ( .A1(n11258), .A2(n11163), .ZN(n11170) );
  NOR2_X1 U12439 ( .A1(n13883), .A2(n13882), .ZN(n13892) );
  INV_X1 U12440 ( .A(n20124), .ZN(n11257) );
  NAND2_X1 U12441 ( .A1(n20124), .A2(n11158), .ZN(n11258) );
  INV_X1 U12442 ( .A(n10400), .ZN(n10179) );
  OR2_X1 U12443 ( .A1(n12755), .A2(n18536), .ZN(n9903) );
  AND4_X1 U12444 ( .A1(n10901), .A2(n10937), .A3(n18122), .A4(n10900), .ZN(
        n10902) );
  AND3_X1 U12445 ( .A1(n14245), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15273), .ZN(n9905) );
  NOR2_X1 U12446 ( .A1(n13201), .A2(n9905), .ZN(n9906) );
  OR2_X1 U12447 ( .A1(n10791), .A2(n12758), .ZN(n9907) );
  NOR2_X1 U12448 ( .A1(n11260), .A2(n11259), .ZN(n9908) );
  INV_X1 U12449 ( .A(n10153), .ZN(n10154) );
  AND2_X1 U12450 ( .A1(n14238), .A2(n13130), .ZN(n9909) );
  AND4_X1 U12451 ( .A1(n12059), .A2(n12058), .A3(n12057), .A4(n12056), .ZN(
        n9910) );
  AND3_X1 U12452 ( .A1(n10866), .A2(n10865), .A3(n10864), .ZN(n9911) );
  AND2_X1 U12453 ( .A1(n16053), .A2(n16052), .ZN(n9912) );
  NAND3_X1 U12454 ( .A1(n10246), .A2(n10245), .A3(n10244), .ZN(n9913) );
  AND3_X1 U12455 ( .A1(n10035), .A2(n10034), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9914) );
  OR2_X2 U12456 ( .A1(n18727), .A2(n10922), .ZN(n9915) );
  AND2_X1 U12457 ( .A1(n15785), .A2(n12650), .ZN(n9916) );
  NAND3_X1 U12458 ( .A1(n10218), .A2(n10217), .A3(n10216), .ZN(n9917) );
  OR2_X1 U12459 ( .A1(n10791), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9918) );
  AND2_X1 U12460 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9919) );
  INV_X1 U12461 ( .A(n11322), .ZN(n11687) );
  INV_X1 U12462 ( .A(n11687), .ZN(n13123) );
  INV_X1 U12463 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19742) );
  INV_X1 U12464 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11330) );
  INV_X1 U12465 ( .A(n17670), .ZN(n10807) );
  INV_X1 U12466 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12335) );
  INV_X1 U12467 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10800) );
  INV_X1 U12468 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10690) );
  AND2_X1 U12469 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .ZN(n9920) );
  NOR2_X1 U12470 ( .A1(n19052), .A2(n18809), .ZN(n12529) );
  INV_X1 U12471 ( .A(n18924), .ZN(n13079) );
  AND4_X1 U12472 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n9921) );
  INV_X1 U12473 ( .A(n17074), .ZN(n10750) );
  AND2_X1 U12474 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9922) );
  AND2_X1 U12475 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9923) );
  INV_X1 U12476 ( .A(n18090), .ZN(n18074) );
  AND4_X1 U12477 ( .A1(n10662), .A2(n10661), .A3(n10660), .A4(n10659), .ZN(
        n9924) );
  OR2_X1 U12478 ( .A1(n16592), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n9925) );
  NOR2_X1 U12479 ( .A1(n16458), .A2(n13108), .ZN(n9926) );
  INV_X1 U12480 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n19998) );
  OR2_X1 U12481 ( .A1(n12836), .A2(n12835), .ZN(n9927) );
  OR2_X1 U12482 ( .A1(n10784), .A2(n15517), .ZN(n9928) );
  INV_X2 U12483 ( .A(n10693), .ZN(n17061) );
  AND2_X1 U12484 ( .A1(n12553), .A2(n12552), .ZN(n9929) );
  INV_X1 U12485 ( .A(n10643), .ZN(n12547) );
  XOR2_X1 U12486 ( .A(n15160), .B(n12304), .Z(n9930) );
  AND4_X1 U12487 ( .A1(n11111), .A2(n11110), .A3(n11109), .A4(n11108), .ZN(
        n9931) );
  AND2_X1 U12488 ( .A1(n12695), .A2(n11134), .ZN(n9932) );
  INV_X1 U12489 ( .A(n11840), .ZN(n11838) );
  NAND2_X1 U12490 ( .A1(n12826), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10015) );
  BUF_X1 U12491 ( .A(n11107), .Z(n11762) );
  AND2_X1 U12492 ( .A1(n10062), .A2(n13011), .ZN(n10063) );
  NAND2_X1 U12493 ( .A1(n12826), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10025) );
  AND2_X1 U12494 ( .A1(n20521), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11825) );
  INV_X1 U12495 ( .A(n14437), .ZN(n11619) );
  INV_X1 U12496 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11305) );
  NOR2_X1 U12497 ( .A1(n11135), .A2(n11136), .ZN(n11137) );
  AOI22_X1 U12498 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11712), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11016) );
  AND3_X1 U12499 ( .A1(n11255), .A2(n11254), .A3(n11253), .ZN(n11262) );
  AOI22_X1 U12500 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n9941) );
  INV_X1 U12501 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U12502 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11106), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11043) );
  OR2_X1 U12503 ( .A1(n11251), .A2(n11250), .ZN(n12566) );
  INV_X1 U12504 ( .A(n13258), .ZN(n11302) );
  INV_X1 U12505 ( .A(n20800), .ZN(n12607) );
  OR2_X1 U12506 ( .A1(n11218), .A2(n11217), .ZN(n12625) );
  INV_X1 U12507 ( .A(n12407), .ZN(n12405) );
  AOI22_X1 U12508 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n9970) );
  INV_X1 U12509 ( .A(n12548), .ZN(n12468) );
  NAND2_X1 U12510 ( .A1(n12422), .A2(n10637), .ZN(n12407) );
  AND2_X1 U12511 ( .A1(n12282), .A2(n12281), .ZN(n12502) );
  INV_X1 U12512 ( .A(n11992), .ZN(n11993) );
  NAND2_X1 U12513 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10736) );
  AND2_X1 U12514 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10862) );
  NOR2_X1 U12515 ( .A1(n11235), .A2(n19998), .ZN(n12622) );
  NOR2_X1 U12516 ( .A1(n14762), .A2(n15771), .ZN(n14750) );
  INV_X1 U12517 ( .A(n13881), .ZN(n11881) );
  AND2_X1 U12518 ( .A1(n11853), .A2(n12621), .ZN(n11848) );
  NOR2_X1 U12519 ( .A1(n10530), .A2(n10545), .ZN(n10531) );
  NAND2_X1 U12520 ( .A1(n12406), .A2(n12405), .ZN(n12416) );
  AOI21_X1 U12521 ( .B1(n10905), .B2(n10906), .A(n12734), .ZN(n10914) );
  OAI21_X1 U12522 ( .B1(n17011), .B2(n17120), .A(n10736), .ZN(n10737) );
  AND2_X1 U12523 ( .A1(n16828), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10671) );
  INV_X1 U12524 ( .A(n11874), .ZN(n11943) );
  OAI211_X1 U12525 ( .C1(n15570), .C2(n20394), .A(n11168), .B(n11167), .ZN(
        n11169) );
  AND2_X1 U12526 ( .A1(n11885), .A2(n11884), .ZN(n13938) );
  NAND2_X1 U12527 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11331) );
  INV_X1 U12528 ( .A(n11481), .ZN(n11495) );
  NAND2_X1 U12529 ( .A1(n15772), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14561) );
  AOI21_X1 U12530 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19734), .A(
        n10531), .ZN(n10544) );
  AND2_X1 U12531 ( .A1(n10475), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10140) );
  NAND2_X1 U12532 ( .A1(n10440), .A2(n10437), .ZN(n10441) );
  AND2_X1 U12533 ( .A1(n13011), .A2(n20926), .ZN(n12882) );
  AND2_X1 U12534 ( .A1(n12361), .A2(n12360), .ZN(n18844) );
  NAND2_X2 U12535 ( .A1(n10038), .A2(n10037), .ZN(n10061) );
  INV_X1 U12536 ( .A(n10738), .ZN(n10739) );
  NOR2_X1 U12537 ( .A1(n10718), .A2(n10717), .ZN(n10719) );
  NOR2_X1 U12538 ( .A1(n10672), .A2(n10671), .ZN(n10682) );
  INV_X1 U12539 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U12540 ( .A1(n10807), .A2(n9928), .ZN(n10786) );
  NOR2_X1 U12541 ( .A1(n10961), .A2(n17728), .ZN(n10964) );
  INV_X1 U12542 ( .A(n19884), .ZN(n19855) );
  NAND2_X1 U12543 ( .A1(n13892), .A2(n13891), .ZN(n19877) );
  NAND2_X1 U12544 ( .A1(n15709), .A2(n15708), .ZN(n14123) );
  AND2_X1 U12546 ( .A1(n11483), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11498) );
  AND2_X1 U12547 ( .A1(n11495), .A2(n11438), .ZN(n14139) );
  NAND2_X1 U12548 ( .A1(n11395), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11420) );
  INV_X1 U12549 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19856) );
  OR2_X1 U12550 ( .A1(n19948), .A2(n12782), .ZN(n14636) );
  INV_X1 U12551 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14550) );
  NAND2_X1 U12552 ( .A1(n12641), .A2(n15785), .ZN(n14601) );
  OR2_X1 U12553 ( .A1(n12709), .A2(n13600), .ZN(n19981) );
  NAND2_X1 U12554 ( .A1(n12680), .A2(n13240), .ZN(n12709) );
  OR2_X1 U12555 ( .A1(n13842), .A2(n14811), .ZN(n20283) );
  INV_X1 U12556 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20482) );
  INV_X1 U12557 ( .A(n12414), .ZN(n13137) );
  NAND2_X1 U12558 ( .A1(n14851), .A2(n15128), .ZN(n13043) );
  NAND2_X1 U12559 ( .A1(n10171), .A2(n9922), .ZN(n13771) );
  AND2_X1 U12560 ( .A1(n13475), .A2(n10143), .ZN(n13519) );
  INV_X1 U12561 ( .A(n10480), .ZN(n10477) );
  AOI21_X1 U12562 ( .B1(n16115), .B2(n18798), .A(n13227), .ZN(n13228) );
  NAND2_X1 U12563 ( .A1(n15605), .A2(n19719), .ZN(n19074) );
  OR2_X1 U12564 ( .A1(n19738), .A2(n19746), .ZN(n19464) );
  INV_X1 U12565 ( .A(n19744), .ZN(n19746) );
  OR2_X1 U12566 ( .A1(n19464), .A2(n19730), .ZN(n19506) );
  INV_X1 U12567 ( .A(n13143), .ZN(n19102) );
  NOR2_X1 U12568 ( .A1(n10918), .A2(n10917), .ZN(n13099) );
  NOR2_X1 U12569 ( .A1(n18111), .A2(n10918), .ZN(n12738) );
  OR2_X1 U12570 ( .A1(n16473), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n13110) );
  INV_X1 U12571 ( .A(n16766), .ZN(n16784) );
  OR2_X1 U12572 ( .A1(n10985), .A2(n17557), .ZN(n16300) );
  INV_X1 U12573 ( .A(n17615), .ZN(n17598) );
  NAND2_X1 U12574 ( .A1(n17520), .A2(n17759), .ZN(n17446) );
  INV_X1 U12575 ( .A(n17770), .ZN(n17416) );
  NAND2_X1 U12576 ( .A1(n9624), .A2(n10794), .ZN(n10795) );
  NOR2_X1 U12577 ( .A1(n17668), .A2(n17997), .ZN(n17667) );
  NAND2_X1 U12578 ( .A1(n17999), .A2(n9624), .ZN(n17669) );
  NOR2_X1 U12579 ( .A1(n17704), .A2(n17703), .ZN(n17702) );
  NOR2_X1 U12580 ( .A1(n17757), .A2(n17751), .ZN(n17750) );
  INV_X1 U12581 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18576) );
  AOI211_X2 U12582 ( .C1(n9592), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n10842), .B(n10841), .ZN(n18115) );
  NAND2_X1 U12583 ( .A1(n13439), .A2(n13534), .ZN(n20795) );
  NAND2_X1 U12584 ( .A1(n11498), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11514) );
  INV_X1 U12585 ( .A(n19877), .ZN(n15642) );
  OR2_X1 U12586 ( .A1(n20795), .A2(n13872), .ZN(n14417) );
  INV_X1 U12587 ( .A(n19839), .ZN(n19868) );
  AND2_X1 U12588 ( .A1(n13892), .A2(n13885), .ZN(n19860) );
  INV_X1 U12589 ( .A(n14470), .ZN(n19900) );
  NOR2_X1 U12590 ( .A1(n14518), .A2(n16338), .ZN(n13260) );
  OR2_X1 U12591 ( .A1(n13534), .A2(n13531), .ZN(n13725) );
  NAND2_X1 U12592 ( .A1(n11646), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11669) );
  NAND2_X1 U12593 ( .A1(n11564), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11598) );
  NAND2_X1 U12594 ( .A1(n11425), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11463) );
  INV_X1 U12595 ( .A(n14636), .ZN(n19941) );
  AND3_X1 U12596 ( .A1(n12777), .A2(n12776), .A3(n13601), .ZN(n19948) );
  INV_X1 U12597 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12654) );
  INV_X1 U12598 ( .A(n19983), .ZN(n19967) );
  AND2_X1 U12599 ( .A1(n12577), .A2(n13842), .ZN(n20121) );
  AND2_X1 U12600 ( .A1(n20121), .A2(n20445), .ZN(n20191) );
  INV_X1 U12601 ( .A(n20283), .ZN(n20286) );
  INV_X1 U12602 ( .A(n20335), .ZN(n20348) );
  INV_X1 U12603 ( .A(n20476), .ZN(n20319) );
  INV_X1 U12604 ( .A(n20427), .ZN(n20420) );
  NOR2_X1 U12605 ( .A1(n12577), .A2(n12555), .ZN(n20446) );
  INV_X1 U12606 ( .A(n20477), .ZN(n20514) );
  INV_X1 U12607 ( .A(n20609), .ZN(n20599) );
  INV_X1 U12608 ( .A(n20395), .ZN(n20617) );
  INV_X1 U12609 ( .A(n20414), .ZN(n20652) );
  INV_X1 U12610 ( .A(n20418), .ZN(n20659) );
  INV_X1 U12611 ( .A(n20666), .ZN(n20681) );
  OR2_X1 U12612 ( .A1(n16259), .A2(n19789), .ZN(n13322) );
  NAND2_X1 U12613 ( .A1(n13075), .A2(n13079), .ZN(n13080) );
  INV_X1 U12614 ( .A(n9691), .ZN(n18921) );
  AND2_X1 U12615 ( .A1(n12355), .A2(n12354), .ZN(n14151) );
  OAI21_X1 U12616 ( .B1(n10646), .B2(n14932), .A(n10645), .ZN(n10647) );
  AND2_X1 U12617 ( .A1(n14938), .A2(n14937), .ZN(n14935) );
  INV_X1 U12618 ( .A(n18978), .ZN(n18998) );
  AND2_X1 U12619 ( .A1(n13424), .A2(n19772), .ZN(n19003) );
  AND2_X1 U12620 ( .A1(n16124), .A2(n13400), .ZN(n16115) );
  INV_X1 U12621 ( .A(n15331), .ZN(n16046) );
  NAND2_X1 U12622 ( .A1(n13158), .A2(n19633), .ZN(n13213) );
  OR2_X1 U12623 ( .A1(n15304), .A2(n13191), .ZN(n15390) );
  INV_X1 U12624 ( .A(n19158), .ZN(n19576) );
  NAND2_X1 U12625 ( .A1(n16263), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19719) );
  OAI21_X1 U12626 ( .B1(n19086), .B2(n19085), .A(n19084), .ZN(n19121) );
  AND2_X1 U12627 ( .A1(n19129), .A2(n19127), .ZN(n19148) );
  NAND2_X1 U12628 ( .A1(n19780), .A2(n19074), .ZN(n19158) );
  INV_X1 U12629 ( .A(n19248), .ZN(n19218) );
  INV_X1 U12630 ( .A(n19278), .ZN(n19271) );
  AND2_X1 U12631 ( .A1(n19249), .A2(n19730), .ZN(n19307) );
  INV_X1 U12632 ( .A(n19366), .ZN(n19331) );
  OAI21_X1 U12633 ( .B1(n19361), .B2(n19341), .A(n19576), .ZN(n19363) );
  INV_X1 U12634 ( .A(n19386), .ZN(n19393) );
  NOR2_X1 U12635 ( .A1(n19368), .A2(n19752), .ZN(n19428) );
  OAI211_X1 U12636 ( .C1(n19498), .C2(n19469), .A(n19468), .B(n19576), .ZN(
        n19501) );
  OAI21_X1 U12637 ( .B1(n19547), .B2(n19546), .A(n19545), .ZN(n19564) );
  NAND2_X1 U12638 ( .A1(n18558), .A2(n13099), .ZN(n18532) );
  NAND2_X2 U12639 ( .A1(n17332), .A2(n17811), .ZN(n18539) );
  INV_X1 U12640 ( .A(n16793), .ZN(n16786) );
  NOR2_X1 U12641 ( .A1(n18596), .A2(n13103), .ZN(n16766) );
  NAND4_X1 U12642 ( .A1(n9600), .A2(n18755), .A3(n18610), .A4(n18601), .ZN(
        n16795) );
  AND2_X1 U12643 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16916), .ZN(n16901) );
  NOR2_X1 U12644 ( .A1(n17259), .A2(n16931), .ZN(n16916) );
  AND2_X1 U12645 ( .A1(n15493), .A2(n17107), .ZN(n17081) );
  NOR2_X1 U12646 ( .A1(n17134), .A2(n17117), .ZN(n17111) );
  NOR2_X1 U12647 ( .A1(n17340), .A2(n17206), .ZN(n17201) );
  OAI211_X1 U12648 ( .C1(n17087), .C2(n16888), .A(n10758), .B(n10757), .ZN(
        n17267) );
  INV_X1 U12649 ( .A(n17329), .ZN(n17293) );
  OAI211_X1 U12650 ( .C1(n16821), .C2(n20927), .A(n10782), .B(n10781), .ZN(
        n15517) );
  NOR2_X1 U12651 ( .A1(n10980), .A2(n17667), .ZN(n17965) );
  INV_X1 U12652 ( .A(n17446), .ZN(n17508) );
  NAND2_X1 U12653 ( .A1(n12764), .A2(n12763), .ZN(n12765) );
  NOR2_X2 U12654 ( .A1(n18767), .A2(n15488), .ZN(n18559) );
  INV_X1 U12655 ( .A(n18546), .ZN(n18574) );
  INV_X1 U12656 ( .A(n17332), .ZN(n18749) );
  OR2_X1 U12657 ( .A1(n13441), .A2(n19796), .ZN(n13439) );
  INV_X1 U12658 ( .A(n19847), .ZN(n14414) );
  INV_X1 U12659 ( .A(n19860), .ZN(n19893) );
  INV_X1 U12660 ( .A(n14468), .ZN(n19904) );
  INV_X1 U12661 ( .A(n19908), .ZN(n19938) );
  INV_X1 U12662 ( .A(n13725), .ZN(n13746) );
  INV_X1 U12663 ( .A(n15781), .ZN(n19953) );
  NAND2_X1 U12664 ( .A1(n12705), .A2(n12689), .ZN(n19977) );
  NAND2_X1 U12665 ( .A1(n20121), .A2(n20319), .ZN(n20077) );
  NAND2_X1 U12666 ( .A1(n20121), .A2(n20362), .ZN(n20115) );
  NAND2_X1 U12667 ( .A1(n20121), .A2(n20572), .ZN(n20151) );
  INV_X1 U12668 ( .A(n20191), .ZN(n20187) );
  NAND2_X1 U12669 ( .A1(n20286), .A2(n20319), .ZN(n20231) );
  NAND2_X1 U12670 ( .A1(n20286), .A2(n20362), .ZN(n20274) );
  NAND2_X1 U12671 ( .A1(n20286), .A2(n20572), .ZN(n20313) );
  NAND2_X1 U12672 ( .A1(n20286), .A2(n20445), .ZN(n20335) );
  NAND2_X1 U12673 ( .A1(n20446), .A2(n20572), .ZN(n20467) );
  NAND2_X1 U12674 ( .A1(n20529), .A2(n20528), .ZN(n20609) );
  NAND2_X1 U12675 ( .A1(n20573), .A2(n20445), .ZN(n20685) );
  INV_X1 U12676 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15944) );
  NOR2_X1 U12677 ( .A1(n13322), .A2(n13329), .ZN(n19786) );
  OR3_X1 U12678 ( .A1(n13078), .A2(n14277), .A3(n13077), .ZN(n18924) );
  INV_X1 U12679 ( .A(n10647), .ZN(n10648) );
  INV_X1 U12680 ( .A(n13608), .ZN(n14915) );
  AND2_X1 U12681 ( .A1(n13015), .A2(n13014), .ZN(n13016) );
  INV_X1 U12682 ( .A(n18995), .ZN(n18973) );
  AND2_X1 U12683 ( .A1(n16003), .A2(n13677), .ZN(n19002) );
  AOI21_X1 U12684 ( .B1(n16154), .B2(n19046), .A(n13229), .ZN(n13230) );
  INV_X1 U12685 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20875) );
  XNOR2_X1 U12686 ( .A(n15121), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16157) );
  OR2_X1 U12687 ( .A1(n13213), .A2(n19761), .ZN(n16191) );
  OR2_X1 U12688 ( .A1(n13213), .A2(n13161), .ZN(n19058) );
  INV_X1 U12689 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19757) );
  OR2_X1 U12690 ( .A1(n19132), .A2(n19507), .ZN(n19152) );
  AOI211_X2 U12691 ( .C1(n19160), .C2(n19159), .A(n19158), .B(n19157), .ZN(
        n19185) );
  OR2_X1 U12692 ( .A1(n19186), .A2(n19507), .ZN(n19216) );
  OR2_X1 U12693 ( .A1(n19186), .A2(n19752), .ZN(n19248) );
  INV_X1 U12694 ( .A(n19307), .ZN(n19285) );
  NAND2_X1 U12695 ( .A1(n19281), .A2(n19752), .ZN(n19335) );
  OR2_X1 U12696 ( .A1(n19731), .A2(n19752), .ZN(n19366) );
  NAND2_X1 U12697 ( .A1(n19428), .A2(n19744), .ZN(n19427) );
  INV_X1 U12698 ( .A(n19465), .ZN(n19504) );
  NAND2_X1 U12699 ( .A1(n19511), .A2(n19507), .ZN(n19535) );
  NAND2_X1 U12700 ( .A1(n19580), .A2(n19752), .ZN(n19568) );
  NAND2_X1 U12701 ( .A1(n19580), .A2(n19507), .ZN(n19631) );
  AOI21_X1 U12702 ( .B1(n18533), .B2(n18532), .A(n17330), .ZN(n18768) );
  NAND2_X1 U12703 ( .A1(n18593), .A2(n18757), .ZN(n16440) );
  INV_X1 U12704 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17626) );
  INV_X1 U12705 ( .A(n16794), .ZN(n16783) );
  INV_X1 U12706 ( .A(n16851), .ZN(n16864) );
  AND2_X1 U12707 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16865), .ZN(n16871) );
  INV_X1 U12708 ( .A(n17121), .ZN(n17114) );
  NAND2_X1 U12709 ( .A1(n17131), .A2(n17259), .ZN(n17121) );
  INV_X1 U12710 ( .A(n15517), .ZN(n17261) );
  INV_X1 U12711 ( .A(n17287), .ZN(n17270) );
  NAND2_X1 U12712 ( .A1(n15613), .A2(n17141), .ZN(n17290) );
  NAND2_X1 U12713 ( .A1(n17331), .A2(n17292), .ZN(n17329) );
  OR2_X1 U12714 ( .A1(n17565), .A2(n17846), .ZN(n17530) );
  NAND2_X1 U12715 ( .A1(n17752), .A2(n15517), .ZN(n17622) );
  NOR2_X1 U12716 ( .A1(n17615), .A2(n17508), .ZN(n17744) );
  INV_X1 U12717 ( .A(n17752), .ZN(n17763) );
  AOI21_X1 U12718 ( .B1(n12767), .B2(n12766), .A(n12765), .ZN(n12768) );
  INV_X1 U12719 ( .A(n18009), .ZN(n17960) );
  OAI21_X2 U12720 ( .B1(n12745), .B2(n12744), .A(n18757), .ZN(n18090) );
  OAI211_X1 U12721 ( .C1(n15194), .C2(n16109), .A(n12515), .B(n12514), .ZN(
        P2_U2985) );
  NAND2_X1 U12722 ( .A1(n13231), .A2(n13230), .ZN(P2_U2995) );
  INV_X1 U12723 ( .A(n13114), .ZN(P3_U2641) );
  AOI22_X1 U12724 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n9937) );
  AND2_X4 U12725 ( .A1(n14075), .A2(n9883), .ZN(n12790) );
  AND2_X4 U12726 ( .A1(n16236), .A2(n10085), .ZN(n10400) );
  AOI22_X1 U12727 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9936) );
  AND2_X4 U12728 ( .A1(n14074), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10183) );
  AOI22_X1 U12729 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n9935) );
  NAND4_X1 U12730 ( .A1(n9937), .A2(n9936), .A3(n9935), .A4(n9934), .ZN(n9938)
         );
  AOI22_X1 U12731 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n9942) );
  AOI22_X1 U12732 ( .A1(n12845), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n9940) );
  NAND4_X1 U12733 ( .A1(n9943), .A2(n9942), .A3(n9941), .A4(n9940), .ZN(n9944)
         );
  NAND2_X1 U12734 ( .A1(n9944), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9945) );
  AOI22_X1 U12735 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U12736 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n9949) );
  AOI22_X1 U12737 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n9948) );
  AOI22_X1 U12738 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n9947) );
  NAND4_X1 U12739 ( .A1(n9950), .A2(n9949), .A3(n9948), .A4(n9947), .ZN(n9951)
         );
  NAND2_X1 U12740 ( .A1(n9951), .A2(n10529), .ZN(n9958) );
  AOI22_X1 U12741 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U12742 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U12743 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n9953) );
  AOI22_X1 U12744 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n9952) );
  NAND4_X1 U12745 ( .A1(n9955), .A2(n9954), .A3(n9953), .A4(n9952), .ZN(n9956)
         );
  NAND2_X2 U12746 ( .A1(n9958), .A2(n9957), .ZN(n13012) );
  AOI22_X1 U12747 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10002), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U12748 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n9961) );
  AOI22_X1 U12749 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U12750 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U12751 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U12752 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n9966) );
  AOI22_X1 U12753 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n9965) );
  AOI22_X1 U12754 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n9964) );
  INV_X2 U12755 ( .A(n10048), .ZN(n13143) );
  AOI22_X1 U12756 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U12757 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n9972) );
  AOI22_X1 U12758 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n9971) );
  NAND4_X1 U12759 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n9974)
         );
  NAND2_X1 U12760 ( .A1(n9974), .A2(n10529), .ZN(n9982) );
  AND2_X1 U12761 ( .A1(n10001), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n9975) );
  AOI21_X1 U12762 ( .B1(n10183), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n9975), .ZN(n9979) );
  AOI22_X1 U12763 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U12764 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U12765 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n9976) );
  NAND4_X1 U12766 ( .A1(n9979), .A2(n9978), .A3(n9977), .A4(n9976), .ZN(n9980)
         );
  NAND2_X1 U12767 ( .A1(n9980), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9981) );
  NAND2_X4 U12768 ( .A1(n9982), .A2(n9981), .ZN(n13011) );
  NOR2_X1 U12769 ( .A1(n13143), .A2(n13011), .ZN(n9983) );
  AOI22_X1 U12770 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U12771 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U12772 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U12773 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9984) );
  NAND4_X1 U12774 ( .A1(n9987), .A2(n9986), .A3(n9985), .A4(n9984), .ZN(n9988)
         );
  AOI22_X1 U12775 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n9992) );
  AOI22_X1 U12776 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U12777 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n9990) );
  AOI22_X1 U12778 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9989) );
  NAND4_X1 U12779 ( .A1(n9992), .A2(n9991), .A3(n9990), .A4(n9989), .ZN(n9993)
         );
  AOI22_X1 U12780 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U12781 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n9999) );
  AOI22_X1 U12782 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n9998) );
  NAND4_X1 U12783 ( .A1(n10000), .A2(n9999), .A3(n9998), .A4(n9997), .ZN(
        n10008) );
  AOI22_X1 U12784 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10006) );
  AOI22_X1 U12785 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10005) );
  AOI22_X1 U12786 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10004) );
  NAND4_X1 U12787 ( .A1(n10006), .A2(n10005), .A3(n10004), .A4(n10003), .ZN(
        n10007) );
  MUX2_X2 U12788 ( .A(n10008), .B(n10007), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n16265) );
  NAND2_X1 U12789 ( .A1(n10092), .A2(n19076), .ZN(n10044) );
  AOI22_X1 U12790 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U12791 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10011) );
  AOI22_X1 U12792 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U12793 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10009) );
  NAND4_X1 U12794 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10013) );
  AOI22_X1 U12795 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10019) );
  AOI22_X1 U12796 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U12797 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9627), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U12798 ( .A1(n10002), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10014) );
  NAND4_X1 U12799 ( .A1(n10019), .A2(n10018), .A3(n10017), .A4(n10016), .ZN(
        n10020) );
  AOI22_X1 U12800 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U12801 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U12802 ( .A1(n10024), .A2(n10023), .ZN(n10029) );
  AOI22_X1 U12803 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U12804 ( .A1(n10002), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10026) );
  NAND3_X1 U12805 ( .A1(n10027), .A2(n10026), .A3(n10025), .ZN(n10028) );
  NOR2_X1 U12806 ( .A1(n10029), .A2(n10028), .ZN(n10030) );
  NAND2_X1 U12807 ( .A1(n10030), .A2(n10529), .ZN(n10038) );
  AOI22_X1 U12808 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10002), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10032) );
  AOI22_X1 U12809 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10400), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10031) );
  AOI22_X1 U12810 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10035) );
  AOI22_X1 U12811 ( .A1(n10183), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10034) );
  NAND4_X1 U12812 ( .A1(n13182), .A2(n10061), .A3(n10048), .A4(n13011), .ZN(
        n10039) );
  NOR2_X2 U12813 ( .A1(n10039), .A2(n10053), .ZN(n12449) );
  INV_X1 U12814 ( .A(n10039), .ZN(n10041) );
  NAND2_X1 U12815 ( .A1(n10553), .A2(n16265), .ZN(n10043) );
  NAND2_X1 U12816 ( .A1(n10044), .A2(n10043), .ZN(n10052) );
  MUX2_X1 U12817 ( .A(n13012), .B(n13011), .S(n13143), .Z(n10046) );
  AND2_X1 U12818 ( .A1(n10053), .A2(n10061), .ZN(n10045) );
  NAND2_X1 U12819 ( .A1(n10056), .A2(n13182), .ZN(n10069) );
  NAND3_X1 U12820 ( .A1(n10046), .A2(n10045), .A3(n10069), .ZN(n10051) );
  NAND4_X1 U12821 ( .A1(n10067), .A2(n10048), .A3(n10047), .A4(n13011), .ZN(
        n10049) );
  NOR2_X2 U12822 ( .A1(n10049), .A2(n10053), .ZN(n13469) );
  INV_X1 U12823 ( .A(n13469), .ZN(n10050) );
  NAND3_X1 U12824 ( .A1(n10051), .A2(n19076), .A3(n10050), .ZN(n13177) );
  AND2_X2 U12825 ( .A1(n10052), .A2(n13177), .ZN(n10096) );
  NAND2_X1 U12826 ( .A1(n10054), .A2(n10053), .ZN(n12862) );
  INV_X1 U12827 ( .A(n12862), .ZN(n10055) );
  NAND2_X1 U12828 ( .A1(n10055), .A2(n19102), .ZN(n12860) );
  NAND2_X1 U12829 ( .A1(n10056), .A2(n13143), .ZN(n12858) );
  AND2_X1 U12830 ( .A1(n12858), .A2(n13011), .ZN(n10057) );
  NAND2_X1 U12831 ( .A1(n13180), .A2(n13182), .ZN(n10059) );
  NAND2_X1 U12832 ( .A1(n10059), .A2(n10058), .ZN(n10094) );
  INV_X2 U12833 ( .A(n12144), .ZN(n10075) );
  NAND2_X1 U12834 ( .A1(n10094), .A2(n10075), .ZN(n10060) );
  NAND2_X1 U12835 ( .A1(n10096), .A2(n10060), .ZN(n10084) );
  AND2_X2 U12836 ( .A1(n10061), .A2(n10067), .ZN(n13175) );
  NAND2_X1 U12837 ( .A1(n12872), .A2(n10063), .ZN(n10064) );
  NOR2_X1 U12838 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U12839 ( .A1(n12883), .A2(n9996), .ZN(n10068) );
  NAND2_X1 U12840 ( .A1(n10068), .A2(n10067), .ZN(n10070) );
  NAND2_X1 U12841 ( .A1(n10070), .A2(n10069), .ZN(n10073) );
  NOR2_X2 U12842 ( .A1(n10073), .A2(n10072), .ZN(n10552) );
  NAND2_X1 U12843 ( .A1(n10153), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10080) );
  AND2_X2 U12844 ( .A1(n13175), .A2(n10075), .ZN(n10087) );
  AND2_X2 U12845 ( .A1(n10087), .A2(n9613), .ZN(n13186) );
  AND2_X4 U12846 ( .A1(n13186), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U12847 ( .A1(n10621), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10078) );
  AOI22_X1 U12848 ( .A1(n10098), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10077) );
  INV_X1 U12849 ( .A(n13186), .ZN(n16224) );
  AOI21_X1 U12850 ( .B1(n16224), .B2(n10085), .A(n19780), .ZN(n10086) );
  OAI21_X1 U12851 ( .B1(n9611), .B2(n10087), .A(n10086), .ZN(n10091) );
  NAND2_X1 U12852 ( .A1(n10099), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10088) );
  NAND2_X1 U12853 ( .A1(n10091), .A2(n10090), .ZN(n10126) );
  INV_X1 U12854 ( .A(n10092), .ZN(n10093) );
  NAND2_X1 U12855 ( .A1(n10094), .A2(n10093), .ZN(n10095) );
  NAND2_X1 U12856 ( .A1(n10096), .A2(n10095), .ZN(n10097) );
  NAND2_X1 U12857 ( .A1(n10097), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10105) );
  INV_X1 U12858 ( .A(n10099), .ZN(n10151) );
  NAND2_X1 U12859 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U12860 ( .A1(n10151), .A2(n10100), .ZN(n10101) );
  AOI21_X1 U12861 ( .B1(n10098), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10101), .ZN(
        n10104) );
  NAND2_X1 U12862 ( .A1(n10153), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10103) );
  NAND2_X1 U12863 ( .A1(n10621), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10102) );
  NAND4_X1 U12864 ( .A1(n10105), .A2(n10104), .A3(n10103), .A4(n10102), .ZN(
        n10127) );
  AOI21_X1 U12865 ( .B1(n19780), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U12866 ( .A1(n10621), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U12867 ( .A1(n10098), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10109) );
  NAND2_X1 U12868 ( .A1(n10153), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10108) );
  NAND3_X1 U12869 ( .A1(n10110), .A2(n10109), .A3(n10108), .ZN(n10111) );
  NAND2_X1 U12870 ( .A1(n10112), .A2(n10111), .ZN(n10113) );
  INV_X1 U12871 ( .A(n10114), .ZN(n10117) );
  INV_X1 U12872 ( .A(n10115), .ZN(n10116) );
  NAND2_X1 U12873 ( .A1(n19780), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15603) );
  INV_X1 U12874 ( .A(n15603), .ZN(n10158) );
  NAND2_X1 U12875 ( .A1(n11973), .A2(n10158), .ZN(n10124) );
  NAND2_X1 U12876 ( .A1(n13012), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U12877 ( .A1(n10120), .A2(n20926), .ZN(n10162) );
  NAND2_X1 U12878 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19429) );
  NAND2_X1 U12879 ( .A1(n19429), .A2(n19742), .ZN(n10121) );
  NAND2_X1 U12880 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19536) );
  INV_X1 U12881 ( .A(n19536), .ZN(n19571) );
  AND2_X1 U12882 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19571), .ZN(
        n10159) );
  INV_X1 U12883 ( .A(n10159), .ZN(n10160) );
  NAND2_X1 U12884 ( .A1(n10121), .A2(n10160), .ZN(n19220) );
  INV_X1 U12885 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19784) );
  NAND2_X1 U12886 ( .A1(n19784), .A2(n20926), .ZN(n19539) );
  NOR2_X1 U12887 ( .A1(n19220), .A2(n19539), .ZN(n10122) );
  AOI21_X1 U12888 ( .B1(n10162), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10122), .ZN(n10123) );
  NOR2_X1 U12889 ( .A1(n13012), .A2(n19780), .ZN(n10125) );
  INV_X1 U12890 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12098) );
  OR2_X1 U12891 ( .A1(n10127), .A2(n10126), .ZN(n10128) );
  NOR2_X1 U12892 ( .A1(n19539), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10129) );
  AOI21_X1 U12893 ( .B1(n10162), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10129), .ZN(n10130) );
  INV_X1 U12894 ( .A(n10517), .ZN(n10475) );
  XNOR2_X1 U12895 ( .A(n10139), .B(n10140), .ZN(n13472) );
  INV_X1 U12896 ( .A(n10134), .ZN(n10135) );
  NAND2_X1 U12897 ( .A1(n11967), .A2(n10135), .ZN(n10136) );
  XNOR2_X1 U12898 ( .A(n19751), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19221) );
  INV_X1 U12899 ( .A(n19539), .ZN(n19724) );
  NAND2_X1 U12900 ( .A1(n19221), .A2(n19724), .ZN(n19401) );
  INV_X1 U12901 ( .A(n19401), .ZN(n10137) );
  AOI21_X1 U12902 ( .B1(n10162), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10137), .ZN(n10138) );
  INV_X1 U12903 ( .A(n10139), .ZN(n10142) );
  INV_X1 U12904 ( .A(n10140), .ZN(n10141) );
  NAND2_X1 U12905 ( .A1(n10142), .A2(n10141), .ZN(n10143) );
  NAND2_X1 U12906 ( .A1(n13520), .A2(n13519), .ZN(n10148) );
  INV_X1 U12907 ( .A(n10144), .ZN(n10145) );
  NAND2_X1 U12908 ( .A1(n10146), .A2(n10145), .ZN(n10147) );
  INV_X1 U12909 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12137) );
  NAND2_X1 U12910 ( .A1(n10098), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U12911 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10155) );
  OAI211_X1 U12912 ( .C1(n13207), .C2(n12137), .A(n10156), .B(n10155), .ZN(
        n10157) );
  NAND2_X1 U12913 ( .A1(n11974), .A2(n10158), .ZN(n10164) );
  NAND2_X1 U12914 ( .A1(n10159), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19569) );
  NAND2_X1 U12915 ( .A1(n19734), .A2(n10160), .ZN(n10161) );
  AND3_X1 U12916 ( .A1(n19724), .A2(n19569), .A3(n10161), .ZN(n19459) );
  AOI21_X1 U12917 ( .B1(n10162), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19459), .ZN(n10163) );
  INV_X1 U12918 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U12919 ( .A1(n13616), .A2(n13615), .ZN(n10170) );
  INV_X1 U12920 ( .A(n10165), .ZN(n10167) );
  AND2_X1 U12921 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13012), .ZN(
        n10166) );
  AOI21_X1 U12922 ( .B1(n10168), .B2(n10167), .A(n10166), .ZN(n10169) );
  INV_X1 U12923 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10237) );
  NOR2_X1 U12924 ( .A1(n10517), .A2(n10237), .ZN(n13605) );
  INV_X1 U12925 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12216) );
  AND2_X2 U12926 ( .A1(n14075), .A2(n10401), .ZN(n12250) );
  AOI22_X1 U12927 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10176) );
  AND2_X2 U12928 ( .A1(n14074), .A2(n10401), .ZN(n12252) );
  AOI22_X1 U12929 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U12930 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10174) );
  NAND2_X1 U12931 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10173) );
  NAND4_X1 U12932 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10178) );
  INV_X1 U12933 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10390) );
  INV_X1 U12934 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10391) );
  OAI22_X1 U12935 ( .A1(n12260), .A2(n10390), .B1(n12258), .B2(n10391), .ZN(
        n10177) );
  NOR2_X1 U12936 ( .A1(n10178), .A2(n10177), .ZN(n10191) );
  INV_X1 U12937 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10385) );
  OR2_X2 U12938 ( .A1(n10179), .A2(n10529), .ZN(n12264) );
  INV_X1 U12939 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10379) );
  OAI22_X1 U12940 ( .A1(n12008), .A2(n10385), .B1(n12264), .B2(n10379), .ZN(
        n10182) );
  INV_X1 U12941 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10180) );
  INV_X1 U12942 ( .A(n9601), .ZN(n12810) );
  INV_X1 U12943 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10383) );
  OAI22_X1 U12944 ( .A1(n12268), .A2(n10180), .B1(n12266), .B2(n10383), .ZN(
        n10181) );
  NOR2_X1 U12945 ( .A1(n10182), .A2(n10181), .ZN(n10190) );
  INV_X1 U12946 ( .A(n10183), .ZN(n12795) );
  INV_X1 U12947 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10186) );
  INV_X1 U12948 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10384) );
  OAI22_X1 U12949 ( .A1(n12170), .A2(n10186), .B1(n12272), .B2(n10384), .ZN(
        n10188) );
  NAND2_X1 U12950 ( .A1(n16235), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12012) );
  INV_X1 U12951 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10380) );
  INV_X1 U12952 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10386) );
  OAI22_X1 U12953 ( .A1(n12275), .A2(n10380), .B1(n12017), .B2(n10386), .ZN(
        n10187) );
  NOR2_X1 U12954 ( .A1(n10188), .A2(n10187), .ZN(n10189) );
  AND3_X1 U12955 ( .A1(n10191), .A2(n10190), .A3(n10189), .ZN(n12930) );
  AOI22_X1 U12956 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U12957 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U12958 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10194) );
  NAND2_X1 U12959 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10193) );
  NAND4_X1 U12960 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10198) );
  INV_X1 U12961 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12026) );
  INV_X1 U12962 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12064) );
  OAI22_X1 U12963 ( .A1(n12026), .A2(n12275), .B1(n12017), .B2(n12064), .ZN(
        n10197) );
  NOR2_X1 U12964 ( .A1(n10198), .A2(n10197), .ZN(n10205) );
  INV_X1 U12965 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12074) );
  INV_X1 U12966 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12070) );
  OAI22_X1 U12967 ( .A1(n12008), .A2(n12074), .B1(n12264), .B2(n12070), .ZN(
        n10200) );
  INV_X1 U12968 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12065) );
  INV_X1 U12969 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12069) );
  OAI22_X1 U12970 ( .A1(n12170), .A2(n12065), .B1(n12266), .B2(n12069), .ZN(
        n10199) );
  NOR2_X1 U12971 ( .A1(n10200), .A2(n10199), .ZN(n10204) );
  INV_X1 U12972 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12076) );
  INV_X1 U12973 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10366) );
  OAI22_X1 U12974 ( .A1(n12268), .A2(n12076), .B1(n12272), .B2(n10366), .ZN(
        n10202) );
  INV_X1 U12975 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20816) );
  INV_X1 U12976 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12068) );
  OAI22_X1 U12977 ( .A1(n20816), .A2(n12260), .B1(n12258), .B2(n12068), .ZN(
        n10201) );
  NOR2_X1 U12978 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NAND3_X1 U12979 ( .A1(n10205), .A2(n10204), .A3(n10203), .ZN(n13799) );
  AOI22_X1 U12980 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U12981 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U12982 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10207) );
  NAND2_X1 U12983 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10206) );
  NAND4_X1 U12984 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10211) );
  INV_X1 U12985 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12093) );
  OAI22_X1 U12986 ( .A1(n12098), .A2(n12260), .B1(n12258), .B2(n12093), .ZN(
        n10210) );
  NOR2_X1 U12987 ( .A1(n10211), .A2(n10210), .ZN(n10218) );
  INV_X1 U12988 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12092) );
  INV_X1 U12989 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12090) );
  OAI22_X1 U12990 ( .A1(n12008), .A2(n12092), .B1(n12264), .B2(n12090), .ZN(
        n10213) );
  INV_X1 U12991 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12099) );
  INV_X1 U12992 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12097) );
  OAI22_X1 U12993 ( .A1(n12268), .A2(n12099), .B1(n12266), .B2(n12097), .ZN(
        n10212) );
  NOR2_X1 U12994 ( .A1(n10213), .A2(n10212), .ZN(n10217) );
  INV_X1 U12995 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12088) );
  INV_X1 U12996 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10350) );
  OAI22_X1 U12997 ( .A1(n12170), .A2(n12088), .B1(n12272), .B2(n10350), .ZN(
        n10215) );
  INV_X1 U12998 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10347) );
  INV_X1 U12999 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12087) );
  OAI22_X1 U13000 ( .A1(n10347), .A2(n12275), .B1(n12017), .B2(n12087), .ZN(
        n10214) );
  NOR2_X1 U13001 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  AOI22_X1 U13002 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U13003 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U13004 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10221) );
  NAND2_X1 U13005 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10220) );
  NAND4_X1 U13006 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10225) );
  INV_X1 U13007 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11968) );
  INV_X1 U13008 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11975) );
  OAI22_X1 U13009 ( .A1(n11968), .A2(n12258), .B1(n12017), .B2(n11975), .ZN(
        n10224) );
  NOR2_X1 U13010 ( .A1(n10225), .A2(n10224), .ZN(n10232) );
  INV_X1 U13011 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12009) );
  INV_X1 U13012 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11986) );
  OAI22_X1 U13013 ( .A1(n12008), .A2(n12009), .B1(n12264), .B2(n11986), .ZN(
        n10227) );
  INV_X1 U13014 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20841) );
  INV_X1 U13015 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11979) );
  OAI22_X1 U13016 ( .A1(n12170), .A2(n20841), .B1(n12272), .B2(n11979), .ZN(
        n10226) );
  NOR2_X1 U13017 ( .A1(n10227), .A2(n10226), .ZN(n10231) );
  INV_X1 U13018 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11970) );
  INV_X1 U13019 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11984) );
  OAI22_X1 U13020 ( .A1(n12268), .A2(n11970), .B1(n12266), .B2(n11984), .ZN(
        n10229) );
  INV_X1 U13021 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11976) );
  OAI22_X1 U13022 ( .A1(n11976), .A2(n12275), .B1(n12260), .B2(n11999), .ZN(
        n10228) );
  NOR2_X1 U13023 ( .A1(n10229), .A2(n10228), .ZN(n10230) );
  AND3_X1 U13024 ( .A1(n10232), .A2(n10231), .A3(n10230), .ZN(n13912) );
  AOI22_X1 U13025 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13026 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10235) );
  NAND2_X1 U13027 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10234) );
  NAND2_X1 U13028 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10233) );
  NAND4_X1 U13029 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10239) );
  INV_X1 U13030 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12162) );
  OAI22_X1 U13031 ( .A1(n10237), .A2(n12260), .B1(n12258), .B2(n12162), .ZN(
        n10238) );
  NOR2_X1 U13032 ( .A1(n10239), .A2(n10238), .ZN(n10246) );
  INV_X1 U13033 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12168) );
  INV_X1 U13034 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12164) );
  OAI22_X1 U13035 ( .A1(n12008), .A2(n12168), .B1(n12264), .B2(n12164), .ZN(
        n10241) );
  INV_X1 U13036 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12171) );
  INV_X1 U13037 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12163) );
  OAI22_X1 U13038 ( .A1(n12268), .A2(n12171), .B1(n12266), .B2(n12163), .ZN(
        n10240) );
  NOR2_X1 U13039 ( .A1(n10241), .A2(n10240), .ZN(n10245) );
  INV_X1 U13040 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12159) );
  INV_X1 U13041 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10321) );
  OAI22_X1 U13042 ( .A1(n12170), .A2(n12159), .B1(n12272), .B2(n10321), .ZN(
        n10243) );
  INV_X1 U13043 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10318) );
  INV_X1 U13044 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12158) );
  OAI22_X1 U13045 ( .A1(n10318), .A2(n12275), .B1(n12017), .B2(n12158), .ZN(
        n10242) );
  NOR2_X1 U13046 ( .A1(n10243), .A2(n10242), .ZN(n10244) );
  INV_X1 U13047 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12806) );
  OAI22_X1 U13048 ( .A1(n12008), .A2(n12806), .B1(n12268), .B2(n9699), .ZN(
        n10248) );
  INV_X1 U13049 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12213) );
  INV_X1 U13050 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12805) );
  OAI22_X1 U13051 ( .A1(n12264), .A2(n12213), .B1(n12266), .B2(n12805), .ZN(
        n10247) );
  NOR2_X1 U13052 ( .A1(n10248), .A2(n10247), .ZN(n10259) );
  AOI22_X1 U13053 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U13054 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10251) );
  NAND2_X1 U13055 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10250) );
  NAND2_X1 U13056 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10249) );
  NAND4_X1 U13057 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10254) );
  INV_X1 U13058 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12212) );
  INV_X1 U13059 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12209) );
  OAI22_X1 U13060 ( .A1(n12258), .A2(n12212), .B1(n12017), .B2(n12209), .ZN(
        n10253) );
  NOR2_X1 U13061 ( .A1(n10254), .A2(n10253), .ZN(n10258) );
  INV_X1 U13062 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12811) );
  INV_X1 U13063 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12809) );
  OAI22_X1 U13064 ( .A1(n12170), .A2(n12811), .B1(n12272), .B2(n12809), .ZN(
        n10256) );
  INV_X1 U13065 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12794) );
  OAI22_X1 U13066 ( .A1(n12260), .A2(n12216), .B1(n12275), .B2(n12794), .ZN(
        n10255) );
  NOR2_X1 U13067 ( .A1(n10256), .A2(n10255), .ZN(n10257) );
  NAND3_X1 U13068 ( .A1(n10259), .A2(n10258), .A3(n10257), .ZN(n14040) );
  AOI22_X1 U13069 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U13070 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U13071 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10261) );
  NAND2_X1 U13072 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10260) );
  NAND4_X1 U13073 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10265) );
  INV_X1 U13074 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13770) );
  INV_X1 U13075 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12263) );
  OAI22_X1 U13076 ( .A1(n12260), .A2(n13770), .B1(n12258), .B2(n12263), .ZN(
        n10264) );
  NOR2_X1 U13077 ( .A1(n10265), .A2(n10264), .ZN(n10272) );
  INV_X1 U13078 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12271) );
  INV_X1 U13079 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12265) );
  OAI22_X1 U13080 ( .A1(n12008), .A2(n12271), .B1(n12264), .B2(n12265), .ZN(
        n10267) );
  INV_X1 U13081 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12274) );
  INV_X1 U13082 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12823) );
  OAI22_X1 U13083 ( .A1(n12268), .A2(n12274), .B1(n12266), .B2(n12823), .ZN(
        n10266) );
  NOR2_X1 U13084 ( .A1(n10267), .A2(n10266), .ZN(n10271) );
  INV_X1 U13085 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12259) );
  INV_X1 U13086 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12242) );
  OAI22_X1 U13087 ( .A1(n12170), .A2(n12259), .B1(n12272), .B2(n12242), .ZN(
        n10269) );
  INV_X1 U13088 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12241) );
  INV_X1 U13089 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12257) );
  OAI22_X1 U13090 ( .A1(n12275), .A2(n12241), .B1(n12017), .B2(n12257), .ZN(
        n10268) );
  NOR2_X1 U13091 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  AND3_X1 U13092 ( .A1(n10272), .A2(n10271), .A3(n10270), .ZN(n12952) );
  INV_X1 U13093 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12114) );
  INV_X1 U13094 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10273) );
  OAI22_X1 U13095 ( .A1(n12114), .A2(n12268), .B1(n12170), .B2(n10273), .ZN(
        n10275) );
  INV_X1 U13096 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10424) );
  INV_X1 U13097 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12115) );
  OAI22_X1 U13098 ( .A1(n10424), .A2(n12275), .B1(n12017), .B2(n12115), .ZN(
        n10274) );
  NOR2_X1 U13099 ( .A1(n10275), .A2(n10274), .ZN(n10287) );
  AOI22_X1 U13100 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13101 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U13102 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10278) );
  NAND2_X1 U13103 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10277) );
  NAND4_X1 U13104 ( .A1(n10280), .A2(n10279), .A3(n10278), .A4(n10277), .ZN(
        n10282) );
  INV_X1 U13105 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10421) );
  INV_X1 U13106 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12118) );
  OAI22_X1 U13107 ( .A1(n12260), .A2(n10421), .B1(n12258), .B2(n12118), .ZN(
        n10281) );
  NOR2_X1 U13108 ( .A1(n10282), .A2(n10281), .ZN(n10286) );
  INV_X1 U13109 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12120) );
  INV_X1 U13110 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n20853) );
  OAI22_X1 U13111 ( .A1(n12008), .A2(n12120), .B1(n12264), .B2(n20853), .ZN(
        n10284) );
  INV_X1 U13112 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12119) );
  INV_X1 U13113 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10417) );
  OAI22_X1 U13114 ( .A1(n12119), .A2(n12266), .B1(n12272), .B2(n10417), .ZN(
        n10283) );
  NOR2_X1 U13115 ( .A1(n10284), .A2(n10283), .ZN(n10285) );
  AND3_X1 U13116 ( .A1(n10287), .A2(n10286), .A3(n10285), .ZN(n14173) );
  AOI22_X1 U13117 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13118 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U13119 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10289) );
  NAND2_X1 U13120 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10288) );
  NAND4_X1 U13121 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10293) );
  OAI22_X1 U13122 ( .A1(n12260), .A2(n12241), .B1(n12258), .B2(n12265), .ZN(
        n10292) );
  NOR2_X1 U13123 ( .A1(n10293), .A2(n10292), .ZN(n10300) );
  OAI22_X1 U13124 ( .A1(n12008), .A2(n12242), .B1(n12264), .B2(n12823), .ZN(
        n10295) );
  OAI22_X1 U13125 ( .A1(n12268), .A2(n12257), .B1(n12266), .B2(n12271), .ZN(
        n10294) );
  NOR2_X1 U13126 ( .A1(n10295), .A2(n10294), .ZN(n10299) );
  INV_X1 U13127 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12273) );
  OAI22_X1 U13128 ( .A1(n12170), .A2(n13770), .B1(n12272), .B2(n12273), .ZN(
        n10297) );
  INV_X1 U13129 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n19178) );
  OAI22_X1 U13130 ( .A1(n19178), .A2(n12275), .B1(n12017), .B2(n12263), .ZN(
        n10296) );
  NOR2_X1 U13131 ( .A1(n10297), .A2(n10296), .ZN(n10298) );
  NAND3_X1 U13132 ( .A1(n10300), .A2(n10299), .A3(n10298), .ZN(n14905) );
  AOI22_X1 U13133 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13134 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U13135 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U13136 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10301) );
  NAND4_X1 U13137 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10306) );
  OAI22_X1 U13138 ( .A1(n12260), .A2(n12794), .B1(n12258), .B2(n12213), .ZN(
        n10305) );
  NOR2_X1 U13139 ( .A1(n10306), .A2(n10305), .ZN(n10313) );
  OAI22_X1 U13140 ( .A1(n12008), .A2(n12809), .B1(n12264), .B2(n12805), .ZN(
        n10308) );
  OAI22_X1 U13141 ( .A1(n12268), .A2(n12209), .B1(n12266), .B2(n12806), .ZN(
        n10307) );
  NOR2_X1 U13142 ( .A1(n10308), .A2(n10307), .ZN(n10312) );
  INV_X1 U13143 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12807) );
  OAI22_X1 U13144 ( .A1(n12170), .A2(n12216), .B1(n12272), .B2(n12807), .ZN(
        n10310) );
  INV_X1 U13145 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12192) );
  OAI22_X1 U13146 ( .A1(n12275), .A2(n12192), .B1(n12017), .B2(n12212), .ZN(
        n10309) );
  NOR2_X1 U13147 ( .A1(n10310), .A2(n10309), .ZN(n10311) );
  NAND3_X1 U13148 ( .A1(n10313), .A2(n10312), .A3(n10311), .ZN(n14914) );
  AOI22_X1 U13149 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13150 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10316) );
  NAND2_X1 U13151 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10315) );
  NAND2_X1 U13152 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10314) );
  NAND4_X1 U13153 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10320) );
  OAI22_X1 U13154 ( .A1(n10318), .A2(n12260), .B1(n12258), .B2(n12164), .ZN(
        n10319) );
  NOR2_X1 U13155 ( .A1(n10320), .A2(n10319), .ZN(n10329) );
  OAI22_X1 U13156 ( .A1(n12008), .A2(n10321), .B1(n12264), .B2(n12163), .ZN(
        n10323) );
  OAI22_X1 U13157 ( .A1(n12268), .A2(n12158), .B1(n12266), .B2(n12168), .ZN(
        n10322) );
  NOR2_X1 U13158 ( .A1(n10323), .A2(n10322), .ZN(n10328) );
  INV_X1 U13159 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12169) );
  OAI22_X1 U13160 ( .A1(n12170), .A2(n10237), .B1(n12272), .B2(n12169), .ZN(
        n10326) );
  INV_X1 U13161 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10324) );
  OAI22_X1 U13162 ( .A1(n10324), .A2(n12275), .B1(n12017), .B2(n12162), .ZN(
        n10325) );
  NOR2_X1 U13163 ( .A1(n10326), .A2(n10325), .ZN(n10327) );
  AND3_X1 U13164 ( .A1(n10329), .A2(n10328), .A3(n10327), .ZN(n14919) );
  AOI22_X1 U13165 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13166 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10332) );
  NAND2_X1 U13167 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10331) );
  NAND2_X1 U13168 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10330) );
  NAND4_X1 U13169 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10335) );
  OAI22_X1 U13170 ( .A1(n11976), .A2(n12260), .B1(n12258), .B2(n11986), .ZN(
        n10334) );
  NOR2_X1 U13171 ( .A1(n10335), .A2(n10334), .ZN(n10342) );
  OAI22_X1 U13172 ( .A1(n12008), .A2(n11979), .B1(n12264), .B2(n11984), .ZN(
        n10337) );
  OAI22_X1 U13173 ( .A1(n12268), .A2(n11975), .B1(n12266), .B2(n12009), .ZN(
        n10336) );
  NOR2_X1 U13174 ( .A1(n10337), .A2(n10336), .ZN(n10341) );
  INV_X1 U13175 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12010) );
  OAI22_X1 U13176 ( .A1(n12170), .A2(n11999), .B1(n12272), .B2(n12010), .ZN(
        n10339) );
  INV_X1 U13177 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12000) );
  OAI22_X1 U13178 ( .A1(n12000), .A2(n12275), .B1(n12017), .B2(n11968), .ZN(
        n10338) );
  NOR2_X1 U13179 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  AND3_X1 U13180 ( .A1(n10342), .A2(n10341), .A3(n10340), .ZN(n14923) );
  NOR2_X1 U13181 ( .A1(n14919), .A2(n14923), .ZN(n10359) );
  AOI22_X1 U13182 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13183 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U13184 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10344) );
  NAND2_X1 U13185 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10343) );
  NAND4_X1 U13186 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10349) );
  OAI22_X1 U13187 ( .A1(n10347), .A2(n12260), .B1(n12258), .B2(n12090), .ZN(
        n10348) );
  NOR2_X1 U13188 ( .A1(n10349), .A2(n10348), .ZN(n10358) );
  OAI22_X1 U13189 ( .A1(n12008), .A2(n10350), .B1(n12264), .B2(n12097), .ZN(
        n10352) );
  OAI22_X1 U13190 ( .A1(n12268), .A2(n12087), .B1(n12266), .B2(n12092), .ZN(
        n10351) );
  NOR2_X1 U13191 ( .A1(n10352), .A2(n10351), .ZN(n10357) );
  INV_X1 U13192 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12096) );
  OAI22_X1 U13193 ( .A1(n12170), .A2(n12098), .B1(n12272), .B2(n12096), .ZN(
        n10355) );
  INV_X1 U13194 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10353) );
  OAI22_X1 U13195 ( .A1(n10353), .A2(n12275), .B1(n12017), .B2(n12093), .ZN(
        n10354) );
  NOR2_X1 U13196 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  NAND3_X1 U13197 ( .A1(n10358), .A2(n10357), .A3(n10356), .ZN(n14930) );
  AND2_X1 U13198 ( .A1(n10359), .A2(n14930), .ZN(n14911) );
  AND2_X1 U13199 ( .A1(n14914), .A2(n14911), .ZN(n14904) );
  AND2_X1 U13200 ( .A1(n14905), .A2(n14904), .ZN(n10374) );
  AOI22_X1 U13201 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13202 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U13203 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10361) );
  NAND2_X1 U13204 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10360) );
  NAND4_X1 U13205 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10365) );
  OAI22_X1 U13206 ( .A1(n12026), .A2(n12260), .B1(n12258), .B2(n12070), .ZN(
        n10364) );
  NOR2_X1 U13207 ( .A1(n10365), .A2(n10364), .ZN(n10373) );
  OAI22_X1 U13208 ( .A1(n12008), .A2(n10366), .B1(n12264), .B2(n12069), .ZN(
        n10368) );
  OAI22_X1 U13209 ( .A1(n12268), .A2(n12064), .B1(n12266), .B2(n12074), .ZN(
        n10367) );
  NOR2_X1 U13210 ( .A1(n10368), .A2(n10367), .ZN(n10372) );
  INV_X1 U13211 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12075) );
  OAI22_X1 U13212 ( .A1(n12170), .A2(n20816), .B1(n12272), .B2(n12075), .ZN(
        n10370) );
  INV_X1 U13213 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12036) );
  OAI22_X1 U13214 ( .A1(n12036), .A2(n12275), .B1(n12017), .B2(n12068), .ZN(
        n10369) );
  NOR2_X1 U13215 ( .A1(n10370), .A2(n10369), .ZN(n10371) );
  NAND3_X1 U13216 ( .A1(n10373), .A2(n10372), .A3(n10371), .ZN(n14937) );
  AND2_X1 U13217 ( .A1(n10374), .A2(n14937), .ZN(n10397) );
  AOI22_X1 U13218 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13219 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10377) );
  NAND2_X1 U13220 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10376) );
  NAND2_X1 U13221 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10375) );
  NAND4_X1 U13222 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10382) );
  OAI22_X1 U13223 ( .A1(n12260), .A2(n10380), .B1(n12258), .B2(n10379), .ZN(
        n10381) );
  NOR2_X1 U13224 ( .A1(n10382), .A2(n10381), .ZN(n10396) );
  OAI22_X1 U13225 ( .A1(n12008), .A2(n10384), .B1(n12264), .B2(n10383), .ZN(
        n10388) );
  OAI22_X1 U13226 ( .A1(n12268), .A2(n10386), .B1(n12266), .B2(n10385), .ZN(
        n10387) );
  NOR2_X1 U13227 ( .A1(n10388), .A2(n10387), .ZN(n10395) );
  INV_X1 U13228 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10389) );
  OAI22_X1 U13229 ( .A1(n12170), .A2(n10390), .B1(n12272), .B2(n10389), .ZN(
        n10393) );
  INV_X1 U13230 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n19165) );
  OAI22_X1 U13231 ( .A1(n19165), .A2(n12275), .B1(n12017), .B2(n10391), .ZN(
        n10392) );
  NOR2_X1 U13232 ( .A1(n10393), .A2(n10392), .ZN(n10394) );
  NAND3_X1 U13233 ( .A1(n10396), .A2(n10395), .A3(n10394), .ZN(n14217) );
  NAND2_X1 U13234 ( .A1(n10397), .A2(n14217), .ZN(n10398) );
  NOR2_X1 U13235 ( .A1(n14173), .A2(n10398), .ZN(n10399) );
  AOI22_X1 U13236 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10408) );
  INV_X1 U13237 ( .A(n12808), .ZN(n12842) );
  AOI22_X1 U13238 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10407) );
  AND2_X1 U13239 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10402) );
  OR2_X1 U13240 ( .A1(n10402), .A2(n10401), .ZN(n12848) );
  INV_X1 U13241 ( .A(n12848), .ZN(n10504) );
  NAND2_X1 U13242 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13243 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10403) );
  AND3_X1 U13244 ( .A1(n10504), .A2(n10404), .A3(n10403), .ZN(n10406) );
  AOI22_X1 U13245 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9963), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10405) );
  NAND4_X1 U13246 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10416) );
  AOI22_X1 U13247 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13248 ( .A1(n12790), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13249 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U13250 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10410) );
  NAND2_X1 U13251 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10409) );
  AND3_X1 U13252 ( .A1(n10410), .A2(n12848), .A3(n10409), .ZN(n10411) );
  NAND4_X1 U13253 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10415) );
  NAND2_X1 U13254 ( .A1(n10416), .A2(n10415), .ZN(n10438) );
  NOR2_X1 U13255 ( .A1(n13146), .A2(n10438), .ZN(n10436) );
  OAI22_X1 U13256 ( .A1(n12008), .A2(n10417), .B1(n12264), .B2(n12119), .ZN(
        n10419) );
  OAI22_X1 U13257 ( .A1(n12268), .A2(n12115), .B1(n12266), .B2(n12120), .ZN(
        n10418) );
  NOR2_X1 U13258 ( .A1(n10419), .A2(n10418), .ZN(n10433) );
  INV_X1 U13259 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10420) );
  OAI22_X1 U13260 ( .A1(n12170), .A2(n10421), .B1(n12272), .B2(n10420), .ZN(
        n10423) );
  INV_X1 U13261 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19184) );
  OAI22_X1 U13262 ( .A1(n19184), .A2(n12275), .B1(n12017), .B2(n12118), .ZN(
        n10422) );
  NOR2_X1 U13263 ( .A1(n10423), .A2(n10422), .ZN(n10432) );
  OAI22_X1 U13264 ( .A1(n10424), .A2(n12260), .B1(n12258), .B2(n20853), .ZN(
        n10425) );
  INV_X1 U13265 ( .A(n10425), .ZN(n10431) );
  AOI22_X1 U13266 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13267 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U13268 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10427) );
  NAND2_X1 U13269 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10426) );
  AND4_X1 U13270 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  NAND4_X1 U13271 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10435) );
  INV_X1 U13272 ( .A(n10438), .ZN(n10434) );
  NAND2_X1 U13273 ( .A1(n10435), .A2(n10434), .ZN(n10457) );
  OAI22_X1 U13274 ( .A1(n10436), .A2(n10435), .B1(n13146), .B2(n10457), .ZN(
        n10460) );
  INV_X1 U13275 ( .A(n10460), .ZN(n10437) );
  NOR2_X1 U13276 ( .A1(n13571), .A2(n10438), .ZN(n14899) );
  INV_X1 U13277 ( .A(n10439), .ZN(n10440) );
  AOI22_X1 U13278 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12842), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13279 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13280 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9627), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U13281 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10443) );
  NAND2_X1 U13282 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10442) );
  AND3_X1 U13283 ( .A1(n10443), .A2(n12848), .A3(n10442), .ZN(n10444) );
  NAND4_X1 U13284 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10455) );
  AOI22_X1 U13285 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13286 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U13287 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10449) );
  NAND2_X1 U13288 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10448) );
  AND3_X1 U13289 ( .A1(n10504), .A2(n10449), .A3(n10448), .ZN(n10451) );
  AOI22_X1 U13290 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10450) );
  NAND4_X1 U13291 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10454) );
  AND2_X1 U13292 ( .A1(n10455), .A2(n10454), .ZN(n14893) );
  INV_X1 U13293 ( .A(n14893), .ZN(n10459) );
  INV_X1 U13294 ( .A(n10457), .ZN(n10456) );
  AND2_X1 U13295 ( .A1(n10456), .A2(n14893), .ZN(n10476) );
  AOI211_X1 U13296 ( .C1(n10459), .C2(n10457), .A(n10517), .B(n10476), .ZN(
        n14892) );
  INV_X1 U13297 ( .A(n14899), .ZN(n10458) );
  AOI22_X1 U13298 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13299 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U13300 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13301 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10461) );
  AND3_X1 U13302 ( .A1(n10504), .A2(n10462), .A3(n10461), .ZN(n10464) );
  AOI22_X1 U13303 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10463) );
  NAND4_X1 U13304 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10474) );
  AOI22_X1 U13305 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13306 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13307 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U13308 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10468) );
  NAND2_X1 U13309 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10467) );
  AND3_X1 U13310 ( .A1(n10468), .A2(n12848), .A3(n10467), .ZN(n10469) );
  NAND4_X1 U13311 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n10473) );
  AND2_X1 U13312 ( .A1(n10474), .A2(n10473), .ZN(n10478) );
  NAND2_X1 U13313 ( .A1(n10476), .A2(n10478), .ZN(n10497) );
  OAI211_X1 U13314 ( .C1(n10476), .C2(n10478), .A(n10475), .B(n10497), .ZN(
        n10480) );
  INV_X1 U13315 ( .A(n10478), .ZN(n10479) );
  NOR2_X1 U13316 ( .A1(n13571), .A2(n10479), .ZN(n14886) );
  AOI22_X1 U13317 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12842), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13318 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13319 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U13320 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10484) );
  NAND2_X1 U13321 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10483) );
  AND3_X1 U13322 ( .A1(n10484), .A2(n12848), .A3(n10483), .ZN(n10485) );
  NAND4_X1 U13323 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10496) );
  AOI22_X1 U13324 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13325 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13326 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16235), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10492) );
  NAND2_X1 U13327 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10490) );
  NAND2_X1 U13328 ( .A1(n9963), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10489) );
  AND3_X1 U13329 ( .A1(n10504), .A2(n10490), .A3(n10489), .ZN(n10491) );
  NAND4_X1 U13330 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10495) );
  NAND2_X1 U13331 ( .A1(n10496), .A2(n10495), .ZN(n10499) );
  AOI21_X1 U13332 ( .B1(n10497), .B2(n10499), .A(n10517), .ZN(n10498) );
  OR2_X1 U13333 ( .A1(n10497), .A2(n10499), .ZN(n10518) );
  NAND2_X1 U13334 ( .A1(n10498), .A2(n10518), .ZN(n10500) );
  NOR2_X1 U13335 ( .A1(n13571), .A2(n10499), .ZN(n14879) );
  INV_X1 U13336 ( .A(n10500), .ZN(n10501) );
  AOI22_X1 U13337 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13338 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10507) );
  NAND2_X1 U13339 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10503) );
  NAND2_X1 U13340 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10502) );
  AND3_X1 U13341 ( .A1(n10504), .A2(n10503), .A3(n10502), .ZN(n10506) );
  AOI22_X1 U13342 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10505) );
  NAND4_X1 U13343 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10516) );
  AOI22_X1 U13344 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13345 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13346 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10512) );
  NAND2_X1 U13347 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10510) );
  NAND2_X1 U13348 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10509) );
  AND3_X1 U13349 ( .A1(n10510), .A2(n10509), .A3(n12848), .ZN(n10511) );
  NAND4_X1 U13350 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10515) );
  NAND2_X1 U13351 ( .A1(n10516), .A2(n10515), .ZN(n10519) );
  AOI21_X1 U13352 ( .B1(n10518), .B2(n10519), .A(n10517), .ZN(n10521) );
  INV_X1 U13353 ( .A(n10518), .ZN(n10520) );
  INV_X1 U13354 ( .A(n10519), .ZN(n10522) );
  NAND2_X1 U13355 ( .A1(n10520), .A2(n10522), .ZN(n12818) );
  NAND2_X1 U13356 ( .A1(n10521), .A2(n12818), .ZN(n12789) );
  XNOR2_X1 U13357 ( .A(n12788), .B(n12789), .ZN(n10524) );
  NAND2_X1 U13358 ( .A1(n13146), .A2(n10522), .ZN(n10523) );
  AOI21_X1 U13359 ( .B1(n10524), .B2(n10523), .A(n12817), .ZN(n14959) );
  XNOR2_X1 U13360 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U13361 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19757), .ZN(
        n10537) );
  INV_X1 U13362 ( .A(n10537), .ZN(n10525) );
  AOI22_X1 U13363 ( .A1(n10538), .A2(n10525), .B1(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19751), .ZN(n10534) );
  INV_X1 U13364 ( .A(n10534), .ZN(n10527) );
  MUX2_X1 U13365 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n19742), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10533) );
  INV_X1 U13366 ( .A(n10533), .ZN(n10526) );
  NAND2_X1 U13367 ( .A1(n10527), .A2(n10526), .ZN(n10535) );
  NAND2_X1 U13368 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19742), .ZN(
        n10528) );
  NAND2_X1 U13369 ( .A1(n10535), .A2(n10528), .ZN(n10546) );
  INV_X1 U13370 ( .A(n10546), .ZN(n10530) );
  XNOR2_X1 U13371 ( .A(n10529), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10545) );
  INV_X1 U13372 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13471) );
  INV_X1 U13373 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15607) );
  NOR2_X1 U13374 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15607), .ZN(
        n10532) );
  AOI221_X1 U13375 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10544), 
        .C1(n13471), .C2(n10544), .A(n10532), .ZN(n12458) );
  INV_X1 U13376 ( .A(n12458), .ZN(n10549) );
  NAND2_X1 U13377 ( .A1(n19076), .A2(n13571), .ZN(n19773) );
  NAND2_X1 U13378 ( .A1(n10534), .A2(n10533), .ZN(n10536) );
  NAND2_X1 U13379 ( .A1(n10536), .A2(n10535), .ZN(n12437) );
  MUX2_X1 U13380 ( .A(n12144), .B(n19773), .S(n12437), .Z(n10543) );
  OAI21_X1 U13381 ( .B1(n19757), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10537), .ZN(n12145) );
  INV_X1 U13382 ( .A(n12145), .ZN(n12441) );
  NAND2_X1 U13383 ( .A1(n10538), .A2(n12441), .ZN(n12451) );
  NAND2_X1 U13384 ( .A1(n10075), .A2(n12451), .ZN(n10540) );
  XNOR2_X1 U13385 ( .A(n10538), .B(n10537), .ZN(n12438) );
  OAI211_X1 U13386 ( .C1(n13571), .C2(n12441), .A(n19076), .B(n12438), .ZN(
        n10539) );
  OAI211_X1 U13387 ( .C1(n10541), .C2(n12437), .A(n10540), .B(n10539), .ZN(
        n10542) );
  NAND2_X1 U13388 ( .A1(n10543), .A2(n10542), .ZN(n10547) );
  NAND3_X1 U13389 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10544), .A3(
        n13471), .ZN(n12153) );
  XNOR2_X1 U13390 ( .A(n10546), .B(n10545), .ZN(n12136) );
  NAND2_X1 U13391 ( .A1(n12153), .A2(n12136), .ZN(n12436) );
  MUX2_X1 U13392 ( .A(n10547), .B(n12144), .S(n12436), .Z(n10548) );
  NAND2_X1 U13393 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  MUX2_X1 U13394 ( .A(n10550), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19780), .Z(n13142) );
  AND2_X1 U13395 ( .A1(n16265), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13425) );
  NAND2_X1 U13396 ( .A1(n12458), .A2(n13425), .ZN(n10551) );
  INV_X1 U13397 ( .A(n16263), .ZN(n10554) );
  NAND2_X1 U13398 ( .A1(n10552), .A2(n10553), .ZN(n16219) );
  INV_X1 U13399 ( .A(n16219), .ZN(n16257) );
  NAND2_X1 U13400 ( .A1(n10554), .A2(n16257), .ZN(n13462) );
  NAND2_X1 U13401 ( .A1(n13462), .A2(n16224), .ZN(n10556) );
  INV_X1 U13402 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15404) );
  NAND2_X1 U13403 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15404), .ZN(n13066) );
  INV_X1 U13404 ( .A(n13066), .ZN(n10555) );
  AND2_X1 U13405 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10555), .ZN(n19633) );
  NAND2_X1 U13406 ( .A1(n10556), .A2(n19633), .ZN(n13608) );
  INV_X1 U13407 ( .A(n13011), .ZN(n19116) );
  INV_X1 U13408 ( .A(n14942), .ZN(n14175) );
  NAND2_X1 U13409 ( .A1(n14959), .A2(n14175), .ZN(n10649) );
  INV_X1 U13410 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13411 ( .A1(n13059), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10557) );
  OAI21_X1 U13412 ( .B1(n13207), .B2(n10558), .A(n10557), .ZN(n10559) );
  AOI21_X1 U13413 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10559), .ZN(n10644) );
  NAND2_X1 U13414 ( .A1(n10561), .A2(n10560), .ZN(n10566) );
  INV_X1 U13415 ( .A(n10562), .ZN(n10563) );
  OR2_X1 U13416 ( .A1(n10564), .A2(n10563), .ZN(n10565) );
  NAND2_X1 U13417 ( .A1(n10566), .A2(n10565), .ZN(n13611) );
  NAND2_X1 U13418 ( .A1(n10621), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13419 ( .A1(n10098), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10567) );
  NAND2_X1 U13420 ( .A1(n10568), .A2(n10567), .ZN(n10569) );
  AOI21_X1 U13421 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n10569), .ZN(n13612) );
  NAND2_X1 U13422 ( .A1(n10621), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13423 ( .A1(n10098), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10571) );
  NAND2_X1 U13424 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  AOI21_X1 U13425 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10573), .ZN(n13739) );
  INV_X1 U13426 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14193) );
  AOI22_X1 U13427 ( .A1(n10098), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10575) );
  NAND2_X1 U13428 ( .A1(n10621), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10574) );
  OAI211_X1 U13429 ( .C1(n10154), .C2(n14193), .A(n10575), .B(n10574), .ZN(
        n13749) );
  NAND2_X1 U13430 ( .A1(n10621), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13431 ( .A1(n10098), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10576) );
  NAND2_X1 U13432 ( .A1(n10577), .A2(n10576), .ZN(n10578) );
  AOI21_X1 U13433 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10578), .ZN(n13766) );
  NAND2_X1 U13434 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10582) );
  NAND2_X1 U13435 ( .A1(n10621), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10580) );
  AOI22_X1 U13436 ( .A1(n10098), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10579) );
  AND2_X1 U13437 ( .A1(n10580), .A2(n10579), .ZN(n10581) );
  NAND2_X1 U13438 ( .A1(n10582), .A2(n10581), .ZN(n13789) );
  NAND2_X1 U13439 ( .A1(n10621), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13440 ( .A1(n13059), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10583) );
  NAND2_X1 U13441 ( .A1(n10584), .A2(n10583), .ZN(n10585) );
  AOI21_X1 U13442 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10585), .ZN(n13800) );
  INV_X1 U13443 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16183) );
  AOI22_X1 U13444 ( .A1(n13059), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10587) );
  NAND2_X1 U13445 ( .A1(n10621), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10586) );
  OAI211_X1 U13446 ( .C1(n10154), .C2(n16183), .A(n10587), .B(n10586), .ZN(
        n13856) );
  NAND2_X1 U13447 ( .A1(n10621), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13448 ( .A1(n13059), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10588) );
  NAND2_X1 U13449 ( .A1(n10589), .A2(n10588), .ZN(n10590) );
  AOI21_X1 U13450 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10590), .ZN(n13909) );
  NAND2_X1 U13451 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10594) );
  NAND2_X1 U13452 ( .A1(n10621), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13453 ( .A1(n13059), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10591) );
  AND2_X1 U13454 ( .A1(n10592), .A2(n10591), .ZN(n10593) );
  NAND2_X1 U13455 ( .A1(n10594), .A2(n10593), .ZN(n14032) );
  INV_X1 U13456 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U13457 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10596) );
  AOI22_X1 U13458 ( .A1(n13059), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10595) );
  OAI211_X1 U13459 ( .C1(n12326), .C2(n13207), .A(n10596), .B(n10595), .ZN(
        n14037) );
  NAND2_X1 U13460 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10600) );
  NAND2_X1 U13461 ( .A1(n10621), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13462 ( .A1(n13059), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10597) );
  AND2_X1 U13463 ( .A1(n10598), .A2(n10597), .ZN(n10599) );
  NAND2_X1 U13464 ( .A1(n10600), .A2(n10599), .ZN(n14108) );
  NAND2_X1 U13465 ( .A1(n10621), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13466 ( .A1(n13059), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10601) );
  NAND2_X1 U13467 ( .A1(n10602), .A2(n10601), .ZN(n10603) );
  AOI21_X1 U13468 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10603), .ZN(n14170) );
  NOR2_X2 U13469 ( .A1(n14171), .A2(n14170), .ZN(n14160) );
  INV_X1 U13470 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12350) );
  NAND2_X1 U13471 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10605) );
  AOI22_X1 U13472 ( .A1(n13059), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10604) );
  OAI211_X1 U13473 ( .C1(n12350), .C2(n13207), .A(n10605), .B(n10604), .ZN(
        n14162) );
  NAND2_X1 U13474 ( .A1(n10621), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13475 ( .A1(n13059), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10606) );
  NAND2_X1 U13476 ( .A1(n10607), .A2(n10606), .ZN(n10608) );
  AOI21_X1 U13477 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10608), .ZN(n14939) );
  NAND2_X1 U13478 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10612) );
  NAND2_X1 U13479 ( .A1(n10621), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13480 ( .A1(n13059), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10609) );
  AND2_X1 U13481 ( .A1(n10610), .A2(n10609), .ZN(n10611) );
  NAND2_X1 U13482 ( .A1(n10612), .A2(n10611), .ZN(n12526) );
  NAND2_X1 U13483 ( .A1(n10621), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13484 ( .A1(n13059), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10613) );
  NAND2_X1 U13485 ( .A1(n10614), .A2(n10613), .ZN(n10615) );
  AOI21_X1 U13486 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10615), .ZN(n13217) );
  NAND2_X1 U13487 ( .A1(n10621), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13488 ( .A1(n13059), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10618) );
  NAND2_X1 U13489 ( .A1(n10619), .A2(n10618), .ZN(n10620) );
  AOI21_X1 U13490 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10620), .ZN(n14852) );
  NAND2_X1 U13491 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13492 ( .A1(n10621), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13493 ( .A1(n13059), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10622) );
  AND2_X1 U13494 ( .A1(n10623), .A2(n10622), .ZN(n10624) );
  NAND2_X1 U13495 ( .A1(n10625), .A2(n10624), .ZN(n14841) );
  NAND2_X1 U13496 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10629) );
  NAND2_X1 U13497 ( .A1(n10621), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13498 ( .A1(n13059), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10626) );
  AND2_X1 U13499 ( .A1(n10627), .A2(n10626), .ZN(n10628) );
  NAND2_X1 U13500 ( .A1(n10629), .A2(n10628), .ZN(n14906) );
  INV_X1 U13501 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U13502 ( .A1(n13059), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10630) );
  OAI21_X1 U13503 ( .B1(n13207), .B2(n12388), .A(n10630), .ZN(n10631) );
  AOI21_X1 U13504 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13204), .A(
        n10631), .ZN(n14901) );
  NAND2_X1 U13505 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10635) );
  NAND2_X1 U13506 ( .A1(n10621), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13507 ( .A1(n13059), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10632) );
  AND2_X1 U13508 ( .A1(n10633), .A2(n10632), .ZN(n10634) );
  NAND2_X1 U13509 ( .A1(n10635), .A2(n10634), .ZN(n13277) );
  NAND2_X1 U13510 ( .A1(n13276), .A2(n13277), .ZN(n13275) );
  INV_X1 U13511 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13512 ( .A1(n13059), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10636) );
  OAI21_X1 U13513 ( .B1(n13207), .B2(n10637), .A(n10636), .ZN(n10638) );
  AOI21_X1 U13514 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10638), .ZN(n14888) );
  NAND2_X1 U13515 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10642) );
  NAND2_X1 U13516 ( .A1(n10621), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10640) );
  AOI22_X1 U13517 ( .A1(n13059), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10639) );
  AND2_X1 U13518 ( .A1(n10640), .A2(n10639), .ZN(n10641) );
  NAND2_X1 U13519 ( .A1(n10642), .A2(n10641), .ZN(n14881) );
  AOI21_X1 U13520 ( .B1(n10644), .B2(n9660), .A(n10643), .ZN(n15959) );
  INV_X1 U13521 ( .A(n15959), .ZN(n10646) );
  NAND2_X1 U13522 ( .A1(n13608), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10645) );
  NAND2_X1 U13523 ( .A1(n10649), .A2(n10648), .ZN(P2_U2860) );
  INV_X1 U13524 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16308) );
  NAND2_X2 U13525 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10650), .ZN(
        n16821) );
  INV_X1 U13526 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U13527 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10654) );
  INV_X2 U13528 ( .A(n9586), .ZN(n17062) );
  AOI22_X1 U13529 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10750), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10653) );
  OAI211_X1 U13530 ( .C1(n16821), .C2(n17084), .A(n10654), .B(n10653), .ZN(
        n10655) );
  INV_X1 U13531 ( .A(n10655), .ZN(n10670) );
  INV_X2 U13532 ( .A(n9587), .ZN(n17014) );
  AOI22_X1 U13533 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13534 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10701), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10661) );
  NAND2_X1 U13535 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10665), .ZN(
        n10844) );
  AOI22_X1 U13536 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10660) );
  INV_X4 U13537 ( .A(n10732), .ZN(n16828) );
  NAND2_X1 U13538 ( .A1(n16828), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10659) );
  INV_X1 U13539 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17100) );
  NOR2_X1 U13540 ( .A1(n9598), .A2(n17100), .ZN(n10664) );
  AOI22_X1 U13541 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U13542 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17758), .ZN(
        n17757) );
  INV_X1 U13543 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U13544 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10681) );
  INV_X1 U13545 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16949) );
  INV_X1 U13546 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10674) );
  INV_X1 U13547 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10673) );
  INV_X1 U13548 ( .A(n10675), .ZN(n10678) );
  AOI22_X1 U13549 ( .A1(n10676), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10677) );
  OAI211_X1 U13550 ( .C1(n16821), .C2(n16949), .A(n10678), .B(n10677), .ZN(
        n10679) );
  INV_X1 U13551 ( .A(n10679), .ZN(n10680) );
  NAND3_X1 U13552 ( .A1(n10682), .A2(n10681), .A3(n10680), .ZN(n10689) );
  AOI22_X1 U13553 ( .A1(n10701), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13554 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10750), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10686) );
  INV_X2 U13555 ( .A(n10699), .ZN(n15473) );
  AOI22_X1 U13556 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10685) );
  NAND2_X1 U13557 ( .A1(n10683), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10684) );
  NAND4_X1 U13558 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10688) );
  NOR2_X1 U13559 ( .A1(n10949), .A2(n10690), .ZN(n10691) );
  INV_X1 U13560 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18071) );
  INV_X1 U13561 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U13562 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10693), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10694) );
  OAI21_X1 U13563 ( .B1(n17011), .B2(n17128), .A(n10694), .ZN(n10696) );
  INV_X1 U13564 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16935) );
  INV_X1 U13565 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17046) );
  OAI22_X1 U13566 ( .A1(n15507), .A2(n16935), .B1(n10844), .B2(n17046), .ZN(
        n10695) );
  AOI22_X1 U13567 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10750), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10697) );
  INV_X1 U13568 ( .A(n10697), .ZN(n10698) );
  AOI22_X1 U13569 ( .A1(n16828), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10706) );
  INV_X1 U13570 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n20883) );
  AOI22_X1 U13571 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13572 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10701), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10702) );
  INV_X1 U13573 ( .A(n10702), .ZN(n10703) );
  XNOR2_X1 U13574 ( .A(n18071), .B(n10709), .ZN(n17739) );
  NOR2_X1 U13575 ( .A1(n18071), .A2(n10709), .ZN(n10710) );
  INV_X1 U13576 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U13577 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13578 ( .A1(n15473), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10711) );
  OAI211_X1 U13579 ( .C1(n16821), .C2(n16919), .A(n10712), .B(n10711), .ZN(
        n10713) );
  AOI22_X1 U13580 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10715) );
  INV_X1 U13581 ( .A(n10715), .ZN(n10718) );
  INV_X1 U13582 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17122) );
  NAND2_X1 U13583 ( .A1(n16828), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10716) );
  OAI21_X1 U13584 ( .B1(n17011), .B2(n17122), .A(n10716), .ZN(n10717) );
  AOI22_X1 U13585 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13586 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13587 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10657), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10723) );
  NAND2_X1 U13588 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10722) );
  NAND4_X1 U13589 ( .A1(n10725), .A2(n10724), .A3(n10723), .A4(n10722), .ZN(
        n10726) );
  INV_X1 U13590 ( .A(n10952), .ZN(n17277) );
  INV_X1 U13591 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13592 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10721), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10731) );
  OAI21_X1 U13593 ( .B1(n10811), .B2(n10892), .A(n10731), .ZN(n10745) );
  AOI22_X1 U13594 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13595 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13596 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16828), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10733) );
  NAND3_X1 U13597 ( .A1(n10735), .A2(n10734), .A3(n10733), .ZN(n10743) );
  AOI22_X1 U13598 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10741) );
  INV_X1 U13599 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17120) );
  INV_X1 U13600 ( .A(n10737), .ZN(n10740) );
  INV_X1 U13601 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17021) );
  INV_X1 U13602 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16905) );
  OAI22_X1 U13603 ( .A1(n16821), .A2(n17021), .B1(n17061), .B2(n16905), .ZN(
        n10738) );
  NAND3_X1 U13604 ( .A1(n10741), .A2(n10740), .A3(n10739), .ZN(n10742) );
  AOI211_X2 U13605 ( .C1(n9599), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n10745), .B(n10744), .ZN(n17273) );
  XOR2_X1 U13606 ( .A(n10747), .B(n17273), .Z(n17719) );
  NAND2_X1 U13607 ( .A1(n9658), .A2(n9785), .ZN(n10746) );
  INV_X1 U13608 ( .A(n17273), .ZN(n10963) );
  INV_X1 U13609 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U13610 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10758) );
  INV_X1 U13611 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U13612 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13613 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10748) );
  OAI211_X1 U13614 ( .C1(n16821), .C2(n15472), .A(n10749), .B(n10748), .ZN(
        n10756) );
  AOI22_X1 U13615 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13616 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13617 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10657), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U13618 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10751) );
  NAND4_X1 U13619 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10755) );
  NOR2_X2 U13620 ( .A1(n17707), .A2(n17706), .ZN(n17705) );
  NAND2_X1 U13621 ( .A1(n17706), .A2(n17707), .ZN(n10759) );
  INV_X1 U13622 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U13623 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n17027), .ZN(n10761) );
  OAI21_X1 U13624 ( .B1(n17109), .B2(n17011), .A(n10761), .ZN(n10771) );
  INV_X1 U13625 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13626 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n9595), .ZN(n10768) );
  INV_X1 U13627 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U13628 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n9596), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10762) );
  OAI21_X1 U13629 ( .B1(n15507), .B2(n16995), .A(n10762), .ZN(n10766) );
  INV_X1 U13630 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16807) );
  AOI22_X1 U13631 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n17066), .ZN(n10764) );
  AOI22_X1 U13632 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n17047), .B1(
        n10701), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10763) );
  OAI211_X1 U13633 ( .C1(n16807), .C2(n16821), .A(n10764), .B(n10763), .ZN(
        n10765) );
  AOI211_X1 U13634 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n10766), .B(n10765), .ZN(n10767) );
  OAI211_X1 U13635 ( .C1(n16957), .C2(n10769), .A(n10768), .B(n10767), .ZN(
        n10770) );
  INV_X1 U13636 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n20927) );
  AOI22_X1 U13637 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10782) );
  INV_X1 U13638 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U13639 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13640 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10773) );
  OAI211_X1 U13641 ( .C1(n10732), .C2(n16987), .A(n10774), .B(n10773), .ZN(
        n10780) );
  AOI22_X1 U13642 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13643 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10777) );
  INV_X2 U13644 ( .A(n17074), .ZN(n17047) );
  AOI22_X1 U13645 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13646 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10775) );
  NAND4_X1 U13647 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10779) );
  AOI211_X1 U13648 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n10780), .B(n10779), .ZN(n10781) );
  INV_X1 U13649 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18015) );
  NOR2_X1 U13650 ( .A1(n17684), .A2(n18015), .ZN(n17683) );
  NOR2_X1 U13651 ( .A1(n10785), .A2(n10786), .ZN(n10787) );
  INV_X1 U13652 ( .A(n10789), .ZN(n10788) );
  INV_X1 U13653 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17997) );
  NAND2_X1 U13654 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17972) );
  INV_X1 U13655 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17946) );
  NOR2_X1 U13656 ( .A1(n17972), .A2(n17946), .ZN(n17953) );
  NAND2_X1 U13657 ( .A1(n17953), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17926) );
  NAND2_X1 U13658 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17575) );
  NOR2_X1 U13659 ( .A1(n17926), .A2(n17575), .ZN(n17902) );
  NAND2_X1 U13660 ( .A1(n17902), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17876) );
  NAND2_X1 U13661 ( .A1(n9654), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10796) );
  NOR2_X1 U13662 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17646) );
  INV_X1 U13663 ( .A(n17646), .ZN(n10793) );
  NAND2_X1 U13664 ( .A1(n17628), .A2(n17946), .ZN(n17604) );
  NOR2_X2 U13665 ( .A1(n17604), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17566) );
  INV_X1 U13666 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17945) );
  NAND2_X1 U13667 ( .A1(n17566), .A2(n17945), .ZN(n17582) );
  INV_X1 U13668 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17932) );
  INV_X1 U13669 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17899) );
  NAND2_X1 U13670 ( .A1(n17932), .A2(n17899), .ZN(n17911) );
  INV_X1 U13671 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17890) );
  NOR2_X1 U13672 ( .A1(n10794), .A2(n17890), .ZN(n17879) );
  INV_X1 U13673 ( .A(n17879), .ZN(n17538) );
  INV_X1 U13674 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17884) );
  INV_X1 U13675 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17850) );
  NAND2_X1 U13676 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17849) );
  NOR3_X1 U13677 ( .A1(n17884), .A2(n17850), .A3(n17849), .ZN(n17475) );
  NAND2_X1 U13678 ( .A1(n17475), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12760) );
  NOR2_X1 U13679 ( .A1(n17538), .A2(n12760), .ZN(n17804) );
  NAND2_X1 U13680 ( .A1(n17804), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17465) );
  NAND2_X1 U13681 ( .A1(n10791), .A2(n17884), .ZN(n17531) );
  NOR2_X1 U13682 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17531), .ZN(
        n10798) );
  INV_X1 U13683 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17861) );
  NAND2_X1 U13684 ( .A1(n10798), .A2(n17861), .ZN(n17501) );
  NOR2_X1 U13685 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17501), .ZN(
        n17476) );
  INV_X1 U13686 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17839) );
  NAND2_X1 U13687 ( .A1(n17476), .A2(n17839), .ZN(n17477) );
  OAI22_X1 U13688 ( .A1(n9631), .A2(n17465), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17477), .ZN(n10799) );
  NAND2_X1 U13689 ( .A1(n17474), .A2(n10799), .ZN(n17457) );
  INV_X1 U13690 ( .A(n12760), .ZN(n10802) );
  AND2_X1 U13691 ( .A1(n10802), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10803) );
  AND3_X2 U13692 ( .A1(n9645), .A2(n17455), .A3(n10803), .ZN(n10805) );
  INV_X1 U13693 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17801) );
  NAND2_X1 U13694 ( .A1(n10791), .A2(n17455), .ZN(n10804) );
  NAND2_X1 U13695 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17767) );
  INV_X1 U13696 ( .A(n17767), .ZN(n10806) );
  NOR2_X1 U13697 ( .A1(n10807), .A2(n10806), .ZN(n10808) );
  INV_X1 U13698 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12758) );
  NAND3_X1 U13699 ( .A1(n12756), .A2(n12758), .A3(n10791), .ZN(n15515) );
  NOR2_X1 U13700 ( .A1(n16288), .A2(n16287), .ZN(n10810) );
  XNOR2_X1 U13701 ( .A(n10810), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15591) );
  INV_X1 U13702 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U13703 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13704 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10812) );
  OAI211_X1 U13705 ( .C1(n16821), .C2(n15448), .A(n10813), .B(n10812), .ZN(
        n10821) );
  INV_X1 U13706 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U13707 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13708 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10814) );
  OAI21_X1 U13709 ( .B1(n15507), .B2(n17130), .A(n10814), .ZN(n10817) );
  AOI22_X1 U13710 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10815) );
  OAI21_X1 U13711 ( .B1(n17065), .B2(n10674), .A(n10815), .ZN(n10816) );
  AOI211_X1 U13712 ( .C1(n9599), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n10817), .B(n10816), .ZN(n10818) );
  OAI211_X1 U13713 ( .C1(n16957), .C2(n17073), .A(n10819), .B(n10818), .ZN(
        n10820) );
  AOI211_X4 U13714 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n10821), .B(n10820), .ZN(n17332) );
  INV_X1 U13715 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U13716 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10831) );
  INV_X1 U13717 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U13718 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13719 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10822) );
  OAI211_X1 U13720 ( .C1(n16821), .C2(n17044), .A(n10823), .B(n10822), .ZN(
        n10829) );
  AOI22_X1 U13721 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13722 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13723 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U13724 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10824) );
  NAND4_X1 U13725 ( .A1(n10827), .A2(n10826), .A3(n10825), .A4(n10824), .ZN(
        n10828) );
  AOI211_X1 U13726 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n10829), .B(n10828), .ZN(n10830) );
  INV_X1 U13727 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13728 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10832) );
  OAI21_X1 U13729 ( .B1(n10811), .B2(n10833), .A(n10832), .ZN(n10842) );
  INV_X1 U13730 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U13731 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13732 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16828), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10834) );
  OAI21_X1 U13733 ( .B1(n15507), .B2(n17122), .A(n10834), .ZN(n10838) );
  INV_X1 U13734 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15460) );
  AOI22_X1 U13735 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13736 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10835) );
  OAI211_X1 U13737 ( .C1(n16821), .C2(n15460), .A(n10836), .B(n10835), .ZN(
        n10837) );
  AOI211_X1 U13738 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n10838), .B(n10837), .ZN(n10839) );
  OAI211_X1 U13739 ( .C1(n9587), .C2(n15459), .A(n10840), .B(n10839), .ZN(
        n10841) );
  INV_X1 U13740 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U13741 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10843) );
  OAI21_X1 U13742 ( .B1(n15507), .B2(n17085), .A(n10843), .ZN(n10854) );
  INV_X1 U13743 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13744 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10851) );
  INV_X1 U13745 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U13746 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10845) );
  OAI21_X1 U13747 ( .B1(n16957), .B2(n15431), .A(n10845), .ZN(n10849) );
  INV_X1 U13748 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U13749 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13750 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10846) );
  OAI211_X1 U13751 ( .C1(n16821), .C2(n17086), .A(n10847), .B(n10846), .ZN(
        n10848) );
  AOI211_X1 U13752 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n10849), .B(n10848), .ZN(n10850) );
  OAI211_X1 U13753 ( .C1(n9587), .C2(n10852), .A(n10851), .B(n10850), .ZN(
        n10853) );
  INV_X1 U13754 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16820) );
  INV_X1 U13755 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16831) );
  OAI22_X1 U13756 ( .A1(n16957), .A2(n16820), .B1(n10732), .B2(n16831), .ZN(
        n10859) );
  AOI22_X1 U13757 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13758 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13759 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10855) );
  NAND3_X1 U13760 ( .A1(n10857), .A2(n10856), .A3(n10855), .ZN(n10858) );
  AOI211_X1 U13761 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n10859), .B(n10858), .ZN(n10867) );
  INV_X1 U13762 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U13763 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10860) );
  OAI21_X1 U13764 ( .B1(n15507), .B2(n16982), .A(n10860), .ZN(n10861) );
  INV_X1 U13765 ( .A(n10861), .ZN(n10866) );
  AOI22_X1 U13766 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10865) );
  INV_X1 U13767 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16979) );
  INV_X1 U13768 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17113) );
  INV_X1 U13769 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20847) );
  OAI22_X1 U13770 ( .A1(n15507), .A2(n17113), .B1(n16957), .B2(n20847), .ZN(
        n10878) );
  AOI22_X1 U13771 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13772 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10875) );
  INV_X1 U13773 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U13774 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16828), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10868) );
  OAI21_X1 U13775 ( .B1(n9644), .B2(n16889), .A(n10868), .ZN(n10873) );
  INV_X1 U13776 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13777 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13778 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10869) );
  OAI211_X1 U13779 ( .C1(n16821), .C2(n10871), .A(n10870), .B(n10869), .ZN(
        n10872) );
  AOI211_X1 U13780 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n10873), .B(n10872), .ZN(n10874) );
  NAND3_X1 U13781 ( .A1(n10876), .A2(n10875), .A3(n10874), .ZN(n10877) );
  INV_X1 U13782 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16808) );
  AOI22_X1 U13783 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10888) );
  INV_X1 U13784 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U13785 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13786 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10879) );
  OAI211_X1 U13787 ( .C1(n16821), .C2(n16997), .A(n10880), .B(n10879), .ZN(
        n10886) );
  AOI22_X1 U13788 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U13789 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U13790 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U13791 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10881) );
  NAND4_X1 U13792 ( .A1(n10884), .A2(n10883), .A3(n10882), .A4(n10881), .ZN(
        n10885) );
  AOI211_X1 U13793 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n10886), .B(n10885), .ZN(n10887) );
  OAI211_X1 U13794 ( .C1(n16957), .C2(n16808), .A(n10888), .B(n10887), .ZN(
        n10921) );
  INV_X1 U13795 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17013) );
  OAI22_X1 U13796 ( .A1(n15507), .A2(n17120), .B1(n10811), .B2(n17013), .ZN(
        n10899) );
  AOI22_X1 U13797 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13798 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10896) );
  INV_X1 U13799 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U13800 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10889) );
  OAI21_X1 U13801 ( .B1(n17065), .B2(n17010), .A(n10889), .ZN(n10894) );
  AOI22_X1 U13802 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13803 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10890) );
  OAI211_X1 U13804 ( .C1(n16821), .C2(n10892), .A(n10891), .B(n10890), .ZN(
        n10893) );
  AOI211_X1 U13805 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n10894), .B(n10893), .ZN(n10895) );
  NAND3_X1 U13806 ( .A1(n10897), .A2(n10896), .A3(n10895), .ZN(n10898) );
  INV_X1 U13807 ( .A(n10906), .ZN(n10900) );
  NOR2_X1 U13808 ( .A1(n18127), .A2(n18122), .ZN(n10910) );
  NAND4_X1 U13809 ( .A1(n18115), .A2(n18119), .A3(n10908), .A4(n10910), .ZN(
        n10918) );
  NAND2_X1 U13810 ( .A1(n16730), .A2(n18749), .ZN(n10920) );
  NOR2_X1 U13811 ( .A1(n16439), .A2(n10920), .ZN(n14227) );
  NOR2_X1 U13812 ( .A1(n10902), .A2(n14227), .ZN(n18533) );
  INV_X1 U13813 ( .A(n18122), .ZN(n17144) );
  NOR2_X1 U13814 ( .A1(n18127), .A2(n17144), .ZN(n10935) );
  NAND2_X1 U13815 ( .A1(n10935), .A2(n18549), .ZN(n15486) );
  INV_X1 U13816 ( .A(n15486), .ZN(n10903) );
  NAND3_X1 U13817 ( .A1(n10908), .A2(n17332), .A3(n10903), .ZN(n10904) );
  INV_X2 U13818 ( .A(n18564), .ZN(n18558) );
  NOR2_X1 U13819 ( .A1(n17332), .A2(n10937), .ZN(n10915) );
  NOR2_X1 U13820 ( .A1(n18122), .A2(n12731), .ZN(n12733) );
  INV_X1 U13821 ( .A(n12733), .ZN(n10905) );
  NOR2_X1 U13822 ( .A1(n18122), .A2(n10921), .ZN(n15613) );
  NOR2_X1 U13823 ( .A1(n18134), .A2(n15613), .ZN(n15612) );
  NAND2_X1 U13824 ( .A1(n17332), .A2(n10901), .ZN(n10919) );
  NAND2_X1 U13825 ( .A1(n18111), .A2(n10910), .ZN(n12743) );
  AOI21_X1 U13826 ( .B1(n10906), .B2(n12743), .A(n10901), .ZN(n10913) );
  INV_X1 U13827 ( .A(n15613), .ZN(n18570) );
  INV_X1 U13828 ( .A(n18119), .ZN(n10936) );
  OAI22_X1 U13829 ( .A1(n10908), .A2(n10907), .B1(n18570), .B2(n10936), .ZN(
        n10912) );
  AND2_X1 U13830 ( .A1(n10920), .A2(n18111), .ZN(n10938) );
  OAI21_X1 U13831 ( .B1(n10910), .B2(n18134), .A(n10936), .ZN(n10909) );
  OAI21_X1 U13832 ( .B1(n10910), .B2(n10938), .A(n10909), .ZN(n10911) );
  NOR3_X2 U13833 ( .A1(n10913), .A2(n10912), .A3(n10911), .ZN(n12736) );
  AOI21_X1 U13834 ( .B1(n18533), .B2(n10915), .A(n10917), .ZN(n10916) );
  INV_X1 U13835 ( .A(n10916), .ZN(n18548) );
  AOI21_X4 U13836 ( .B1(n18549), .B2(n18558), .A(n18548), .ZN(n18571) );
  NAND2_X1 U13837 ( .A1(n10920), .A2(n10919), .ZN(n18767) );
  NOR2_X1 U13838 ( .A1(n18119), .A2(n10921), .ZN(n18550) );
  NAND3_X1 U13839 ( .A1(n10937), .A2(n12733), .A3(n18550), .ZN(n15488) );
  NOR2_X2 U13840 ( .A1(n17768), .A2(n18559), .ZN(n17811) );
  OAI22_X1 U13841 ( .A1(n18727), .A2(n18576), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10942) );
  NOR2_X1 U13842 ( .A1(n18733), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10941) );
  INV_X1 U13843 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18545) );
  INV_X1 U13844 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18411) );
  AND2_X1 U13845 ( .A1(n10942), .A2(n10941), .ZN(n10923) );
  AOI21_X1 U13846 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18576), .A(
        n10923), .ZN(n10928) );
  OAI22_X1 U13847 ( .A1(n10651), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18411), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10927) );
  NOR2_X1 U13848 ( .A1(n10928), .A2(n10927), .ZN(n10924) );
  AOI21_X1 U13849 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18411), .A(
        n10924), .ZN(n10925) );
  AOI22_X1 U13850 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18545), .B1(
        n10925), .B2(n18711), .ZN(n10929) );
  INV_X1 U13851 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18585) );
  NOR2_X1 U13852 ( .A1(n10925), .A2(n18711), .ZN(n10930) );
  NAND2_X1 U13853 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18545), .ZN(
        n10926) );
  OAI22_X1 U13854 ( .A1(n10929), .A2(n18585), .B1(n10930), .B2(n10926), .ZN(
        n10933) );
  AOI211_X1 U13855 ( .C1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n18733), .A(
        n10941), .B(n10933), .ZN(n10940) );
  XNOR2_X1 U13856 ( .A(n10928), .B(n10927), .ZN(n10947) );
  OAI21_X1 U13857 ( .B1(n18585), .B2(n10930), .A(n10929), .ZN(n10931) );
  OAI21_X1 U13858 ( .B1(n18545), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n10931), .ZN(n10945) );
  INV_X1 U13859 ( .A(n10945), .ZN(n10932) );
  OAI21_X1 U13860 ( .B1(n10933), .B2(n10947), .A(n10932), .ZN(n10943) );
  AOI21_X1 U13861 ( .B1(n10942), .B2(n10940), .A(n10943), .ZN(n18541) );
  NAND2_X1 U13862 ( .A1(n18111), .A2(n18749), .ZN(n10934) );
  NOR2_X1 U13863 ( .A1(n18127), .A2(n10934), .ZN(n12741) );
  OAI21_X1 U13864 ( .B1(n10936), .B2(n10935), .A(n18570), .ZN(n10939) );
  AND3_X1 U13865 ( .A1(n10939), .A2(n10938), .A3(n10937), .ZN(n12737) );
  NAND2_X1 U13866 ( .A1(n12741), .A2(n12737), .ZN(n12755) );
  INV_X1 U13867 ( .A(n10940), .ZN(n10946) );
  XOR2_X1 U13868 ( .A(n10942), .B(n10941), .Z(n10944) );
  OAI21_X1 U13869 ( .B1(n10945), .B2(n10944), .A(n10943), .ZN(n13100) );
  OAI21_X1 U13870 ( .B1(n10947), .B2(n10946), .A(n13100), .ZN(n18536) );
  INV_X1 U13871 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18753) );
  NOR2_X1 U13872 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18753), .ZN(n17760) );
  NAND2_X1 U13873 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n17760), .ZN(n18603) );
  INV_X1 U13874 ( .A(n18603), .ZN(n18757) );
  NAND2_X1 U13875 ( .A1(n15591), .A2(n17671), .ZN(n10993) );
  NAND3_X1 U13876 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17789) );
  INV_X1 U13877 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10948) );
  NOR2_X1 U13878 ( .A1(n17789), .A2(n10948), .ZN(n12759) );
  INV_X1 U13879 ( .A(n12759), .ZN(n17765) );
  NAND2_X1 U13880 ( .A1(n10949), .A2(n17758), .ZN(n10953) );
  NAND2_X1 U13881 ( .A1(n17280), .A2(n10953), .ZN(n10951) );
  NAND2_X1 U13882 ( .A1(n10952), .A2(n10951), .ZN(n10962) );
  NOR2_X1 U13883 ( .A1(n17273), .A2(n10962), .ZN(n10950) );
  NAND2_X1 U13884 ( .A1(n10950), .A2(n17267), .ZN(n10969) );
  NOR2_X1 U13885 ( .A1(n17264), .A2(n10969), .ZN(n10973) );
  NAND2_X1 U13886 ( .A1(n10973), .A2(n15517), .ZN(n10974) );
  XOR2_X1 U13887 ( .A(n17267), .B(n10950), .Z(n10967) );
  AND2_X1 U13888 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10967), .ZN(
        n10968) );
  INV_X1 U13889 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18041) );
  XNOR2_X1 U13890 ( .A(n10952), .B(n10951), .ZN(n10960) );
  NOR2_X1 U13891 ( .A1(n18041), .A2(n10960), .ZN(n10961) );
  XOR2_X1 U13892 ( .A(n17280), .B(n10953), .Z(n10954) );
  NOR2_X1 U13893 ( .A1(n10954), .A2(n18071), .ZN(n10959) );
  XNOR2_X1 U13894 ( .A(n18071), .B(n10954), .ZN(n17742) );
  INV_X1 U13895 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18730) );
  NOR2_X1 U13896 ( .A1(n17291), .A2(n18730), .ZN(n10957) );
  INV_X1 U13897 ( .A(n17758), .ZN(n10956) );
  NAND3_X1 U13898 ( .A1(n10956), .A2(n17291), .A3(n18730), .ZN(n10955) );
  OAI221_X1 U13899 ( .B1(n10957), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n10956), .C2(n17291), .A(n10955), .ZN(n17741) );
  NOR2_X1 U13900 ( .A1(n17742), .A2(n17741), .ZN(n10958) );
  NOR2_X1 U13901 ( .A1(n10959), .A2(n10958), .ZN(n17730) );
  XNOR2_X1 U13902 ( .A(n18041), .B(n10960), .ZN(n17729) );
  NOR2_X1 U13903 ( .A1(n17730), .A2(n17729), .ZN(n17728) );
  XOR2_X1 U13904 ( .A(n10963), .B(n10962), .Z(n10965) );
  NOR2_X1 U13905 ( .A1(n10964), .A2(n10965), .ZN(n10966) );
  XNOR2_X1 U13906 ( .A(n10965), .B(n10964), .ZN(n17715) );
  XNOR2_X1 U13907 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n10967), .ZN(
        n17703) );
  XNOR2_X1 U13908 ( .A(n17264), .B(n10969), .ZN(n10971) );
  NOR2_X1 U13909 ( .A1(n10970), .A2(n10971), .ZN(n10972) );
  INV_X1 U13910 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18026) );
  XNOR2_X1 U13911 ( .A(n10971), .B(n10970), .ZN(n17696) );
  XOR2_X1 U13912 ( .A(n17261), .B(n10973), .Z(n10976) );
  NAND2_X1 U13913 ( .A1(n10975), .A2(n10976), .ZN(n17680) );
  NOR2_X1 U13914 ( .A1(n10974), .A2(n10978), .ZN(n10980) );
  INV_X1 U13915 ( .A(n10974), .ZN(n10979) );
  OR2_X1 U13916 ( .A1(n10976), .A2(n10975), .ZN(n17681) );
  OAI21_X1 U13917 ( .B1(n10979), .B2(n10978), .A(n17681), .ZN(n10977) );
  INV_X1 U13918 ( .A(n17965), .ZN(n12757) );
  NAND2_X1 U13919 ( .A1(n17804), .A2(n17549), .ZN(n17483) );
  NOR2_X1 U13920 ( .A1(n17765), .A2(n17483), .ZN(n17426) );
  NAND2_X1 U13921 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15522) );
  NOR2_X1 U13922 ( .A1(n15522), .A2(n16308), .ZN(n16327) );
  INV_X1 U13923 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n20944) );
  NAND2_X1 U13924 ( .A1(n16327), .A2(n20944), .ZN(n15595) );
  INV_X1 U13925 ( .A(n15595), .ZN(n10981) );
  INV_X1 U13926 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18714) );
  NAND2_X1 U13927 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17721) );
  INV_X1 U13928 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18765) );
  INV_X1 U13929 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18704) );
  OAI21_X1 U13930 ( .B1(n18765), .B2(n18714), .A(n18704), .ZN(n18756) );
  NAND4_X1 U13931 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17623) );
  INV_X1 U13932 ( .A(n17623), .ZN(n10982) );
  NAND2_X1 U13933 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16607) );
  INV_X1 U13934 ( .A(n16607), .ZN(n17600) );
  INV_X1 U13935 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17586) );
  INV_X1 U13936 ( .A(n17558), .ZN(n10984) );
  INV_X1 U13937 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17543) );
  INV_X1 U13938 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17506) );
  NAND3_X1 U13939 ( .A1(n17487), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17470) );
  INV_X1 U13940 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17469) );
  INV_X1 U13941 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17432) );
  INV_X1 U13942 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17403) );
  INV_X1 U13943 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16469) );
  XOR2_X1 U13944 ( .A(n13088), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16457) );
  NAND2_X1 U13945 ( .A1(n16310), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10985) );
  NOR2_X1 U13946 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18765), .ZN(n17520) );
  INV_X1 U13947 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17755) );
  NAND2_X1 U13948 ( .A1(n18765), .A2(n18714), .ZN(n18752) );
  NAND2_X1 U13949 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18094) );
  NOR2_X1 U13950 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18704), .ZN(
        n18728) );
  AOI21_X1 U13951 ( .B1(n18752), .B2(n18094), .A(n18728), .ZN(n18103) );
  NOR2_X1 U13952 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18103), .ZN(n18385) );
  INV_X1 U13953 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16436) );
  NOR3_X1 U13954 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16436), .ZN(n18441) );
  NAND2_X1 U13955 ( .A1(n18385), .A2(n18441), .ZN(n18201) );
  INV_X1 U13956 ( .A(n17612), .ZN(n17557) );
  INV_X1 U13957 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13107) );
  NOR2_X1 U13958 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17446), .ZN(
        n16311) );
  INV_X1 U13959 ( .A(n13098), .ZN(n13084) );
  INV_X1 U13960 ( .A(n17520), .ZN(n17593) );
  INV_X1 U13961 ( .A(n18201), .ZN(n18477) );
  NAND2_X1 U13962 ( .A1(n18477), .A2(n10985), .ZN(n16314) );
  OAI211_X1 U13963 ( .C1(n13084), .C2(n17593), .A(n17759), .B(n16314), .ZN(
        n16317) );
  NOR2_X1 U13964 ( .A1(n16311), .A2(n16317), .ZN(n16298) );
  NAND2_X1 U13965 ( .A1(n18714), .A2(n18704), .ZN(n18708) );
  NOR3_X1 U13966 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18708), .ZN(n13104) );
  NAND2_X1 U13967 ( .A1(n18050), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n15592) );
  OAI221_X1 U13968 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16300), .C1(
        n13107), .C2(n16298), .A(n15592), .ZN(n10986) );
  AOI21_X1 U13969 ( .B1(n17615), .B2(n16457), .A(n10986), .ZN(n10989) );
  NAND2_X1 U13970 ( .A1(n17804), .A2(n12759), .ZN(n15520) );
  INV_X1 U13971 ( .A(n15520), .ZN(n12749) );
  NAND2_X1 U13972 ( .A1(n12749), .A2(n17827), .ZN(n17772) );
  INV_X1 U13973 ( .A(n16327), .ZN(n15587) );
  NOR2_X1 U13974 ( .A1(n17772), .A2(n15587), .ZN(n16302) );
  INV_X1 U13975 ( .A(n17876), .ZN(n17553) );
  NAND2_X1 U13976 ( .A1(n17969), .A2(n17553), .ZN(n17909) );
  NOR2_X1 U13977 ( .A1(n17909), .A2(n15520), .ZN(n17770) );
  OAI22_X1 U13978 ( .A1(n16302), .A2(n17764), .B1(n16307), .B2(n17674), .ZN(
        n10987) );
  NAND2_X1 U13979 ( .A1(n10987), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U13980 ( .A1(n10993), .A2(n10992), .ZN(P3_U2800) );
  AND2_X2 U13981 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10997), .ZN(
        n10996) );
  AND2_X2 U13982 ( .A1(n13811), .A2(n13824), .ZN(n11106) );
  AOI22_X1 U13983 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11106), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11003) );
  INV_X1 U13984 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10994) );
  NOR2_X2 U13985 ( .A1(n10995), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11007) );
  AND2_X2 U13986 ( .A1(n10996), .A2(n13811), .ZN(n11172) );
  AND2_X2 U13987 ( .A1(n10999), .A2(n13811), .ZN(n11212) );
  AND2_X2 U13988 ( .A1(n11006), .A2(n10999), .ZN(n11219) );
  AOI22_X1 U13989 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11053), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13990 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U13991 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11036), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11010) );
  AND2_X2 U13992 ( .A1(n13811), .A2(n13581), .ZN(n11227) );
  AOI22_X1 U13993 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11009) );
  AND2_X2 U13994 ( .A1(n11007), .A2(n13581), .ZN(n11100) );
  AOI22_X1 U13995 ( .A1(n11205), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U13996 ( .A1(n11205), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U13997 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U13998 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U13999 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11106), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14000 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U14001 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11053), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14002 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11212), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11018) );
  INV_X1 U14003 ( .A(n11121), .ZN(n11034) );
  AOI22_X1 U14004 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14005 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11026) );
  CLKBUF_X3 U14006 ( .A(n11036), .Z(n11788) );
  AOI22_X1 U14007 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U14008 ( .A1(n11205), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11053), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U14009 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11106), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U14010 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11212), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14011 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14012 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U14013 ( .A1(n11034), .A2(n12686), .ZN(n11045) );
  NAND2_X1 U14014 ( .A1(n11826), .A2(n11116), .ZN(n11862) );
  AOI22_X1 U14015 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11107), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U14016 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U14017 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U14018 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14019 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11212), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U14020 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U14021 ( .A1(n11053), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n11210), .ZN(n11041) );
  NAND2_X1 U14022 ( .A1(n11045), .A2(n11152), .ZN(n12656) );
  NAND2_X1 U14023 ( .A1(n11047), .A2(n12686), .ZN(n12660) );
  NAND2_X1 U14024 ( .A1(n11046), .A2(n11129), .ZN(n11117) );
  OR2_X2 U14025 ( .A1(n13671), .A2(n11117), .ZN(n13649) );
  AND2_X2 U14026 ( .A1(n11131), .A2(n11135), .ZN(n12775) );
  AOI21_X1 U14027 ( .B1(n11105), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n11048), .ZN(n11052) );
  AOI22_X1 U14028 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11049) );
  NAND4_X1 U14029 ( .A1(n11052), .A2(n11051), .A3(n11050), .A4(n11049), .ZN(
        n11059) );
  AOI22_X1 U14030 ( .A1(n11106), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_13__3__SCAN_IN), .B2(n11107), .ZN(n11056) );
  AOI22_X1 U14031 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11212), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14032 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11053), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11054) );
  NAND4_X1 U14033 ( .A1(n11057), .A2(n11056), .A3(n11055), .A4(n11054), .ZN(
        n11058) );
  OR2_X2 U14034 ( .A1(n11059), .A2(n11058), .ZN(n11120) );
  NAND2_X1 U14035 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11063) );
  NAND2_X1 U14036 ( .A1(n11205), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11062) );
  NAND2_X1 U14037 ( .A1(n11712), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11061) );
  NAND2_X1 U14038 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11060) );
  NAND2_X1 U14039 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11067) );
  NAND2_X1 U14040 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11066) );
  NAND2_X1 U14041 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11065) );
  NAND2_X1 U14042 ( .A1(n11106), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11064) );
  NAND2_X1 U14043 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11071) );
  NAND2_X1 U14044 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11070) );
  NAND2_X1 U14045 ( .A1(n11212), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11069) );
  NAND2_X1 U14046 ( .A1(n11053), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11068) );
  NAND2_X1 U14047 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11075) );
  NAND2_X1 U14048 ( .A1(n11105), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11074) );
  NAND2_X1 U14049 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11073) );
  NAND2_X1 U14050 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11072) );
  NAND4_X4 U14051 ( .A1(n11079), .A2(n11078), .A3(n11077), .A4(n11076), .ZN(
        n11136) );
  NAND2_X2 U14052 ( .A1(n11120), .A2(n11136), .ZN(n11892) );
  NAND2_X1 U14053 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11083) );
  NAND2_X1 U14054 ( .A1(n11205), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11082) );
  NAND2_X1 U14055 ( .A1(n11712), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11081) );
  NAND2_X1 U14056 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11080) );
  NAND2_X1 U14057 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U14058 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11086) );
  NAND2_X1 U14059 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11085) );
  NAND2_X1 U14060 ( .A1(n11106), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11084) );
  NAND2_X1 U14061 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11091) );
  NAND2_X1 U14062 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11090) );
  NAND2_X1 U14063 ( .A1(n11212), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U14064 ( .A1(n11053), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11088) );
  NAND2_X1 U14065 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U14066 ( .A1(n11105), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11094) );
  NAND2_X1 U14067 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11093) );
  NAND2_X1 U14068 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11092) );
  AOI22_X1 U14069 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11103) );
  AOI22_X1 U14070 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11212), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14071 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U14072 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11106), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14073 ( .A1(n11241), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11108) );
  OAI22_X1 U14074 ( .A1(n11818), .A2(n11892), .B1(n13882), .B2(n9594), .ZN(
        n12702) );
  INV_X1 U14075 ( .A(n12702), .ZN(n13576) );
  NAND2_X1 U14076 ( .A1(n13882), .A2(n11136), .ZN(n13595) );
  OAI21_X1 U14077 ( .B1(n20800), .B2(n12686), .A(n13595), .ZN(n11113) );
  INV_X1 U14078 ( .A(n11113), .ZN(n11114) );
  INV_X1 U14079 ( .A(n11120), .ZN(n11115) );
  NAND2_X1 U14080 ( .A1(n11115), .A2(n19999), .ZN(n11867) );
  NAND2_X2 U14081 ( .A1(n11892), .A2(n11867), .ZN(n13622) );
  NAND2_X1 U14082 ( .A1(n13622), .A2(n11130), .ZN(n12695) );
  NAND3_X1 U14083 ( .A1(n11150), .A2(n9647), .A3(n9932), .ZN(n11805) );
  NAND2_X1 U14084 ( .A1(n12567), .A2(n11121), .ZN(n11119) );
  NAND2_X1 U14085 ( .A1(n11117), .A2(n13258), .ZN(n11118) );
  NAND2_X1 U14086 ( .A1(n11119), .A2(n11118), .ZN(n11128) );
  NAND2_X1 U14087 ( .A1(n11818), .A2(n11123), .ZN(n11124) );
  NAND2_X1 U14088 ( .A1(n11126), .A2(n11124), .ZN(n11125) );
  AOI22_X1 U14089 ( .A1(n11805), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11252), 
        .B2(n11156), .ZN(n11141) );
  NAND2_X1 U14090 ( .A1(n11126), .A2(n12775), .ZN(n11127) );
  NOR2_X1 U14091 ( .A1(n11128), .A2(n11127), .ZN(n12661) );
  NAND2_X1 U14092 ( .A1(n12661), .A2(n13875), .ZN(n13232) );
  NAND2_X1 U14093 ( .A1(n13232), .A2(n9657), .ZN(n12687) );
  INV_X1 U14094 ( .A(n12673), .ZN(n11133) );
  XNOR2_X1 U14095 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12670) );
  NAND2_X1 U14096 ( .A1(n13241), .A2(n11137), .ZN(n13577) );
  INV_X1 U14097 ( .A(n13577), .ZN(n11138) );
  OAI21_X1 U14098 ( .B1(n13235), .B2(n12670), .A(n12684), .ZN(n11139) );
  OR2_X2 U14099 ( .A1(n12687), .A2(n11139), .ZN(n11140) );
  NAND2_X2 U14100 ( .A1(n11140), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U14101 ( .A1(n11141), .A2(n11159), .ZN(n11164) );
  NAND2_X1 U14102 ( .A1(n11164), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11146) );
  AND2_X1 U14103 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11166) );
  INV_X1 U14104 ( .A(n11166), .ZN(n11143) );
  NAND2_X1 U14105 ( .A1(n20521), .A2(n20482), .ZN(n11142) );
  NAND2_X1 U14106 ( .A1(n11143), .A2(n11142), .ZN(n20392) );
  NOR2_X1 U14107 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15934) );
  NAND2_X1 U14108 ( .A1(n15934), .A2(n19998), .ZN(n12781) );
  NAND2_X1 U14109 ( .A1(n15944), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20687) );
  NAND2_X1 U14110 ( .A1(n20687), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11160) );
  OAI21_X1 U14111 ( .B1(n20392), .B2(n12781), .A(n11160), .ZN(n11144) );
  INV_X1 U14112 ( .A(n11144), .ZN(n11145) );
  NAND2_X1 U14113 ( .A1(n11146), .A2(n11145), .ZN(n11147) );
  NAND2_X1 U14114 ( .A1(n11164), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11149) );
  INV_X1 U14115 ( .A(n20687), .ZN(n15570) );
  MUX2_X1 U14116 ( .A(n15570), .B(n12781), .S(n20521), .Z(n11148) );
  NAND2_X1 U14117 ( .A1(n11149), .A2(n11148), .ZN(n11203) );
  INV_X1 U14118 ( .A(n11152), .ZN(n11153) );
  NAND2_X1 U14119 ( .A1(n15934), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19799) );
  AOI21_X1 U14120 ( .B1(n11153), .B2(n12607), .A(n19799), .ZN(n11155) );
  INV_X1 U14121 ( .A(n13875), .ZN(n12681) );
  NAND2_X1 U14122 ( .A1(n13440), .A2(n11126), .ZN(n11154) );
  OR2_X1 U14123 ( .A1(n11134), .A2(n11116), .ZN(n12703) );
  NAND2_X1 U14124 ( .A1(n11156), .A2(n13875), .ZN(n12699) );
  INV_X1 U14125 ( .A(n11256), .ZN(n11158) );
  INV_X1 U14126 ( .A(n11159), .ZN(n11162) );
  NAND2_X1 U14127 ( .A1(n11160), .A2(n10997), .ZN(n11161) );
  NAND2_X1 U14128 ( .A1(n11162), .A2(n11161), .ZN(n11163) );
  NAND2_X1 U14129 ( .A1(n11165), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11168) );
  NAND2_X1 U14130 ( .A1(n11166), .A2(n20394), .ZN(n20434) );
  OAI21_X1 U14131 ( .B1(n11166), .B2(n20394), .A(n20434), .ZN(n20007) );
  INV_X1 U14132 ( .A(n12781), .ZN(n11186) );
  NAND2_X1 U14133 ( .A1(n20007), .A2(n11186), .ZN(n11167) );
  NAND2_X1 U14134 ( .A1(n11171), .A2(n13825), .ZN(n13582) );
  INV_X1 U14135 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U14136 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14137 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11175) );
  AOI22_X1 U14138 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11174) );
  AOI22_X1 U14139 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11173) );
  NAND4_X1 U14140 ( .A1(n11176), .A2(n11175), .A3(n11174), .A4(n11173), .ZN(
        n11182) );
  AOI22_X1 U14141 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14142 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14143 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U14144 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11177) );
  NAND4_X1 U14145 ( .A1(n11180), .A2(n11179), .A3(n11178), .A4(n11177), .ZN(
        n11181) );
  INV_X1 U14146 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11183) );
  OAI22_X1 U14147 ( .A1(n11845), .A2(n11183), .B1(n11189), .B2(n12578), .ZN(
        n11184) );
  NAND2_X1 U14148 ( .A1(n11165), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11188) );
  NOR3_X1 U14149 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20394), .A3(
        n20482), .ZN(n20285) );
  NAND2_X1 U14150 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20285), .ZN(
        n20276) );
  INV_X1 U14151 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20435) );
  NAND3_X1 U14152 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20614) );
  NOR2_X1 U14153 ( .A1(n20521), .A2(n20614), .ZN(n20658) );
  AOI21_X1 U14154 ( .B1(n20276), .B2(n20435), .A(n20658), .ZN(n20316) );
  AOI22_X1 U14155 ( .A1(n20316), .A2(n11186), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20687), .ZN(n11187) );
  NAND2_X1 U14156 ( .A1(n13808), .A2(n19998), .ZN(n11201) );
  AOI22_X1 U14157 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14158 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11762), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14159 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14160 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11190) );
  NAND4_X1 U14161 ( .A1(n11193), .A2(n11192), .A3(n11191), .A4(n11190), .ZN(
        n11199) );
  AOI22_X1 U14162 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14163 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14164 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14165 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11194) );
  NAND4_X1 U14166 ( .A1(n11197), .A2(n11196), .A3(n11195), .A4(n11194), .ZN(
        n11198) );
  OR2_X1 U14167 ( .A1(n11199), .A2(n11198), .ZN(n12585) );
  AOI22_X1 U14168 ( .A1(n11840), .A2(n12585), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11853), .ZN(n11200) );
  AOI22_X1 U14169 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11712), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14170 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14171 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14172 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11206) );
  NAND4_X1 U14173 ( .A1(n11209), .A2(n11208), .A3(n11207), .A4(n11206), .ZN(
        n11218) );
  BUF_X1 U14174 ( .A(n11210), .Z(n11221) );
  AOI22_X1 U14175 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14176 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14177 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14178 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11213) );
  NAND4_X1 U14179 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(
        n11217) );
  NAND2_X1 U14180 ( .A1(n12686), .A2(n12625), .ZN(n11235) );
  NOR2_X1 U14181 ( .A1(n11260), .A2(n12625), .ZN(n11240) );
  AOI22_X1 U14182 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11220), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14183 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n11221), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14184 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14185 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11222) );
  NAND4_X1 U14186 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11233) );
  AOI22_X1 U14187 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11784), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14188 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11211), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14189 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14190 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11228) );
  NAND4_X1 U14191 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n11232) );
  MUX2_X1 U14192 ( .A(n12622), .B(n11240), .S(n12565), .Z(n11234) );
  INV_X1 U14193 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11237) );
  AOI21_X1 U14194 ( .B1(n13882), .B2(n12565), .A(n19998), .ZN(n11236) );
  OAI211_X1 U14195 ( .C1(n11845), .C2(n11237), .A(n11236), .B(n11235), .ZN(
        n11318) );
  NAND2_X1 U14196 ( .A1(n11319), .A2(n11318), .ZN(n11239) );
  INV_X1 U14197 ( .A(n12622), .ZN(n11238) );
  INV_X1 U14198 ( .A(n11240), .ZN(n11255) );
  NAND2_X1 U14199 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11254) );
  AOI22_X1 U14200 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11786), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14201 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11762), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14202 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14203 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11242) );
  NAND4_X1 U14204 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n11251) );
  AOI22_X1 U14205 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14206 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14207 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14208 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11246) );
  NAND4_X1 U14209 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n11250) );
  NAND2_X1 U14210 ( .A1(n11252), .A2(n12566), .ZN(n11253) );
  NAND2_X1 U14211 ( .A1(n11257), .A2(n11256), .ZN(n20522) );
  INV_X1 U14212 ( .A(n14423), .ZN(n11261) );
  INV_X1 U14213 ( .A(n12566), .ZN(n11259) );
  AOI21_X2 U14214 ( .B1(n11261), .B2(n19998), .A(n9908), .ZN(n12564) );
  NAND2_X1 U14215 ( .A1(n11308), .A2(n12564), .ZN(n11311) );
  INV_X1 U14216 ( .A(n11262), .ZN(n11263) );
  AOI22_X1 U14217 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14218 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14219 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14220 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11266) );
  NAND4_X1 U14221 ( .A1(n11269), .A2(n11268), .A3(n11267), .A4(n11266), .ZN(
        n11275) );
  AOI22_X1 U14222 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14223 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14224 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14225 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11270) );
  NAND4_X1 U14226 ( .A1(n11273), .A2(n11272), .A3(n11271), .A4(n11270), .ZN(
        n11274) );
  OR2_X1 U14227 ( .A1(n11275), .A2(n11274), .ZN(n12593) );
  NAND2_X1 U14228 ( .A1(n11840), .A2(n12593), .ZN(n11277) );
  NAND2_X1 U14229 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14230 ( .A1(n11277), .A2(n11276), .ZN(n11339) );
  AOI22_X1 U14231 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11786), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14232 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14233 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14234 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11278) );
  NAND4_X1 U14235 ( .A1(n11281), .A2(n11280), .A3(n11279), .A4(n11278), .ZN(
        n11287) );
  AOI22_X1 U14236 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14237 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14238 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14239 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11282) );
  NAND4_X1 U14240 ( .A1(n11285), .A2(n11284), .A3(n11283), .A4(n11282), .ZN(
        n11286) );
  OR2_X1 U14241 ( .A1(n11287), .A2(n11286), .ZN(n12604) );
  NAND2_X1 U14242 ( .A1(n11840), .A2(n12604), .ZN(n11289) );
  NAND2_X1 U14243 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11288) );
  NAND2_X1 U14244 ( .A1(n11289), .A2(n11288), .ZN(n11384) );
  NAND2_X1 U14245 ( .A1(n11387), .A2(n11384), .ZN(n11361) );
  NAND2_X1 U14246 ( .A1(n11290), .A2(n11361), .ZN(n12592) );
  NAND2_X1 U14247 ( .A1(n11291), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11481) );
  AND2_X1 U14248 ( .A1(n20689), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13122) );
  INV_X1 U14249 ( .A(n13122), .ZN(n11368) );
  INV_X1 U14250 ( .A(n11331), .ZN(n11292) );
  AND2_X1 U14251 ( .A1(n11345), .A2(n19856), .ZN(n11293) );
  OR2_X1 U14252 ( .A1(n11293), .A2(n11362), .ZN(n19852) );
  OR2_X1 U14253 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n11800) );
  NAND2_X1 U14254 ( .A1(n19852), .A2(n9602), .ZN(n11294) );
  OAI21_X1 U14255 ( .B1(n19856), .B2(n11368), .A(n11294), .ZN(n11295) );
  AOI21_X1 U14256 ( .B1(n13123), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11295), .ZN(
        n11296) );
  INV_X1 U14257 ( .A(n11296), .ZN(n11297) );
  NAND2_X1 U14258 ( .A1(n11300), .A2(n11299), .ZN(n11301) );
  NAND2_X1 U14259 ( .A1(n11302), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11343) );
  XNOR2_X1 U14260 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13666) );
  AOI21_X1 U14261 ( .B1(n9602), .B2(n13666), .A(n13122), .ZN(n11304) );
  NAND2_X1 U14262 ( .A1(n13123), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11303) );
  OAI211_X1 U14263 ( .C1(n11343), .C2(n11305), .A(n11304), .B(n11303), .ZN(
        n11306) );
  INV_X1 U14264 ( .A(n11306), .ZN(n11307) );
  INV_X1 U14265 ( .A(n12564), .ZN(n11310) );
  INV_X1 U14266 ( .A(n11308), .ZN(n11309) );
  NAND2_X1 U14267 ( .A1(n11310), .A2(n11309), .ZN(n11312) );
  NAND2_X1 U14268 ( .A1(n13840), .A2(n11495), .ZN(n11317) );
  INV_X1 U14269 ( .A(n11343), .ZN(n11313) );
  NAND2_X1 U14270 ( .A1(n11313), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11315) );
  AOI22_X1 U14271 ( .A1(n13123), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20689), .ZN(n11314) );
  AND2_X1 U14272 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  NAND2_X1 U14273 ( .A1(n11317), .A2(n11316), .ZN(n13524) );
  NAND2_X1 U14274 ( .A1(n12563), .A2(n11291), .ZN(n11320) );
  NAND2_X1 U14275 ( .A1(n11320), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13486) );
  INV_X1 U14276 ( .A(n13963), .ZN(n20123) );
  NAND2_X1 U14277 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20689), .ZN(
        n11324) );
  NAND2_X1 U14278 ( .A1(n11322), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11323) );
  OAI211_X1 U14279 ( .C1(n11343), .C2(n13652), .A(n11324), .B(n11323), .ZN(
        n11325) );
  AOI21_X1 U14280 ( .B1(n20123), .B2(n11495), .A(n11325), .ZN(n13487) );
  OR2_X1 U14281 ( .A1(n13486), .A2(n13487), .ZN(n13488) );
  NAND2_X1 U14282 ( .A1(n13487), .A2(n9602), .ZN(n11326) );
  NAND2_X1 U14283 ( .A1(n13488), .A2(n11326), .ZN(n13523) );
  NAND2_X1 U14284 ( .A1(n13524), .A2(n13523), .ZN(n13658) );
  INV_X1 U14285 ( .A(n13658), .ZN(n11327) );
  NAND2_X1 U14286 ( .A1(n13656), .A2(n11327), .ZN(n13661) );
  NAND2_X1 U14287 ( .A1(n13122), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13657) );
  NAND2_X1 U14288 ( .A1(n13661), .A2(n13657), .ZN(n13731) );
  INV_X1 U14289 ( .A(n11346), .ZN(n11334) );
  INV_X1 U14290 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14291 ( .A1(n11332), .A2(n11331), .ZN(n11333) );
  NAND2_X1 U14292 ( .A1(n11334), .A2(n11333), .ZN(n13896) );
  AOI22_X1 U14293 ( .A1(n13896), .A2(n9602), .B1(n13122), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11336) );
  NAND2_X1 U14294 ( .A1(n13123), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11335) );
  OAI211_X1 U14295 ( .C1(n11343), .C2(n11330), .A(n11336), .B(n11335), .ZN(
        n11337) );
  INV_X1 U14296 ( .A(n11337), .ZN(n11338) );
  XNOR2_X1 U14297 ( .A(n11340), .B(n11339), .ZN(n12583) );
  INV_X1 U14298 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13828) );
  NAND2_X1 U14299 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14300 ( .A1(n13123), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11341) );
  OAI211_X1 U14301 ( .C1(n11343), .C2(n13828), .A(n11342), .B(n11341), .ZN(
        n11344) );
  NAND2_X1 U14302 ( .A1(n11344), .A2(n11800), .ZN(n11348) );
  OAI21_X1 U14303 ( .B1(n11346), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11345), .ZN(n19952) );
  NAND2_X1 U14304 ( .A1(n19952), .A2(n9602), .ZN(n11347) );
  NAND2_X1 U14305 ( .A1(n11348), .A2(n11347), .ZN(n11349) );
  NAND2_X1 U14306 ( .A1(n13795), .A2(n13796), .ZN(n13794) );
  AOI22_X1 U14307 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14308 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14309 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14310 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11350) );
  NAND4_X1 U14311 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n11360) );
  AOI22_X1 U14312 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11358) );
  INV_X1 U14313 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U14314 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14315 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14316 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11354), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11355) );
  NAND4_X1 U14317 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11359) );
  OR2_X1 U14318 ( .A1(n11360), .A2(n11359), .ZN(n12612) );
  AOI22_X1 U14319 ( .A1(n11840), .A2(n12612), .B1(n11853), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11383) );
  INV_X1 U14320 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13868) );
  NOR2_X1 U14321 ( .A1(n11362), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11363) );
  OR2_X1 U14322 ( .A1(n11391), .A2(n11363), .ZN(n19843) );
  AOI22_X1 U14323 ( .A1(n19843), .A2(n9602), .B1(n13122), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11364) );
  OAI21_X1 U14324 ( .B1(n11687), .B2(n13868), .A(n11364), .ZN(n11365) );
  INV_X1 U14325 ( .A(n13865), .ZN(n11366) );
  INV_X1 U14326 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11367) );
  NOR2_X1 U14327 ( .A1(n11368), .A2(n11367), .ZN(n11369) );
  AOI21_X1 U14328 ( .B1(n13123), .B2(P1_EAX_REG_8__SCAN_IN), .A(n11369), .ZN(
        n11382) );
  XNOR2_X1 U14329 ( .A(n11395), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14655) );
  NAND2_X1 U14330 ( .A1(n14655), .A2(n9602), .ZN(n11381) );
  AOI22_X1 U14331 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11786), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14332 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11756), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14333 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11788), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14334 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11370) );
  NAND4_X1 U14335 ( .A1(n11373), .A2(n11372), .A3(n11371), .A4(n11370), .ZN(
        n11379) );
  AOI22_X1 U14336 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11220), .B1(
        n11762), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14337 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11211), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14338 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11221), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14339 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11374) );
  NAND4_X1 U14340 ( .A1(n11377), .A2(n11376), .A3(n11375), .A4(n11374), .ZN(
        n11378) );
  OAI21_X1 U14341 ( .B1(n11379), .B2(n11378), .A(n11495), .ZN(n11380) );
  AND3_X1 U14342 ( .A1(n11382), .A2(n11381), .A3(n11380), .ZN(n14403) );
  INV_X1 U14343 ( .A(n11383), .ZN(n11385) );
  AND2_X1 U14344 ( .A1(n11385), .A2(n11384), .ZN(n11386) );
  NAND2_X1 U14345 ( .A1(n11840), .A2(n12625), .ZN(n11389) );
  NAND2_X1 U14346 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U14347 ( .A1(n11389), .A2(n11388), .ZN(n11390) );
  INV_X1 U14348 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14540) );
  NOR2_X1 U14349 ( .A1(n11391), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11392) );
  OR2_X1 U14350 ( .A1(n11395), .A2(n11392), .ZN(n19830) );
  AOI22_X1 U14351 ( .A1(n19830), .A2(n9602), .B1(n13122), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11393) );
  OAI21_X1 U14352 ( .B1(n11687), .B2(n14540), .A(n11393), .ZN(n11394) );
  XNOR2_X1 U14353 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11420), .ZN(
        n19819) );
  AOI22_X1 U14354 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14355 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14356 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11712), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14357 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11396) );
  NAND4_X1 U14358 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(
        n11405) );
  AOI22_X1 U14359 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14360 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14361 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14362 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11400) );
  NAND4_X1 U14363 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n11404) );
  OR2_X1 U14364 ( .A1(n11405), .A2(n11404), .ZN(n11406) );
  AOI22_X1 U14365 ( .A1(n11495), .A2(n11406), .B1(n13122), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11408) );
  NAND2_X1 U14366 ( .A1(n13123), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11407) );
  OAI211_X1 U14367 ( .C1(n19819), .C2(n11800), .A(n11408), .B(n11407), .ZN(
        n13862) );
  AOI22_X1 U14368 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14369 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14370 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14371 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11409) );
  NAND4_X1 U14372 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n11418) );
  AOI22_X1 U14373 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14374 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14375 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14376 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11413) );
  NAND4_X1 U14377 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11417) );
  NOR2_X1 U14378 ( .A1(n11418), .A2(n11417), .ZN(n11423) );
  INV_X1 U14379 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11419) );
  XNOR2_X1 U14380 ( .A(n11424), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14647) );
  NAND2_X1 U14381 ( .A1(n14647), .A2(n9602), .ZN(n11422) );
  AOI22_X1 U14382 ( .A1(n13123), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13122), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11421) );
  OAI211_X1 U14383 ( .C1(n11423), .C2(n11481), .A(n11422), .B(n11421), .ZN(
        n13971) );
  NAND2_X1 U14384 ( .A1(n11322), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11427) );
  OAI21_X1 U14385 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11425), .A(
        n11463), .ZN(n15792) );
  AOI22_X1 U14386 ( .A1(n9602), .A2(n15792), .B1(n13122), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11426) );
  NAND2_X1 U14387 ( .A1(n11427), .A2(n11426), .ZN(n14117) );
  AOI22_X1 U14388 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14389 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14390 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14391 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11428) );
  NAND4_X1 U14392 ( .A1(n11431), .A2(n11430), .A3(n11429), .A4(n11428), .ZN(
        n11437) );
  AOI22_X1 U14393 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14394 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14395 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14396 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11432) );
  NAND4_X1 U14397 ( .A1(n11435), .A2(n11434), .A3(n11433), .A4(n11432), .ZN(
        n11436) );
  OR2_X1 U14398 ( .A1(n11437), .A2(n11436), .ZN(n11438) );
  INV_X1 U14399 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15702) );
  XNOR2_X1 U14400 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11478), .ZN(
        n14638) );
  AOI22_X1 U14401 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11762), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14402 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14403 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14404 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11439) );
  NAND4_X1 U14405 ( .A1(n11442), .A2(n11441), .A3(n11440), .A4(n11439), .ZN(
        n11448) );
  AOI22_X1 U14406 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14407 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14408 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14409 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11443) );
  NAND4_X1 U14410 ( .A1(n11446), .A2(n11445), .A3(n11444), .A4(n11443), .ZN(
        n11447) );
  OR2_X1 U14411 ( .A1(n11448), .A2(n11447), .ZN(n11449) );
  AOI22_X1 U14412 ( .A1(n11495), .A2(n11449), .B1(n13122), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11451) );
  NAND2_X1 U14413 ( .A1(n13123), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11450) );
  OAI211_X1 U14414 ( .C1(n14638), .C2(n11800), .A(n11451), .B(n11450), .ZN(
        n14122) );
  INV_X1 U14415 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14183) );
  AOI22_X1 U14416 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14417 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14418 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14419 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11452) );
  NAND4_X1 U14420 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11461) );
  AOI22_X1 U14421 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14422 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14423 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14424 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11456) );
  NAND4_X1 U14425 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11460) );
  OR2_X1 U14426 ( .A1(n11461), .A2(n11460), .ZN(n11462) );
  NAND2_X1 U14427 ( .A1(n11495), .A2(n11462), .ZN(n11466) );
  XNOR2_X1 U14428 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11463), .ZN(
        n15780) );
  INV_X1 U14429 ( .A(n15780), .ZN(n11464) );
  AOI22_X1 U14430 ( .A1(n13122), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n9602), .B2(n11464), .ZN(n11465) );
  OAI211_X1 U14431 ( .C1(n11687), .C2(n14183), .A(n11466), .B(n11465), .ZN(
        n14121) );
  NAND2_X1 U14432 ( .A1(n14122), .A2(n14121), .ZN(n11467) );
  AOI22_X1 U14433 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11762), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14434 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14435 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14436 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11468) );
  NAND4_X1 U14437 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11477) );
  AOI22_X1 U14438 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14439 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14440 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14441 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11472) );
  NAND4_X1 U14442 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n11476) );
  NOR2_X1 U14443 ( .A1(n11477), .A2(n11476), .ZN(n11482) );
  INV_X1 U14444 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14129) );
  XNOR2_X1 U14445 ( .A(n11483), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15692) );
  NAND2_X1 U14446 ( .A1(n15692), .A2(n9602), .ZN(n11480) );
  AOI22_X1 U14447 ( .A1(n13123), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n13122), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11479) );
  OAI211_X1 U14448 ( .C1(n11482), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        n14066) );
  XOR2_X1 U14449 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11498), .Z(
        n15775) );
  AOI22_X1 U14450 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14451 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14452 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14453 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11484) );
  NAND4_X1 U14454 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(
        n11493) );
  AOI22_X1 U14455 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11762), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14456 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14457 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14458 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11488) );
  NAND4_X1 U14459 ( .A1(n11491), .A2(n11490), .A3(n11489), .A4(n11488), .ZN(
        n11492) );
  OR2_X1 U14460 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  AOI22_X1 U14461 ( .A1(n11495), .A2(n11494), .B1(n13122), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U14462 ( .A1(n11322), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11496) );
  OAI211_X1 U14463 ( .C1(n15775), .C2(n11800), .A(n11497), .B(n11496), .ZN(
        n14143) );
  INV_X1 U14464 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11499) );
  XNOR2_X1 U14465 ( .A(n11514), .B(n11499), .ZN(n15765) );
  INV_X1 U14466 ( .A(n13649), .ZN(n15542) );
  NAND2_X1 U14467 ( .A1(n15542), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14468 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11786), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14469 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14470 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11785), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14471 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11500) );
  NAND4_X1 U14472 ( .A1(n11503), .A2(n11502), .A3(n11501), .A4(n11500), .ZN(
        n11509) );
  AOI22_X1 U14473 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11221), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14474 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n11756), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14475 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n11784), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14476 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11504) );
  NAND4_X1 U14477 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n11508) );
  NOR2_X1 U14478 ( .A1(n11509), .A2(n11508), .ZN(n11512) );
  AOI21_X1 U14479 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n11499), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11510) );
  AOI21_X1 U14480 ( .B1(n11322), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11510), .ZN(
        n11511) );
  OAI21_X1 U14481 ( .B1(n11773), .B2(n11512), .A(n11511), .ZN(n11513) );
  OAI21_X1 U14482 ( .B1(n15765), .B2(n11800), .A(n11513), .ZN(n14207) );
  XNOR2_X1 U14483 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11531), .ZN(
        n15760) );
  INV_X1 U14484 ( .A(n15760), .ZN(n11528) );
  AOI22_X1 U14485 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11107), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14486 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14487 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14488 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11515) );
  NAND4_X1 U14489 ( .A1(n11518), .A2(n11517), .A3(n11516), .A4(n11515), .ZN(
        n11524) );
  AOI22_X1 U14490 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11786), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14491 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14492 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14493 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11519) );
  NAND4_X1 U14494 ( .A1(n11522), .A2(n11521), .A3(n11520), .A4(n11519), .ZN(
        n11523) );
  NOR2_X1 U14495 ( .A1(n11524), .A2(n11523), .ZN(n11526) );
  AOI22_X1 U14496 ( .A1(n13123), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13122), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11525) );
  OAI21_X1 U14497 ( .B1(n11773), .B2(n11526), .A(n11525), .ZN(n11527) );
  AOI21_X1 U14498 ( .B1(n11528), .B2(n9602), .A(n11527), .ZN(n14389) );
  NAND2_X1 U14499 ( .A1(n14386), .A2(n11529), .ZN(n14373) );
  INV_X1 U14500 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11530) );
  INV_X1 U14501 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11532) );
  XNOR2_X1 U14502 ( .A(n11563), .B(n11532), .ZN(n14611) );
  NAND2_X1 U14503 ( .A1(n14611), .A2(n9602), .ZN(n11548) );
  AOI22_X1 U14504 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14505 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14506 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14507 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11533) );
  NAND4_X1 U14508 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11544) );
  AOI22_X1 U14509 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14510 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11541) );
  AOI21_X1 U14511 ( .B1(n11739), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A(n9602), .ZN(n11538) );
  NAND2_X1 U14512 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11537) );
  AND2_X1 U14513 ( .A1(n11538), .A2(n11537), .ZN(n11540) );
  AOI22_X1 U14514 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11539) );
  NAND4_X1 U14515 ( .A1(n11542), .A2(n11541), .A3(n11540), .A4(n11539), .ZN(
        n11543) );
  NAND2_X1 U14516 ( .A1(n11773), .A2(n11800), .ZN(n11612) );
  OAI21_X1 U14517 ( .B1(n11544), .B2(n11543), .A(n11612), .ZN(n11546) );
  AOI22_X1 U14518 ( .A1(n13123), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20689), .ZN(n11545) );
  NAND2_X1 U14519 ( .A1(n11546), .A2(n11545), .ZN(n11547) );
  NAND2_X1 U14520 ( .A1(n11548), .A2(n11547), .ZN(n14374) );
  AOI22_X1 U14521 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14522 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11107), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14523 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14524 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11549) );
  NAND4_X1 U14525 ( .A1(n11552), .A2(n11551), .A3(n11550), .A4(n11549), .ZN(
        n11558) );
  AOI22_X1 U14526 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14527 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14528 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14529 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11553) );
  NAND4_X1 U14530 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n11557) );
  NOR2_X1 U14531 ( .A1(n11558), .A2(n11557), .ZN(n11562) );
  INV_X1 U14532 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20359) );
  OAI21_X1 U14533 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20359), .A(
        n20689), .ZN(n11559) );
  INV_X1 U14534 ( .A(n11559), .ZN(n11560) );
  AOI21_X1 U14535 ( .B1(n11322), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11560), .ZN(
        n11561) );
  OAI21_X1 U14536 ( .B1(n11773), .B2(n11562), .A(n11561), .ZN(n11566) );
  OAI21_X1 U14537 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11564), .A(
        n11598), .ZN(n15759) );
  OR2_X1 U14538 ( .A1(n11800), .A2(n15759), .ZN(n11565) );
  AND2_X1 U14539 ( .A1(n11566), .A2(n11565), .ZN(n14456) );
  AOI22_X1 U14540 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14541 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14542 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11570) );
  AOI21_X1 U14543 ( .B1(n11787), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A(n9602), .ZN(n11568) );
  NAND2_X1 U14544 ( .A1(n11620), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11567) );
  AND2_X1 U14545 ( .A1(n11568), .A2(n11567), .ZN(n11569) );
  NAND4_X1 U14546 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(
        n11578) );
  AOI22_X1 U14547 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11784), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14548 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14549 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14550 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11573) );
  NAND4_X1 U14551 ( .A1(n11576), .A2(n11575), .A3(n11574), .A4(n11573), .ZN(
        n11577) );
  OR2_X1 U14552 ( .A1(n11578), .A2(n11577), .ZN(n11579) );
  NAND2_X1 U14553 ( .A1(n11612), .A2(n11579), .ZN(n11582) );
  AOI22_X1 U14554 ( .A1(n13123), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20689), .ZN(n11581) );
  XNOR2_X1 U14555 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11598), .ZN(
        n15750) );
  AND2_X1 U14556 ( .A1(n9602), .A2(n15750), .ZN(n11580) );
  AOI21_X1 U14557 ( .B1(n11582), .B2(n11581), .A(n11580), .ZN(n14454) );
  AOI22_X1 U14558 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14559 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14560 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14561 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11583) );
  NAND4_X1 U14562 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n11592) );
  AOI22_X1 U14563 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14564 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14565 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14566 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11587) );
  NAND4_X1 U14567 ( .A1(n11590), .A2(n11589), .A3(n11588), .A4(n11587), .ZN(
        n11591) );
  NOR2_X1 U14568 ( .A1(n11592), .A2(n11591), .ZN(n11596) );
  NAND2_X1 U14569 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U14570 ( .A1(n11800), .A2(n11593), .ZN(n11594) );
  AOI21_X1 U14571 ( .B1(n11322), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11594), .ZN(
        n11595) );
  OAI21_X1 U14572 ( .B1(n11773), .B2(n11596), .A(n11595), .ZN(n11601) );
  INV_X1 U14573 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11597) );
  OAI21_X1 U14574 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11599), .A(
        n11645), .ZN(n15749) );
  OR2_X1 U14575 ( .A1(n11800), .A2(n15749), .ZN(n11600) );
  NAND2_X1 U14576 ( .A1(n11601), .A2(n11600), .ZN(n14444) );
  AOI22_X1 U14577 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11107), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14578 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14579 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14580 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14581 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11614) );
  AOI22_X1 U14582 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14583 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14584 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11609) );
  AOI21_X1 U14585 ( .B1(n11787), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A(n9602), .ZN(n11607) );
  NAND2_X1 U14586 ( .A1(n11620), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11606) );
  AND2_X1 U14587 ( .A1(n11607), .A2(n11606), .ZN(n11608) );
  NAND4_X1 U14588 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11613) );
  OAI21_X1 U14589 ( .B1(n11614), .B2(n11613), .A(n11612), .ZN(n11616) );
  AOI22_X1 U14590 ( .A1(n13123), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20689), .ZN(n11615) );
  NAND2_X1 U14591 ( .A1(n11616), .A2(n11615), .ZN(n11618) );
  XNOR2_X1 U14592 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n11645), .ZN(
        n15634) );
  NAND2_X1 U14593 ( .A1(n15634), .A2(n9602), .ZN(n11617) );
  NAND2_X1 U14594 ( .A1(n11618), .A2(n11617), .ZN(n14437) );
  AOI22_X1 U14595 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11107), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14596 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14597 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13810), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14598 ( .A1(n11620), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11621) );
  NAND4_X1 U14599 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11630) );
  AOI22_X1 U14600 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11786), .B1(
        n11784), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14601 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n11220), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U14602 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n11221), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14603 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11625) );
  NAND4_X1 U14604 ( .A1(n11628), .A2(n11627), .A3(n11626), .A4(n11625), .ZN(
        n11629) );
  NOR2_X1 U14605 ( .A1(n11630), .A2(n11629), .ZN(n11650) );
  AOI22_X1 U14606 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14607 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14608 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14609 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11631) );
  NAND4_X1 U14610 ( .A1(n11634), .A2(n11633), .A3(n11632), .A4(n11631), .ZN(
        n11640) );
  AOI22_X1 U14611 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11712), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14612 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14613 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14614 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11635) );
  NAND4_X1 U14615 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11639) );
  NOR2_X1 U14616 ( .A1(n11640), .A2(n11639), .ZN(n11649) );
  XNOR2_X1 U14617 ( .A(n11650), .B(n11649), .ZN(n11644) );
  NAND2_X1 U14618 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11641) );
  NAND2_X1 U14619 ( .A1(n11800), .A2(n11641), .ZN(n11642) );
  AOI21_X1 U14620 ( .B1(n11322), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11642), .ZN(
        n11643) );
  OAI21_X1 U14621 ( .B1(n11644), .B2(n11773), .A(n11643), .ZN(n11648) );
  INV_X1 U14622 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15630) );
  OAI21_X1 U14623 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n11646), .A(
        n11669), .ZN(n15744) );
  OR2_X1 U14624 ( .A1(n11800), .A2(n15744), .ZN(n11647) );
  NAND2_X1 U14625 ( .A1(n11648), .A2(n11647), .ZN(n14359) );
  NOR2_X1 U14626 ( .A1(n11650), .A2(n11649), .ZN(n11684) );
  AOI22_X1 U14627 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14628 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14629 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14630 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14631 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11660) );
  AOI22_X1 U14632 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11712), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14633 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14634 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11656) );
  INV_X1 U14635 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n20886) );
  AOI22_X1 U14636 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11655) );
  NAND4_X1 U14637 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(
        n11659) );
  OR2_X1 U14638 ( .A1(n11660), .A2(n11659), .ZN(n11683) );
  INV_X1 U14639 ( .A(n11683), .ZN(n11661) );
  XNOR2_X1 U14640 ( .A(n11684), .B(n11661), .ZN(n11662) );
  INV_X1 U14641 ( .A(n11773), .ZN(n11797) );
  NAND2_X1 U14642 ( .A1(n11662), .A2(n11797), .ZN(n11667) );
  NAND2_X1 U14643 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11663) );
  NAND2_X1 U14644 ( .A1(n11800), .A2(n11663), .ZN(n11664) );
  AOI21_X1 U14645 ( .B1(n11322), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11664), .ZN(
        n11666) );
  XNOR2_X1 U14646 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n11669), .ZN(
        n14594) );
  AND2_X1 U14647 ( .A1(n9602), .A2(n14594), .ZN(n11665) );
  AOI21_X1 U14648 ( .B1(n11667), .B2(n11666), .A(n11665), .ZN(n14349) );
  NAND2_X1 U14649 ( .A1(n14348), .A2(n14349), .ZN(n14347) );
  INV_X1 U14650 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11668) );
  OR2_X1 U14651 ( .A1(n11670), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11671) );
  NAND2_X1 U14652 ( .A1(n11670), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U14653 ( .A1(n11671), .A2(n11725), .ZN(n15735) );
  AOI22_X1 U14654 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14655 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11105), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14656 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14657 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11673) );
  NAND4_X1 U14658 ( .A1(n11676), .A2(n11675), .A3(n11674), .A4(n11673), .ZN(
        n11682) );
  AOI22_X1 U14659 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11786), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14660 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14661 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14662 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14663 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11681) );
  NOR2_X1 U14664 ( .A1(n11682), .A2(n11681), .ZN(n11691) );
  NAND2_X1 U14665 ( .A1(n11684), .A2(n11683), .ZN(n11690) );
  XNOR2_X1 U14666 ( .A(n11691), .B(n11690), .ZN(n11685) );
  NOR2_X1 U14667 ( .A1(n11685), .A2(n11773), .ZN(n11689) );
  INV_X1 U14668 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14492) );
  NAND2_X1 U14669 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11686) );
  OAI211_X1 U14670 ( .C1(n11687), .C2(n14492), .A(n11800), .B(n11686), .ZN(
        n11688) );
  OAI22_X1 U14671 ( .A1(n15735), .A2(n11800), .B1(n11689), .B2(n11688), .ZN(
        n14491) );
  NOR2_X1 U14672 ( .A1(n11691), .A2(n11690), .ZN(n11720) );
  INV_X1 U14673 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20823) );
  AOI22_X1 U14674 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14675 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14676 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14677 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11692) );
  NAND4_X1 U14678 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11701) );
  AOI22_X1 U14679 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11712), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14680 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14681 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14682 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11696) );
  NAND4_X1 U14683 ( .A1(n11699), .A2(n11698), .A3(n11697), .A4(n11696), .ZN(
        n11700) );
  OR2_X1 U14684 ( .A1(n11701), .A2(n11700), .ZN(n11719) );
  XNOR2_X1 U14685 ( .A(n11720), .B(n11719), .ZN(n11705) );
  NAND2_X1 U14686 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11702) );
  NAND2_X1 U14687 ( .A1(n11800), .A2(n11702), .ZN(n11703) );
  AOI21_X1 U14688 ( .B1(n11322), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11703), .ZN(
        n11704) );
  OAI21_X1 U14689 ( .B1(n11705), .B2(n11773), .A(n11704), .ZN(n11707) );
  XNOR2_X1 U14690 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(n11725), .ZN(
        n14586) );
  NAND2_X1 U14691 ( .A1(n9602), .A2(n14586), .ZN(n11706) );
  NAND2_X1 U14692 ( .A1(n11707), .A2(n11706), .ZN(n14334) );
  AOI22_X1 U14693 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14694 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14695 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14696 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11708) );
  NAND4_X1 U14697 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11718) );
  AOI22_X1 U14698 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14699 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11712), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14700 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14701 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U14702 ( .A1(n11716), .A2(n11715), .A3(n11714), .A4(n11713), .ZN(
        n11717) );
  NOR2_X1 U14703 ( .A1(n11718), .A2(n11717), .ZN(n11733) );
  NAND2_X1 U14704 ( .A1(n11720), .A2(n11719), .ZN(n11732) );
  XNOR2_X1 U14705 ( .A(n11733), .B(n11732), .ZN(n11724) );
  NAND2_X1 U14706 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14707 ( .A1(n11800), .A2(n11721), .ZN(n11722) );
  AOI21_X1 U14708 ( .B1(n11322), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11722), .ZN(
        n11723) );
  OAI21_X1 U14709 ( .B1(n11724), .B2(n11773), .A(n11723), .ZN(n11731) );
  INV_X1 U14710 ( .A(n11725), .ZN(n11726) );
  INV_X1 U14711 ( .A(n11727), .ZN(n11728) );
  INV_X1 U14712 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14576) );
  NAND2_X1 U14713 ( .A1(n11728), .A2(n14576), .ZN(n11729) );
  AND2_X1 U14714 ( .A1(n11752), .A2(n11729), .ZN(n14580) );
  NAND2_X1 U14715 ( .A1(n14580), .A2(n9602), .ZN(n11730) );
  NOR2_X1 U14716 ( .A1(n11733), .A2(n11732), .ZN(n11770) );
  AOI22_X1 U14717 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14718 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14719 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14720 ( .A1(n11219), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14721 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11745) );
  INV_X1 U14722 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20813) );
  AOI22_X1 U14723 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14724 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13810), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14725 ( .A1(n11785), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14726 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11740) );
  NAND4_X1 U14727 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11744) );
  OR2_X1 U14728 ( .A1(n11745), .A2(n11744), .ZN(n11769) );
  XNOR2_X1 U14729 ( .A(n11770), .B(n11769), .ZN(n11749) );
  NAND2_X1 U14730 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11746) );
  NAND2_X1 U14731 ( .A1(n11800), .A2(n11746), .ZN(n11747) );
  AOI21_X1 U14732 ( .B1(n13123), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11747), .ZN(
        n11748) );
  OAI21_X1 U14733 ( .B1(n11749), .B2(n11773), .A(n11748), .ZN(n11751) );
  XNOR2_X1 U14734 ( .A(n11752), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14566) );
  NAND2_X1 U14735 ( .A1(n14566), .A2(n9602), .ZN(n11750) );
  NAND2_X1 U14736 ( .A1(n11751), .A2(n11750), .ZN(n14311) );
  INV_X1 U14737 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14568) );
  NAND2_X1 U14738 ( .A1(n11753), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13115) );
  INV_X1 U14739 ( .A(n11753), .ZN(n11754) );
  INV_X1 U14740 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14297) );
  NAND2_X1 U14741 ( .A1(n11754), .A2(n14297), .ZN(n11755) );
  NAND2_X1 U14742 ( .A1(n13115), .A2(n11755), .ZN(n14296) );
  AOI22_X1 U14743 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11756), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14744 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14745 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14746 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11757) );
  NAND4_X1 U14747 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n11768) );
  AOI22_X1 U14748 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14749 ( .A1(n11762), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U14750 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14751 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11779), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11763) );
  NAND4_X1 U14752 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n11767) );
  NOR2_X1 U14753 ( .A1(n11768), .A2(n11767), .ZN(n11778) );
  NAND2_X1 U14754 ( .A1(n11770), .A2(n11769), .ZN(n11777) );
  XNOR2_X1 U14755 ( .A(n11778), .B(n11777), .ZN(n11774) );
  AOI21_X1 U14756 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20689), .A(
        n9602), .ZN(n11772) );
  NAND2_X1 U14757 ( .A1(n13123), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11771) );
  OAI211_X1 U14758 ( .C1(n11774), .C2(n11773), .A(n11772), .B(n11771), .ZN(
        n11775) );
  OAI21_X1 U14759 ( .B1(n11800), .B2(n14296), .A(n11775), .ZN(n12779) );
  INV_X1 U14760 ( .A(n12779), .ZN(n11776) );
  NOR2_X1 U14761 ( .A1(n11778), .A2(n11777), .ZN(n11796) );
  AOI22_X1 U14762 ( .A1(n11210), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11219), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14763 ( .A1(n13810), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14764 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11620), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14765 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11672), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11780) );
  NAND4_X1 U14766 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11794) );
  AOI22_X1 U14767 ( .A1(n11784), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11762), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14768 ( .A1(n11756), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14769 ( .A1(n11786), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11785), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14770 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11787), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11789) );
  NAND4_X1 U14771 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11793) );
  NOR2_X1 U14772 ( .A1(n11794), .A2(n11793), .ZN(n11795) );
  XNOR2_X1 U14773 ( .A(n11796), .B(n11795), .ZN(n11798) );
  NAND2_X1 U14774 ( .A1(n11798), .A2(n11797), .ZN(n11804) );
  NAND2_X1 U14775 ( .A1(n20689), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U14776 ( .A1(n11800), .A2(n11799), .ZN(n11801) );
  AOI21_X1 U14777 ( .B1(n13123), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11801), .ZN(
        n11803) );
  XNOR2_X1 U14778 ( .A(n13115), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14547) );
  AND2_X1 U14779 ( .A1(n14547), .A2(n9602), .ZN(n11802) );
  OR2_X1 U14780 ( .A1(n13671), .A2(n13532), .ZN(n12658) );
  OR2_X1 U14781 ( .A1(n11805), .A2(n12658), .ZN(n13600) );
  XNOR2_X1 U14782 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U14783 ( .A1(n11825), .A2(n11824), .ZN(n11807) );
  NAND2_X1 U14784 ( .A1(n20482), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11806) );
  NAND2_X1 U14785 ( .A1(n11807), .A2(n11806), .ZN(n11836) );
  XNOR2_X1 U14786 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11835) );
  NAND2_X1 U14787 ( .A1(n11836), .A2(n11835), .ZN(n11809) );
  NAND2_X1 U14788 ( .A1(n20394), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U14789 ( .A1(n11809), .A2(n11808), .ZN(n11816) );
  XNOR2_X1 U14790 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11815) );
  NAND2_X1 U14791 ( .A1(n11816), .A2(n11815), .ZN(n11811) );
  NAND2_X1 U14792 ( .A1(n20435), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U14793 ( .A1(n11811), .A2(n11810), .ZN(n11849) );
  NOR2_X1 U14794 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13828), .ZN(
        n11812) );
  OR2_X1 U14795 ( .A1(n11849), .A2(n11812), .ZN(n11814) );
  INV_X1 U14796 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19993) );
  OR2_X1 U14797 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19993), .ZN(
        n11813) );
  AND2_X1 U14798 ( .A1(n11814), .A2(n11813), .ZN(n12669) );
  NAND2_X1 U14799 ( .A1(n11848), .A2(n12669), .ZN(n11861) );
  NAND2_X1 U14800 ( .A1(n12669), .A2(n11840), .ZN(n11859) );
  XNOR2_X1 U14801 ( .A(n11816), .B(n11815), .ZN(n12665) );
  INV_X1 U14802 ( .A(n11825), .ZN(n11817) );
  OAI21_X1 U14803 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20521), .A(
        n11817), .ZN(n11819) );
  NOR2_X1 U14804 ( .A1(n11838), .A2(n11819), .ZN(n11823) );
  INV_X1 U14805 ( .A(n11819), .ZN(n11821) );
  NAND2_X1 U14806 ( .A1(n11826), .A2(n19999), .ZN(n11820) );
  NAND2_X1 U14807 ( .A1(n11820), .A2(n13532), .ZN(n11837) );
  OAI211_X1 U14808 ( .C1(n13882), .C2(n11818), .A(n11821), .B(n11837), .ZN(
        n11822) );
  OAI21_X1 U14809 ( .B1(n11848), .B2(n11823), .A(n11822), .ZN(n11830) );
  INV_X1 U14810 ( .A(n11830), .ZN(n11834) );
  XNOR2_X1 U14811 ( .A(n11825), .B(n11824), .ZN(n12666) );
  NAND2_X1 U14812 ( .A1(n11826), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11828) );
  OAI21_X1 U14813 ( .B1(n11838), .B2(n13532), .A(n11828), .ZN(n11827) );
  AOI21_X1 U14814 ( .B1(n11853), .B2(n12666), .A(n11827), .ZN(n11831) );
  INV_X1 U14815 ( .A(n11831), .ZN(n11833) );
  AND2_X1 U14816 ( .A1(n11828), .A2(n11136), .ZN(n11829) );
  NAND2_X1 U14817 ( .A1(n11838), .A2(n11829), .ZN(n11850) );
  AOI22_X1 U14818 ( .A1(n12666), .A2(n11850), .B1(n11831), .B2(n11830), .ZN(
        n11832) );
  AOI21_X1 U14819 ( .B1(n11834), .B2(n11833), .A(n11832), .ZN(n11844) );
  XNOR2_X1 U14820 ( .A(n11836), .B(n11835), .ZN(n12664) );
  INV_X1 U14821 ( .A(n11837), .ZN(n11841) );
  NOR2_X1 U14822 ( .A1(n11838), .A2(n12664), .ZN(n11839) );
  AOI211_X1 U14823 ( .C1(n11853), .C2(n12664), .A(n11841), .B(n11839), .ZN(
        n11843) );
  NAND2_X1 U14824 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  OAI22_X1 U14825 ( .A1(n11844), .A2(n11843), .B1(n12664), .B2(n11842), .ZN(
        n11847) );
  NAND2_X1 U14826 ( .A1(n11845), .A2(n12665), .ZN(n11846) );
  AOI22_X1 U14827 ( .A1(n11848), .A2(n12665), .B1(n11847), .B2(n11846), .ZN(
        n11856) );
  OR3_X1 U14828 ( .A1(n11849), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n19993), .ZN(n11851) );
  NOR2_X1 U14829 ( .A1(n11853), .A2(n11851), .ZN(n11855) );
  INV_X1 U14830 ( .A(n11850), .ZN(n11852) );
  INV_X1 U14831 ( .A(n11851), .ZN(n12667) );
  NAND3_X1 U14832 ( .A1(n11853), .A2(n11852), .A3(n12667), .ZN(n11854) );
  OAI21_X1 U14833 ( .B1(n11856), .B2(n11855), .A(n11854), .ZN(n11857) );
  AOI21_X1 U14834 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19998), .A(
        n11857), .ZN(n11858) );
  NAND2_X1 U14835 ( .A1(n11859), .A2(n11858), .ZN(n11860) );
  OR2_X1 U14836 ( .A1(n20687), .A2(n19998), .ZN(n19796) );
  OR2_X1 U14837 ( .A1(n13601), .A2(n19796), .ZN(n11866) );
  INV_X1 U14838 ( .A(n19796), .ZN(n13240) );
  NAND3_X1 U14839 ( .A1(n14210), .A2(n12686), .A3(n13240), .ZN(n11863) );
  NOR2_X1 U14840 ( .A1(n11863), .A2(n11862), .ZN(n13242) );
  NAND3_X1 U14841 ( .A1(n13242), .A2(n13901), .A3(n11864), .ZN(n11865) );
  NAND2_X1 U14842 ( .A1(n19904), .A2(n11129), .ZN(n14470) );
  OR2_X1 U14843 ( .A1(n13901), .A2(n11867), .ZN(n11933) );
  NAND2_X1 U14844 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n9625), .ZN(
        n11868) );
  AND2_X1 U14845 ( .A1(n11933), .A2(n11868), .ZN(n11869) );
  NAND2_X1 U14846 ( .A1(n11870), .A2(n11869), .ZN(n11873) );
  NAND2_X1 U14847 ( .A1(n11867), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11872) );
  INV_X1 U14848 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13859) );
  NAND2_X1 U14849 ( .A1(n11928), .A2(n13859), .ZN(n11871) );
  NAND2_X1 U14850 ( .A1(n11872), .A2(n11871), .ZN(n13623) );
  MUX2_X1 U14851 ( .A(n11874), .B(n11867), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11877) );
  NAND2_X1 U14852 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n9625), .ZN(
        n11875) );
  AND2_X1 U14853 ( .A1(n11933), .A2(n11875), .ZN(n11876) );
  NAND2_X1 U14854 ( .A1(n11877), .A2(n11876), .ZN(n13933) );
  NAND2_X1 U14855 ( .A1(n13901), .A2(n11928), .ZN(n11952) );
  MUX2_X1 U14856 ( .A(n11952), .B(n11928), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11880) );
  OR2_X1 U14857 ( .A1(n13622), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11879) );
  NAND2_X1 U14858 ( .A1(n11880), .A2(n11879), .ZN(n13881) );
  INV_X1 U14859 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13942) );
  NAND2_X1 U14860 ( .A1(n11943), .A2(n13942), .ZN(n11885) );
  INV_X1 U14861 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19963) );
  NAND2_X1 U14862 ( .A1(n11867), .A2(n19963), .ZN(n11883) );
  OAI211_X1 U14863 ( .C1(n9625), .C2(P1_EBX_REG_4__SCAN_IN), .A(n11883), .B(
        n11928), .ZN(n11884) );
  OR2_X1 U14864 ( .A1(n13622), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11887) );
  MUX2_X1 U14865 ( .A(n11952), .B(n11928), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n11886) );
  AND2_X1 U14866 ( .A1(n11887), .A2(n11886), .ZN(n13850) );
  OR2_X1 U14867 ( .A1(n11952), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U14868 ( .A1(n11928), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11889) );
  OAI211_X1 U14869 ( .C1(n9625), .C2(P1_EBX_REG_7__SCAN_IN), .A(n11956), .B(
        n11889), .ZN(n11890) );
  AND2_X1 U14870 ( .A1(n11891), .A2(n11890), .ZN(n15903) );
  OR2_X1 U14871 ( .A1(n11874), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n11895) );
  INV_X1 U14872 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15900) );
  NAND2_X1 U14873 ( .A1(n11956), .A2(n15900), .ZN(n11893) );
  OAI211_X1 U14874 ( .C1(n9625), .C2(P1_EBX_REG_6__SCAN_IN), .A(n11893), .B(
        n11892), .ZN(n11894) );
  NAND2_X1 U14875 ( .A1(n11895), .A2(n11894), .ZN(n15915) );
  MUX2_X1 U14876 ( .A(n11874), .B(n11956), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11898) );
  NAND2_X1 U14877 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n9625), .ZN(
        n11897) );
  AND3_X1 U14878 ( .A1(n11898), .A2(n11933), .A3(n11897), .ZN(n14404) );
  MUX2_X1 U14879 ( .A(n11952), .B(n11928), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n11899) );
  OAI21_X1 U14880 ( .B1(n13622), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11899), .ZN(n13905) );
  INV_X1 U14881 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14049) );
  NAND2_X1 U14882 ( .A1(n11943), .A2(n14049), .ZN(n11903) );
  INV_X1 U14883 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11900) );
  NAND2_X1 U14884 ( .A1(n11956), .A2(n11900), .ZN(n11901) );
  OAI211_X1 U14885 ( .C1(n9625), .C2(P1_EBX_REG_10__SCAN_IN), .A(n11901), .B(
        n11928), .ZN(n11902) );
  AND2_X1 U14886 ( .A1(n11903), .A2(n11902), .ZN(n13975) );
  OR2_X1 U14887 ( .A1(n11952), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U14888 ( .A1(n11928), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11904) );
  OAI211_X1 U14889 ( .C1(n9625), .C2(P1_EBX_REG_11__SCAN_IN), .A(n11956), .B(
        n11904), .ZN(n11905) );
  AND2_X1 U14890 ( .A1(n11906), .A2(n11905), .ZN(n15708) );
  MUX2_X1 U14891 ( .A(n11952), .B(n11928), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11908) );
  OR2_X1 U14892 ( .A1(n13622), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11907) );
  AND2_X1 U14893 ( .A1(n11908), .A2(n11907), .ZN(n14126) );
  OR2_X1 U14894 ( .A1(n11874), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n11911) );
  INV_X1 U14895 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U14896 ( .A1(n11956), .A2(n14791), .ZN(n11909) );
  OAI211_X1 U14897 ( .C1(n9625), .C2(P1_EBX_REG_12__SCAN_IN), .A(n11909), .B(
        n11928), .ZN(n11910) );
  NAND2_X1 U14898 ( .A1(n11911), .A2(n11910), .ZN(n14793) );
  NAND2_X1 U14899 ( .A1(n14126), .A2(n14793), .ZN(n11912) );
  MUX2_X1 U14900 ( .A(n11874), .B(n11956), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11915) );
  INV_X1 U14901 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15852) );
  OAI21_X1 U14902 ( .B1(n13901), .B2(n15852), .A(n11933), .ZN(n11913) );
  INV_X1 U14903 ( .A(n11913), .ZN(n11914) );
  AND2_X1 U14904 ( .A1(n11915), .A2(n11914), .ZN(n14114) );
  OR2_X1 U14905 ( .A1(n11952), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n11918) );
  NAND2_X1 U14906 ( .A1(n11928), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11916) );
  OAI211_X1 U14907 ( .C1(n9625), .C2(P1_EBX_REG_15__SCAN_IN), .A(n11956), .B(
        n11916), .ZN(n11917) );
  AND2_X1 U14908 ( .A1(n11918), .A2(n11917), .ZN(n15681) );
  INV_X1 U14909 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15672) );
  NAND2_X1 U14910 ( .A1(n11943), .A2(n15672), .ZN(n11922) );
  INV_X1 U14911 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11919) );
  NAND2_X1 U14912 ( .A1(n11956), .A2(n11919), .ZN(n11920) );
  OAI211_X1 U14913 ( .C1(n9625), .C2(P1_EBX_REG_16__SCAN_IN), .A(n11920), .B(
        n11928), .ZN(n11921) );
  NAND2_X1 U14914 ( .A1(n11922), .A2(n11921), .ZN(n14208) );
  MUX2_X1 U14915 ( .A(n11952), .B(n11928), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11924) );
  OR2_X1 U14916 ( .A1(n13622), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U14917 ( .A1(n11924), .A2(n11923), .ZN(n14390) );
  INV_X1 U14918 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U14919 ( .A1(n11943), .A2(n14465), .ZN(n11927) );
  INV_X1 U14920 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15831) );
  NAND2_X1 U14921 ( .A1(n11956), .A2(n15831), .ZN(n11925) );
  OAI211_X1 U14922 ( .C1(n9625), .C2(P1_EBX_REG_18__SCAN_IN), .A(n11925), .B(
        n11928), .ZN(n11926) );
  AND2_X1 U14923 ( .A1(n11927), .A2(n11926), .ZN(n14380) );
  OR2_X1 U14924 ( .A1(n11952), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n11931) );
  NAND2_X1 U14925 ( .A1(n11928), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11929) );
  OAI211_X1 U14926 ( .C1(n9625), .C2(P1_EBX_REG_19__SCAN_IN), .A(n11956), .B(
        n11929), .ZN(n11930) );
  AND2_X1 U14927 ( .A1(n11931), .A2(n11930), .ZN(n14458) );
  MUX2_X1 U14928 ( .A(n11874), .B(n11956), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11935) );
  NAND2_X1 U14929 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n9625), .ZN(
        n11932) );
  AND2_X1 U14930 ( .A1(n11933), .A2(n11932), .ZN(n11934) );
  NAND2_X1 U14931 ( .A1(n11935), .A2(n11934), .ZN(n14451) );
  MUX2_X1 U14932 ( .A(n11952), .B(n11928), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11937) );
  OR2_X1 U14933 ( .A1(n13622), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U14934 ( .A1(n11937), .A2(n11936), .ZN(n14447) );
  INV_X1 U14935 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15631) );
  NAND2_X1 U14936 ( .A1(n11943), .A2(n15631), .ZN(n11940) );
  INV_X1 U14937 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14602) );
  NAND2_X1 U14938 ( .A1(n11956), .A2(n14602), .ZN(n11938) );
  OAI211_X1 U14939 ( .C1(n9625), .C2(P1_EBX_REG_22__SCAN_IN), .A(n11938), .B(
        n11928), .ZN(n11939) );
  AND2_X1 U14940 ( .A1(n11940), .A2(n11939), .ZN(n14438) );
  MUX2_X1 U14941 ( .A(n11952), .B(n11892), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11942) );
  OR2_X1 U14942 ( .A1(n13622), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U14943 ( .A1(n11942), .A2(n11941), .ZN(n14361) );
  INV_X1 U14944 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14352) );
  NAND2_X1 U14945 ( .A1(n11943), .A2(n14352), .ZN(n11946) );
  INV_X1 U14946 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U14947 ( .A1(n11956), .A2(n12646), .ZN(n11944) );
  OAI211_X1 U14948 ( .C1(n9625), .C2(P1_EBX_REG_24__SCAN_IN), .A(n11944), .B(
        n11928), .ZN(n11945) );
  NAND2_X1 U14949 ( .A1(n11946), .A2(n11945), .ZN(n14346) );
  OR2_X1 U14950 ( .A1(n11952), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n11949) );
  NAND2_X1 U14951 ( .A1(n11928), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11947) );
  OAI211_X1 U14952 ( .C1(n9625), .C2(P1_EBX_REG_25__SCAN_IN), .A(n11956), .B(
        n11947), .ZN(n11948) );
  NAND2_X1 U14953 ( .A1(n11949), .A2(n11948), .ZN(n15622) );
  MUX2_X1 U14954 ( .A(n11874), .B(n11956), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n11951) );
  NAND2_X1 U14955 ( .A1(n9625), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11950) );
  AND2_X1 U14956 ( .A1(n11951), .A2(n11950), .ZN(n14335) );
  OR2_X1 U14957 ( .A1(n11952), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U14958 ( .A1(n11928), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11953) );
  OAI211_X1 U14959 ( .C1(n9625), .C2(P1_EBX_REG_27__SCAN_IN), .A(n11956), .B(
        n11953), .ZN(n11954) );
  AND2_X1 U14960 ( .A1(n11955), .A2(n11954), .ZN(n14326) );
  AND2_X2 U14961 ( .A1(n14336), .A2(n14326), .ZN(n14328) );
  MUX2_X1 U14962 ( .A(n11874), .B(n11956), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11958) );
  NAND2_X1 U14963 ( .A1(n9625), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11957) );
  NAND2_X1 U14964 ( .A1(n11958), .A2(n11957), .ZN(n14307) );
  OR2_X1 U14965 ( .A1(n13622), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11960) );
  INV_X1 U14966 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14430) );
  NAND2_X1 U14967 ( .A1(n13901), .A2(n14430), .ZN(n11959) );
  NAND2_X1 U14968 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  OAI22_X1 U14969 ( .A1(n11961), .A2(n11878), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11874), .ZN(n14302) );
  INV_X1 U14970 ( .A(n11961), .ZN(n11962) );
  AND2_X1 U14971 ( .A1(n9625), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11963) );
  AOI21_X1 U14972 ( .B1(n13622), .B2(P1_EBX_REG_30__SCAN_IN), .A(n11963), .ZN(
        n12690) );
  NAND2_X1 U14973 ( .A1(n14210), .A2(n19904), .ZN(n14472) );
  NOR2_X1 U14974 ( .A1(n14287), .A2(n14472), .ZN(n11965) );
  INV_X1 U14975 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14292) );
  NOR2_X1 U14976 ( .A1(n19904), .A2(n14292), .ZN(n11964) );
  NOR2_X1 U14977 ( .A1(n11965), .A2(n11964), .ZN(n11966) );
  OAI21_X1 U14978 ( .B1(n14553), .B2(n14470), .A(n11966), .ZN(P1_U2842) );
  INV_X1 U14979 ( .A(n15402), .ZN(n13574) );
  NAND2_X1 U14980 ( .A1(n15393), .A2(n13574), .ZN(n11996) );
  NAND2_X1 U14981 ( .A1(n11967), .A2(n15402), .ZN(n11990) );
  OAI22_X1 U14983 ( .A1(n12010), .A2(n19543), .B1(n12196), .B2(n11968), .ZN(
        n11972) );
  INV_X1 U14984 ( .A(n11974), .ZN(n13617) );
  NAND2_X1 U14985 ( .A1(n11969), .A2(n15402), .ZN(n11992) );
  OR2_X2 U14986 ( .A1(n11991), .A2(n11992), .ZN(n12185) );
  OAI22_X1 U14987 ( .A1(n11970), .A2(n12185), .B1(n12198), .B2(n20841), .ZN(
        n11971) );
  NOR2_X1 U14988 ( .A1(n11972), .A2(n11971), .ZN(n12006) );
  OR2_X2 U14989 ( .A1(n11998), .A2(n11990), .ZN(n19126) );
  OAI22_X1 U14990 ( .A1(n11976), .A2(n19126), .B1(n12186), .B2(n11975), .ZN(
        n11982) );
  OR2_X2 U14991 ( .A1(n9607), .A2(n11996), .ZN(n12187) );
  INV_X1 U14992 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11980) );
  INV_X1 U14993 ( .A(n11983), .ZN(n11978) );
  OAI22_X1 U14994 ( .A1(n12187), .A2(n11980), .B1(n19508), .B2(n11979), .ZN(
        n11981) );
  NOR2_X1 U14995 ( .A1(n11982), .A2(n11981), .ZN(n12005) );
  OR2_X2 U14996 ( .A1(n9607), .A2(n11997), .ZN(n12181) );
  INV_X1 U14997 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11987) );
  OAI22_X1 U14998 ( .A1(n12181), .A2(n11987), .B1(n12190), .B2(n11986), .ZN(
        n11988) );
  NOR2_X1 U14999 ( .A1(n11989), .A2(n11988), .ZN(n12004) );
  INV_X1 U15000 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11995) );
  OR2_X2 U15001 ( .A1(n11991), .A2(n11990), .ZN(n12182) );
  INV_X1 U15002 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11994) );
  OAI22_X1 U15003 ( .A1(n11995), .A2(n12182), .B1(n12195), .B2(n11994), .ZN(
        n12002) );
  NOR2_X1 U15004 ( .A1(n12002), .A2(n12001), .ZN(n12003) );
  NAND4_X1 U15005 ( .A1(n12006), .A2(n12004), .A3(n12005), .A4(n12003), .ZN(
        n12007) );
  NAND2_X1 U15006 ( .A1(n12007), .A2(n13571), .ZN(n12025) );
  INV_X1 U15007 ( .A(n12008), .ZN(n12045) );
  INV_X1 U15008 ( .A(n12268), .ZN(n12123) );
  AOI22_X1 U15009 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12045), .B1(
        n12123), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12016) );
  INV_X1 U15010 ( .A(n12264), .ZN(n12054) );
  INV_X1 U15011 ( .A(n12266), .ZN(n12055) );
  AOI22_X1 U15012 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n12054), .B1(
        n12055), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12015) );
  OAI22_X1 U15013 ( .A1(n12170), .A2(n12010), .B1(n12272), .B2(n12009), .ZN(
        n12011) );
  INV_X1 U15014 ( .A(n12011), .ZN(n12014) );
  INV_X1 U15015 ( .A(n12012), .ZN(n12126) );
  INV_X1 U15016 ( .A(n12260), .ZN(n12125) );
  AOI22_X1 U15017 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12126), .B1(
        n12125), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12013) );
  NAND4_X1 U15018 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(
        n12023) );
  AOI22_X1 U15019 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10276), .B1(
        n10192), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12021) );
  INV_X1 U15020 ( .A(n12017), .ZN(n12048) );
  AOI22_X1 U15021 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12048), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15022 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15023 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12018) );
  NAND4_X1 U15024 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12022) );
  INV_X1 U15025 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12071) );
  OAI22_X1 U15026 ( .A1(n12071), .A2(n12187), .B1(n19126), .B2(n12026), .ZN(
        n12030) );
  NAND2_X1 U15027 ( .A1(n12027), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12028) );
  OAI211_X1 U15028 ( .C1(n12069), .C2(n19431), .A(n12028), .B(n13571), .ZN(
        n12029) );
  NOR2_X1 U15029 ( .A1(n12030), .A2(n12029), .ZN(n12044) );
  OAI22_X1 U15030 ( .A1(n12075), .A2(n19543), .B1(n12185), .B2(n12076), .ZN(
        n12032) );
  OAI22_X1 U15031 ( .A1(n12065), .A2(n12198), .B1(n12186), .B2(n12064), .ZN(
        n12031) );
  NOR2_X1 U15032 ( .A1(n12032), .A2(n12031), .ZN(n12043) );
  OAI22_X1 U15033 ( .A1(n12074), .A2(n19463), .B1(n12190), .B2(n12070), .ZN(
        n12035) );
  INV_X1 U15034 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12033) );
  NOR2_X1 U15035 ( .A1(n12035), .A2(n12034), .ZN(n12042) );
  INV_X1 U15036 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12037) );
  OAI22_X1 U15037 ( .A1(n12037), .A2(n12182), .B1(n12191), .B2(n12036), .ZN(
        n12040) );
  INV_X1 U15038 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12038) );
  OAI22_X1 U15039 ( .A1(n12038), .A2(n12195), .B1(n12196), .B2(n12068), .ZN(
        n12039) );
  NOR2_X1 U15040 ( .A1(n12040), .A2(n12039), .ZN(n12041) );
  NAND4_X1 U15041 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n12108) );
  AOI22_X1 U15042 ( .A1(n12045), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12125), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12053) );
  INV_X1 U15043 ( .A(n12046), .ZN(n12124) );
  AOI22_X1 U15044 ( .A1(n12124), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10192), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12052) );
  INV_X1 U15045 ( .A(n12272), .ZN(n12047) );
  AOI22_X1 U15046 ( .A1(n12048), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12047), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15047 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12049), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15048 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15049 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15050 ( .A1(n12123), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12054), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15051 ( .A1(n12055), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12126), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12056) );
  OR2_X1 U15052 ( .A1(n13315), .A2(n13571), .ZN(n12478) );
  INV_X1 U15053 ( .A(n12478), .ZN(n12082) );
  AOI22_X1 U15054 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15055 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12062) );
  NAND2_X1 U15056 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12061) );
  NAND2_X1 U15057 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12060) );
  NAND4_X1 U15058 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(
        n12067) );
  OAI22_X1 U15059 ( .A1(n12065), .A2(n12260), .B1(n12258), .B2(n12064), .ZN(
        n12066) );
  NOR2_X1 U15060 ( .A1(n12067), .A2(n12066), .ZN(n12081) );
  OAI22_X1 U15061 ( .A1(n12008), .A2(n12069), .B1(n12264), .B2(n12068), .ZN(
        n12073) );
  OAI22_X1 U15062 ( .A1(n12268), .A2(n12071), .B1(n12266), .B2(n12070), .ZN(
        n12072) );
  NOR2_X1 U15063 ( .A1(n12073), .A2(n12072), .ZN(n12080) );
  OAI22_X1 U15064 ( .A1(n12170), .A2(n12075), .B1(n12272), .B2(n12074), .ZN(
        n12078) );
  OAI22_X1 U15065 ( .A1(n20816), .A2(n12275), .B1(n12017), .B2(n12076), .ZN(
        n12077) );
  NOR2_X1 U15066 ( .A1(n12078), .A2(n12077), .ZN(n12079) );
  INV_X1 U15067 ( .A(n12479), .ZN(n12892) );
  NAND2_X1 U15068 ( .A1(n12082), .A2(n12892), .ZN(n12482) );
  AOI22_X1 U15069 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15070 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12085) );
  NAND2_X1 U15071 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12084) );
  NAND2_X1 U15072 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12083) );
  NAND4_X1 U15073 ( .A1(n12086), .A2(n12085), .A3(n12084), .A4(n12083), .ZN(
        n12106) );
  OAI22_X1 U15074 ( .A1(n12088), .A2(n12260), .B1(n12258), .B2(n12087), .ZN(
        n12089) );
  INV_X1 U15075 ( .A(n12089), .ZN(n12104) );
  INV_X1 U15076 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12091) );
  OAI22_X1 U15077 ( .A1(n12268), .A2(n12091), .B1(n12266), .B2(n12090), .ZN(
        n12095) );
  OAI22_X1 U15078 ( .A1(n12093), .A2(n12264), .B1(n12272), .B2(n12092), .ZN(
        n12094) );
  NOR2_X1 U15079 ( .A1(n12095), .A2(n12094), .ZN(n12103) );
  OAI22_X1 U15080 ( .A1(n12097), .A2(n12008), .B1(n12170), .B2(n12096), .ZN(
        n12101) );
  OAI22_X1 U15081 ( .A1(n12099), .A2(n12017), .B1(n12275), .B2(n12098), .ZN(
        n12100) );
  NOR2_X1 U15082 ( .A1(n12101), .A2(n12100), .ZN(n12102) );
  NAND3_X1 U15083 ( .A1(n12104), .A2(n12103), .A3(n12102), .ZN(n12105) );
  NOR2_X1 U15084 ( .A1(n12106), .A2(n12105), .ZN(n12899) );
  NAND2_X1 U15085 ( .A1(n12482), .A2(n12899), .ZN(n12107) );
  AOI22_X1 U15086 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15087 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12112) );
  NAND2_X1 U15088 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12111) );
  NAND2_X1 U15089 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12110) );
  NAND4_X1 U15090 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12117) );
  OAI22_X1 U15091 ( .A1(n12258), .A2(n12115), .B1(n12017), .B2(n12114), .ZN(
        n12116) );
  NOR2_X1 U15092 ( .A1(n12117), .A2(n12116), .ZN(n12133) );
  OAI22_X1 U15093 ( .A1(n12008), .A2(n12119), .B1(n12264), .B2(n12118), .ZN(
        n12122) );
  OAI22_X1 U15094 ( .A1(n20853), .A2(n12266), .B1(n12272), .B2(n12120), .ZN(
        n12121) );
  NOR2_X1 U15095 ( .A1(n12122), .A2(n12121), .ZN(n12132) );
  NAND2_X1 U15096 ( .A1(n12123), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12130) );
  NAND2_X1 U15097 ( .A1(n12124), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12129) );
  NAND2_X1 U15098 ( .A1(n12125), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12128) );
  NAND2_X1 U15099 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12127) );
  AND4_X1 U15100 ( .A1(n12130), .A2(n12129), .A3(n12128), .A4(n12127), .ZN(
        n12131) );
  INV_X1 U15101 ( .A(n12419), .ZN(n13138) );
  MUX2_X1 U15102 ( .A(n12899), .B(n12437), .S(n12144), .Z(n12452) );
  INV_X1 U15103 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12146) );
  INV_X1 U15104 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13476) );
  NAND2_X1 U15105 ( .A1(n12146), .A2(n13476), .ZN(n12135) );
  MUX2_X1 U15106 ( .A(n12907), .B(n12136), .S(n12144), .Z(n12455) );
  MUX2_X1 U15107 ( .A(n12455), .B(n12137), .S(n9593), .Z(n12138) );
  OAI21_X1 U15108 ( .B1(n12140), .B2(n12138), .A(n12226), .ZN(n13924) );
  INV_X1 U15109 ( .A(n12140), .ZN(n12143) );
  NAND2_X1 U15110 ( .A1(n12141), .A2(n12149), .ZN(n12142) );
  NAND2_X1 U15111 ( .A1(n12143), .A2(n12142), .ZN(n14020) );
  INV_X1 U15112 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13512) );
  MUX2_X1 U15113 ( .A(n13315), .B(n12145), .S(n12144), .Z(n12147) );
  MUX2_X1 U15114 ( .A(n12147), .B(n12146), .S(n9593), .Z(n13946) );
  INV_X1 U15115 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13308) );
  OR2_X1 U15116 ( .A1(n13946), .A2(n13308), .ZN(n15170) );
  NAND3_X1 U15117 ( .A1(n9593), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n12148) );
  NAND2_X1 U15118 ( .A1(n12149), .A2(n12148), .ZN(n15171) );
  NOR2_X1 U15119 ( .A1(n15170), .A2(n15171), .ZN(n12150) );
  NAND2_X1 U15120 ( .A1(n15170), .A2(n15171), .ZN(n15169) );
  OAI21_X1 U15121 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12150), .A(
        n15169), .ZN(n13419) );
  XNOR2_X1 U15122 ( .A(n14020), .B(n13512), .ZN(n13418) );
  OR2_X1 U15123 ( .A1(n13419), .A2(n13418), .ZN(n13505) );
  OAI21_X1 U15124 ( .B1(n14020), .B2(n13512), .A(n13505), .ZN(n16116) );
  NAND2_X1 U15125 ( .A1(n16118), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12151) );
  NAND2_X1 U15126 ( .A1(n12152), .A2(n12151), .ZN(n19044) );
  INV_X1 U15127 ( .A(n12153), .ZN(n12177) );
  AOI22_X1 U15128 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12250), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15129 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12252), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12156) );
  NAND2_X1 U15130 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12155) );
  NAND2_X1 U15131 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12154) );
  NAND4_X1 U15132 ( .A1(n12157), .A2(n12156), .A3(n12155), .A4(n12154), .ZN(
        n12161) );
  OAI22_X1 U15133 ( .A1(n12159), .A2(n12260), .B1(n12258), .B2(n12158), .ZN(
        n12160) );
  NOR2_X1 U15134 ( .A1(n12161), .A2(n12160), .ZN(n12176) );
  OAI22_X1 U15135 ( .A1(n12008), .A2(n12163), .B1(n12264), .B2(n12162), .ZN(
        n12167) );
  INV_X1 U15136 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12165) );
  OAI22_X1 U15137 ( .A1(n12268), .A2(n12165), .B1(n12266), .B2(n12164), .ZN(
        n12166) );
  NOR2_X1 U15138 ( .A1(n12167), .A2(n12166), .ZN(n12175) );
  OAI22_X1 U15139 ( .A1(n12170), .A2(n12169), .B1(n12272), .B2(n12168), .ZN(
        n12173) );
  OAI22_X1 U15140 ( .A1(n10237), .A2(n12275), .B1(n12017), .B2(n12171), .ZN(
        n12172) );
  NOR2_X1 U15141 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  MUX2_X1 U15142 ( .A(n12177), .B(n12180), .S(n10075), .Z(n12450) );
  XNOR2_X1 U15143 ( .A(n12226), .B(n12225), .ZN(n12178) );
  XNOR2_X1 U15144 ( .A(n12178), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19045) );
  INV_X1 U15145 ( .A(n12178), .ZN(n18948) );
  NAND2_X1 U15146 ( .A1(n18948), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12179) );
  INV_X1 U15147 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12791) );
  OAI22_X1 U15148 ( .A1(n12791), .A2(n12181), .B1(n19431), .B2(n12805), .ZN(
        n12184) );
  INV_X1 U15149 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12793) );
  OAI22_X1 U15150 ( .A1(n12793), .A2(n12182), .B1(n19543), .B2(n12807), .ZN(
        n12183) );
  NOR2_X1 U15151 ( .A1(n12184), .A2(n12183), .ZN(n12204) );
  OAI22_X1 U15152 ( .A1(n9699), .A2(n12185), .B1(n12186), .B2(n12209), .ZN(
        n12189) );
  INV_X1 U15153 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12792) );
  OAI22_X1 U15154 ( .A1(n12792), .A2(n12187), .B1(n19508), .B2(n12809), .ZN(
        n12188) );
  NOR2_X1 U15155 ( .A1(n12189), .A2(n12188), .ZN(n12203) );
  OAI22_X1 U15156 ( .A1(n12806), .A2(n19463), .B1(n12190), .B2(n12213), .ZN(
        n12194) );
  OAI22_X1 U15157 ( .A1(n12192), .A2(n12191), .B1(n19082), .B2(n12216), .ZN(
        n12193) );
  NOR2_X1 U15158 ( .A1(n12194), .A2(n12193), .ZN(n12202) );
  INV_X1 U15159 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12197) );
  OAI22_X1 U15160 ( .A1(n12197), .A2(n19191), .B1(n12196), .B2(n12212), .ZN(
        n12200) );
  OAI22_X1 U15161 ( .A1(n12794), .A2(n19126), .B1(n12198), .B2(n12811), .ZN(
        n12199) );
  NOR2_X1 U15162 ( .A1(n12200), .A2(n12199), .ZN(n12201) );
  NAND4_X1 U15163 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12224) );
  AOI22_X1 U15164 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15165 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12207) );
  NAND2_X1 U15166 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12206) );
  NAND2_X1 U15167 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12205) );
  NAND4_X1 U15168 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12211) );
  OAI22_X1 U15169 ( .A1(n12260), .A2(n12811), .B1(n12258), .B2(n12209), .ZN(
        n12210) );
  NOR2_X1 U15170 ( .A1(n12211), .A2(n12210), .ZN(n12221) );
  OAI22_X1 U15171 ( .A1(n12008), .A2(n12805), .B1(n12264), .B2(n12212), .ZN(
        n12215) );
  OAI22_X1 U15172 ( .A1(n12268), .A2(n12792), .B1(n12266), .B2(n12213), .ZN(
        n12214) );
  NOR2_X1 U15173 ( .A1(n12215), .A2(n12214), .ZN(n12220) );
  OAI22_X1 U15174 ( .A1(n12170), .A2(n12807), .B1(n12272), .B2(n12806), .ZN(
        n12218) );
  OAI22_X1 U15175 ( .A1(n12275), .A2(n12216), .B1(n12017), .B2(n9699), .ZN(
        n12217) );
  NOR2_X1 U15176 ( .A1(n12218), .A2(n12217), .ZN(n12219) );
  NAND3_X1 U15177 ( .A1(n12221), .A2(n12220), .A3(n12219), .ZN(n12916) );
  INV_X1 U15178 ( .A(n12916), .ZN(n12222) );
  NAND2_X1 U15179 ( .A1(n12222), .A2(n13146), .ZN(n12223) );
  NAND2_X1 U15180 ( .A1(n12494), .A2(n12419), .ZN(n12228) );
  INV_X1 U15181 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13743) );
  OAI21_X1 U15182 ( .B1(n9677), .B2(n12227), .A(n12287), .ZN(n18923) );
  INV_X1 U15183 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U15184 ( .A1(n12229), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12230) );
  OAI22_X1 U15185 ( .A1(n12271), .A2(n19463), .B1(n19431), .B2(n12823), .ZN(
        n12234) );
  INV_X1 U15186 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12232) );
  OAI22_X1 U15187 ( .A1(n12232), .A2(n12181), .B1(n12190), .B2(n12265), .ZN(
        n12233) );
  NOR2_X1 U15188 ( .A1(n12234), .A2(n12233), .ZN(n12248) );
  OAI22_X1 U15189 ( .A1(n19178), .A2(n12191), .B1(n19082), .B2(n13770), .ZN(
        n12238) );
  INV_X1 U15190 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12236) );
  INV_X1 U15191 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12235) );
  OAI22_X1 U15192 ( .A1(n12236), .A2(n12182), .B1(n19191), .B2(n12235), .ZN(
        n12237) );
  NOR2_X1 U15193 ( .A1(n12238), .A2(n12237), .ZN(n12247) );
  OAI22_X1 U15194 ( .A1(n12273), .A2(n19543), .B1(n12196), .B2(n12263), .ZN(
        n12240) );
  OAI22_X1 U15195 ( .A1(n12274), .A2(n12185), .B1(n12198), .B2(n12259), .ZN(
        n12239) );
  NOR2_X1 U15196 ( .A1(n12240), .A2(n12239), .ZN(n12246) );
  OAI22_X1 U15197 ( .A1(n12241), .A2(n19126), .B1(n12186), .B2(n12257), .ZN(
        n12244) );
  INV_X1 U15198 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12267) );
  OAI22_X1 U15199 ( .A1(n12267), .A2(n12187), .B1(n19508), .B2(n12242), .ZN(
        n12243) );
  NOR2_X1 U15200 ( .A1(n12244), .A2(n12243), .ZN(n12245) );
  NAND4_X1 U15201 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(
        n12282) );
  AOI22_X1 U15202 ( .A1(n12250), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12249), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15203 ( .A1(n12252), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12251), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12255) );
  NAND2_X1 U15204 ( .A1(n10192), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12254) );
  NAND2_X1 U15205 ( .A1(n10276), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12253) );
  NAND4_X1 U15206 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12253), .ZN(
        n12262) );
  OAI22_X1 U15207 ( .A1(n12260), .A2(n12259), .B1(n12258), .B2(n12257), .ZN(
        n12261) );
  NOR2_X1 U15208 ( .A1(n12262), .A2(n12261), .ZN(n12280) );
  OAI22_X1 U15209 ( .A1(n12008), .A2(n12823), .B1(n12264), .B2(n12263), .ZN(
        n12270) );
  OAI22_X1 U15210 ( .A1(n12268), .A2(n12267), .B1(n12266), .B2(n12265), .ZN(
        n12269) );
  NOR2_X1 U15211 ( .A1(n12270), .A2(n12269), .ZN(n12279) );
  OAI22_X1 U15212 ( .A1(n12170), .A2(n12273), .B1(n12272), .B2(n12271), .ZN(
        n12277) );
  OAI22_X1 U15213 ( .A1(n12275), .A2(n13770), .B1(n12017), .B2(n12274), .ZN(
        n12276) );
  NOR2_X1 U15214 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  NAND2_X1 U15215 ( .A1(n12920), .A2(n13146), .ZN(n12281) );
  NAND2_X1 U15216 ( .A1(n12495), .A2(n12419), .ZN(n12283) );
  XNOR2_X1 U15217 ( .A(n12287), .B(n12286), .ZN(n14012) );
  NAND2_X1 U15218 ( .A1(n12284), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12285) );
  NAND2_X1 U15219 ( .A1(n9593), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12288) );
  NOR2_X1 U15220 ( .A1(n12292), .A2(n12288), .ZN(n12289) );
  OR2_X1 U15221 ( .A1(n12307), .A2(n12289), .ZN(n13983) );
  NOR2_X1 U15222 ( .A1(n13983), .A2(n12419), .ZN(n12301) );
  AND2_X1 U15223 ( .A1(n12301), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16098) );
  XNOR2_X1 U15224 ( .A(n12291), .B(n12290), .ZN(n18909) );
  AND2_X1 U15225 ( .A1(n18909), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16095) );
  INV_X1 U15226 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13806) );
  INV_X1 U15227 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13997) );
  INV_X1 U15228 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18883) );
  NAND2_X1 U15229 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12299), .ZN(n12293) );
  OR2_X1 U15230 ( .A1(n12322), .A2(n12294), .ZN(n18884) );
  OR2_X1 U15231 ( .A1(n18884), .A2(n12419), .ZN(n12295) );
  INV_X1 U15232 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12317) );
  AND2_X1 U15233 ( .A1(n12295), .A2(n12317), .ZN(n16067) );
  INV_X1 U15234 ( .A(n16067), .ZN(n12312) );
  NAND2_X1 U15235 ( .A1(n12306), .A2(n13997), .ZN(n12299) );
  NOR2_X1 U15236 ( .A1(n12306), .A2(n13997), .ZN(n12296) );
  NAND2_X1 U15237 ( .A1(n9593), .A2(n12296), .ZN(n12297) );
  AND2_X1 U15238 ( .A1(n12420), .A2(n12297), .ZN(n12298) );
  NAND2_X1 U15239 ( .A1(n12299), .A2(n12298), .ZN(n13994) );
  OR2_X1 U15240 ( .A1(n13994), .A2(n12419), .ZN(n12300) );
  NAND2_X1 U15241 ( .A1(n12300), .A2(n16183), .ZN(n16078) );
  INV_X1 U15242 ( .A(n12301), .ZN(n12303) );
  INV_X1 U15243 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U15244 ( .A1(n12303), .A2(n12302), .ZN(n16097) );
  INV_X1 U15245 ( .A(n18909), .ZN(n12305) );
  INV_X1 U15246 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12304) );
  NAND2_X1 U15247 ( .A1(n12305), .A2(n12304), .ZN(n16096) );
  AND2_X1 U15248 ( .A1(n16097), .A2(n16096), .ZN(n15369) );
  INV_X1 U15249 ( .A(n12306), .ZN(n12310) );
  NAND2_X1 U15250 ( .A1(n9593), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12308) );
  MUX2_X1 U15251 ( .A(n12308), .B(n9593), .S(n12307), .Z(n12309) );
  AND2_X1 U15252 ( .A1(n12310), .A2(n12309), .ZN(n12314) );
  AOI21_X1 U15253 ( .B1(n12314), .B2(n13138), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15371) );
  INV_X1 U15254 ( .A(n15371), .ZN(n12311) );
  AND2_X1 U15255 ( .A1(n15369), .A2(n12311), .ZN(n16074) );
  AND2_X1 U15256 ( .A1(n16078), .A2(n16074), .ZN(n16062) );
  AND2_X1 U15257 ( .A1(n12312), .A2(n16062), .ZN(n12313) );
  INV_X1 U15258 ( .A(n12314), .ZN(n18895) );
  INV_X1 U15259 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12315) );
  OR2_X1 U15260 ( .A1(n12419), .A2(n12315), .ZN(n12316) );
  OR2_X1 U15261 ( .A1(n18895), .A2(n12316), .ZN(n15370) );
  OR3_X1 U15262 ( .A1(n13994), .A2(n12419), .A3(n16183), .ZN(n16077) );
  NAND2_X1 U15263 ( .A1(n15370), .A2(n16077), .ZN(n16063) );
  OR2_X1 U15264 ( .A1(n12419), .A2(n12317), .ZN(n12318) );
  NOR2_X1 U15265 ( .A1(n18884), .A2(n12318), .ZN(n16066) );
  NOR2_X1 U15266 ( .A1(n16063), .A2(n16066), .ZN(n12319) );
  NAND2_X1 U15267 ( .A1(n9593), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12321) );
  NAND3_X1 U15268 ( .A1(n9593), .A2(n12323), .A3(P2_EBX_REG_12__SCAN_IN), .ZN(
        n12324) );
  NAND2_X1 U15269 ( .A1(n12328), .A2(n12324), .ZN(n18871) );
  OR2_X1 U15270 ( .A1(n18871), .A2(n12419), .ZN(n15363) );
  NAND2_X1 U15271 ( .A1(n12328), .A2(n12327), .ZN(n12329) );
  NAND2_X1 U15272 ( .A1(n12358), .A2(n12329), .ZN(n18855) );
  OR2_X1 U15273 ( .A1(n18855), .A2(n12419), .ZN(n12330) );
  INV_X1 U15274 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12377) );
  NAND2_X1 U15275 ( .A1(n12330), .A2(n12377), .ZN(n15148) );
  NAND2_X1 U15276 ( .A1(n9593), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12346) );
  INV_X1 U15277 ( .A(n12344), .ZN(n12332) );
  INV_X1 U15278 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12334) );
  NOR2_X2 U15279 ( .A1(n12343), .A2(n12341), .ZN(n12339) );
  INV_X1 U15280 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14921) );
  AND3_X1 U15281 ( .A1(n12336), .A2(n9593), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n12337) );
  NOR2_X1 U15282 ( .A1(n12383), .A2(n12337), .ZN(n12366) );
  INV_X1 U15283 ( .A(n12366), .ZN(n14848) );
  INV_X1 U15284 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12364) );
  OAI21_X1 U15285 ( .B1(n14848), .B2(n12419), .A(n12364), .ZN(n15106) );
  NAND2_X1 U15286 ( .A1(n9593), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12338) );
  XNOR2_X1 U15287 ( .A(n12339), .B(n12338), .ZN(n12379) );
  INV_X1 U15288 ( .A(n12379), .ZN(n14861) );
  NAND2_X1 U15289 ( .A1(n14861), .A2(n13138), .ZN(n12340) );
  INV_X1 U15290 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15287) );
  NAND2_X1 U15291 ( .A1(n12340), .A2(n15287), .ZN(n15118) );
  INV_X1 U15292 ( .A(n12341), .ZN(n12342) );
  XNOR2_X1 U15293 ( .A(n12343), .B(n12342), .ZN(n18799) );
  NAND2_X1 U15294 ( .A1(n18799), .A2(n13138), .ZN(n12367) );
  INV_X1 U15295 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16151) );
  NAND2_X1 U15296 ( .A1(n12367), .A2(n16151), .ZN(n13223) );
  XNOR2_X1 U15297 ( .A(n12348), .B(n12344), .ZN(n12368) );
  INV_X1 U15298 ( .A(n12368), .ZN(n18810) );
  NAND2_X1 U15299 ( .A1(n18810), .A2(n13138), .ZN(n12345) );
  INV_X1 U15300 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n20842) );
  NAND2_X1 U15301 ( .A1(n12345), .A2(n20842), .ZN(n13220) );
  AND2_X1 U15302 ( .A1(n13223), .A2(n13220), .ZN(n15115) );
  AND2_X1 U15303 ( .A1(n15118), .A2(n15115), .ZN(n15104) );
  OR2_X1 U15304 ( .A1(n9669), .A2(n12346), .ZN(n12347) );
  AND2_X1 U15305 ( .A1(n12348), .A2(n12347), .ZN(n12370) );
  INV_X1 U15306 ( .A(n12370), .ZN(n18819) );
  INV_X1 U15307 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15135) );
  OAI21_X1 U15308 ( .B1(n18819), .B2(n12419), .A(n15135), .ZN(n12521) );
  INV_X1 U15309 ( .A(n12349), .ZN(n12351) );
  NAND2_X1 U15310 ( .A1(n12351), .A2(n12350), .ZN(n12355) );
  INV_X1 U15311 ( .A(n12420), .ZN(n12352) );
  AOI21_X1 U15312 ( .B1(n12349), .B2(n12353), .A(n12352), .ZN(n12354) );
  NAND2_X1 U15313 ( .A1(n14151), .A2(n13138), .ZN(n12356) );
  XNOR2_X1 U15314 ( .A(n12356), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15317) );
  OR2_X1 U15315 ( .A1(n12358), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12360) );
  NAND3_X1 U15316 ( .A1(n12360), .A2(n9593), .A3(P2_EBX_REG_15__SCAN_IN), .ZN(
        n12357) );
  AND2_X1 U15317 ( .A1(n12357), .A2(n12349), .ZN(n12375) );
  INV_X1 U15318 ( .A(n12375), .ZN(n18831) );
  INV_X1 U15319 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12373) );
  OAI21_X1 U15320 ( .B1(n18831), .B2(n12419), .A(n12373), .ZN(n15327) );
  NAND2_X1 U15321 ( .A1(n9593), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12359) );
  MUX2_X1 U15322 ( .A(n9593), .B(n12359), .S(n12358), .Z(n12361) );
  NAND2_X1 U15323 ( .A1(n18844), .A2(n13138), .ZN(n12362) );
  INV_X1 U15324 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12371) );
  NAND2_X1 U15325 ( .A1(n12362), .A2(n12371), .ZN(n16049) );
  AND4_X1 U15326 ( .A1(n12521), .A2(n15317), .A3(n15327), .A4(n16049), .ZN(
        n12363) );
  NAND3_X1 U15327 ( .A1(n15106), .A2(n15104), .A3(n12363), .ZN(n12382) );
  NOR2_X1 U15328 ( .A1(n12419), .A2(n12364), .ZN(n12365) );
  NAND2_X1 U15329 ( .A1(n12366), .A2(n12365), .ZN(n15105) );
  OR2_X1 U15330 ( .A1(n12367), .A2(n16151), .ZN(n13224) );
  OR3_X1 U15331 ( .A1(n12368), .A2(n12419), .A3(n20842), .ZN(n13222) );
  AND2_X1 U15332 ( .A1(n13224), .A2(n13222), .ZN(n15101) );
  NOR2_X1 U15333 ( .A1(n12419), .A2(n15135), .ZN(n12369) );
  NAND2_X1 U15334 ( .A1(n12370), .A2(n12369), .ZN(n12520) );
  NOR2_X1 U15335 ( .A1(n12419), .A2(n12371), .ZN(n12372) );
  NAND2_X1 U15336 ( .A1(n18844), .A2(n12372), .ZN(n16048) );
  NOR2_X1 U15337 ( .A1(n12419), .A2(n12373), .ZN(n12374) );
  NAND2_X1 U15338 ( .A1(n12375), .A2(n12374), .ZN(n15326) );
  AND2_X1 U15339 ( .A1(n16048), .A2(n15326), .ZN(n12518) );
  INV_X1 U15340 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15307) );
  NOR2_X1 U15341 ( .A1(n12419), .A2(n15307), .ZN(n12376) );
  NAND2_X1 U15342 ( .A1(n14151), .A2(n12376), .ZN(n12519) );
  OR2_X1 U15343 ( .A1(n12419), .A2(n12377), .ZN(n12378) );
  OR2_X1 U15344 ( .A1(n18855), .A2(n12378), .ZN(n15147) );
  AND4_X1 U15345 ( .A1(n12520), .A2(n12518), .A3(n12519), .A4(n15147), .ZN(
        n12380) );
  OR3_X1 U15346 ( .A1(n12379), .A2(n12419), .A3(n15287), .ZN(n15117) );
  AND4_X1 U15347 ( .A1(n15105), .A2(n15101), .A3(n12380), .A4(n15117), .ZN(
        n12381) );
  NAND2_X1 U15348 ( .A1(n9593), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12384) );
  INV_X1 U15349 ( .A(n12384), .ZN(n12385) );
  NAND2_X1 U15350 ( .A1(n12386), .A2(n12385), .ZN(n12387) );
  NAND2_X1 U15351 ( .A1(n12399), .A2(n12387), .ZN(n15528) );
  OR2_X1 U15352 ( .A1(n15528), .A2(n12419), .ZN(n12391) );
  INV_X1 U15353 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15243) );
  NAND2_X1 U15354 ( .A1(n12391), .A2(n15243), .ZN(n15255) );
  INV_X1 U15355 ( .A(n12398), .ZN(n12389) );
  XNOR2_X1 U15356 ( .A(n12399), .B(n12389), .ZN(n15993) );
  NAND2_X1 U15357 ( .A1(n15993), .A2(n13138), .ZN(n12395) );
  XNOR2_X1 U15358 ( .A(n12395), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15091) );
  AND2_X1 U15359 ( .A1(n15255), .A2(n15091), .ZN(n12390) );
  NAND2_X1 U15360 ( .A1(n15086), .A2(n12390), .ZN(n15089) );
  INV_X1 U15361 ( .A(n15091), .ZN(n12393) );
  INV_X1 U15362 ( .A(n12391), .ZN(n12392) );
  NAND2_X1 U15363 ( .A1(n12392), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15256) );
  INV_X1 U15364 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12394) );
  OR2_X1 U15365 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  AND2_X1 U15366 ( .A1(n15088), .A2(n12396), .ZN(n12397) );
  NAND3_X1 U15367 ( .A1(n12401), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n9593), .ZN(
        n12400) );
  NAND2_X1 U15368 ( .A1(n12400), .A2(n12420), .ZN(n12402) );
  OR2_X1 U15369 ( .A1(n12402), .A2(n12422), .ZN(n13274) );
  AND2_X1 U15370 ( .A1(n12403), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15231) );
  INV_X1 U15371 ( .A(n12403), .ZN(n12404) );
  INV_X1 U15372 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13196) );
  NAND2_X1 U15373 ( .A1(n12404), .A2(n13196), .ZN(n15230) );
  INV_X1 U15374 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12406) );
  NAND3_X1 U15375 ( .A1(n9593), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n12407), .ZN(
        n12408) );
  AND2_X1 U15376 ( .A1(n13137), .A2(n12408), .ZN(n15972) );
  INV_X1 U15377 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15069) );
  NOR2_X1 U15378 ( .A1(n12419), .A2(n15069), .ZN(n12409) );
  NAND2_X1 U15379 ( .A1(n15972), .A2(n12409), .ZN(n12430) );
  INV_X1 U15380 ( .A(n15972), .ZN(n12410) );
  OAI21_X1 U15381 ( .B1(n12410), .B2(n12419), .A(n15069), .ZN(n12411) );
  NAND2_X1 U15382 ( .A1(n12430), .A2(n12411), .ZN(n15068) );
  NAND2_X1 U15383 ( .A1(n9593), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12415) );
  INV_X1 U15384 ( .A(n12415), .ZN(n12417) );
  NAND2_X1 U15385 ( .A1(n12417), .A2(n12416), .ZN(n12418) );
  NAND2_X1 U15386 ( .A1(n12425), .A2(n12418), .ZN(n15964) );
  INV_X1 U15387 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15062) );
  NAND2_X1 U15388 ( .A1(n12540), .A2(n15062), .ZN(n12423) );
  AOI21_X1 U15389 ( .B1(n12422), .B2(n10637), .A(n12421), .ZN(n15982) );
  INV_X1 U15390 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12424) );
  NAND2_X1 U15391 ( .A1(n12424), .A2(n15062), .ZN(n12428) );
  INV_X1 U15392 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12466) );
  AOI21_X1 U15393 ( .B1(n12426), .B2(n12425), .A(n13073), .ZN(n14823) );
  NAND2_X1 U15394 ( .A1(n14823), .A2(n13138), .ZN(n12541) );
  INV_X1 U15395 ( .A(n12541), .ZN(n12427) );
  OAI21_X1 U15396 ( .B1(n12431), .B2(n12428), .A(n12427), .ZN(n12433) );
  INV_X1 U15397 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16129) );
  NAND2_X1 U15398 ( .A1(n15082), .A2(n12430), .ZN(n12537) );
  NAND2_X1 U15399 ( .A1(n9593), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13072) );
  XNOR2_X1 U15400 ( .A(n13073), .B(n13072), .ZN(n12435) );
  INV_X1 U15401 ( .A(n12435), .ZN(n15946) );
  NAND3_X1 U15402 ( .A1(n15946), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13138), .ZN(n14238) );
  INV_X1 U15403 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12434) );
  OAI21_X1 U15404 ( .B1(n12435), .B2(n12419), .A(n12434), .ZN(n13130) );
  NOR2_X1 U15405 ( .A1(n12437), .A2(n12436), .ZN(n12440) );
  AND2_X1 U15406 ( .A1(n12438), .A2(n12440), .ZN(n12439) );
  OR2_X1 U15407 ( .A1(n12458), .A2(n12439), .ZN(n16259) );
  AOI21_X1 U15408 ( .B1(n12441), .B2(n12440), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n12442) );
  INV_X1 U15409 ( .A(n12442), .ZN(n12443) );
  OR2_X1 U15410 ( .A1(n16259), .A2(n12443), .ZN(n12448) );
  AOI21_X1 U15411 ( .B1(n12445), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16269) );
  NAND2_X1 U15412 ( .A1(n12170), .A2(n16269), .ZN(n12446) );
  INV_X1 U15413 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13466) );
  AOI21_X1 U15414 ( .B1(n12446), .B2(n13466), .A(n15404), .ZN(n19754) );
  INV_X1 U15415 ( .A(n19754), .ZN(n12447) );
  AND2_X1 U15416 ( .A1(n12448), .A2(n12447), .ZN(n19766) );
  NAND2_X1 U15417 ( .A1(n12449), .A2(n13571), .ZN(n12460) );
  INV_X1 U15418 ( .A(n12450), .ZN(n12454) );
  NAND2_X1 U15419 ( .A1(n12452), .A2(n12451), .ZN(n12453) );
  NAND2_X1 U15420 ( .A1(n12454), .A2(n12453), .ZN(n12457) );
  INV_X1 U15421 ( .A(n12455), .ZN(n12456) );
  NOR2_X1 U15422 ( .A1(n12457), .A2(n12456), .ZN(n12459) );
  OR2_X1 U15423 ( .A1(n12459), .A2(n12458), .ZN(n19763) );
  AND2_X1 U15424 ( .A1(n13146), .A2(n16265), .ZN(n19776) );
  NAND2_X1 U15425 ( .A1(n12449), .A2(n19776), .ZN(n19762) );
  OAI22_X1 U15426 ( .A1(n19766), .A2(n12460), .B1(n19763), .B2(n19762), .ZN(
        n13154) );
  AND2_X1 U15427 ( .A1(n16265), .A2(n19633), .ZN(n12461) );
  NAND2_X1 U15428 ( .A1(n13154), .A2(n12461), .ZN(n13331) );
  OR2_X1 U15429 ( .A1(n13331), .A2(n13146), .ZN(n16109) );
  INV_X1 U15430 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12462) );
  INV_X1 U15431 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15164) );
  INV_X1 U15432 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18894) );
  INV_X1 U15433 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16073) );
  INV_X1 U15434 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15151) );
  INV_X1 U15435 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18830) );
  INV_X1 U15436 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15139) );
  INV_X1 U15437 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20810) );
  INV_X1 U15438 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20815) );
  INV_X1 U15439 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15095) );
  INV_X1 U15440 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15078) );
  NOR2_X2 U15441 ( .A1(n13046), .A2(n15078), .ZN(n13048) );
  INV_X1 U15442 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15059) );
  INV_X1 U15443 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12550) );
  AOI21_X1 U15444 ( .B1(n12462), .B2(n12544), .A(n13054), .ZN(n15952) );
  NOR2_X1 U15445 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19635) );
  INV_X1 U15446 ( .A(n19635), .ZN(n19726) );
  AND2_X1 U15447 ( .A1(n19539), .A2(n19726), .ZN(n19782) );
  OR2_X1 U15448 ( .A1(n19782), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12463) );
  NAND2_X1 U15449 ( .A1(n13331), .A2(n12463), .ZN(n16124) );
  INV_X1 U15450 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19725) );
  NAND2_X1 U15451 ( .A1(n19725), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12464) );
  NAND2_X1 U15452 ( .A1(n15603), .A2(n12464), .ZN(n13400) );
  AOI22_X1 U15453 ( .A1(n13059), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12465) );
  OAI21_X1 U15454 ( .B1(n13207), .B2(n12466), .A(n12465), .ZN(n12467) );
  AOI21_X1 U15455 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12467), .ZN(n12548) );
  INV_X1 U15456 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15457 ( .A1(n13059), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12470) );
  OAI21_X1 U15458 ( .B1(n13207), .B2(n12471), .A(n12470), .ZN(n12472) );
  AOI21_X1 U15459 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12472), .ZN(n12474) );
  OR2_X2 U15460 ( .A1(n12473), .A2(n12474), .ZN(n13203) );
  NAND2_X1 U15461 ( .A1(n12473), .A2(n12474), .ZN(n12475) );
  NAND2_X1 U15462 ( .A1(n13203), .A2(n12475), .ZN(n15947) );
  AND2_X1 U15463 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19743) );
  INV_X1 U15464 ( .A(n19047), .ZN(n16034) );
  NOR2_X1 U15465 ( .A1(n19539), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n18774) );
  NAND2_X1 U15466 ( .A1(n19040), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15184) );
  INV_X1 U15467 ( .A(n16124), .ZN(n19041) );
  NAND2_X1 U15468 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12476) );
  OAI211_X1 U15469 ( .C1(n15947), .C2(n16034), .A(n15184), .B(n12476), .ZN(
        n12477) );
  AOI21_X1 U15470 ( .B1(n15952), .B2(n16115), .A(n12477), .ZN(n12515) );
  NAND2_X1 U15471 ( .A1(n12478), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13317) );
  XNOR2_X1 U15472 ( .A(n13315), .B(n12479), .ZN(n12480) );
  NOR2_X1 U15473 ( .A1(n13317), .A2(n12480), .ZN(n12481) );
  INV_X1 U15474 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15176) );
  XNOR2_X1 U15475 ( .A(n13317), .B(n12480), .ZN(n15175) );
  NOR2_X1 U15476 ( .A1(n15176), .A2(n15175), .ZN(n15174) );
  NOR2_X1 U15477 ( .A1(n12481), .A2(n15174), .ZN(n12483) );
  NOR2_X1 U15478 ( .A1(n12483), .A2(n13512), .ZN(n12484) );
  XOR2_X1 U15479 ( .A(n12899), .B(n12482), .Z(n13414) );
  XNOR2_X1 U15480 ( .A(n13512), .B(n12483), .ZN(n13413) );
  NOR2_X1 U15481 ( .A1(n13414), .A2(n13413), .ZN(n13412) );
  NOR2_X1 U15482 ( .A1(n12484), .A2(n13412), .ZN(n12485) );
  XOR2_X1 U15483 ( .A(n9705), .B(n12485), .Z(n16119) );
  OR2_X1 U15484 ( .A1(n12485), .A2(n9705), .ZN(n12491) );
  NAND2_X1 U15485 ( .A1(n12490), .A2(n12491), .ZN(n12489) );
  INV_X1 U15486 ( .A(n12486), .ZN(n12488) );
  NAND2_X1 U15487 ( .A1(n12488), .A2(n12487), .ZN(n12492) );
  XNOR2_X1 U15488 ( .A(n12489), .B(n12492), .ZN(n19043) );
  INV_X1 U15489 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19059) );
  NAND3_X1 U15490 ( .A1(n12492), .A2(n12490), .A3(n12491), .ZN(n12493) );
  NAND2_X1 U15491 ( .A1(n14186), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12500) );
  NAND2_X1 U15492 ( .A1(n12498), .A2(n12496), .ZN(n12499) );
  INV_X1 U15493 ( .A(n15158), .ZN(n12505) );
  INV_X1 U15494 ( .A(n12502), .ZN(n12503) );
  XNOR2_X1 U15495 ( .A(n12507), .B(n12419), .ZN(n15159) );
  NAND2_X1 U15496 ( .A1(n15158), .A2(n15159), .ZN(n12506) );
  NAND2_X1 U15497 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n12508), .ZN(
        n12509) );
  NAND2_X1 U15498 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15272) );
  NOR2_X1 U15499 ( .A1(n12315), .A2(n15272), .ZN(n15342) );
  NAND4_X1 U15500 ( .A1(n15342), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12523) );
  NOR3_X1 U15501 ( .A1(n15307), .A2(n12373), .A3(n15135), .ZN(n15294) );
  NAND4_X1 U15502 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15294), .A3(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15093) );
  NOR2_X1 U15503 ( .A1(n12523), .A2(n15093), .ZN(n15260) );
  NAND2_X1 U15504 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15260), .ZN(
        n15248) );
  NAND2_X1 U15505 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16136) );
  NOR2_X1 U15506 ( .A1(n15248), .A2(n16136), .ZN(n13193) );
  INV_X1 U15507 ( .A(n12511), .ZN(n12510) );
  AOI21_X1 U15508 ( .B1(n12510), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12512) );
  NAND2_X1 U15509 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14244) );
  NOR2_X1 U15510 ( .A1(n12512), .A2(n14243), .ZN(n15192) );
  INV_X1 U15511 ( .A(n13331), .ZN(n12513) );
  AND2_X1 U15512 ( .A1(n12513), .A2(n13146), .ZN(n19048) );
  NAND2_X1 U15513 ( .A1(n15192), .A2(n19048), .ZN(n12514) );
  NAND2_X1 U15514 ( .A1(n13220), .A2(n13222), .ZN(n12522) );
  INV_X1 U15515 ( .A(n15327), .ZN(n12517) );
  NAND2_X1 U15516 ( .A1(n15318), .A2(n15317), .ZN(n15316) );
  NAND2_X1 U15517 ( .A1(n12521), .A2(n12520), .ZN(n15131) );
  XOR2_X1 U15518 ( .A(n12522), .B(n15102), .Z(n15292) );
  INV_X1 U15519 ( .A(n16109), .ZN(n19046) );
  NAND2_X1 U15520 ( .A1(n15292), .A2(n19046), .ZN(n12536) );
  INV_X1 U15521 ( .A(n12523), .ZN(n15293) );
  NOR2_X2 U15522 ( .A1(n16032), .A2(n15307), .ZN(n16031) );
  NOR2_X2 U15523 ( .A1(n15133), .A2(n20842), .ZN(n15121) );
  AOI21_X1 U15524 ( .B1(n20842), .B2(n15133), .A(n15121), .ZN(n15299) );
  OR2_X1 U15525 ( .A1(n12526), .A2(n12525), .ZN(n12527) );
  AND2_X1 U15526 ( .A1(n12524), .A2(n12527), .ZN(n14931) );
  NAND2_X1 U15527 ( .A1(n14931), .A2(n19047), .ZN(n12533) );
  INV_X1 U15528 ( .A(n16115), .ZN(n19052) );
  OAI21_X1 U15529 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12528), .A(
        n13023), .ZN(n18809) );
  AOI22_X1 U15530 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19040), .ZN(n12530) );
  INV_X1 U15531 ( .A(n12530), .ZN(n12531) );
  NOR2_X1 U15532 ( .A1(n12529), .A2(n12531), .ZN(n12532) );
  NAND2_X1 U15533 ( .A1(n12533), .A2(n12532), .ZN(n12534) );
  AOI21_X1 U15534 ( .B1(n15299), .B2(n19048), .A(n12534), .ZN(n12535) );
  NAND2_X1 U15535 ( .A1(n12536), .A2(n12535), .ZN(P2_U2996) );
  INV_X1 U15536 ( .A(n12537), .ZN(n12538) );
  XNOR2_X1 U15537 ( .A(n12541), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12542) );
  XNOR2_X1 U15538 ( .A(n12543), .B(n12542), .ZN(n15208) );
  XNOR2_X1 U15539 ( .A(n12511), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15206) );
  NAND2_X1 U15540 ( .A1(n15206), .A2(n19048), .ZN(n12553) );
  INV_X1 U15541 ( .A(n12544), .ZN(n12545) );
  AOI21_X1 U15542 ( .B1(n12550), .B2(n13052), .A(n12545), .ZN(n14826) );
  INV_X1 U15543 ( .A(n12473), .ZN(n12546) );
  AOI21_X1 U15544 ( .B1(n12548), .B2(n12547), .A(n12546), .ZN(n15201) );
  NAND2_X1 U15545 ( .A1(n15201), .A2(n19047), .ZN(n12549) );
  NAND2_X1 U15546 ( .A1(n19040), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15197) );
  OAI211_X1 U15547 ( .C1(n16124), .C2(n12550), .A(n12549), .B(n15197), .ZN(
        n12551) );
  AOI21_X1 U15548 ( .B1(n14826), .B2(n16115), .A(n12551), .ZN(n12552) );
  OAI21_X1 U15549 ( .B1(n15208), .B2(n16109), .A(n9929), .ZN(P2_U2986) );
  NOR2_X1 U15550 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14630) );
  AND2_X1 U15551 ( .A1(n14630), .A2(n14791), .ZN(n14618) );
  NOR2_X1 U15552 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12554) );
  INV_X1 U15553 ( .A(n13841), .ZN(n12555) );
  NAND2_X1 U15554 ( .A1(n12566), .A2(n12565), .ZN(n12579) );
  XNOR2_X1 U15555 ( .A(n12579), .B(n12578), .ZN(n12557) );
  NAND2_X1 U15556 ( .A1(n13882), .A2(n11120), .ZN(n12560) );
  INV_X1 U15557 ( .A(n12560), .ZN(n12556) );
  AOI21_X1 U15558 ( .B1(n12557), .B2(n12607), .A(n12556), .ZN(n12558) );
  NAND2_X1 U15559 ( .A1(n12559), .A2(n12558), .ZN(n13662) );
  INV_X1 U15560 ( .A(n12621), .ZN(n12591) );
  OAI21_X1 U15561 ( .B1(n20800), .B2(n12565), .A(n12560), .ZN(n12561) );
  INV_X1 U15562 ( .A(n12561), .ZN(n12562) );
  NAND2_X2 U15563 ( .A1(n13494), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13493) );
  NAND2_X1 U15564 ( .A1(n12564), .A2(n11136), .ZN(n12571) );
  OAI21_X1 U15565 ( .B1(n12566), .B2(n12565), .A(n12579), .ZN(n12568) );
  OAI21_X1 U15566 ( .B1(n12568), .B2(n20800), .A(n12567), .ZN(n12569) );
  INV_X1 U15567 ( .A(n12569), .ZN(n12570) );
  NAND2_X1 U15568 ( .A1(n12571), .A2(n12570), .ZN(n12572) );
  XNOR2_X1 U15569 ( .A(n13493), .B(n12572), .ZN(n13527) );
  NAND2_X1 U15570 ( .A1(n13527), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13528) );
  INV_X1 U15571 ( .A(n13493), .ZN(n12573) );
  NAND2_X1 U15572 ( .A1(n12573), .A2(n12572), .ZN(n12574) );
  INV_X1 U15573 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19990) );
  NAND2_X1 U15574 ( .A1(n13662), .A2(n13663), .ZN(n13664) );
  NAND2_X1 U15575 ( .A1(n12575), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12576) );
  INV_X1 U15576 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19955) );
  NAND2_X1 U15577 ( .A1(n12579), .A2(n12578), .ZN(n12584) );
  XNOR2_X1 U15578 ( .A(n12584), .B(n12585), .ZN(n12580) );
  OAI22_X1 U15579 ( .A1(n12577), .A2(n12591), .B1(n20800), .B2(n12580), .ZN(
        n13776) );
  NAND2_X1 U15580 ( .A1(n12581), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12582) );
  NAND2_X1 U15581 ( .A1(n13775), .A2(n12582), .ZN(n19943) );
  NAND2_X1 U15582 ( .A1(n12583), .A2(n12621), .ZN(n12588) );
  NAND2_X1 U15583 ( .A1(n12585), .A2(n12584), .ZN(n12594) );
  XNOR2_X1 U15584 ( .A(n12593), .B(n12594), .ZN(n12586) );
  NAND2_X1 U15585 ( .A1(n12607), .A2(n12586), .ZN(n12587) );
  NAND2_X1 U15586 ( .A1(n12588), .A2(n12587), .ZN(n12589) );
  XNOR2_X1 U15587 ( .A(n12589), .B(n19963), .ZN(n19942) );
  NAND2_X1 U15588 ( .A1(n19943), .A2(n19942), .ZN(n19945) );
  NAND2_X1 U15589 ( .A1(n12589), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12590) );
  NAND2_X1 U15590 ( .A1(n19945), .A2(n12590), .ZN(n15806) );
  OR2_X1 U15591 ( .A1(n12592), .A2(n12591), .ZN(n12599) );
  INV_X1 U15592 ( .A(n12593), .ZN(n12595) );
  NOR2_X1 U15593 ( .A1(n12595), .A2(n12594), .ZN(n12605) );
  INV_X1 U15594 ( .A(n12605), .ZN(n12596) );
  XNOR2_X1 U15595 ( .A(n12604), .B(n12596), .ZN(n12597) );
  NAND2_X1 U15596 ( .A1(n12607), .A2(n12597), .ZN(n12598) );
  NAND2_X1 U15597 ( .A1(n12599), .A2(n12598), .ZN(n12600) );
  INV_X1 U15598 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15926) );
  XNOR2_X1 U15599 ( .A(n12600), .B(n15926), .ZN(n15805) );
  NAND2_X1 U15600 ( .A1(n12600), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12601) );
  NAND3_X1 U15601 ( .A1(n12602), .A2(n12603), .A3(n12621), .ZN(n12609) );
  NAND2_X1 U15602 ( .A1(n12605), .A2(n12604), .ZN(n12613) );
  XNOR2_X1 U15603 ( .A(n12612), .B(n12613), .ZN(n12606) );
  NAND2_X1 U15604 ( .A1(n12607), .A2(n12606), .ZN(n12608) );
  NAND2_X1 U15605 ( .A1(n15800), .A2(n15900), .ZN(n12610) );
  INV_X1 U15606 ( .A(n15800), .ZN(n12611) );
  INV_X1 U15607 ( .A(n12612), .ZN(n12614) );
  NOR2_X1 U15608 ( .A1(n12614), .A2(n12613), .ZN(n12624) );
  XNOR2_X1 U15609 ( .A(n12625), .B(n12624), .ZN(n12615) );
  NOR2_X1 U15610 ( .A1(n20800), .A2(n12615), .ZN(n12616) );
  AOI21_X1 U15611 ( .B1(n12617), .B2(n12621), .A(n12616), .ZN(n12618) );
  INV_X1 U15612 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15912) );
  NAND2_X1 U15613 ( .A1(n12618), .A2(n15912), .ZN(n15795) );
  NAND2_X1 U15614 ( .A1(n15793), .A2(n15795), .ZN(n12620) );
  INV_X1 U15615 ( .A(n12618), .ZN(n12619) );
  NAND2_X1 U15616 ( .A1(n12619), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15794) );
  NAND2_X1 U15617 ( .A1(n12620), .A2(n15794), .ZN(n14651) );
  AND2_X1 U15618 ( .A1(n12622), .A2(n12621), .ZN(n12623) );
  AND2_X4 U15619 ( .A1(n12602), .A2(n12623), .ZN(n15785) );
  NAND2_X1 U15620 ( .A1(n12625), .A2(n12624), .ZN(n12626) );
  NOR2_X1 U15621 ( .A1(n20800), .A2(n12626), .ZN(n12627) );
  INV_X1 U15622 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12628) );
  NAND2_X1 U15623 ( .A1(n14652), .A2(n12628), .ZN(n12629) );
  INV_X1 U15624 ( .A(n14652), .ZN(n12630) );
  NAND2_X1 U15625 ( .A1(n12630), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12631) );
  INV_X1 U15626 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12632) );
  NAND2_X1 U15627 ( .A1(n9588), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14622) );
  NAND2_X1 U15628 ( .A1(n15785), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12633) );
  NAND2_X1 U15629 ( .A1(n14622), .A2(n12633), .ZN(n14762) );
  AOI21_X1 U15630 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n15785), .ZN(n14631) );
  NOR2_X1 U15631 ( .A1(n15785), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14633) );
  OAI21_X1 U15632 ( .B1(n15785), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n14622), .ZN(n14634) );
  NOR3_X1 U15633 ( .A1(n14631), .A2(n14633), .A3(n14634), .ZN(n14621) );
  NAND2_X1 U15634 ( .A1(n15772), .A2(n15852), .ZN(n12634) );
  NAND2_X1 U15635 ( .A1(n14621), .A2(n12634), .ZN(n14764) );
  NAND2_X1 U15636 ( .A1(n14764), .A2(n14750), .ZN(n12636) );
  MUX2_X1 U15637 ( .A(n11919), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .S(
        n15785), .Z(n14766) );
  NOR2_X1 U15638 ( .A1(n15785), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12635) );
  NOR2_X1 U15639 ( .A1(n14766), .A2(n12635), .ZN(n14767) );
  NAND2_X1 U15640 ( .A1(n12636), .A2(n14767), .ZN(n14751) );
  INV_X1 U15641 ( .A(n14751), .ZN(n12637) );
  INV_X1 U15642 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14732) );
  NAND2_X1 U15643 ( .A1(n15831), .A2(n14732), .ZN(n12638) );
  INV_X1 U15644 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14733) );
  INV_X1 U15645 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12639) );
  AND2_X1 U15646 ( .A1(n14733), .A2(n12639), .ZN(n12640) );
  NAND2_X1 U15647 ( .A1(n14723), .A2(n12640), .ZN(n12641) );
  XNOR2_X1 U15648 ( .A(n15785), .B(n15831), .ZN(n14609) );
  NAND3_X1 U15649 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12708) );
  OAI21_X2 U15650 ( .B1(n14608), .B2(n12708), .A(n15772), .ZN(n14599) );
  NAND2_X1 U15651 ( .A1(n14599), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12642) );
  NAND2_X1 U15652 ( .A1(n14601), .A2(n12642), .ZN(n14555) );
  NAND3_X1 U15653 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12718) );
  NAND2_X1 U15654 ( .A1(n14555), .A2(n12718), .ZN(n12644) );
  NAND2_X1 U15655 ( .A1(n12642), .A2(n15772), .ZN(n14589) );
  NAND2_X1 U15656 ( .A1(n12644), .A2(n12643), .ZN(n12649) );
  NAND2_X1 U15657 ( .A1(n14555), .A2(n15785), .ZN(n14554) );
  INV_X1 U15658 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12645) );
  INV_X1 U15659 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15739) );
  NAND3_X1 U15660 ( .A1(n12646), .A2(n12645), .A3(n15739), .ZN(n14557) );
  NAND2_X1 U15661 ( .A1(n15785), .A2(n14557), .ZN(n12647) );
  NAND2_X1 U15662 ( .A1(n14554), .A2(n12647), .ZN(n14572) );
  INV_X1 U15663 ( .A(n14572), .ZN(n12648) );
  INV_X1 U15664 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14687) );
  INV_X1 U15665 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14564) );
  NAND2_X1 U15666 ( .A1(n14687), .A2(n14564), .ZN(n14679) );
  INV_X1 U15667 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12650) );
  NAND2_X1 U15668 ( .A1(n14549), .A2(n14550), .ZN(n12653) );
  AND2_X1 U15669 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U15670 ( .A1(n14670), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12719) );
  NOR2_X1 U15671 ( .A1(n9588), .A2(n12719), .ZN(n12651) );
  NAND2_X1 U15672 ( .A1(n14548), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12652) );
  NOR2_X1 U15673 ( .A1(n12697), .A2(n11130), .ZN(n12657) );
  NAND2_X1 U15674 ( .A1(n13649), .A2(n13882), .ZN(n12683) );
  AND2_X1 U15675 ( .A1(n12657), .A2(n12683), .ZN(n12777) );
  AND2_X1 U15676 ( .A1(n12658), .A2(n19999), .ZN(n12659) );
  NAND2_X1 U15677 ( .A1(n12660), .A2(n12659), .ZN(n12701) );
  NAND2_X1 U15678 ( .A1(n12777), .A2(n12701), .ZN(n12663) );
  NAND2_X1 U15679 ( .A1(n12662), .A2(n13882), .ZN(n13451) );
  NAND2_X1 U15680 ( .A1(n12663), .A2(n13451), .ZN(n13593) );
  NOR4_X1 U15681 ( .A1(n12667), .A2(n12666), .A3(n12665), .A4(n12664), .ZN(
        n12668) );
  NOR2_X1 U15682 ( .A1(n12669), .A2(n12668), .ZN(n13450) );
  NAND2_X1 U15683 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20797) );
  NAND2_X1 U15684 ( .A1(n13450), .A2(n20797), .ZN(n13234) );
  INV_X1 U15685 ( .A(n12670), .ZN(n12671) );
  INV_X1 U15686 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20701) );
  NAND2_X1 U15687 ( .A1(n12671), .A2(n20701), .ZN(n15597) );
  AND2_X1 U15688 ( .A1(n11136), .A2(n15597), .ZN(n12672) );
  OR2_X1 U15689 ( .A1(n13234), .A2(n12672), .ZN(n12677) );
  INV_X1 U15690 ( .A(n15597), .ZN(n13591) );
  OAI21_X1 U15691 ( .B1(n11136), .B2(n13591), .A(n20797), .ZN(n13888) );
  OAI211_X1 U15692 ( .C1(n12674), .C2(n13888), .A(n19999), .B(n13258), .ZN(
        n12675) );
  NAND2_X1 U15693 ( .A1(n12675), .A2(n13601), .ZN(n12676) );
  MUX2_X1 U15694 ( .A(n12677), .B(n12676), .S(n9594), .Z(n12679) );
  INV_X1 U15695 ( .A(n13601), .ZN(n15574) );
  NAND3_X1 U15696 ( .A1(n15574), .A2(n15542), .A3(n11136), .ZN(n12678) );
  NAND3_X1 U15697 ( .A1(n13593), .A2(n12679), .A3(n12678), .ZN(n12680) );
  INV_X1 U15698 ( .A(n12709), .ZN(n12705) );
  NAND2_X1 U15699 ( .A1(n12777), .A2(n12775), .ZN(n15560) );
  NOR2_X1 U15700 ( .A1(n12681), .A2(n11130), .ZN(n12682) );
  NAND2_X1 U15701 ( .A1(n12683), .A2(n12682), .ZN(n13584) );
  NAND2_X1 U15702 ( .A1(n15560), .A2(n13584), .ZN(n13448) );
  NOR2_X1 U15703 ( .A1(n12685), .A2(n12686), .ZN(n12688) );
  OR3_X1 U15704 ( .A1(n13448), .A2(n12688), .A3(n12687), .ZN(n12689) );
  AOI22_X1 U15705 ( .A1(n13622), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n9625), .ZN(n12691) );
  INV_X1 U15706 ( .A(n14429), .ZN(n12724) );
  OR2_X1 U15707 ( .A1(n12674), .A2(n20800), .ZN(n15568) );
  OAI21_X1 U15708 ( .B1(n12685), .B2(n11046), .A(n15568), .ZN(n12693) );
  INV_X1 U15709 ( .A(n12693), .ZN(n12694) );
  INV_X1 U15710 ( .A(n12718), .ZN(n14556) );
  INV_X1 U15711 ( .A(n13595), .ZN(n13873) );
  NAND2_X1 U15712 ( .A1(n12662), .A2(n13873), .ZN(n15544) );
  NAND2_X1 U15713 ( .A1(n11818), .A2(n13873), .ZN(n12696) );
  AND2_X1 U15714 ( .A1(n12696), .A2(n12695), .ZN(n12700) );
  INV_X1 U15715 ( .A(n11134), .ZN(n13241) );
  OAI21_X1 U15716 ( .B1(n12697), .B2(n13241), .A(n11136), .ZN(n12698) );
  NAND4_X1 U15717 ( .A1(n12701), .A2(n12700), .A3(n12699), .A4(n12698), .ZN(
        n13580) );
  OAI21_X1 U15718 ( .B1(n13882), .B2(n11123), .A(n12702), .ZN(n12704) );
  NAND2_X1 U15719 ( .A1(n12704), .A2(n12703), .ZN(n12706) );
  OAI21_X1 U15720 ( .B1(n13580), .B2(n12706), .A(n12705), .ZN(n14731) );
  NAND2_X1 U15721 ( .A1(n14731), .A2(n19981), .ZN(n13625) );
  INV_X1 U15722 ( .A(n13625), .ZN(n12707) );
  INV_X1 U15723 ( .A(n19981), .ZN(n15890) );
  NOR2_X1 U15724 ( .A1(n14602), .A2(n12708), .ZN(n14706) );
  INV_X1 U15725 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14757) );
  NAND3_X1 U15726 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14758) );
  NOR2_X1 U15727 ( .A1(n14757), .A2(n14758), .ZN(n15832) );
  NAND2_X1 U15728 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15832), .ZN(
        n12717) );
  INV_X1 U15729 ( .A(n12717), .ZN(n14707) );
  NAND2_X1 U15730 ( .A1(n13630), .A2(n14731), .ZN(n15888) );
  INV_X1 U15731 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15889) );
  NOR2_X1 U15732 ( .A1(n19963), .A2(n19955), .ZN(n19954) );
  NAND2_X1 U15733 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19954), .ZN(
        n15891) );
  NOR3_X1 U15734 ( .A1(n19990), .A2(n15889), .A3(n15891), .ZN(n15871) );
  NAND3_X1 U15735 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15877) );
  NOR3_X1 U15736 ( .A1(n11900), .A2(n12632), .A3(n15877), .ZN(n14788) );
  AND2_X1 U15737 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14788), .ZN(
        n14783) );
  NAND2_X1 U15738 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14783), .ZN(
        n15845) );
  INV_X1 U15739 ( .A(n15845), .ZN(n12710) );
  AND2_X1 U15740 ( .A1(n15871), .A2(n12710), .ZN(n15855) );
  NAND2_X1 U15741 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15855), .ZN(
        n12715) );
  OR2_X1 U15742 ( .A1(n12781), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19957) );
  NAND2_X1 U15743 ( .A1(n12709), .A2(n19957), .ZN(n14801) );
  OAI21_X1 U15744 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14731), .A(
        n14801), .ZN(n15887) );
  AOI21_X1 U15745 ( .B1(n15888), .B2(n12715), .A(n15887), .ZN(n12713) );
  INV_X1 U15746 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15846) );
  AOI21_X1 U15747 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15921) );
  NOR2_X1 U15748 ( .A1(n15921), .A2(n15891), .ZN(n15872) );
  NAND2_X1 U15749 ( .A1(n12710), .A2(n15872), .ZN(n14729) );
  NOR2_X1 U15750 ( .A1(n15846), .A2(n14729), .ZN(n12716) );
  INV_X1 U15751 ( .A(n12716), .ZN(n12711) );
  NAND2_X1 U15752 ( .A1(n15890), .A2(n12711), .ZN(n12712) );
  NAND2_X1 U15753 ( .A1(n12713), .A2(n12712), .ZN(n15860) );
  INV_X1 U15754 ( .A(n15860), .ZN(n15853) );
  OAI21_X1 U15755 ( .B1(n14772), .B2(n14707), .A(n15853), .ZN(n14746) );
  INV_X1 U15756 ( .A(n14746), .ZN(n14735) );
  OAI21_X1 U15757 ( .B1(n14772), .B2(n14706), .A(n14735), .ZN(n15818) );
  AOI21_X1 U15758 ( .B1(n15739), .B2(n15890), .A(n15818), .ZN(n14708) );
  OAI21_X1 U15759 ( .B1(n14556), .B2(n14772), .A(n14708), .ZN(n15815) );
  INV_X1 U15760 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14696) );
  NAND2_X1 U15761 ( .A1(n14708), .A2(n14772), .ZN(n14668) );
  OAI21_X1 U15762 ( .B1(n15815), .B2(n14696), .A(n14668), .ZN(n14678) );
  NAND2_X1 U15763 ( .A1(n14678), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14667) );
  INV_X1 U15764 ( .A(n14670), .ZN(n14680) );
  OAI21_X1 U15765 ( .B1(n14667), .B2(n14680), .A(n14668), .ZN(n12714) );
  NAND2_X1 U15766 ( .A1(n12714), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14662) );
  NAND3_X1 U15767 ( .A1(n14662), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14668), .ZN(n12722) );
  INV_X1 U15768 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20755) );
  NOR2_X1 U15769 ( .A1(n19957), .A2(n20755), .ZN(n13117) );
  INV_X1 U15770 ( .A(n13117), .ZN(n12721) );
  INV_X1 U15771 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13626) );
  NAND2_X1 U15772 ( .A1(n13626), .A2(n13630), .ZN(n14799) );
  NAND2_X1 U15773 ( .A1(n15888), .A2(n14799), .ZN(n14790) );
  NOR2_X1 U15774 ( .A1(n12715), .A2(n14790), .ZN(n14705) );
  AOI21_X1 U15775 ( .B1(n12716), .B2(n15890), .A(n14705), .ZN(n15821) );
  NOR2_X1 U15776 ( .A1(n15821), .A2(n12717), .ZN(n14740) );
  NAND2_X1 U15777 ( .A1(n14706), .A2(n14740), .ZN(n15810) );
  NOR2_X1 U15778 ( .A1(n15810), .A2(n12718), .ZN(n14697) );
  NAND2_X1 U15779 ( .A1(n14697), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14669) );
  NOR2_X1 U15780 ( .A1(n14669), .A2(n12719), .ZN(n14663) );
  NAND3_X1 U15781 ( .A1(n14663), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12654), .ZN(n12720) );
  NAND3_X1 U15782 ( .A1(n12722), .A2(n12721), .A3(n12720), .ZN(n12723) );
  OAI21_X1 U15783 ( .B1(n13129), .B2(n19977), .A(n12725), .ZN(P1_U3000) );
  NAND2_X1 U15784 ( .A1(n12726), .A2(n12728), .ZN(n17420) );
  NOR2_X1 U15785 ( .A1(n17419), .A2(n12756), .ZN(n17401) );
  AOI22_X1 U15786 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n10791), .B1(
        n9624), .B2(n12758), .ZN(n17402) );
  AND2_X1 U15787 ( .A1(n12729), .A2(n15517), .ZN(n12730) );
  NOR2_X1 U15788 ( .A1(n15522), .A2(n17772), .ZN(n16319) );
  OR2_X1 U15789 ( .A1(n17416), .A2(n15522), .ZN(n16309) );
  NOR2_X1 U15790 ( .A1(n12755), .A2(n15517), .ZN(n18000) );
  INV_X1 U15791 ( .A(n18559), .ZN(n18540) );
  NAND2_X1 U15792 ( .A1(n18546), .A2(n18540), .ZN(n17898) );
  NOR3_X1 U15793 ( .A1(n9785), .A2(n18041), .A3(n9789), .ZN(n18027) );
  NOR2_X1 U15794 ( .A1(n18071), .A2(n10690), .ZN(n18040) );
  AND2_X1 U15795 ( .A1(n18027), .A2(n18040), .ZN(n18003) );
  NAND4_X1 U15796 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n18003), .ZN(n17939) );
  NOR2_X1 U15797 ( .A1(n17876), .A2(n17939), .ZN(n17829) );
  INV_X1 U15798 ( .A(n18571), .ZN(n17987) );
  NOR2_X1 U15799 ( .A1(n18730), .A2(n17939), .ZN(n17963) );
  NAND2_X1 U15800 ( .A1(n17553), .A2(n17963), .ZN(n17900) );
  NAND2_X1 U15801 ( .A1(n17879), .A2(n17475), .ZN(n17832) );
  NOR2_X1 U15802 ( .A1(n17900), .A2(n17832), .ZN(n17835) );
  NAND4_X1 U15803 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n12759), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A4(n17835), .ZN(n12747) );
  INV_X1 U15804 ( .A(n9600), .ZN(n17892) );
  INV_X1 U15805 ( .A(n18536), .ZN(n12740) );
  INV_X1 U15806 ( .A(n13100), .ZN(n18535) );
  INV_X1 U15807 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18626) );
  NAND2_X1 U15808 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18626), .ZN(n18763) );
  INV_X1 U15809 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18629) );
  NOR2_X1 U15810 ( .A1(n18763), .A2(n18629), .ZN(n18628) );
  NOR2_X1 U15811 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18613) );
  NOR3_X1 U15812 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18628), .A3(n18613), 
        .ZN(n18748) );
  XOR2_X1 U15813 ( .A(n12731), .B(n18749), .Z(n12732) );
  NAND2_X1 U15814 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18759) );
  OAI21_X1 U15815 ( .B1(n18748), .B2(n12732), .A(n18759), .ZN(n16437) );
  NOR3_X1 U15816 ( .A1(n12733), .A2(n18535), .A3(n16437), .ZN(n12739) );
  INV_X1 U15817 ( .A(n12734), .ZN(n12735) );
  OAI211_X1 U15818 ( .C1(n12738), .C2(n12737), .A(n12736), .B(n12735), .ZN(
        n14229) );
  AOI211_X1 U15819 ( .C1(n12741), .C2(n12740), .A(n12739), .B(n14229), .ZN(
        n12742) );
  INV_X1 U15820 ( .A(n12742), .ZN(n12745) );
  AOI21_X1 U15821 ( .B1(n12743), .B2(n18119), .A(n15487), .ZN(n12744) );
  OAI21_X1 U15822 ( .B1(n10690), .B2(n18730), .A(n18071), .ZN(n18066) );
  NAND2_X1 U15823 ( .A1(n18027), .A2(n18066), .ZN(n18001) );
  NAND3_X1 U15824 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12746) );
  NOR2_X1 U15825 ( .A1(n18001), .A2(n12746), .ZN(n17923) );
  NAND2_X1 U15826 ( .A1(n17553), .A2(n17923), .ZN(n17831) );
  NAND2_X1 U15827 ( .A1(n18559), .A2(n17831), .ZN(n17878) );
  OAI21_X1 U15828 ( .B1(n12749), .B2(n18540), .A(n17878), .ZN(n17766) );
  AOI211_X1 U15829 ( .C1(n17987), .C2(n12747), .A(n18052), .B(n17766), .ZN(
        n12748) );
  OAI221_X1 U15830 ( .B1(n18546), .B2(n12749), .C1(n18546), .C2(n17829), .A(
        n12748), .ZN(n15586) );
  AOI21_X1 U15831 ( .B1(n9795), .B2(n17898), .A(n15586), .ZN(n15519) );
  INV_X1 U15832 ( .A(n15519), .ZN(n12750) );
  AOI21_X1 U15833 ( .B1(n16309), .B2(n18000), .A(n12750), .ZN(n12751) );
  OAI21_X1 U15834 ( .B1(n16319), .B2(n18539), .A(n12751), .ZN(n12752) );
  OAI21_X1 U15835 ( .B1(n12753), .B2(n12752), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12769) );
  NOR2_X1 U15836 ( .A1(n18090), .A2(n12754), .ZN(n12766) );
  INV_X1 U15837 ( .A(n12755), .ZN(n18537) );
  NAND2_X1 U15838 ( .A1(n18537), .A2(n18074), .ZN(n18083) );
  NOR2_X2 U15839 ( .A1(n17261), .A2(n18083), .ZN(n18009) );
  NAND3_X1 U15840 ( .A1(n12756), .A2(n18009), .A3(n17402), .ZN(n12764) );
  INV_X1 U15841 ( .A(n18539), .ZN(n17966) );
  AOI22_X1 U15842 ( .A1(n18000), .A2(n17969), .B1(n17966), .B2(n12757), .ZN(
        n17875) );
  INV_X1 U15843 ( .A(n17831), .ZN(n17787) );
  INV_X1 U15844 ( .A(n17768), .ZN(n18039) );
  NOR2_X1 U15845 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18574), .ZN(
        n18077) );
  NOR2_X1 U15846 ( .A1(n18039), .A2(n18077), .ZN(n17873) );
  AOI22_X1 U15847 ( .A1(n18559), .A2(n17787), .B1(n17829), .B2(n17873), .ZN(
        n17786) );
  OAI21_X1 U15848 ( .B1(n17875), .B2(n17876), .A(n17786), .ZN(n17825) );
  NAND3_X1 U15849 ( .A1(n18074), .A2(n17879), .A3(n17825), .ZN(n17802) );
  NAND3_X1 U15850 ( .A1(n12759), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n12758), .ZN(n17418) );
  NOR3_X1 U15851 ( .A1(n12760), .A2(n17802), .A3(n17418), .ZN(n12762) );
  AND2_X1 U15852 ( .A1(n18050), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n12761) );
  OAI21_X1 U15853 ( .B1(n12769), .B2(n18050), .A(n12768), .ZN(P3_U2834) );
  AOI21_X1 U15854 ( .B1(n12770), .B2(n14670), .A(n15785), .ZN(n12772) );
  OR2_X2 U15855 ( .A1(n12772), .A2(n12771), .ZN(n12774) );
  XNOR2_X1 U15856 ( .A(n9588), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12773) );
  XNOR2_X1 U15857 ( .A(n12774), .B(n12773), .ZN(n14677) );
  AND2_X1 U15858 ( .A1(n12775), .A2(n13240), .ZN(n12776) );
  INV_X1 U15859 ( .A(n12778), .ZN(n14310) );
  AOI21_X1 U15860 ( .B1(n12779), .B2(n14310), .A(n13121), .ZN(n14295) );
  NAND3_X1 U15861 ( .A1(n19998), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15939) );
  INV_X1 U15862 ( .A(n15939), .ZN(n12780) );
  OR2_X1 U15863 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20567) );
  INV_X2 U15864 ( .A(n20567), .ZN(n20625) );
  NAND2_X1 U15865 ( .A1(n20567), .A2(n12781), .ZN(n20796) );
  AND2_X1 U15866 ( .A1(n20796), .A2(n19998), .ZN(n12782) );
  NAND2_X1 U15867 ( .A1(n19998), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15565) );
  NAND2_X1 U15868 ( .A1(n20359), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12783) );
  AND2_X1 U15869 ( .A1(n15565), .A2(n12783), .ZN(n13491) );
  INV_X1 U15870 ( .A(n13491), .ZN(n12784) );
  INV_X1 U15871 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20753) );
  NOR2_X1 U15872 ( .A1(n19957), .A2(n20753), .ZN(n14674) );
  AOI21_X1 U15873 ( .B1(n19941), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14674), .ZN(n12785) );
  OAI21_X1 U15874 ( .B1(n19953), .B2(n14296), .A(n12785), .ZN(n12786) );
  AOI21_X1 U15875 ( .B1(n14295), .B2(n19947), .A(n12786), .ZN(n12787) );
  OAI21_X1 U15876 ( .B1(n14677), .B2(n19803), .A(n12787), .ZN(P1_U2970) );
  INV_X1 U15877 ( .A(n12790), .ZN(n12808) );
  OAI22_X1 U15878 ( .A1(n12808), .A2(n12792), .B1(n10179), .B2(n12791), .ZN(
        n12801) );
  OAI22_X1 U15879 ( .A1(n12795), .A2(n12794), .B1(n12810), .B2(n12793), .ZN(
        n12800) );
  AOI22_X1 U15880 ( .A1(n12826), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12798) );
  NAND2_X1 U15881 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12797) );
  NAND2_X1 U15882 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12796) );
  NAND4_X1 U15883 ( .A1(n12798), .A2(n12848), .A3(n12797), .A4(n12796), .ZN(
        n12799) );
  NOR3_X1 U15884 ( .A1(n12801), .A2(n12800), .A3(n12799), .ZN(n12816) );
  AOI22_X1 U15885 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12804) );
  AOI21_X1 U15886 ( .B1(n12845), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n12848), .ZN(n12803) );
  OAI211_X1 U15887 ( .C1(n12802), .C2(n12805), .A(n12804), .B(n12803), .ZN(
        n12814) );
  OAI22_X1 U15888 ( .A1(n12808), .A2(n12807), .B1(n10179), .B2(n12806), .ZN(
        n12813) );
  OAI22_X1 U15889 ( .A1(n9628), .A2(n12811), .B1(n12810), .B2(n12809), .ZN(
        n12812) );
  NOR3_X1 U15890 ( .A1(n12814), .A2(n12813), .A3(n12812), .ZN(n12815) );
  NOR2_X1 U15891 ( .A1(n12816), .A2(n12815), .ZN(n14875) );
  INV_X1 U15892 ( .A(n12818), .ZN(n14872) );
  NAND3_X1 U15893 ( .A1(n14872), .A2(n14875), .A3(n13571), .ZN(n12836) );
  AOI22_X1 U15894 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U15895 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12819) );
  NAND2_X1 U15896 ( .A1(n12820), .A2(n12819), .ZN(n12834) );
  AOI22_X1 U15897 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12822) );
  AOI21_X1 U15898 ( .B1(n12845), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n12848), .ZN(n12821) );
  OAI211_X1 U15899 ( .C1(n12802), .C2(n12823), .A(n12822), .B(n12821), .ZN(
        n12833) );
  AOI22_X1 U15900 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U15901 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12824) );
  NAND2_X1 U15902 ( .A1(n12825), .A2(n12824), .ZN(n12832) );
  AOI22_X1 U15903 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12826), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12830) );
  NAND2_X1 U15904 ( .A1(n16235), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12829) );
  NAND2_X1 U15905 ( .A1(n12827), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12828) );
  NAND4_X1 U15906 ( .A1(n12830), .A2(n12848), .A3(n12829), .A4(n12828), .ZN(
        n12831) );
  OAI22_X1 U15907 ( .A1(n12834), .A2(n12833), .B1(n12832), .B2(n12831), .ZN(
        n12835) );
  XNOR2_X1 U15908 ( .A(n12836), .B(n12835), .ZN(n14869) );
  OAI21_X1 U15909 ( .B1(n14868), .B2(n14869), .A(n9927), .ZN(n12856) );
  AOI22_X1 U15910 ( .A1(n9610), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U15911 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10185), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U15912 ( .A1(n12838), .A2(n12837), .ZN(n12853) );
  AOI22_X1 U15913 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16235), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12840) );
  AOI21_X1 U15914 ( .B1(n12845), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n12848), .ZN(n12839) );
  OAI211_X1 U15915 ( .C1(n12841), .C2(n20853), .A(n12840), .B(n12839), .ZN(
        n12852) );
  AOI22_X1 U15916 ( .A1(n10400), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12844) );
  AOI22_X1 U15917 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9627), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U15918 ( .A1(n12844), .A2(n12843), .ZN(n12851) );
  AOI22_X1 U15919 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16235), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12849) );
  NAND2_X1 U15920 ( .A1(n12826), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12847) );
  NAND2_X1 U15921 ( .A1(n12845), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12846) );
  NAND4_X1 U15922 ( .A1(n12849), .A2(n12848), .A3(n12847), .A4(n12846), .ZN(
        n12850) );
  OAI22_X1 U15923 ( .A1(n12853), .A2(n12852), .B1(n12851), .B2(n12850), .ZN(
        n12854) );
  INV_X1 U15924 ( .A(n12854), .ZN(n12855) );
  XNOR2_X1 U15925 ( .A(n12856), .B(n12855), .ZN(n14286) );
  NAND2_X1 U15926 ( .A1(n12858), .A2(n10061), .ZN(n12859) );
  NAND2_X1 U15927 ( .A1(n12857), .A2(n12859), .ZN(n12866) );
  INV_X1 U15928 ( .A(n13175), .ZN(n13170) );
  AND2_X1 U15929 ( .A1(n12860), .A2(n13170), .ZN(n12865) );
  NOR2_X1 U15930 ( .A1(n19102), .A2(n13571), .ZN(n12867) );
  OAI21_X1 U15931 ( .B1(n12867), .B2(n16265), .A(n13011), .ZN(n12861) );
  NAND2_X1 U15932 ( .A1(n12861), .A2(n10061), .ZN(n12864) );
  NAND2_X1 U15933 ( .A1(n12862), .A2(n13011), .ZN(n12863) );
  NAND2_X1 U15934 ( .A1(n12863), .A2(n19776), .ZN(n13181) );
  AND4_X1 U15935 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n13181), .ZN(
        n13150) );
  NAND2_X1 U15936 ( .A1(n13150), .A2(n12867), .ZN(n16262) );
  INV_X1 U15937 ( .A(n16262), .ZN(n12871) );
  NAND2_X1 U15938 ( .A1(n10066), .A2(n12857), .ZN(n16258) );
  NAND2_X1 U15939 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n15600) );
  AND2_X1 U15940 ( .A1(n12868), .A2(n15600), .ZN(n13330) );
  NAND2_X1 U15941 ( .A1(n16258), .A2(n13330), .ZN(n12869) );
  NOR2_X1 U15942 ( .A1(n16259), .A2(n12869), .ZN(n12870) );
  AOI21_X1 U15943 ( .B1(n16263), .B2(n12871), .A(n12870), .ZN(n13464) );
  NAND2_X1 U15944 ( .A1(n9613), .A2(n12872), .ZN(n13176) );
  NAND2_X1 U15945 ( .A1(n13464), .A2(n13176), .ZN(n12873) );
  OR2_X1 U15946 ( .A1(n18995), .A2(n10056), .ZN(n18978) );
  NAND2_X1 U15947 ( .A1(n12876), .A2(n12956), .ZN(n12881) );
  INV_X1 U15948 ( .A(n10056), .ZN(n12878) );
  NAND2_X1 U15949 ( .A1(n12878), .A2(n12901), .ZN(n12897) );
  MUX2_X1 U15950 ( .A(n13011), .B(n19757), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12879) );
  AND2_X1 U15951 ( .A1(n12897), .A2(n12879), .ZN(n12880) );
  NAND2_X1 U15952 ( .A1(n12881), .A2(n12880), .ZN(n13311) );
  NAND2_X4 U15953 ( .A1(n12883), .A2(n12882), .ZN(n13167) );
  INV_X1 U15954 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18789) );
  INV_X1 U15955 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12885) );
  NAND2_X1 U15956 ( .A1(n13571), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12884) );
  OAI211_X1 U15957 ( .C1(n13011), .C2(n12885), .A(n12884), .B(n20926), .ZN(
        n12886) );
  INV_X1 U15958 ( .A(n12886), .ZN(n12887) );
  NAND2_X1 U15959 ( .A1(n13311), .A2(n13310), .ZN(n12895) );
  INV_X1 U15960 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19659) );
  NOR2_X1 U15961 ( .A1(n13011), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U15962 ( .A1(n12900), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12901), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12888) );
  XNOR2_X1 U15963 ( .A(n12895), .B(n12890), .ZN(n13687) );
  NAND2_X1 U15964 ( .A1(n10056), .A2(n13011), .ZN(n12891) );
  MUX2_X1 U15965 ( .A(n12891), .B(n19751), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12894) );
  NAND2_X1 U15966 ( .A1(n12956), .A2(n12892), .ZN(n12893) );
  NAND2_X1 U15967 ( .A1(n12894), .A2(n12893), .ZN(n13686) );
  INV_X1 U15968 ( .A(n12895), .ZN(n13313) );
  OAI21_X1 U15969 ( .B1(n13687), .B2(n13686), .A(n9659), .ZN(n12896) );
  INV_X1 U15970 ( .A(n12896), .ZN(n12905) );
  NAND2_X1 U15971 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12898) );
  OAI211_X1 U15972 ( .C1(n12944), .C2(n12899), .A(n12898), .B(n12897), .ZN(
        n12904) );
  XNOR2_X1 U15973 ( .A(n12905), .B(n12904), .ZN(n13499) );
  INV_X1 U15974 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19661) );
  OR2_X1 U15975 ( .A1(n13167), .A2(n19661), .ZN(n12903) );
  AOI22_X1 U15976 ( .A1(n13164), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13163), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12902) );
  NAND2_X1 U15977 ( .A1(n12903), .A2(n12902), .ZN(n13498) );
  NOR2_X1 U15978 ( .A1(n13499), .A2(n13498), .ZN(n13500) );
  NOR2_X1 U15979 ( .A1(n12905), .A2(n12904), .ZN(n12906) );
  INV_X1 U15980 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U15981 ( .A1(n12956), .A2(n12907), .B1(n13164), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U15982 ( .A1(n12901), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12908) );
  OAI211_X1 U15983 ( .C1(n13167), .C2(n12910), .A(n12909), .B(n12908), .ZN(
        n13922) );
  NAND2_X1 U15984 ( .A1(n13921), .A2(n13922), .ZN(n18941) );
  INV_X1 U15985 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12911) );
  OR2_X1 U15986 ( .A1(n13167), .A2(n12911), .ZN(n12915) );
  AOI22_X1 U15987 ( .A1(n13164), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13163), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12914) );
  NAND2_X1 U15988 ( .A1(n12956), .A2(n12912), .ZN(n12913) );
  INV_X1 U15989 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U15990 ( .A1(n13164), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13163), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12918) );
  NAND2_X1 U15991 ( .A1(n12956), .A2(n12916), .ZN(n12917) );
  OAI211_X1 U15992 ( .C1(n13167), .C2(n12919), .A(n12918), .B(n12917), .ZN(
        n14097) );
  INV_X1 U15993 ( .A(n12920), .ZN(n12921) );
  NAND2_X1 U15994 ( .A1(n12956), .A2(n12921), .ZN(n12922) );
  INV_X1 U15995 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19666) );
  OR2_X1 U15996 ( .A1(n13167), .A2(n19666), .ZN(n12924) );
  AOI22_X1 U15997 ( .A1(n13164), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13163), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12923) );
  NAND2_X1 U15998 ( .A1(n12924), .A2(n12923), .ZN(n13683) );
  NAND2_X1 U15999 ( .A1(n12956), .A2(n13138), .ZN(n12925) );
  INV_X1 U16000 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19668) );
  OR2_X1 U16001 ( .A1(n13167), .A2(n19668), .ZN(n12928) );
  AOI22_X1 U16002 ( .A1(n13164), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13163), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12927) );
  NAND2_X1 U16003 ( .A1(n12928), .A2(n12927), .ZN(n13685) );
  INV_X1 U16004 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12929) );
  OR2_X1 U16005 ( .A1(n13167), .A2(n12929), .ZN(n12933) );
  AOI22_X1 U16006 ( .A1(n13164), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13163), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12932) );
  INV_X1 U16007 ( .A(n12930), .ZN(n13787) );
  NAND2_X1 U16008 ( .A1(n12956), .A2(n13787), .ZN(n12931) );
  INV_X1 U16009 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U16010 ( .A1(n13164), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13163), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U16011 ( .A1(n12956), .A2(n13799), .ZN(n12934) );
  OAI211_X1 U16012 ( .C1(n13167), .C2(n12936), .A(n12935), .B(n12934), .ZN(
        n13680) );
  INV_X1 U16013 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12937) );
  OR2_X1 U16014 ( .A1(n13167), .A2(n12937), .ZN(n12940) );
  AOI22_X1 U16015 ( .A1(n13164), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12939) );
  NAND2_X1 U16016 ( .A1(n12956), .A2(n9917), .ZN(n12938) );
  AND3_X1 U16017 ( .A1(n12940), .A2(n12939), .A3(n12938), .ZN(n13764) );
  INV_X1 U16018 ( .A(n13167), .ZN(n12941) );
  NAND2_X1 U16019 ( .A1(n12941), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16020 ( .A1(n13164), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12942) );
  OAI211_X1 U16021 ( .C1(n12944), .C2(n13912), .A(n12943), .B(n12942), .ZN(
        n13784) );
  INV_X1 U16022 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12945) );
  OR2_X1 U16023 ( .A1(n13167), .A2(n12945), .ZN(n12948) );
  AOI22_X1 U16024 ( .A1(n13164), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12947) );
  NAND2_X1 U16025 ( .A1(n12956), .A2(n9913), .ZN(n12946) );
  AND3_X1 U16026 ( .A1(n12948), .A2(n12947), .A3(n12946), .ZN(n15360) );
  INV_X1 U16027 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15152) );
  AOI22_X1 U16028 ( .A1(n13164), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12950) );
  NAND2_X1 U16029 ( .A1(n12956), .A2(n14040), .ZN(n12949) );
  OAI211_X1 U16030 ( .C1(n13167), .C2(n15152), .A(n12950), .B(n12949), .ZN(
        n13849) );
  INV_X1 U16031 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12951) );
  OR2_X1 U16032 ( .A1(n13167), .A2(n12951), .ZN(n12955) );
  AOI22_X1 U16033 ( .A1(n13164), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12954) );
  INV_X1 U16034 ( .A(n12952), .ZN(n14105) );
  NAND2_X1 U16035 ( .A1(n12956), .A2(n14105), .ZN(n12953) );
  AND3_X1 U16036 ( .A1(n12955), .A2(n12954), .A3(n12953), .ZN(n16165) );
  INV_X1 U16037 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U16038 ( .A1(n13164), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12958) );
  INV_X1 U16039 ( .A(n14173), .ZN(n14177) );
  NAND2_X1 U16040 ( .A1(n12956), .A2(n14177), .ZN(n12957) );
  OAI211_X1 U16041 ( .C1(n13167), .C2(n12959), .A(n12958), .B(n12957), .ZN(
        n13957) );
  INV_X1 U16042 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n14159) );
  OR2_X1 U16043 ( .A1(n13167), .A2(n14159), .ZN(n12961) );
  AOI22_X1 U16044 ( .A1(n13164), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12960) );
  AND2_X1 U16045 ( .A1(n12961), .A2(n12960), .ZN(n14157) );
  INV_X1 U16046 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19680) );
  OR2_X1 U16047 ( .A1(n13167), .A2(n19680), .ZN(n12963) );
  AOI22_X1 U16048 ( .A1(n13164), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12962) );
  NAND2_X1 U16049 ( .A1(n12963), .A2(n12962), .ZN(n15037) );
  NAND2_X1 U16050 ( .A1(n14155), .A2(n15037), .ZN(n15027) );
  INV_X1 U16051 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n12964) );
  OR2_X1 U16052 ( .A1(n13167), .A2(n12964), .ZN(n12966) );
  AOI22_X1 U16053 ( .A1(n13164), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12965) );
  AND2_X1 U16054 ( .A1(n12966), .A2(n12965), .ZN(n15028) );
  NOR2_X2 U16055 ( .A1(n15027), .A2(n15028), .ZN(n16006) );
  INV_X1 U16056 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20940) );
  OR2_X1 U16057 ( .A1(n13167), .A2(n20940), .ZN(n12968) );
  AOI22_X1 U16058 ( .A1(n13164), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12967) );
  NAND2_X1 U16059 ( .A1(n12968), .A2(n12967), .ZN(n16008) );
  INV_X1 U16060 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19684) );
  OR2_X1 U16061 ( .A1(n13167), .A2(n19684), .ZN(n12970) );
  AOI22_X1 U16062 ( .A1(n13164), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12969) );
  NAND2_X1 U16063 ( .A1(n12970), .A2(n12969), .ZN(n14855) );
  INV_X1 U16064 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19686) );
  OR2_X1 U16065 ( .A1(n13167), .A2(n19686), .ZN(n12972) );
  AOI22_X1 U16066 ( .A1(n13164), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12971) );
  NAND2_X1 U16067 ( .A1(n12972), .A2(n12971), .ZN(n14844) );
  INV_X1 U16068 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12973) );
  OR2_X1 U16069 ( .A1(n13167), .A2(n12973), .ZN(n12975) );
  AOI22_X1 U16070 ( .A1(n13164), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12974) );
  AND2_X1 U16071 ( .A1(n12975), .A2(n12974), .ZN(n15005) );
  INV_X1 U16072 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19688) );
  OR2_X1 U16073 ( .A1(n13167), .A2(n19688), .ZN(n12977) );
  AOI22_X1 U16074 ( .A1(n13164), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12976) );
  NAND2_X1 U16075 ( .A1(n12977), .A2(n12976), .ZN(n14996) );
  INV_X1 U16076 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n12978) );
  OR2_X1 U16077 ( .A1(n13167), .A2(n12978), .ZN(n12980) );
  AOI22_X1 U16078 ( .A1(n13164), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12979) );
  AND2_X1 U16079 ( .A1(n12980), .A2(n12979), .ZN(n13280) );
  NOR2_X2 U16080 ( .A1(n13279), .A2(n13280), .ZN(n14978) );
  INV_X1 U16081 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19691) );
  OR2_X1 U16082 ( .A1(n13167), .A2(n19691), .ZN(n12982) );
  AOI22_X1 U16083 ( .A1(n13164), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12981) );
  NAND2_X1 U16084 ( .A1(n12982), .A2(n12981), .ZN(n14979) );
  NAND2_X1 U16085 ( .A1(n14978), .A2(n14979), .ZN(n14969) );
  INV_X1 U16086 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n12983) );
  OR2_X1 U16087 ( .A1(n13167), .A2(n12983), .ZN(n12985) );
  AOI22_X1 U16088 ( .A1(n13164), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12984) );
  AND2_X1 U16089 ( .A1(n12985), .A2(n12984), .ZN(n14971) );
  NOR2_X2 U16090 ( .A1(n14969), .A2(n14971), .ZN(n14960) );
  INV_X1 U16091 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19694) );
  OR2_X1 U16092 ( .A1(n13167), .A2(n19694), .ZN(n12987) );
  AOI22_X1 U16093 ( .A1(n13164), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U16094 ( .A1(n12987), .A2(n12986), .ZN(n14961) );
  INV_X1 U16095 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19695) );
  OR2_X1 U16096 ( .A1(n13167), .A2(n19695), .ZN(n12989) );
  AOI22_X1 U16097 ( .A1(n13164), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12988) );
  NAND2_X1 U16098 ( .A1(n12989), .A2(n12988), .ZN(n14829) );
  INV_X1 U16099 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19697) );
  OR2_X1 U16100 ( .A1(n13167), .A2(n19697), .ZN(n12991) );
  AOI22_X1 U16101 ( .A1(n13164), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12990) );
  NAND2_X1 U16102 ( .A1(n12991), .A2(n12990), .ZN(n14943) );
  NAND2_X1 U16103 ( .A1(n14944), .A2(n14943), .ZN(n14946) );
  INV_X1 U16104 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12992) );
  OR2_X1 U16105 ( .A1(n13167), .A2(n12992), .ZN(n12994) );
  AOI22_X1 U16106 ( .A1(n13164), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12901), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12993) );
  AND2_X1 U16107 ( .A1(n12994), .A2(n12993), .ZN(n12995) );
  NOR2_X2 U16108 ( .A1(n14946), .A2(n12995), .ZN(n13162) );
  AOI21_X1 U16109 ( .B1(n14946), .B2(n12995), .A(n13162), .ZN(n14247) );
  NAND2_X1 U16110 ( .A1(n9593), .A2(n13011), .ZN(n12996) );
  NOR4_X1 U16111 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13000) );
  NOR4_X1 U16112 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12999) );
  NOR4_X1 U16113 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12998) );
  NOR4_X1 U16114 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12997) );
  NAND4_X1 U16115 ( .A1(n13000), .A2(n12999), .A3(n12998), .A4(n12997), .ZN(
        n13005) );
  NOR4_X1 U16116 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13003) );
  NOR4_X1 U16117 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13002) );
  NOR4_X1 U16118 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13001) );
  INV_X1 U16119 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19663) );
  NAND4_X1 U16120 ( .A1(n13003), .A2(n13002), .A3(n13001), .A4(n19663), .ZN(
        n13004) );
  OAI21_X1 U16121 ( .B1(n13005), .B2(n13004), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13380) );
  INV_X1 U16122 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13006) );
  OR2_X1 U16123 ( .A1(n19071), .A2(n13006), .ZN(n13008) );
  NAND2_X1 U16124 ( .A1(n19071), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13007) );
  AND2_X1 U16125 ( .A1(n13008), .A2(n13007), .ZN(n13355) );
  INV_X1 U16126 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13009) );
  OAI22_X1 U16127 ( .A1(n16003), .A2(n13355), .B1(n18973), .B2(n13009), .ZN(
        n13010) );
  AOI21_X1 U16128 ( .B1(n14247), .B2(n18996), .A(n13010), .ZN(n13015) );
  NAND2_X1 U16129 ( .A1(n13012), .A2(n13011), .ZN(n13013) );
  OR2_X1 U16130 ( .A1(n18995), .A2(n13013), .ZN(n13677) );
  INV_X1 U16131 ( .A(n13380), .ZN(n19070) );
  NOR2_X1 U16132 ( .A1(n13677), .A2(n19070), .ZN(n18963) );
  NOR2_X1 U16133 ( .A1(n13677), .A2(n19071), .ZN(n18962) );
  AOI22_X1 U16134 ( .A1(n18963), .A2(BUF2_REG_30__SCAN_IN), .B1(n18962), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n13014) );
  OAI21_X1 U16135 ( .B1(n14286), .B2(n18978), .A(n13016), .ZN(P2_U2889) );
  INV_X1 U16136 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13017) );
  INV_X1 U16137 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13019) );
  OAI22_X4 U16138 ( .A1(n14267), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19780), 
        .B2(n13019), .ZN(n13949) );
  INV_X4 U16139 ( .A(n13949), .ZN(n18939) );
  AOI21_X1 U16140 ( .B1(n13042), .B2(n20815), .A(n13021), .ZN(n15113) );
  AOI21_X1 U16141 ( .B1(n20810), .B2(n13023), .A(n13022), .ZN(n18798) );
  AOI21_X1 U16142 ( .B1(n15139), .B2(n13041), .A(n12528), .ZN(n15138) );
  AOI21_X1 U16143 ( .B1(n18830), .B2(n13040), .A(n13026), .ZN(n18836) );
  AOI21_X1 U16144 ( .B1(n15151), .B2(n13027), .A(n13028), .ZN(n15150) );
  AOI21_X1 U16145 ( .B1(n16073), .B2(n13039), .A(n13030), .ZN(n18890) );
  AOI21_X1 U16146 ( .B1(n18894), .B2(n13031), .A(n13032), .ZN(n18900) );
  AOI21_X1 U16147 ( .B1(n15164), .B2(n13033), .A(n13034), .ZN(n18908) );
  AOI21_X1 U16148 ( .B1(n20875), .B2(n13035), .A(n13036), .ZN(n18930) );
  AOI21_X1 U16149 ( .B1(n16125), .B2(n13037), .A(n13038), .ZN(n16114) );
  INV_X1 U16150 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13950) );
  AOI22_X1 U16151 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13308), .B1(n13950), 
        .B2(n19780), .ZN(n14057) );
  AOI22_X1 U16152 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15176), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19780), .ZN(n14056) );
  NOR2_X1 U16153 ( .A1(n14057), .A2(n14056), .ZN(n14055) );
  OAI21_X1 U16154 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13037), .ZN(n14017) );
  NAND2_X1 U16155 ( .A1(n14055), .A2(n14017), .ZN(n13919) );
  NOR2_X1 U16156 ( .A1(n16114), .A2(n13919), .ZN(n18938) );
  OAI21_X1 U16157 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13038), .A(
        n13035), .ZN(n19051) );
  NAND2_X1 U16158 ( .A1(n18938), .A2(n19051), .ZN(n18928) );
  NOR2_X1 U16159 ( .A1(n18930), .A2(n18928), .ZN(n14006) );
  OAI21_X1 U16160 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13036), .A(
        n13033), .ZN(n14199) );
  NAND2_X1 U16161 ( .A1(n14006), .A2(n14199), .ZN(n18906) );
  NOR2_X1 U16162 ( .A1(n18908), .A2(n18906), .ZN(n13980) );
  OAI21_X1 U16163 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13034), .A(
        n13031), .ZN(n16106) );
  NAND2_X1 U16164 ( .A1(n13980), .A2(n16106), .ZN(n18898) );
  NOR2_X1 U16165 ( .A1(n18900), .A2(n18898), .ZN(n13992) );
  OAI21_X1 U16166 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13032), .A(
        n13039), .ZN(n16086) );
  NAND2_X1 U16167 ( .A1(n13992), .A2(n16086), .ZN(n18880) );
  NOR2_X1 U16168 ( .A1(n18890), .A2(n18880), .ZN(n18879) );
  OAI21_X1 U16169 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13030), .A(
        n13027), .ZN(n18870) );
  NAND2_X1 U16170 ( .A1(n18879), .A2(n18870), .ZN(n18862) );
  NOR2_X1 U16171 ( .A1(n15150), .A2(n18862), .ZN(n18842) );
  OAI21_X1 U16172 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13028), .A(
        n13040), .ZN(n18843) );
  NAND2_X1 U16173 ( .A1(n18842), .A2(n18843), .ZN(n18834) );
  NOR2_X1 U16174 ( .A1(n18836), .A2(n18834), .ZN(n14152) );
  OAI21_X1 U16175 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13026), .A(
        n13041), .ZN(n16040) );
  NAND2_X1 U16176 ( .A1(n14152), .A2(n16040), .ZN(n18822) );
  NOR2_X1 U16177 ( .A1(n15138), .A2(n18822), .ZN(n18807) );
  NAND2_X1 U16178 ( .A1(n18807), .A2(n18809), .ZN(n18796) );
  NOR2_X1 U16179 ( .A1(n18798), .A2(n18796), .ZN(n14851) );
  OAI21_X1 U16180 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13022), .A(
        n13042), .ZN(n15128) );
  OAI21_X1 U16181 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13021), .A(
        n13044), .ZN(n16030) );
  INV_X1 U16182 ( .A(n16030), .ZN(n15533) );
  AOI21_X1 U16183 ( .B1(n15095), .B2(n13044), .A(n13047), .ZN(n15997) );
  NOR2_X1 U16184 ( .A1(n15996), .A2(n15997), .ZN(n15995) );
  NOR2_X1 U16185 ( .A1(n18939), .A2(n15995), .ZN(n13269) );
  OAI21_X1 U16186 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n13047), .A(
        n13046), .ZN(n16021) );
  INV_X1 U16187 ( .A(n16021), .ZN(n13271) );
  NOR2_X1 U16188 ( .A1(n13269), .A2(n13271), .ZN(n13270) );
  NOR2_X1 U16189 ( .A1(n18939), .A2(n13270), .ZN(n15986) );
  AOI21_X1 U16190 ( .B1(n15078), .B2(n13046), .A(n13049), .ZN(n15987) );
  NOR2_X1 U16191 ( .A1(n15986), .A2(n15987), .ZN(n15985) );
  NOR2_X1 U16192 ( .A1(n18939), .A2(n15985), .ZN(n15969) );
  OR2_X1 U16193 ( .A1(n13049), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13051) );
  NAND2_X1 U16194 ( .A1(n13053), .A2(n13051), .ZN(n15074) );
  INV_X1 U16195 ( .A(n15074), .ZN(n15971) );
  NOR2_X1 U16196 ( .A1(n15969), .A2(n15971), .ZN(n15970) );
  NOR2_X1 U16197 ( .A1(n18939), .A2(n15970), .ZN(n15960) );
  AOI21_X1 U16198 ( .B1(n15059), .B2(n13053), .A(n9713), .ZN(n15962) );
  NOR2_X1 U16199 ( .A1(n15950), .A2(n15952), .ZN(n15951) );
  NOR2_X1 U16200 ( .A1(n18939), .A2(n15951), .ZN(n13056) );
  XOR2_X1 U16201 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n13054), .Z(
        n15048) );
  NOR2_X1 U16202 ( .A1(n13056), .A2(n15048), .ZN(n14275) );
  INV_X1 U16203 ( .A(n14275), .ZN(n13058) );
  NOR4_X1 U16204 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n15404), .ZN(n13055) );
  INV_X1 U16205 ( .A(n18933), .ZN(n19638) );
  AOI21_X1 U16206 ( .B1(n13056), .B2(n15048), .A(n19638), .ZN(n13057) );
  NAND2_X1 U16207 ( .A1(n13058), .A2(n13057), .ZN(n13083) );
  INV_X1 U16208 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U16209 ( .A1(n13059), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13060) );
  OAI21_X1 U16210 ( .B1(n13207), .B2(n13061), .A(n13060), .ZN(n13062) );
  AOI21_X1 U16211 ( .B1(n13204), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n13062), .ZN(n13202) );
  INV_X1 U16212 ( .A(n15052), .ZN(n13071) );
  INV_X1 U16213 ( .A(n19633), .ZN(n19789) );
  INV_X1 U16214 ( .A(n16258), .ZN(n13329) );
  AND2_X1 U16215 ( .A1(n19786), .A2(n10075), .ZN(n13076) );
  NAND2_X1 U16216 ( .A1(n19725), .A2(n15600), .ZN(n13064) );
  INV_X1 U16217 ( .A(n13064), .ZN(n13077) );
  INV_X1 U16218 ( .A(n14247), .ZN(n13069) );
  INV_X1 U16219 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19642) );
  NOR2_X1 U16220 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19709) );
  INV_X1 U16221 ( .A(n19709), .ZN(n19651) );
  NAND2_X1 U16222 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19642), .ZN(n19793) );
  INV_X2 U16223 ( .A(n19793), .ZN(n19792) );
  NAND2_X2 U16224 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19792), .ZN(n19700) );
  NAND3_X1 U16225 ( .A1(n19642), .A2(n19651), .A3(n19700), .ZN(n19774) );
  INV_X1 U16226 ( .A(n19774), .ZN(n19772) );
  NAND2_X1 U16227 ( .A1(n19772), .A2(n15600), .ZN(n13148) );
  NOR2_X1 U16228 ( .A1(n13148), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16215) );
  AND2_X1 U16229 ( .A1(n16215), .A2(n19776), .ZN(n13063) );
  AND2_X1 U16230 ( .A1(n19786), .A2(n13063), .ZN(n18958) );
  INV_X1 U16231 ( .A(n18958), .ZN(n18937) );
  NOR2_X1 U16232 ( .A1(n13322), .A2(n10066), .ZN(n13332) );
  NAND2_X1 U16233 ( .A1(n13332), .A2(n13146), .ZN(n13423) );
  OR2_X1 U16234 ( .A1(n13423), .A2(n16215), .ZN(n14278) );
  INV_X1 U16235 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14277) );
  NAND3_X1 U16236 ( .A1(n13332), .A2(n13064), .A3(n14277), .ZN(n13065) );
  NAND2_X1 U16237 ( .A1(n14278), .A2(n13065), .ZN(n18927) );
  NAND2_X1 U16238 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18927), .ZN(n13068) );
  NOR3_X1 U16239 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13066), .A3(n20926), 
        .ZN(n16218) );
  NOR2_X1 U16240 ( .A1(n9691), .A2(n20926), .ZN(n18912) );
  AOI22_X1 U16241 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n9691), .ZN(n13067) );
  OAI211_X1 U16242 ( .C1(n13069), .C2(n18937), .A(n13068), .B(n13067), .ZN(
        n13070) );
  AOI21_X1 U16243 ( .B1(n13071), .B2(n18932), .A(n13070), .ZN(n13081) );
  NAND2_X1 U16244 ( .A1(n13073), .A2(n13072), .ZN(n13135) );
  NAND2_X1 U16245 ( .A1(n9593), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13074) );
  XNOR2_X1 U16246 ( .A(n13135), .B(n13074), .ZN(n13075) );
  INV_X1 U16247 ( .A(n13075), .ZN(n13132) );
  INV_X1 U16248 ( .A(n13076), .ZN(n13078) );
  AND2_X1 U16249 ( .A1(n13081), .A2(n13080), .ZN(n13082) );
  NAND2_X1 U16250 ( .A1(n13083), .A2(n13082), .ZN(P2_U2825) );
  NAND2_X1 U16251 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17458), .ZN(
        n13085) );
  INV_X1 U16252 ( .A(n13085), .ZN(n13094) );
  NAND3_X1 U16253 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n13094), .ZN(n17406) );
  NOR2_X1 U16254 ( .A1(n17432), .A2(n17406), .ZN(n13097) );
  NAND2_X1 U16255 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n13097), .ZN(
        n13096) );
  AOI21_X1 U16256 ( .B1(n17403), .B2(n13096), .A(n13084), .ZN(n17411) );
  AOI21_X1 U16257 ( .B1(n17432), .B2(n17406), .A(n13097), .ZN(n17434) );
  INV_X1 U16258 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17463) );
  NOR2_X1 U16259 ( .A1(n17463), .A2(n13085), .ZN(n13095) );
  AOI21_X1 U16260 ( .B1(n17463), .B2(n13085), .A(n13095), .ZN(n17459) );
  INV_X1 U16261 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17490) );
  NOR2_X1 U16262 ( .A1(n17755), .A2(n17507), .ZN(n13091) );
  INV_X1 U16263 ( .A(n13091), .ZN(n17485) );
  NOR2_X1 U16264 ( .A1(n17506), .A2(n17485), .ZN(n13093) );
  NAND2_X1 U16265 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13093), .ZN(
        n13087) );
  NAND3_X1 U16266 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(n13093), .ZN(n17445) );
  INV_X1 U16267 ( .A(n17445), .ZN(n13086) );
  AOI21_X1 U16268 ( .B1(n17490), .B2(n13087), .A(n13086), .ZN(n17488) );
  NAND2_X1 U16269 ( .A1(n13088), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13089) );
  INV_X1 U16270 ( .A(n13090), .ZN(n17556) );
  NOR2_X1 U16271 ( .A1(n17755), .A2(n17556), .ZN(n17555) );
  NAND2_X1 U16272 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17555), .ZN(
        n16592) );
  AOI21_X1 U16273 ( .B1(n17506), .B2(n17485), .A(n13093), .ZN(n17509) );
  NOR2_X1 U16274 ( .A1(n13286), .A2(n16717), .ZN(n16539) );
  INV_X1 U16275 ( .A(n13093), .ZN(n13092) );
  INV_X1 U16276 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U16277 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13093), .B1(
        n13092), .B2(n17496), .ZN(n17499) );
  AOI21_X1 U16278 ( .B1(n17469), .B2(n17445), .A(n13094), .ZN(n17473) );
  NOR2_X1 U16279 ( .A1(n16527), .A2(n9763), .ZN(n16522) );
  NOR2_X1 U16280 ( .A1(n17459), .A2(n16522), .ZN(n16521) );
  NOR2_X1 U16281 ( .A1(n16521), .A2(n9763), .ZN(n16507) );
  OAI21_X1 U16282 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13095), .A(
        n17406), .ZN(n17447) );
  INV_X1 U16283 ( .A(n17447), .ZN(n16508) );
  NOR2_X1 U16284 ( .A1(n16506), .A2(n9763), .ZN(n16500) );
  NOR2_X1 U16285 ( .A1(n17434), .A2(n16500), .ZN(n16499) );
  NOR2_X1 U16286 ( .A1(n16499), .A2(n9763), .ZN(n16487) );
  OAI21_X1 U16287 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n13097), .A(
        n13096), .ZN(n17421) );
  INV_X1 U16288 ( .A(n17421), .ZN(n16488) );
  AOI21_X1 U16289 ( .B1(n13098), .B2(n16469), .A(n13088), .ZN(n16468) );
  NOR2_X1 U16290 ( .A1(n16466), .A2(n9763), .ZN(n16456) );
  XOR2_X1 U16291 ( .A(n16457), .B(n16456), .Z(n13113) );
  NAND3_X1 U16292 ( .A1(n18753), .A2(n18765), .A3(n16436), .ZN(n18612) );
  NOR2_X1 U16293 ( .A1(n18714), .A2(n18612), .ZN(n16743) );
  OAI211_X1 U16294 ( .C1(n18749), .C2(n18748), .A(n18759), .B(n16436), .ZN(
        n18596) );
  INV_X1 U16295 ( .A(n18596), .ZN(n13101) );
  NAND2_X1 U16296 ( .A1(n18757), .A2(n13100), .ZN(n17330) );
  NAND2_X1 U16297 ( .A1(n18768), .A2(n10901), .ZN(n13103) );
  AOI211_X4 U16298 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18749), .A(n13101), .B(
        n13103), .ZN(n16794) );
  NAND2_X1 U16299 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18749), .ZN(n13102) );
  AOI211_X4 U16300 ( .C1(n18759), .C2(n16436), .A(n13103), .B(n13102), .ZN(
        n16793) );
  NOR3_X1 U16301 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16760) );
  INV_X1 U16302 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16758) );
  NAND2_X1 U16303 ( .A1(n16760), .A2(n16758), .ZN(n16755) );
  NOR2_X1 U16304 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16755), .ZN(n16738) );
  INV_X1 U16305 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16729) );
  NAND2_X1 U16306 ( .A1(n16738), .A2(n16729), .ZN(n16720) );
  NOR2_X1 U16307 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16720), .ZN(n16703) );
  INV_X1 U16308 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17105) );
  NAND2_X1 U16309 ( .A1(n16703), .A2(n17105), .ZN(n16694) );
  NOR2_X1 U16310 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16694), .ZN(n16677) );
  INV_X1 U16311 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16669) );
  NAND2_X1 U16312 ( .A1(n16677), .A2(n16669), .ZN(n16667) );
  NOR2_X1 U16313 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16667), .ZN(n16656) );
  INV_X1 U16314 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16651) );
  NAND2_X1 U16315 ( .A1(n16656), .A2(n16651), .ZN(n16650) );
  NOR2_X1 U16316 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16650), .ZN(n16634) );
  INV_X1 U16317 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20860) );
  NAND2_X1 U16318 ( .A1(n16634), .A2(n20860), .ZN(n16623) );
  NOR2_X1 U16319 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16623), .ZN(n16604) );
  INV_X1 U16320 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16972) );
  NAND2_X1 U16321 ( .A1(n16604), .A2(n16972), .ZN(n16594) );
  NOR2_X1 U16322 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16594), .ZN(n16583) );
  INV_X1 U16323 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16572) );
  NAND2_X1 U16324 ( .A1(n16583), .A2(n16572), .ZN(n16570) );
  NOR2_X1 U16325 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16570), .ZN(n16562) );
  INV_X1 U16326 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16918) );
  NAND2_X1 U16327 ( .A1(n16562), .A2(n16918), .ZN(n16550) );
  NOR2_X1 U16328 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16550), .ZN(n16541) );
  INV_X1 U16329 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16900) );
  NAND2_X1 U16330 ( .A1(n16541), .A2(n16900), .ZN(n16540) );
  NOR2_X1 U16331 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16540), .ZN(n16533) );
  INV_X1 U16332 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16532) );
  NAND2_X1 U16333 ( .A1(n16533), .A2(n16532), .ZN(n16531) );
  NOR2_X1 U16334 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16531), .ZN(n16520) );
  INV_X1 U16335 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16852) );
  NAND2_X1 U16336 ( .A1(n16520), .A2(n16852), .ZN(n16514) );
  NOR2_X1 U16337 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16514), .ZN(n16498) );
  INV_X1 U16338 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16846) );
  NAND2_X1 U16339 ( .A1(n16498), .A2(n16846), .ZN(n16492) );
  NOR2_X1 U16340 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16492), .ZN(n16478) );
  INV_X1 U16341 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16835) );
  NAND2_X1 U16342 ( .A1(n16478), .A2(n16835), .ZN(n13109) );
  NOR2_X1 U16343 ( .A1(n16786), .A2(n13109), .ZN(n16462) );
  OAI21_X1 U16344 ( .B1(n16794), .B2(n16462), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n13111) );
  INV_X1 U16345 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18675) );
  INV_X1 U16346 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18671) );
  INV_X1 U16347 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18653) );
  INV_X1 U16348 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18635) );
  NAND3_X1 U16349 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16746) );
  NOR2_X1 U16350 ( .A1(n18635), .A2(n16746), .ZN(n16715) );
  NAND2_X1 U16351 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16715), .ZN(n16616) );
  INV_X1 U16352 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18647) );
  INV_X1 U16353 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18645) );
  NAND3_X1 U16354 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n16661) );
  NOR3_X1 U16355 ( .A1(n18647), .A2(n18645), .A3(n16661), .ZN(n16643) );
  NAND2_X1 U16356 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16643), .ZN(n16617) );
  NOR2_X1 U16357 ( .A1(n16616), .A2(n16617), .ZN(n16635) );
  NAND2_X1 U16358 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16635), .ZN(n16621) );
  NOR2_X1 U16359 ( .A1(n18653), .A2(n16621), .ZN(n13289) );
  NAND2_X1 U16360 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n13289), .ZN(n13292) );
  INV_X1 U16361 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18666) );
  NAND3_X1 U16362 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16552) );
  NAND2_X1 U16363 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n13291) );
  NOR3_X1 U16364 ( .A1(n18666), .A2(n16552), .A3(n13291), .ZN(n13302) );
  NAND3_X1 U16365 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(n13302), .ZN(n16536) );
  NOR3_X1 U16366 ( .A1(n18671), .A2(n13292), .A3(n16536), .ZN(n16519) );
  NAND2_X1 U16367 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16519), .ZN(n16509) );
  NOR2_X1 U16368 ( .A1(n18675), .A2(n16509), .ZN(n16497) );
  NAND2_X1 U16369 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16497), .ZN(n13105) );
  NOR2_X1 U16370 ( .A1(n16784), .A2(n13105), .ZN(n16491) );
  NAND4_X1 U16371 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16491), .ZN(n16454) );
  NOR2_X1 U16372 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16454), .ZN(n16458) );
  NAND3_X1 U16373 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n13106) );
  INV_X1 U16374 ( .A(n18768), .ZN(n18755) );
  INV_X1 U16375 ( .A(n16743), .ZN(n18610) );
  NOR2_X1 U16376 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18704), .ZN(n18605) );
  NAND2_X1 U16377 ( .A1(n17760), .A2(n18605), .ZN(n18601) );
  INV_X1 U16378 ( .A(n16795), .ZN(n16764) );
  AND2_X1 U16379 ( .A1(n16766), .A2(n13105), .ZN(n16496) );
  NOR2_X1 U16380 ( .A1(n16764), .A2(n16496), .ZN(n16495) );
  INV_X1 U16381 ( .A(n16495), .ZN(n16503) );
  AOI21_X1 U16382 ( .B1(n16766), .B2(n13106), .A(n16503), .ZN(n16477) );
  INV_X1 U16383 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18686) );
  OAI22_X1 U16384 ( .A1(n16477), .A2(n18686), .B1(n13107), .B2(n16724), .ZN(
        n13108) );
  NAND2_X1 U16385 ( .A1(n16793), .A2(n13109), .ZN(n16473) );
  NAND3_X1 U16386 ( .A1(n13111), .A2(n9926), .A3(n13110), .ZN(n13112) );
  INV_X1 U16387 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14545) );
  INV_X1 U16388 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14258) );
  XNOR2_X1 U16389 ( .A(n13116), .B(n14258), .ZN(n13886) );
  AOI21_X1 U16390 ( .B1(n19941), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13117), .ZN(n13118) );
  OAI21_X1 U16391 ( .B1(n19953), .B2(n13886), .A(n13118), .ZN(n13119) );
  INV_X1 U16392 ( .A(n13119), .ZN(n13128) );
  NAND2_X1 U16393 ( .A1(n13121), .A2(n13120), .ZN(n13126) );
  AOI22_X1 U16394 ( .A1(n13123), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n13122), .ZN(n13124) );
  INV_X1 U16395 ( .A(n13124), .ZN(n13125) );
  XNOR2_X2 U16396 ( .A(n13126), .B(n13125), .ZN(n14252) );
  NAND2_X1 U16397 ( .A1(n14252), .A2(n19947), .ZN(n13127) );
  OAI211_X1 U16398 ( .C1(n13129), .C2(n19803), .A(n13128), .B(n13127), .ZN(
        P1_U2968) );
  NAND2_X1 U16399 ( .A1(n13131), .A2(n13130), .ZN(n14239) );
  AOI21_X1 U16400 ( .B1(n13075), .B2(n13138), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14240) );
  INV_X1 U16401 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13190) );
  INV_X1 U16402 ( .A(n14238), .ZN(n13133) );
  NOR2_X1 U16403 ( .A1(n9646), .A2(n13133), .ZN(n13134) );
  NOR2_X1 U16404 ( .A1(n13135), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13136) );
  MUX2_X1 U16405 ( .A(n13137), .B(n13136), .S(n9593), .Z(n14274) );
  NAND2_X1 U16406 ( .A1(n14274), .A2(n13138), .ZN(n13139) );
  XNOR2_X1 U16407 ( .A(n13139), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13140) );
  XNOR2_X1 U16408 ( .A(n13141), .B(n13140), .ZN(n14273) );
  OAI22_X1 U16409 ( .A1(n16263), .A2(n19076), .B1(n13571), .B2(n13142), .ZN(
        n13144) );
  NAND2_X1 U16410 ( .A1(n13144), .A2(n13143), .ZN(n13157) );
  MUX2_X1 U16411 ( .A(n13145), .B(n10047), .S(n13146), .Z(n13147) );
  NAND2_X1 U16412 ( .A1(n13147), .A2(n15600), .ZN(n13152) );
  INV_X1 U16413 ( .A(n13148), .ZN(n13460) );
  NAND2_X1 U16414 ( .A1(n13460), .A2(n13145), .ZN(n13149) );
  OR2_X1 U16415 ( .A1(n16259), .A2(n13149), .ZN(n13151) );
  AND2_X1 U16416 ( .A1(n13151), .A2(n13150), .ZN(n13463) );
  OAI21_X1 U16417 ( .B1(n16259), .B2(n13152), .A(n13463), .ZN(n13153) );
  NOR2_X1 U16418 ( .A1(n13154), .A2(n13153), .ZN(n13156) );
  NAND3_X1 U16419 ( .A1(n16263), .A2(n13460), .A3(n10047), .ZN(n13155) );
  NAND3_X1 U16420 ( .A1(n13157), .A2(n13156), .A3(n13155), .ZN(n13158) );
  NAND2_X1 U16421 ( .A1(n12449), .A2(n10075), .ZN(n19761) );
  OR2_X1 U16422 ( .A1(n13213), .A2(n19762), .ZN(n16207) );
  NAND2_X1 U16423 ( .A1(n16258), .A2(n13571), .ZN(n13160) );
  AND2_X1 U16424 ( .A1(n16219), .A2(n13160), .ZN(n13161) );
  INV_X1 U16425 ( .A(n19058), .ZN(n16199) );
  INV_X1 U16426 ( .A(n13162), .ZN(n13169) );
  INV_X1 U16427 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n13166) );
  AOI22_X1 U16428 ( .A1(n13164), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n13163), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13165) );
  OAI21_X1 U16429 ( .B1(n13167), .B2(n13166), .A(n13165), .ZN(n13168) );
  AND2_X1 U16430 ( .A1(n19040), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14268) );
  AOI21_X1 U16431 ( .B1(n16199), .B2(n18961), .A(n14268), .ZN(n13215) );
  INV_X1 U16432 ( .A(n15248), .ZN(n13189) );
  NAND2_X1 U16433 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16193) );
  NOR2_X1 U16434 ( .A1(n14093), .A2(n19059), .ZN(n14190) );
  NOR2_X1 U16435 ( .A1(n13213), .A2(n16262), .ZN(n15304) );
  NAND2_X1 U16436 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15389) );
  NOR2_X1 U16437 ( .A1(n13512), .A2(n15389), .ZN(n13188) );
  NAND2_X1 U16438 ( .A1(n13512), .A2(n15389), .ZN(n13517) );
  INV_X1 U16439 ( .A(n12868), .ZN(n13326) );
  NAND2_X1 U16440 ( .A1(n13170), .A2(n19102), .ZN(n13172) );
  NOR2_X1 U16441 ( .A1(n19076), .A2(n10061), .ZN(n13171) );
  AOI21_X1 U16442 ( .B1(n13326), .B2(n13172), .A(n13171), .ZN(n13179) );
  INV_X1 U16443 ( .A(n13173), .ZN(n13174) );
  NAND3_X1 U16444 ( .A1(n10074), .A2(n13175), .A3(n13174), .ZN(n13178) );
  AND4_X1 U16445 ( .A1(n13179), .A2(n13178), .A3(n13177), .A4(n13176), .ZN(
        n13185) );
  NAND2_X1 U16446 ( .A1(n13180), .A2(n13571), .ZN(n14072) );
  NAND2_X1 U16447 ( .A1(n14072), .A2(n13181), .ZN(n13183) );
  NAND2_X1 U16448 ( .A1(n13183), .A2(n13182), .ZN(n13184) );
  NAND2_X1 U16449 ( .A1(n13185), .A2(n13184), .ZN(n16243) );
  NOR2_X1 U16450 ( .A1(n16243), .A2(n13186), .ZN(n13187) );
  NOR2_X1 U16451 ( .A1(n13213), .A2(n13187), .ZN(n13191) );
  OAI211_X1 U16452 ( .C1(n15304), .C2(n13188), .A(n13517), .B(n15390), .ZN(
        n16213) );
  NOR2_X1 U16453 ( .A1(n9705), .A2(n16213), .ZN(n19055) );
  NAND3_X1 U16454 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14190), .A3(
        n19055), .ZN(n16195) );
  NAND2_X1 U16455 ( .A1(n13189), .A2(n16172), .ZN(n16139) );
  NOR2_X1 U16456 ( .A1(n16136), .A2(n16139), .ZN(n15234) );
  AND2_X1 U16457 ( .A1(n15234), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16130) );
  AND2_X1 U16458 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U16459 ( .A1(n16130), .A2(n13198), .ZN(n15195) );
  OR2_X1 U16460 ( .A1(n15195), .A2(n15062), .ZN(n15204) );
  NOR4_X1 U16461 ( .A1(n15204), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14244), .A4(n13190), .ZN(n13201) );
  INV_X1 U16462 ( .A(n15390), .ZN(n15277) );
  NOR2_X1 U16463 ( .A1(n15062), .A2(n14244), .ZN(n15182) );
  INV_X1 U16464 ( .A(n15389), .ZN(n13508) );
  INV_X1 U16465 ( .A(n13191), .ZN(n15306) );
  AOI21_X1 U16466 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13508), .A(
        n15306), .ZN(n13516) );
  INV_X2 U16467 ( .A(n19040), .ZN(n18920) );
  AND2_X1 U16468 ( .A1(n13213), .A2(n18920), .ZN(n15394) );
  INV_X1 U16469 ( .A(n15304), .ZN(n13192) );
  NOR2_X1 U16470 ( .A1(n13192), .A2(n13517), .ZN(n13509) );
  NOR4_X1 U16471 ( .A1(n13516), .A2(n15394), .A3(n13509), .A4(n9705), .ZN(
        n16214) );
  NAND3_X1 U16472 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16214), .A3(
        n14190), .ZN(n14191) );
  OR2_X1 U16473 ( .A1(n14191), .A2(n16193), .ZN(n15274) );
  OR2_X1 U16474 ( .A1(n15390), .A2(n15394), .ZN(n15273) );
  NAND2_X1 U16475 ( .A1(n15274), .A2(n15273), .ZN(n15374) );
  INV_X1 U16476 ( .A(n13193), .ZN(n13194) );
  NAND2_X1 U16477 ( .A1(n15273), .A2(n13194), .ZN(n13195) );
  AND2_X1 U16478 ( .A1(n15374), .A2(n13195), .ZN(n15240) );
  NAND2_X1 U16479 ( .A1(n15390), .A2(n13196), .ZN(n13197) );
  NAND2_X1 U16480 ( .A1(n15240), .A2(n13197), .ZN(n16128) );
  INV_X1 U16481 ( .A(n13198), .ZN(n13199) );
  AND2_X1 U16482 ( .A1(n15390), .A2(n13199), .ZN(n13200) );
  NOR2_X1 U16483 ( .A1(n16128), .A2(n13200), .ZN(n15196) );
  OAI211_X1 U16484 ( .C1(n15277), .C2(n15182), .A(n15196), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U16485 ( .A1(n13204), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13206) );
  AOI22_X1 U16486 ( .A1(n13059), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13205) );
  OAI211_X1 U16487 ( .C1(n13207), .C2(n14277), .A(n13206), .B(n13205), .ZN(
        n13208) );
  NAND2_X1 U16488 ( .A1(n13210), .A2(n13146), .ZN(n13211) );
  AND2_X1 U16489 ( .A1(n13209), .A2(n13211), .ZN(n13212) );
  OR2_X1 U16490 ( .A1(n13213), .A2(n13212), .ZN(n15384) );
  NAND2_X1 U16491 ( .A1(n12524), .A2(n13217), .ZN(n13218) );
  AND2_X1 U16492 ( .A1(n14853), .A2(n13218), .ZN(n18803) );
  INV_X1 U16493 ( .A(n18803), .ZN(n14926) );
  INV_X1 U16494 ( .A(n19048), .ZN(n16108) );
  OAI22_X1 U16495 ( .A1(n16034), .A2(n14926), .B1(n16108), .B2(n16157), .ZN(
        n13219) );
  INV_X1 U16496 ( .A(n13219), .ZN(n13231) );
  INV_X1 U16497 ( .A(n13220), .ZN(n13221) );
  NAND2_X1 U16498 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  XNOR2_X1 U16499 ( .A(n13226), .B(n13225), .ZN(n16154) );
  OAI22_X1 U16500 ( .A1(n16124), .A2(n20810), .B1(n20940), .B2(n18920), .ZN(
        n13227) );
  INV_X1 U16501 ( .A(n13228), .ZN(n13229) );
  OR2_X1 U16502 ( .A1(n13233), .A2(n13234), .ZN(n13239) );
  NAND2_X1 U16503 ( .A1(n11136), .A2(n20797), .ZN(n13533) );
  OAI21_X1 U16504 ( .B1(n13236), .B2(n13533), .A(n13584), .ZN(n13237) );
  NAND2_X1 U16505 ( .A1(n13237), .A2(n13601), .ZN(n13238) );
  NAND2_X1 U16506 ( .A1(n13239), .A2(n13238), .ZN(n13597) );
  NAND2_X1 U16507 ( .A1(n13597), .A2(n13240), .ZN(n13244) );
  NAND3_X1 U16508 ( .A1(n13242), .A2(n13532), .A3(n13241), .ZN(n13243) );
  AND2_X1 U16509 ( .A1(n14539), .A2(n14210), .ZN(n13245) );
  NAND2_X1 U16510 ( .A1(n14252), .A2(n13245), .ZN(n13263) );
  NOR4_X1 U16511 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13249) );
  NOR4_X1 U16512 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13248) );
  NOR4_X1 U16513 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13247) );
  NOR4_X1 U16514 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13246) );
  AND4_X1 U16515 ( .A1(n13249), .A2(n13248), .A3(n13247), .A4(n13246), .ZN(
        n13254) );
  NOR4_X1 U16516 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13252) );
  NOR4_X1 U16517 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13251) );
  NOR4_X1 U16518 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13250) );
  INV_X1 U16519 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20708) );
  AND4_X1 U16520 ( .A1(n13252), .A2(n13251), .A3(n13250), .A4(n20708), .ZN(
        n13253) );
  NAND2_X1 U16521 ( .A1(n13254), .A2(n13253), .ZN(n13255) );
  NOR3_X1 U16522 ( .A1(n14532), .A2(n19996), .A3(n13258), .ZN(n13256) );
  AOI22_X1 U16523 ( .A1(n14527), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14532), .ZN(n13257) );
  INV_X1 U16524 ( .A(n13257), .ZN(n13261) );
  INV_X1 U16525 ( .A(n19996), .ZN(n19994) );
  NOR2_X1 U16526 ( .A1(n13258), .A2(n19994), .ZN(n13259) );
  NAND2_X1 U16527 ( .A1(n14539), .A2(n13259), .ZN(n14518) );
  INV_X1 U16528 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16338) );
  NOR2_X1 U16529 ( .A1(n13261), .A2(n13260), .ZN(n13262) );
  NAND2_X1 U16530 ( .A1(n13263), .A2(n13262), .ZN(P1_U2873) );
  INV_X1 U16531 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20793) );
  NOR3_X1 U16532 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20793), .ZN(n13265) );
  NOR4_X1 U16533 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13264) );
  NAND4_X1 U16534 ( .A1(n19996), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13265), .A4(
        n13264), .ZN(U214) );
  NOR2_X1 U16535 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13267) );
  NOR4_X1 U16536 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13266) );
  NAND4_X1 U16537 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13267), .A4(n13266), .ZN(n13268) );
  NOR2_X1 U16538 ( .A1(n13380), .A2(n13268), .ZN(n16337) );
  NAND2_X1 U16539 ( .A1(n16337), .A2(U214), .ZN(U212) );
  NOR2_X1 U16540 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13268), .ZN(n16420)
         );
  AOI211_X1 U16541 ( .C1(n13271), .C2(n13269), .A(n13270), .B(n19638), .ZN(
        n13285) );
  INV_X1 U16542 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13272) );
  OAI22_X1 U16543 ( .A1(n13272), .A2(n18922), .B1(n12978), .B2(n18921), .ZN(
        n13284) );
  INV_X1 U16544 ( .A(n18927), .ZN(n18952) );
  INV_X1 U16545 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n13273) );
  OAI22_X1 U16546 ( .A1(n13274), .A2(n18924), .B1(n18952), .B2(n13273), .ZN(
        n13283) );
  INV_X1 U16547 ( .A(n18932), .ZN(n18954) );
  OR2_X1 U16548 ( .A1(n13277), .A2(n13276), .ZN(n13278) );
  AND2_X1 U16549 ( .A1(n13275), .A2(n13278), .ZN(n16014) );
  INV_X1 U16550 ( .A(n16014), .ZN(n13281) );
  XNOR2_X1 U16551 ( .A(n13280), .B(n14995), .ZN(n15235) );
  OAI22_X1 U16552 ( .A1(n18954), .A2(n13281), .B1(n18937), .B2(n15235), .ZN(
        n13282) );
  OR4_X1 U16553 ( .A1(n13285), .A2(n13284), .A3(n13283), .A4(n13282), .ZN(
        P2_U2831) );
  AOI211_X1 U16554 ( .C1(n17509), .C2(n13287), .A(n13286), .B(n18610), .ZN(
        n13299) );
  AOI211_X1 U16555 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16550), .A(n16541), .B(
        n16786), .ZN(n13298) );
  INV_X1 U16556 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n13288) );
  OAI22_X1 U16557 ( .A1(n17506), .A2(n16724), .B1(n16783), .B2(n13288), .ZN(
        n13297) );
  INV_X1 U16558 ( .A(n16552), .ZN(n13290) );
  INV_X1 U16559 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18656) );
  NAND2_X1 U16560 ( .A1(n16766), .A2(n13289), .ZN(n16614) );
  NOR2_X1 U16561 ( .A1(n18656), .A2(n16614), .ZN(n16591) );
  NAND2_X1 U16562 ( .A1(n13290), .A2(n16591), .ZN(n16568) );
  NOR2_X1 U16563 ( .A1(n13291), .A2(n16568), .ZN(n13295) );
  INV_X1 U16564 ( .A(n13302), .ZN(n13293) );
  OR2_X1 U16565 ( .A1(n13292), .A2(n16764), .ZN(n16603) );
  NAND2_X1 U16566 ( .A1(n16795), .A2(n16784), .ZN(n16792) );
  OAI21_X1 U16567 ( .B1(n13293), .B2(n16603), .A(n16792), .ZN(n16546) );
  INV_X1 U16568 ( .A(n16546), .ZN(n13294) );
  MUX2_X1 U16569 ( .A(n13295), .B(n13294), .S(P3_REIP_REG_20__SCAN_IN), .Z(
        n13296) );
  OR4_X1 U16570 ( .A1(n13299), .A2(n13298), .A3(n13297), .A4(n13296), .ZN(
        P3_U2651) );
  AOI211_X1 U16571 ( .C1(n17488), .C2(n13301), .A(n13300), .B(n18610), .ZN(
        n13307) );
  AOI211_X1 U16572 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16540), .A(n16533), .B(
        n16786), .ZN(n13306) );
  INV_X1 U16573 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n15490) );
  OAI22_X1 U16574 ( .A1(n17490), .A2(n16724), .B1(n16783), .B2(n15490), .ZN(
        n13305) );
  NAND2_X1 U16575 ( .A1(n13302), .A2(n16591), .ZN(n16547) );
  INV_X1 U16576 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18669) );
  XOR2_X1 U16577 ( .A(n18669), .B(P3_REIP_REG_21__SCAN_IN), .Z(n13303) );
  OAI22_X1 U16578 ( .A1(n16547), .A2(n13303), .B1(n16546), .B2(n18669), .ZN(
        n13304) );
  OR4_X1 U16579 ( .A1(n13307), .A2(n13306), .A3(n13305), .A4(n13304), .ZN(
        P3_U2649) );
  MUX2_X1 U16580 ( .A(n15390), .B(n15394), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13321) );
  NAND2_X1 U16581 ( .A1(n13946), .A2(n13308), .ZN(n13309) );
  NAND2_X1 U16582 ( .A1(n15170), .A2(n13309), .ZN(n13395) );
  NOR2_X1 U16583 ( .A1(n13311), .A2(n13310), .ZN(n13312) );
  NOR2_X1 U16584 ( .A1(n13313), .A2(n13312), .ZN(n18999) );
  INV_X1 U16585 ( .A(n18999), .ZN(n13314) );
  OAI22_X1 U16586 ( .A1(n16191), .A2(n13395), .B1(n19058), .B2(n13314), .ZN(
        n13320) );
  OR2_X1 U16587 ( .A1(n13315), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13316) );
  NAND2_X1 U16588 ( .A1(n13317), .A2(n13316), .ZN(n13397) );
  NAND2_X1 U16589 ( .A1(n19053), .A2(n15402), .ZN(n13318) );
  NAND2_X1 U16590 ( .A1(n19040), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13396) );
  OAI211_X1 U16591 ( .C1(n13397), .C2(n16207), .A(n13318), .B(n13396), .ZN(
        n13319) );
  OR3_X1 U16592 ( .A1(n13321), .A2(n13320), .A3(n13319), .ZN(P2_U3046) );
  INV_X1 U16593 ( .A(n13322), .ZN(n13324) );
  INV_X1 U16594 ( .A(n12857), .ZN(n13323) );
  NAND2_X1 U16595 ( .A1(n13324), .A2(n13323), .ZN(n18955) );
  INV_X1 U16596 ( .A(n18955), .ZN(n13953) );
  INV_X1 U16597 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13325) );
  NOR2_X1 U16598 ( .A1(n13332), .A2(n18774), .ZN(n13327) );
  OAI21_X1 U16599 ( .B1(n13953), .B2(n13325), .A(n13327), .ZN(P2_U2814) );
  NOR2_X1 U16600 ( .A1(n13953), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13328)
         );
  AOI22_X1 U16601 ( .A1(n13328), .A2(n13327), .B1(n13326), .B2(n19786), .ZN(
        P2_U3612) );
  NOR4_X1 U16602 ( .A1(n16259), .A2(n13330), .A3(n13329), .A4(n13460), .ZN(
        n16264) );
  NOR2_X1 U16603 ( .A1(n16264), .A2(n19789), .ZN(n19760) );
  OAI21_X1 U16604 ( .B1(n19760), .B2(n13466), .A(n13331), .ZN(P2_U2819) );
  INV_X2 U16605 ( .A(n13423), .ZN(n13405) );
  OAI21_X1 U16606 ( .B1(n13146), .B2(n15600), .A(n13332), .ZN(n13356) );
  AOI22_X1 U16607 ( .A1(n13405), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13356), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13334) );
  AND3_X1 U16608 ( .A1(n13332), .A2(n15600), .A3(n13571), .ZN(n13403) );
  AOI22_X1 U16609 ( .A1(n19070), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n13380), .ZN(n14981) );
  INV_X1 U16610 ( .A(n14981), .ZN(n13333) );
  NAND2_X1 U16611 ( .A1(n13403), .A2(n13333), .ZN(n13372) );
  NAND2_X1 U16612 ( .A1(n13334), .A2(n13372), .ZN(P2_U2976) );
  AOI22_X1 U16613 ( .A1(n13405), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13356), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13336) );
  AOI22_X1 U16614 ( .A1(n19070), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19071), .ZN(n14973) );
  INV_X1 U16615 ( .A(n14973), .ZN(n13335) );
  NAND2_X1 U16616 ( .A1(n13403), .A2(n13335), .ZN(n13376) );
  NAND2_X1 U16617 ( .A1(n13336), .A2(n13376), .ZN(P2_U2977) );
  AOI22_X1 U16618 ( .A1(n13405), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13356), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U16619 ( .A1(n19070), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19071), .ZN(n14988) );
  INV_X1 U16620 ( .A(n14988), .ZN(n13337) );
  NAND2_X1 U16621 ( .A1(n13403), .A2(n13337), .ZN(n13374) );
  NAND2_X1 U16622 ( .A1(n13338), .A2(n13374), .ZN(P2_U2975) );
  AOI22_X1 U16623 ( .A1(n13405), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13356), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13340) );
  AOI22_X1 U16624 ( .A1(n19070), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n13380), .ZN(n14948) );
  INV_X1 U16625 ( .A(n14948), .ZN(n13339) );
  NAND2_X1 U16626 ( .A1(n13403), .A2(n13339), .ZN(n13383) );
  NAND2_X1 U16627 ( .A1(n13340), .A2(n13383), .ZN(P2_U2980) );
  AOI22_X1 U16628 ( .A1(n13405), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13356), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U16629 ( .A1(n19070), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13380), .ZN(n19081) );
  INV_X1 U16630 ( .A(n19081), .ZN(n13341) );
  NAND2_X1 U16631 ( .A1(n13403), .A2(n13341), .ZN(n13387) );
  NAND2_X1 U16632 ( .A1(n13342), .A2(n13387), .ZN(P2_U2952) );
  AOI22_X1 U16633 ( .A1(n13405), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13356), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U16634 ( .A1(n19070), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19071), .ZN(n14964) );
  INV_X1 U16635 ( .A(n14964), .ZN(n13343) );
  NAND2_X1 U16636 ( .A1(n13403), .A2(n13343), .ZN(n13369) );
  NAND2_X1 U16637 ( .A1(n13344), .A2(n13369), .ZN(P2_U2978) );
  AOI22_X1 U16638 ( .A1(n13405), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13356), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U16639 ( .A1(n19070), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13380), .ZN(n19120) );
  INV_X1 U16640 ( .A(n19120), .ZN(n13345) );
  NAND2_X1 U16641 ( .A1(n13403), .A2(n13345), .ZN(n13347) );
  NAND2_X1 U16642 ( .A1(n13346), .A2(n13347), .ZN(P2_U2974) );
  AOI22_X1 U16643 ( .A1(n13405), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13356), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13348) );
  NAND2_X1 U16644 ( .A1(n13348), .A2(n13347), .ZN(P2_U2959) );
  AOI22_X1 U16645 ( .A1(n13405), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13356), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U16646 ( .A1(n19070), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13380), .ZN(n19109) );
  INV_X1 U16647 ( .A(n19109), .ZN(n13349) );
  NAND2_X1 U16648 ( .A1(n13403), .A2(n13349), .ZN(n13351) );
  NAND2_X1 U16649 ( .A1(n13350), .A2(n13351), .ZN(P2_U2958) );
  AOI22_X1 U16650 ( .A1(n13405), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13356), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13352) );
  NAND2_X1 U16651 ( .A1(n13352), .A2(n13351), .ZN(P2_U2973) );
  AOI22_X1 U16652 ( .A1(n13405), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13356), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13354) );
  AOI22_X1 U16653 ( .A1(n19070), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13380), .ZN(n19106) );
  INV_X1 U16654 ( .A(n19106), .ZN(n13353) );
  NAND2_X1 U16655 ( .A1(n13403), .A2(n13353), .ZN(n13365) );
  NAND2_X1 U16656 ( .A1(n13354), .A2(n13365), .ZN(P2_U2957) );
  INV_X1 U16657 ( .A(n13355), .ZN(n18966) );
  NAND2_X1 U16658 ( .A1(n13403), .A2(n18966), .ZN(n13359) );
  NAND2_X1 U16659 ( .A1(n13404), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13357) );
  OAI211_X1 U16660 ( .C1(n13009), .C2(n13423), .A(n13359), .B(n13357), .ZN(
        P2_U2966) );
  INV_X1 U16661 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19007) );
  NAND2_X1 U16662 ( .A1(n13404), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13358) );
  OAI211_X1 U16663 ( .C1(n19007), .C2(n13423), .A(n13359), .B(n13358), .ZN(
        P2_U2981) );
  INV_X1 U16664 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19011) );
  INV_X1 U16665 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16365) );
  OR2_X1 U16666 ( .A1(n19071), .A2(n16365), .ZN(n13361) );
  NAND2_X1 U16667 ( .A1(n19071), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13360) );
  AND2_X1 U16668 ( .A1(n13361), .A2(n13360), .ZN(n14953) );
  INV_X1 U16669 ( .A(n14953), .ZN(n18969) );
  NAND2_X1 U16670 ( .A1(n13403), .A2(n18969), .ZN(n13364) );
  NAND2_X1 U16671 ( .A1(n13404), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13362) );
  OAI211_X1 U16672 ( .C1(n19011), .C2(n13423), .A(n13364), .B(n13362), .ZN(
        P2_U2979) );
  INV_X1 U16673 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13432) );
  NAND2_X1 U16674 ( .A1(n13404), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13363) );
  OAI211_X1 U16675 ( .C1(n13432), .C2(n13423), .A(n13364), .B(n13363), .ZN(
        P2_U2964) );
  AOI22_X1 U16676 ( .A1(n13405), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13404), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13366) );
  NAND2_X1 U16677 ( .A1(n13366), .A2(n13365), .ZN(P2_U2972) );
  AOI22_X1 U16678 ( .A1(n13405), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13368) );
  AOI22_X1 U16679 ( .A1(n19070), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19071), .ZN(n19103) );
  INV_X1 U16680 ( .A(n19103), .ZN(n13367) );
  NAND2_X1 U16681 ( .A1(n13403), .A2(n13367), .ZN(n13385) );
  NAND2_X1 U16682 ( .A1(n13368), .A2(n13385), .ZN(P2_U2956) );
  AOI22_X1 U16683 ( .A1(n13405), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U16684 ( .A1(n13370), .A2(n13369), .ZN(P2_U2963) );
  AOI22_X1 U16685 ( .A1(n13405), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13404), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13371) );
  OAI22_X1 U16686 ( .A1(n19071), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19070), .ZN(n19098) );
  INV_X1 U16687 ( .A(n19098), .ZN(n16004) );
  NAND2_X1 U16688 ( .A1(n13403), .A2(n16004), .ZN(n13393) );
  NAND2_X1 U16689 ( .A1(n13371), .A2(n13393), .ZN(P2_U2970) );
  AOI22_X1 U16690 ( .A1(n13405), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13373) );
  NAND2_X1 U16691 ( .A1(n13373), .A2(n13372), .ZN(P2_U2961) );
  AOI22_X1 U16692 ( .A1(n13405), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13375) );
  NAND2_X1 U16693 ( .A1(n13375), .A2(n13374), .ZN(P2_U2960) );
  AOI22_X1 U16694 ( .A1(n13405), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13377) );
  NAND2_X1 U16695 ( .A1(n13377), .A2(n13376), .ZN(P2_U2962) );
  AOI22_X1 U16696 ( .A1(n13405), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U16697 ( .A1(n19070), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13380), .ZN(n19094) );
  INV_X1 U16698 ( .A(n19094), .ZN(n13378) );
  NAND2_X1 U16699 ( .A1(n13403), .A2(n13378), .ZN(n13391) );
  NAND2_X1 U16700 ( .A1(n13379), .A2(n13391), .ZN(P2_U2954) );
  AOI22_X1 U16701 ( .A1(n13405), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13382) );
  AOI22_X1 U16702 ( .A1(n19070), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13380), .ZN(n19089) );
  INV_X1 U16703 ( .A(n19089), .ZN(n13381) );
  NAND2_X1 U16704 ( .A1(n13403), .A2(n13381), .ZN(n13389) );
  NAND2_X1 U16705 ( .A1(n13382), .A2(n13389), .ZN(P2_U2953) );
  AOI22_X1 U16706 ( .A1(n13405), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13384) );
  NAND2_X1 U16707 ( .A1(n13384), .A2(n13383), .ZN(P2_U2965) );
  AOI22_X1 U16708 ( .A1(n13405), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13404), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13386) );
  NAND2_X1 U16709 ( .A1(n13386), .A2(n13385), .ZN(P2_U2971) );
  AOI22_X1 U16710 ( .A1(n13405), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13404), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U16711 ( .A1(n13388), .A2(n13387), .ZN(P2_U2967) );
  AOI22_X1 U16712 ( .A1(n13405), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13404), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13390) );
  NAND2_X1 U16713 ( .A1(n13390), .A2(n13389), .ZN(P2_U2968) );
  AOI22_X1 U16714 ( .A1(n13405), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13404), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13392) );
  NAND2_X1 U16715 ( .A1(n13392), .A2(n13391), .ZN(P2_U2969) );
  AOI22_X1 U16716 ( .A1(n13405), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13404), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13394) );
  NAND2_X1 U16717 ( .A1(n13394), .A2(n13393), .ZN(P2_U2955) );
  INV_X1 U16718 ( .A(n13395), .ZN(n13399) );
  OAI21_X1 U16719 ( .B1(n16108), .B2(n13397), .A(n13396), .ZN(n13398) );
  AOI21_X1 U16720 ( .B1(n19046), .B2(n13399), .A(n13398), .ZN(n13402) );
  OAI21_X1 U16721 ( .B1(n19041), .B2(n13400), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13401) );
  OAI211_X1 U16722 ( .C1(n16034), .C2(n13574), .A(n13402), .B(n13401), .ZN(
        P2_U3014) );
  AOI22_X1 U16723 ( .A1(n19070), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19071), .ZN(n13960) );
  INV_X1 U16724 ( .A(n13403), .ZN(n13407) );
  AOI22_X1 U16725 ( .A1(n13405), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13404), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n13406) );
  OAI21_X1 U16726 ( .B1(n13960), .B2(n13407), .A(n13406), .ZN(P2_U2982) );
  INV_X1 U16727 ( .A(n13450), .ZN(n13408) );
  OR2_X1 U16728 ( .A1(n13451), .A2(n13408), .ZN(n13441) );
  NOR2_X1 U16729 ( .A1(n13236), .A2(n19796), .ZN(n13409) );
  AND2_X1 U16730 ( .A1(n20625), .A2(n15944), .ZN(n14044) );
  INV_X1 U16731 ( .A(n14044), .ZN(n13410) );
  NAND2_X1 U16732 ( .A1(n13534), .A2(n13410), .ZN(n13435) );
  AOI21_X1 U16733 ( .B1(n13439), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13435), 
        .ZN(n13411) );
  INV_X1 U16734 ( .A(n13411), .ZN(P1_U2801) );
  AOI21_X1 U16735 ( .B1(n13414), .B2(n13413), .A(n13412), .ZN(n13503) );
  INV_X1 U16736 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14024) );
  AND2_X1 U16737 ( .A1(n19040), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13510) );
  INV_X1 U16738 ( .A(n13510), .ZN(n13415) );
  OAI21_X1 U16739 ( .B1(n16124), .B2(n14024), .A(n13415), .ZN(n13417) );
  NOR2_X1 U16740 ( .A1(n19052), .A2(n14017), .ZN(n13416) );
  AOI211_X1 U16741 ( .C1(n13503), .C2(n19048), .A(n13417), .B(n13416), .ZN(
        n13421) );
  NAND2_X1 U16742 ( .A1(n13419), .A2(n13418), .ZN(n13504) );
  NAND3_X1 U16743 ( .A1(n13505), .A2(n19046), .A3(n13504), .ZN(n13420) );
  OAI211_X1 U16744 ( .C1(n14023), .C2(n16034), .A(n13421), .B(n13420), .ZN(
        P2_U3012) );
  INV_X1 U16745 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14963) );
  NOR2_X1 U16746 ( .A1(n12857), .A2(n13146), .ZN(n13422) );
  NAND2_X1 U16747 ( .A1(n16263), .A2(n13422), .ZN(n13459) );
  OAI21_X1 U16748 ( .B1(n13459), .B2(n19789), .A(n13423), .ZN(n13424) );
  NAND2_X1 U16749 ( .A1(n19003), .A2(n13425), .ZN(n13570) );
  NAND2_X1 U16750 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n15604) );
  NOR2_X1 U16751 ( .A1(n15604), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19018) );
  INV_X1 U16752 ( .A(n19018), .ZN(n16278) );
  INV_X1 U16753 ( .A(n16278), .ZN(n19037) );
  AOI22_X1 U16754 ( .A1(n19037), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13426) );
  OAI21_X1 U16755 ( .B1(n14963), .B2(n13570), .A(n13426), .ZN(P2_U2924) );
  INV_X1 U16756 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U16757 ( .A1(n19037), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13427) );
  OAI21_X1 U16758 ( .B1(n14987), .B2(n13570), .A(n13427), .ZN(P2_U2927) );
  AOI22_X1 U16759 ( .A1(n19037), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13428) );
  OAI21_X1 U16760 ( .B1(n13009), .B2(n13570), .A(n13428), .ZN(P2_U2921) );
  INV_X1 U16761 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U16762 ( .A1(n19037), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13429) );
  OAI21_X1 U16763 ( .B1(n13430), .B2(n13570), .A(n13429), .ZN(P2_U2926) );
  AOI22_X1 U16764 ( .A1(n19037), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13431) );
  OAI21_X1 U16765 ( .B1(n13432), .B2(n13570), .A(n13431), .ZN(P2_U2923) );
  INV_X1 U16766 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U16767 ( .A1(n19037), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13433) );
  OAI21_X1 U16768 ( .B1(n14972), .B2(n13570), .A(n13433), .ZN(P2_U2925) );
  INV_X1 U16769 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14947) );
  AOI22_X1 U16770 ( .A1(n19037), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13434) );
  OAI21_X1 U16771 ( .B1(n14947), .B2(n13570), .A(n13434), .ZN(P2_U2922) );
  INV_X1 U16772 ( .A(n20795), .ZN(n13437) );
  INV_X1 U16773 ( .A(n13440), .ZN(n13436) );
  OAI22_X1 U16774 ( .A1(n13437), .A2(n13436), .B1(P1_READREQUEST_REG_SCAN_IN), 
        .B2(n13435), .ZN(n13438) );
  OAI21_X1 U16775 ( .B1(n13440), .B2(n13439), .A(n13438), .ZN(P1_U3487) );
  INV_X1 U16776 ( .A(n13441), .ZN(n13443) );
  INV_X1 U16777 ( .A(n13236), .ZN(n13442) );
  OAI22_X1 U16778 ( .A1(n13443), .A2(n13442), .B1(n13875), .B2(n13601), .ZN(
        n19797) );
  NOR3_X1 U16779 ( .A1(n13875), .A2(n13901), .A3(n13591), .ZN(n13444) );
  INV_X1 U16780 ( .A(n20797), .ZN(n20691) );
  NOR2_X1 U16781 ( .A1(n13444), .A2(n20691), .ZN(n20799) );
  NOR2_X1 U16782 ( .A1(n19797), .A2(n20799), .ZN(n15557) );
  NOR2_X1 U16783 ( .A1(n15557), .A2(n19796), .ZN(n19805) );
  INV_X1 U16784 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13458) );
  INV_X1 U16785 ( .A(n11130), .ZN(n13445) );
  AND3_X1 U16786 ( .A1(n13446), .A2(n13445), .A3(n19999), .ZN(n13447) );
  OAI21_X1 U16787 ( .B1(n13448), .B2(n13447), .A(n15574), .ZN(n13454) );
  INV_X1 U16788 ( .A(n13600), .ZN(n13449) );
  NAND2_X1 U16789 ( .A1(n13449), .A2(n13601), .ZN(n13453) );
  OR2_X1 U16790 ( .A1(n13451), .A2(n13450), .ZN(n13452) );
  NAND3_X1 U16791 ( .A1(n13454), .A2(n13453), .A3(n13452), .ZN(n13455) );
  NAND2_X1 U16792 ( .A1(n13455), .A2(n11129), .ZN(n15558) );
  INV_X1 U16793 ( .A(n15558), .ZN(n13456) );
  NAND2_X1 U16794 ( .A1(n19805), .A2(n13456), .ZN(n13457) );
  OAI21_X1 U16795 ( .B1(n19805), .B2(n13458), .A(n13457), .ZN(P1_U3484) );
  NOR2_X1 U16796 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20926), .ZN(n19075) );
  INV_X1 U16797 ( .A(n13459), .ZN(n13461) );
  NAND2_X1 U16798 ( .A1(n13461), .A2(n13460), .ZN(n13465) );
  AND4_X1 U16799 ( .A1(n13465), .A2(n13464), .A3(n13463), .A4(n13462), .ZN(
        n16271) );
  NOR2_X1 U16800 ( .A1(n19780), .A2(n15604), .ZN(n15606) );
  INV_X1 U16801 ( .A(n15606), .ZN(n16285) );
  OAI22_X1 U16802 ( .A1(n16271), .A2(n19789), .B1(n13466), .B2(n16285), .ZN(
        n13467) );
  NOR2_X1 U16803 ( .A1(n19075), .A2(n13467), .ZN(n19720) );
  INV_X1 U16804 ( .A(n19720), .ZN(n19714) );
  NAND2_X1 U16805 ( .A1(n13469), .A2(n13468), .ZN(n16268) );
  OR4_X1 U16806 ( .A1(n19720), .A2(n16269), .A3(n19726), .A4(n16268), .ZN(
        n13470) );
  OAI21_X1 U16807 ( .B1(n19714), .B2(n13471), .A(n13470), .ZN(P2_U3595) );
  NAND2_X1 U16808 ( .A1(n13473), .A2(n13472), .ZN(n13474) );
  INV_X1 U16809 ( .A(n15393), .ZN(n14060) );
  MUX2_X1 U16810 ( .A(n14060), .B(n13476), .S(n14932), .Z(n13477) );
  OAI21_X1 U16811 ( .B1(n19744), .B2(n14942), .A(n13477), .ZN(P2_U2886) );
  INV_X1 U16812 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13546) );
  NAND2_X1 U16813 ( .A1(n15544), .A2(n15568), .ZN(n13479) );
  NOR2_X1 U16814 ( .A1(n15597), .A2(n19796), .ZN(n13478) );
  NAND2_X1 U16815 ( .A1(n19908), .A2(n19999), .ZN(n13647) );
  NOR2_X1 U16816 ( .A1(n20689), .A2(n15944), .ZN(n13835) );
  INV_X1 U16817 ( .A(n13835), .ZN(n15940) );
  OR2_X1 U16818 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15940), .ZN(n19907) );
  INV_X1 U16819 ( .A(n19907), .ZN(n20798) );
  INV_X1 U16820 ( .A(n19907), .ZN(n19936) );
  AOI22_X1 U16821 ( .A1(n20798), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13480) );
  OAI21_X1 U16822 ( .B1(n13546), .B2(n13647), .A(n13480), .ZN(P1_U2912) );
  INV_X1 U16823 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13549) );
  AOI22_X1 U16824 ( .A1(n20798), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13481) );
  OAI21_X1 U16825 ( .B1(n13549), .B2(n13647), .A(n13481), .ZN(P1_U2913) );
  INV_X1 U16826 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U16827 ( .A1(n20798), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13482) );
  OAI21_X1 U16828 ( .B1(n13541), .B2(n13647), .A(n13482), .ZN(P1_U2907) );
  AOI22_X1 U16829 ( .A1(n20798), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13483) );
  OAI21_X1 U16830 ( .B1(n14492), .B2(n13647), .A(n13483), .ZN(P1_U2911) );
  INV_X1 U16831 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13536) );
  AOI22_X1 U16832 ( .A1(n20798), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13484) );
  OAI21_X1 U16833 ( .B1(n13536), .B2(n13647), .A(n13484), .ZN(P1_U2909) );
  INV_X1 U16834 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U16835 ( .A1(n20798), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13485) );
  OAI21_X1 U16836 ( .B1(n13705), .B2(n13647), .A(n13485), .ZN(P1_U2908) );
  INV_X1 U16837 ( .A(n13486), .ZN(n13490) );
  INV_X1 U16838 ( .A(n13487), .ZN(n13489) );
  OAI21_X1 U16839 ( .B1(n13490), .B2(n13489), .A(n13488), .ZN(n13961) );
  NAND2_X1 U16840 ( .A1(n13491), .A2(n14636), .ZN(n13496) );
  INV_X1 U16841 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13492) );
  NOR2_X1 U16842 ( .A1(n19957), .A2(n13492), .ZN(n13628) );
  OAI21_X1 U16843 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13494), .A(
        n13493), .ZN(n13634) );
  NOR2_X1 U16844 ( .A1(n13634), .A2(n19803), .ZN(n13495) );
  AOI211_X1 U16845 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13496), .A(
        n13628), .B(n13495), .ZN(n13497) );
  OAI21_X1 U16846 ( .B1(n19995), .B2(n13961), .A(n13497), .ZN(P1_U2999) );
  NAND2_X1 U16847 ( .A1(n13499), .A2(n13498), .ZN(n13502) );
  INV_X1 U16848 ( .A(n13500), .ZN(n13501) );
  NAND2_X1 U16849 ( .A1(n13502), .A2(n13501), .ZN(n14027) );
  INV_X1 U16850 ( .A(n14027), .ZN(n19736) );
  INV_X1 U16851 ( .A(n13503), .ZN(n13507) );
  NAND3_X1 U16852 ( .A1(n19064), .A2(n13505), .A3(n13504), .ZN(n13506) );
  OAI21_X1 U16853 ( .B1(n13507), .B2(n16207), .A(n13506), .ZN(n13515) );
  AOI21_X1 U16854 ( .B1(n15304), .B2(n13508), .A(n15394), .ZN(n13513) );
  AOI211_X1 U16855 ( .C1(n19053), .C2(n11973), .A(n13510), .B(n13509), .ZN(
        n13511) );
  OAI21_X1 U16856 ( .B1(n13513), .B2(n13512), .A(n13511), .ZN(n13514) );
  AOI211_X1 U16857 ( .C1(n13517), .C2(n13516), .A(n13515), .B(n13514), .ZN(
        n13518) );
  OAI21_X1 U16858 ( .B1(n19736), .B2(n19058), .A(n13518), .ZN(P2_U3044) );
  INV_X1 U16859 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13521) );
  MUX2_X1 U16860 ( .A(n14023), .B(n13521), .S(n14932), .Z(n13522) );
  OAI21_X1 U16861 ( .B1(n19738), .B2(n14942), .A(n13522), .ZN(P2_U2885) );
  OAI21_X1 U16862 ( .B1(n13524), .B2(n13523), .A(n13658), .ZN(n14415) );
  INV_X1 U16863 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14418) );
  INV_X1 U16864 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13525) );
  OAI22_X1 U16865 ( .A1(n14636), .A2(n14418), .B1(n19957), .B2(n13525), .ZN(
        n13526) );
  AOI21_X1 U16866 ( .B1(n15781), .B2(n14418), .A(n13526), .ZN(n13530) );
  OR2_X1 U16867 ( .A1(n13527), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14805) );
  NAND3_X1 U16868 ( .A1(n14805), .A2(n19948), .A3(n13528), .ZN(n13529) );
  OAI211_X1 U16869 ( .C1(n14415), .C2(n19995), .A(n13530), .B(n13529), .ZN(
        P1_U2998) );
  AND2_X1 U16870 ( .A1(n20800), .A2(n20691), .ZN(n13531) );
  NAND2_X1 U16871 ( .A1(n13725), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13535) );
  OR2_X1 U16872 ( .A1(n13534), .A2(n13533), .ZN(n13747) );
  INV_X1 U16873 ( .A(n13747), .ZN(n13542) );
  MUX2_X1 U16874 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n19996), .Z(
        n14484) );
  NAND2_X1 U16875 ( .A1(n13542), .A2(n14484), .ZN(n13722) );
  OAI211_X1 U16876 ( .C1(n13694), .C2(n13536), .A(n13535), .B(n13722), .ZN(
        P1_U2948) );
  INV_X1 U16877 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19922) );
  MUX2_X1 U16878 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n19996), .Z(
        n14533) );
  NAND2_X1 U16879 ( .A1(n13542), .A2(n14533), .ZN(n13544) );
  NAND2_X1 U16880 ( .A1(n13725), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13537) );
  OAI211_X1 U16881 ( .C1(n13694), .C2(n19922), .A(n13544), .B(n13537), .ZN(
        P1_U2960) );
  NAND2_X1 U16882 ( .A1(n13725), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13538) );
  MUX2_X1 U16883 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n19996), .Z(
        n14494) );
  NAND2_X1 U16884 ( .A1(n13542), .A2(n14494), .ZN(n13724) );
  OAI211_X1 U16885 ( .C1(n13694), .C2(n14492), .A(n13538), .B(n13724), .ZN(
        P1_U2946) );
  INV_X1 U16886 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13621) );
  NAND2_X1 U16887 ( .A1(n13725), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13539) );
  MUX2_X1 U16888 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n19996), .Z(
        n14473) );
  NAND2_X1 U16889 ( .A1(n13542), .A2(n14473), .ZN(n13727) );
  OAI211_X1 U16890 ( .C1(n13694), .C2(n13621), .A(n13539), .B(n13727), .ZN(
        P1_U2951) );
  NAND2_X1 U16891 ( .A1(n13728), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13540) );
  MUX2_X1 U16892 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n19996), .Z(
        n14476) );
  NAND2_X1 U16893 ( .A1(n13542), .A2(n14476), .ZN(n13730) );
  OAI211_X1 U16894 ( .C1(n13694), .C2(n13541), .A(n13540), .B(n13730), .ZN(
        P1_U2950) );
  INV_X1 U16895 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19917) );
  MUX2_X1 U16896 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n19996), .Z(
        n14487) );
  NAND2_X1 U16897 ( .A1(n13542), .A2(n14487), .ZN(n13718) );
  NAND2_X1 U16898 ( .A1(n13728), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n13543) );
  OAI211_X1 U16899 ( .C1(n13694), .C2(n19917), .A(n13718), .B(n13543), .ZN(
        P1_U2962) );
  NAND2_X1 U16900 ( .A1(n13728), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13545) );
  OAI211_X1 U16901 ( .C1(n13694), .C2(n13546), .A(n13545), .B(n13544), .ZN(
        P1_U2945) );
  INV_X1 U16902 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13639) );
  MUX2_X1 U16903 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n19996), .Z(
        n20017) );
  INV_X1 U16904 ( .A(n20017), .ZN(n13693) );
  NOR2_X1 U16905 ( .A1(n13747), .A2(n13693), .ZN(n13702) );
  AOI21_X1 U16906 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n13725), .A(n13702), 
        .ZN(n13547) );
  OAI21_X1 U16907 ( .B1(n13639), .B2(n13694), .A(n13547), .ZN(P1_U2939) );
  MUX2_X1 U16908 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n19996), .Z(
        n20042) );
  INV_X1 U16909 ( .A(n20042), .ZN(n14541) );
  NOR2_X1 U16910 ( .A1(n13747), .A2(n14541), .ZN(n13697) );
  AOI21_X1 U16911 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n13728), .A(n13697), 
        .ZN(n13548) );
  OAI21_X1 U16912 ( .B1(n13549), .B2(n13694), .A(n13548), .ZN(P1_U2944) );
  INV_X1 U16913 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13642) );
  NAND2_X1 U16914 ( .A1(n19994), .A2(DATAI_5_), .ZN(n13551) );
  NAND2_X1 U16915 ( .A1(n19996), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13550) );
  AND2_X1 U16916 ( .A1(n13551), .A2(n13550), .ZN(n20029) );
  NOR2_X1 U16917 ( .A1(n13747), .A2(n20029), .ZN(n13706) );
  AOI21_X1 U16918 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n13728), .A(n13706), 
        .ZN(n13552) );
  OAI21_X1 U16919 ( .B1(n13642), .B2(n13694), .A(n13552), .ZN(P1_U2942) );
  INV_X1 U16920 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13648) );
  NAND2_X1 U16921 ( .A1(n19994), .A2(DATAI_4_), .ZN(n13554) );
  NAND2_X1 U16922 ( .A1(n19996), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13553) );
  AND2_X1 U16923 ( .A1(n13554), .A2(n13553), .ZN(n20025) );
  NOR2_X1 U16924 ( .A1(n13747), .A2(n20025), .ZN(n13695) );
  AOI21_X1 U16925 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n13725), .A(n13695), 
        .ZN(n13555) );
  OAI21_X1 U16926 ( .B1(n13648), .B2(n13694), .A(n13555), .ZN(P1_U2941) );
  INV_X1 U16927 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13637) );
  MUX2_X1 U16928 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n19996), .Z(
        n20013) );
  INV_X1 U16929 ( .A(n20013), .ZN(n13692) );
  NOR2_X1 U16930 ( .A1(n13747), .A2(n13692), .ZN(n13716) );
  AOI21_X1 U16931 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n13725), .A(n13716), 
        .ZN(n13556) );
  OAI21_X1 U16932 ( .B1(n13637), .B2(n13694), .A(n13556), .ZN(P1_U2938) );
  INV_X1 U16933 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13644) );
  MUX2_X1 U16934 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n19996), .Z(
        n20033) );
  INV_X1 U16935 ( .A(n20033), .ZN(n13867) );
  NOR2_X1 U16936 ( .A1(n13747), .A2(n13867), .ZN(n13712) );
  AOI21_X1 U16937 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n13728), .A(n13712), 
        .ZN(n13557) );
  OAI21_X1 U16938 ( .B1(n13644), .B2(n13694), .A(n13557), .ZN(P1_U2943) );
  INV_X1 U16939 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13559) );
  AOI22_X1 U16940 ( .A1(n19037), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13558) );
  OAI21_X1 U16941 ( .B1(n13559), .B2(n13570), .A(n13558), .ZN(P2_U2928) );
  INV_X1 U16942 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U16943 ( .A1(n19037), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13560) );
  OAI21_X1 U16944 ( .B1(n15006), .B2(n13570), .A(n13560), .ZN(P2_U2929) );
  INV_X1 U16945 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13562) );
  AOI22_X1 U16946 ( .A1(n19018), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13561) );
  OAI21_X1 U16947 ( .B1(n13562), .B2(n13570), .A(n13561), .ZN(P2_U2934) );
  INV_X1 U16948 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13564) );
  AOI22_X1 U16949 ( .A1(n19018), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13563) );
  OAI21_X1 U16950 ( .B1(n13564), .B2(n13570), .A(n13563), .ZN(P2_U2930) );
  INV_X1 U16951 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U16952 ( .A1(n19018), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13565) );
  OAI21_X1 U16953 ( .B1(n15021), .B2(n13570), .A(n13565), .ZN(P2_U2931) );
  INV_X1 U16954 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U16955 ( .A1(n19018), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13566) );
  OAI21_X1 U16956 ( .B1(n13567), .B2(n13570), .A(n13566), .ZN(P2_U2932) );
  INV_X1 U16957 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14220) );
  AOI22_X1 U16958 ( .A1(n19018), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13568) );
  OAI21_X1 U16959 ( .B1(n14220), .B2(n13570), .A(n13568), .ZN(P2_U2935) );
  INV_X1 U16960 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15029) );
  AOI22_X1 U16961 ( .A1(n19018), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13569) );
  OAI21_X1 U16962 ( .B1(n15029), .B2(n13570), .A(n13569), .ZN(P2_U2933) );
  NAND2_X1 U16963 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13572) );
  AND4_X1 U16964 ( .A1(n9996), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13572), 
        .A4(n20926), .ZN(n13573) );
  MUX2_X1 U16965 ( .A(n13574), .B(n12146), .S(n13608), .Z(n13575) );
  OAI21_X1 U16966 ( .B1(n19752), .B2(n14942), .A(n13575), .ZN(P2_U2887) );
  AND3_X1 U16967 ( .A1(n13577), .A2(n12674), .A3(n13576), .ZN(n13578) );
  NAND2_X1 U16968 ( .A1(n13233), .A2(n13578), .ZN(n13579) );
  NOR2_X1 U16969 ( .A1(n13580), .A2(n13579), .ZN(n13650) );
  NAND2_X1 U16970 ( .A1(n13650), .A2(n11864), .ZN(n13819) );
  XNOR2_X1 U16971 ( .A(n15541), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13589) );
  INV_X1 U16972 ( .A(n13583), .ZN(n20002) );
  INV_X1 U16973 ( .A(n13650), .ZN(n15546) );
  NAND2_X1 U16974 ( .A1(n20002), .A2(n15546), .ZN(n13588) );
  NAND2_X1 U16975 ( .A1(n13600), .A2(n13584), .ZN(n13817) );
  XNOR2_X1 U16976 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13585) );
  NOR2_X1 U16977 ( .A1(n15544), .A2(n13585), .ZN(n13586) );
  AOI21_X1 U16978 ( .B1(n13817), .B2(n13589), .A(n13586), .ZN(n13587) );
  OAI211_X1 U16979 ( .C1(n13819), .C2(n13589), .A(n13588), .B(n13587), .ZN(
        n13807) );
  AOI22_X1 U16980 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n15889), .B2(n12654), .ZN(
        n20780) );
  NOR2_X1 U16981 ( .A1(n15944), .A2(n13626), .ZN(n20771) );
  INV_X1 U16982 ( .A(n14819), .ZN(n20774) );
  INV_X1 U16983 ( .A(n13589), .ZN(n13590) );
  AOI222_X1 U16984 ( .A1(n13807), .A2(n15934), .B1(n20780), .B2(n20771), .C1(
        n20774), .C2(n13590), .ZN(n13603) );
  NAND2_X1 U16985 ( .A1(n15544), .A2(n12674), .ZN(n13592) );
  NAND4_X1 U16986 ( .A1(n13592), .A2(n13591), .A3(n20797), .A4(n13601), .ZN(
        n13594) );
  OAI211_X1 U16987 ( .C1(n13595), .C2(n11123), .A(n13594), .B(n13593), .ZN(
        n13596) );
  INV_X1 U16988 ( .A(n13596), .ZN(n13599) );
  INV_X1 U16989 ( .A(n13597), .ZN(n13598) );
  OAI211_X1 U16990 ( .C1(n13601), .C2(n13600), .A(n13599), .B(n13598), .ZN(
        n15548) );
  INV_X1 U16991 ( .A(n15548), .ZN(n13829) );
  NAND2_X1 U16992 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13835), .ZN(n15945) );
  INV_X1 U16993 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19804) );
  OAI22_X1 U16994 ( .A1(n13829), .A2(n19796), .B1(n15945), .B2(n19804), .ZN(
        n15933) );
  AOI21_X1 U16995 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n19998), .A(n15933), 
        .ZN(n20781) );
  NAND2_X1 U16996 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20781), .ZN(
        n13602) );
  OAI21_X1 U16997 ( .B1(n13603), .B2(n20781), .A(n13602), .ZN(P1_U3472) );
  OR2_X1 U16998 ( .A1(n13606), .A2(n13605), .ZN(n13607) );
  NAND2_X1 U16999 ( .A1(n13604), .A2(n13607), .ZN(n18984) );
  INV_X1 U17000 ( .A(n13609), .ZN(n13610) );
  AOI21_X1 U17001 ( .B1(n13612), .B2(n13611), .A(n13610), .ZN(n19054) );
  INV_X1 U17002 ( .A(n19054), .ZN(n18953) );
  NOR2_X1 U17003 ( .A1(n18953), .A2(n13608), .ZN(n13613) );
  AOI21_X1 U17004 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n13608), .A(n13613), .ZN(
        n13614) );
  OAI21_X1 U17005 ( .B1(n14942), .B2(n18984), .A(n13614), .ZN(P2_U2883) );
  XNOR2_X2 U17006 ( .A(n13615), .B(n13616), .ZN(n19730) );
  NOR2_X1 U17007 ( .A1(n13617), .A2(n13608), .ZN(n13618) );
  AOI21_X1 U17008 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n13608), .A(n13618), .ZN(
        n13619) );
  OAI21_X1 U17009 ( .B1(n19730), .B2(n14942), .A(n13619), .ZN(P2_U2884) );
  AOI22_X1 U17010 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n19935), .B1(n20798), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13620) );
  OAI21_X1 U17011 ( .B1(n13621), .B2(n13647), .A(n13620), .ZN(P1_U2906) );
  OR2_X1 U17012 ( .A1(n13622), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13624) );
  NAND2_X1 U17013 ( .A1(n13624), .A2(n13623), .ZN(n13967) );
  INV_X1 U17014 ( .A(n13967), .ZN(n13629) );
  NAND2_X1 U17015 ( .A1(n13626), .A2(n13625), .ZN(n14800) );
  INV_X1 U17016 ( .A(n14800), .ZN(n13627) );
  AOI211_X1 U17017 ( .C1(n19967), .C2(n13629), .A(n13628), .B(n13627), .ZN(
        n13633) );
  INV_X1 U17018 ( .A(n13630), .ZN(n15856) );
  INV_X1 U17019 ( .A(n14801), .ZN(n13631) );
  OAI21_X1 U17020 ( .B1(n15856), .B2(n13631), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13632) );
  OAI211_X1 U17021 ( .C1(n13634), .C2(n19977), .A(n13633), .B(n13632), .ZN(
        P1_U3031) );
  INV_X1 U17022 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13709) );
  AOI22_X1 U17023 ( .A1(n20798), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13635) );
  OAI21_X1 U17024 ( .B1(n13709), .B2(n13647), .A(n13635), .ZN(P1_U2920) );
  AOI22_X1 U17025 ( .A1(n20798), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13636) );
  OAI21_X1 U17026 ( .B1(n13637), .B2(n13647), .A(n13636), .ZN(P1_U2919) );
  AOI22_X1 U17027 ( .A1(n20798), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13638) );
  OAI21_X1 U17028 ( .B1(n13639), .B2(n13647), .A(n13638), .ZN(P1_U2918) );
  INV_X1 U17029 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14516) );
  AOI22_X1 U17030 ( .A1(n20798), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13640) );
  OAI21_X1 U17031 ( .B1(n14516), .B2(n13647), .A(n13640), .ZN(P1_U2917) );
  AOI22_X1 U17032 ( .A1(n20798), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13641) );
  OAI21_X1 U17033 ( .B1(n13642), .B2(n13647), .A(n13641), .ZN(P1_U2915) );
  AOI22_X1 U17034 ( .A1(n20798), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13643) );
  OAI21_X1 U17035 ( .B1(n13644), .B2(n13647), .A(n13643), .ZN(P1_U2914) );
  INV_X1 U17036 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13720) );
  AOI22_X1 U17037 ( .A1(n20798), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13645) );
  OAI21_X1 U17038 ( .B1(n13720), .B2(n13647), .A(n13645), .ZN(P1_U2910) );
  AOI22_X1 U17039 ( .A1(n20798), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13646) );
  OAI21_X1 U17040 ( .B1(n13648), .B2(n13647), .A(n13646), .ZN(P1_U2916) );
  OAI22_X1 U17041 ( .A1(n13963), .A2(n13650), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13649), .ZN(n15540) );
  OAI22_X1 U17042 ( .A1(n15944), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14819), .ZN(n13651) );
  AOI21_X1 U17043 ( .B1(n15540), .B2(n15934), .A(n13651), .ZN(n13655) );
  NOR2_X1 U17044 ( .A1(n15544), .A2(n13652), .ZN(n15539) );
  AOI22_X1 U17045 ( .A1(n15539), .A2(n15934), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20781), .ZN(n13654) );
  OAI21_X1 U17046 ( .B1(n13655), .B2(n20781), .A(n13654), .ZN(P1_U3474) );
  NAND2_X1 U17047 ( .A1(n13656), .A2(n13657), .ZN(n13659) );
  NAND2_X1 U17048 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  AND2_X1 U17049 ( .A1(n13661), .A2(n13660), .ZN(n19890) );
  INV_X1 U17050 ( .A(n19890), .ZN(n13936) );
  NOR2_X1 U17051 ( .A1(n13663), .A2(n13662), .ZN(n19978) );
  INV_X1 U17052 ( .A(n19978), .ZN(n13665) );
  NAND3_X1 U17053 ( .A1(n13665), .A2(n19948), .A3(n13664), .ZN(n13670) );
  INV_X1 U17054 ( .A(n13666), .ZN(n19882) );
  INV_X1 U17055 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13667) );
  INV_X2 U17056 ( .A(n19957), .ZN(n19940) );
  NAND2_X1 U17057 ( .A1(n19940), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n19979) );
  OAI21_X1 U17058 ( .B1(n14636), .B2(n13667), .A(n19979), .ZN(n13668) );
  AOI21_X1 U17059 ( .B1(n19882), .B2(n15781), .A(n13668), .ZN(n13669) );
  OAI211_X1 U17060 ( .C1(n19995), .C2(n13936), .A(n13670), .B(n13669), .ZN(
        P1_U2997) );
  NAND2_X1 U17061 ( .A1(n13671), .A2(n11129), .ZN(n13672) );
  NAND2_X1 U17062 ( .A1(n19994), .A2(DATAI_0_), .ZN(n13674) );
  NAND2_X1 U17063 ( .A1(n19996), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13673) );
  AND2_X1 U17064 ( .A1(n13674), .A2(n13673), .ZN(n20005) );
  INV_X1 U17065 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19939) );
  OAI222_X1 U17066 ( .A1(n13961), .A2(n14543), .B1(n14542), .B2(n20005), .C1(
        n14539), .C2(n19939), .ZN(P1_U2904) );
  AOI21_X1 U17067 ( .B1(n13676), .B2(n13675), .A(n13679), .ZN(n16200) );
  INV_X1 U17068 ( .A(n16200), .ZN(n13678) );
  NOR2_X1 U17069 ( .A1(n18998), .A2(n18996), .ZN(n18982) );
  INV_X1 U17070 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19020) );
  OAI222_X1 U17071 ( .A1(n13678), .A2(n18982), .B1(n14988), .B2(n19002), .C1(
        n19020), .C2(n18973), .ZN(P2_U2911) );
  OR2_X1 U17072 ( .A1(n13680), .A2(n13679), .ZN(n13681) );
  NAND2_X1 U17073 ( .A1(n13681), .A2(n13763), .ZN(n18905) );
  INV_X1 U17074 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19017) );
  OAI222_X1 U17075 ( .A1(n18905), .A2(n18982), .B1(n14981), .B2(n19002), .C1(
        n19017), .C2(n18973), .ZN(P2_U2910) );
  XNOR2_X1 U17076 ( .A(n13682), .B(n13683), .ZN(n14195) );
  INV_X1 U17077 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19024) );
  OAI222_X1 U17078 ( .A1(n14195), .A2(n18982), .B1(n18973), .B2(n19024), .C1(
        n19002), .C2(n19109), .ZN(P2_U2913) );
  XNOR2_X1 U17079 ( .A(n13684), .B(n13685), .ZN(n18914) );
  INV_X1 U17080 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19022) );
  OAI222_X1 U17081 ( .A1(n18914), .A2(n18982), .B1(n18973), .B2(n19022), .C1(
        n19002), .C2(n19120), .ZN(P2_U2912) );
  XNOR2_X1 U17082 ( .A(n13687), .B(n13686), .ZN(n19749) );
  XNOR2_X1 U17083 ( .A(n19744), .B(n19749), .ZN(n13688) );
  NAND2_X1 U17084 ( .A1(n19507), .A2(n18999), .ZN(n18997) );
  NAND2_X1 U17085 ( .A1(n13688), .A2(n18997), .ZN(n13754) );
  OAI21_X1 U17086 ( .B1(n13688), .B2(n18997), .A(n13754), .ZN(n13689) );
  NAND2_X1 U17087 ( .A1(n13689), .A2(n18998), .ZN(n13691) );
  AOI22_X1 U17088 ( .A1(n18996), .A2(n19749), .B1(n18995), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13690) );
  OAI211_X1 U17089 ( .C1(n19089), .C2(n19002), .A(n13691), .B(n13690), .ZN(
        P2_U2918) );
  INV_X1 U17090 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19934) );
  OAI222_X1 U17091 ( .A1(n14415), .A2(n14543), .B1(n14542), .B2(n13692), .C1(
        n14539), .C2(n19934), .ZN(P1_U2903) );
  INV_X1 U17092 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19932) );
  OAI222_X1 U17093 ( .A1(n13936), .A2(n14543), .B1(n14542), .B2(n13693), .C1(
        n14539), .C2(n19932), .ZN(P1_U2902) );
  INV_X1 U17094 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19928) );
  AOI21_X1 U17095 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n13728), .A(n13695), 
        .ZN(n13696) );
  OAI21_X1 U17096 ( .B1(n19928), .B2(n13694), .A(n13696), .ZN(P1_U2956) );
  AOI21_X1 U17097 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n13728), .A(n13697), 
        .ZN(n13698) );
  OAI21_X1 U17098 ( .B1(n14540), .B2(n13694), .A(n13698), .ZN(P1_U2959) );
  MUX2_X1 U17099 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n19996), .Z(
        n20021) );
  INV_X1 U17100 ( .A(n20021), .ZN(n13734) );
  NOR2_X1 U17101 ( .A1(n13747), .A2(n13734), .ZN(n13700) );
  AOI21_X1 U17102 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n13725), .A(n13700), 
        .ZN(n13699) );
  OAI21_X1 U17103 ( .B1(n14516), .B2(n13694), .A(n13699), .ZN(P1_U2940) );
  INV_X1 U17104 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19930) );
  AOI21_X1 U17105 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n13728), .A(n13700), 
        .ZN(n13701) );
  OAI21_X1 U17106 ( .B1(n19930), .B2(n13694), .A(n13701), .ZN(P1_U2955) );
  AOI21_X1 U17107 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n13728), .A(n13702), 
        .ZN(n13703) );
  OAI21_X1 U17108 ( .B1(n19932), .B2(n13694), .A(n13703), .ZN(P1_U2954) );
  MUX2_X1 U17109 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n19996), .Z(
        n14480) );
  INV_X1 U17110 ( .A(n14480), .ZN(n14184) );
  NOR2_X1 U17111 ( .A1(n13747), .A2(n14184), .ZN(n13714) );
  AOI21_X1 U17112 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n13728), .A(n13714), 
        .ZN(n13704) );
  OAI21_X1 U17113 ( .B1(n13705), .B2(n13694), .A(n13704), .ZN(P1_U2949) );
  INV_X1 U17114 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19926) );
  AOI21_X1 U17115 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n13728), .A(n13706), 
        .ZN(n13707) );
  OAI21_X1 U17116 ( .B1(n19926), .B2(n13694), .A(n13707), .ZN(P1_U2957) );
  NOR2_X1 U17117 ( .A1(n13747), .A2(n20005), .ZN(n13710) );
  AOI21_X1 U17118 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n13725), .A(n13710), 
        .ZN(n13708) );
  OAI21_X1 U17119 ( .B1(n13709), .B2(n13694), .A(n13708), .ZN(P1_U2937) );
  AOI21_X1 U17120 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n13728), .A(n13710), 
        .ZN(n13711) );
  OAI21_X1 U17121 ( .B1(n19939), .B2(n13694), .A(n13711), .ZN(P1_U2952) );
  AOI21_X1 U17122 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n13728), .A(n13712), 
        .ZN(n13713) );
  OAI21_X1 U17123 ( .B1(n13868), .B2(n13694), .A(n13713), .ZN(P1_U2958) );
  AOI21_X1 U17124 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n13728), .A(n13714), 
        .ZN(n13715) );
  OAI21_X1 U17125 ( .B1(n14183), .B2(n13694), .A(n13715), .ZN(P1_U2964) );
  AOI21_X1 U17126 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n13728), .A(n13716), 
        .ZN(n13717) );
  OAI21_X1 U17127 ( .B1(n19934), .B2(n13694), .A(n13717), .ZN(P1_U2953) );
  NAND2_X1 U17128 ( .A1(n13728), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13719) );
  OAI211_X1 U17129 ( .C1(n13694), .C2(n13720), .A(n13719), .B(n13718), .ZN(
        P1_U2947) );
  INV_X1 U17130 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19915) );
  NAND2_X1 U17131 ( .A1(n13725), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13721) );
  OAI211_X1 U17132 ( .C1(n13694), .C2(n19915), .A(n13722), .B(n13721), .ZN(
        P1_U2963) );
  INV_X1 U17133 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19919) );
  NAND2_X1 U17134 ( .A1(n13728), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n13723) );
  OAI211_X1 U17135 ( .C1(n13694), .C2(n19919), .A(n13724), .B(n13723), .ZN(
        P1_U2961) );
  INV_X1 U17136 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19910) );
  NAND2_X1 U17137 ( .A1(n13725), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13726) );
  OAI211_X1 U17138 ( .C1(n13694), .C2(n19910), .A(n13727), .B(n13726), .ZN(
        P1_U2966) );
  INV_X1 U17139 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19912) );
  NAND2_X1 U17140 ( .A1(n13728), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n13729) );
  OAI211_X1 U17141 ( .C1(n13694), .C2(n19912), .A(n13730), .B(n13729), .ZN(
        P1_U2965) );
  OAI21_X1 U17142 ( .B1(n13731), .B2(n13733), .A(n13732), .ZN(n13908) );
  OAI222_X1 U17143 ( .A1(n13908), .A2(n14543), .B1(n14542), .B2(n13734), .C1(
        n14539), .C2(n19930), .ZN(P1_U2901) );
  INV_X1 U17144 ( .A(n13604), .ZN(n13737) );
  OAI211_X1 U17145 ( .C1(n13737), .C2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n14175), .B(n13736), .ZN(n13742) );
  AND2_X1 U17146 ( .A1(n13609), .A2(n13739), .ZN(n13740) );
  OR2_X1 U17147 ( .A1(n13738), .A2(n13740), .ZN(n14098) );
  INV_X1 U17148 ( .A(n14098), .ZN(n18931) );
  NAND2_X1 U17149 ( .A1(n18931), .A2(n14915), .ZN(n13741) );
  OAI211_X1 U17150 ( .C1(n14915), .C2(n13743), .A(n13742), .B(n13741), .ZN(
        P2_U2882) );
  INV_X1 U17151 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20885) );
  INV_X1 U17152 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13744) );
  NOR2_X1 U17153 ( .A1(n19994), .A2(n13744), .ZN(n13745) );
  AOI21_X1 U17154 ( .B1(DATAI_15_), .B2(n19994), .A(n13745), .ZN(n14144) );
  INV_X1 U17155 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19906) );
  OAI222_X1 U17156 ( .A1(n13694), .A2(n20885), .B1(n13747), .B2(n14144), .C1(
        n13746), .C2(n19906), .ZN(P1_U2967) );
  XOR2_X1 U17157 ( .A(n13736), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .Z(n13752)
         );
  INV_X1 U17158 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13750) );
  OAI21_X1 U17159 ( .B1(n13738), .B2(n13749), .A(n13748), .ZN(n14202) );
  MUX2_X1 U17160 ( .A(n13750), .B(n14202), .S(n14915), .Z(n13751) );
  OAI21_X1 U17161 ( .B1(n13752), .B2(n14942), .A(n13751), .ZN(P2_U2881) );
  XNOR2_X1 U17162 ( .A(n19738), .B(n14027), .ZN(n13757) );
  INV_X1 U17163 ( .A(n19749), .ZN(n13753) );
  NAND2_X1 U17164 ( .A1(n19744), .A2(n13753), .ZN(n13755) );
  NAND2_X1 U17165 ( .A1(n13755), .A2(n13754), .ZN(n13756) );
  NAND2_X1 U17166 ( .A1(n13757), .A2(n13756), .ZN(n18975) );
  OAI21_X1 U17167 ( .B1(n13757), .B2(n13756), .A(n18975), .ZN(n13758) );
  NAND2_X1 U17168 ( .A1(n13758), .A2(n18998), .ZN(n13761) );
  INV_X1 U17169 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19033) );
  OAI22_X1 U17170 ( .A1(n19002), .A2(n19094), .B1(n18973), .B2(n19033), .ZN(
        n13759) );
  AOI21_X1 U17171 ( .B1(n14027), .B2(n18996), .A(n13759), .ZN(n13760) );
  NAND2_X1 U17172 ( .A1(n13761), .A2(n13760), .ZN(P2_U2917) );
  AOI21_X1 U17173 ( .B1(n13764), .B2(n13763), .A(n13762), .ZN(n16186) );
  INV_X1 U17174 ( .A(n16186), .ZN(n13765) );
  INV_X1 U17175 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19015) );
  OAI222_X1 U17176 ( .A1(n13765), .A2(n18982), .B1(n14973), .B2(n19002), .C1(
        n19015), .C2(n18973), .ZN(P2_U2909) );
  NAND2_X1 U17177 ( .A1(n13766), .A2(n13748), .ZN(n13769) );
  INV_X1 U17178 ( .A(n13767), .ZN(n13768) );
  NAND2_X1 U17179 ( .A1(n13769), .A2(n13768), .ZN(n18913) );
  NOR2_X1 U17180 ( .A1(n13736), .A2(n13770), .ZN(n13772) );
  OAI211_X1 U17181 ( .C1(n13772), .C2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n14175), .B(n13771), .ZN(n13774) );
  INV_X1 U17182 ( .A(n14915), .ZN(n14932) );
  NAND2_X1 U17183 ( .A1(n14932), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n13773) );
  OAI211_X1 U17184 ( .C1(n18913), .C2(n14932), .A(n13774), .B(n13773), .ZN(
        P2_U2880) );
  OAI21_X1 U17185 ( .B1(n13777), .B2(n13776), .A(n13775), .ZN(n19969) );
  INV_X1 U17186 ( .A(n13908), .ZN(n13878) );
  NAND2_X1 U17187 ( .A1(n19940), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n19965) );
  NAND2_X1 U17188 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13778) );
  OAI211_X1 U17189 ( .C1(n19953), .C2(n13896), .A(n19965), .B(n13778), .ZN(
        n13779) );
  AOI21_X1 U17190 ( .B1(n13878), .B2(n19947), .A(n13779), .ZN(n13780) );
  OAI21_X1 U17191 ( .B1(n19969), .B2(n19803), .A(n13780), .ZN(P1_U2996) );
  INV_X1 U17192 ( .A(n13781), .ZN(n13782) );
  XNOR2_X1 U17193 ( .A(n13732), .B(n13782), .ZN(n19946) );
  INV_X1 U17194 ( .A(n19946), .ZN(n13783) );
  OAI222_X1 U17195 ( .A1(n14543), .A2(n13783), .B1(n14542), .B2(n20025), .C1(
        n14539), .C2(n19928), .ZN(P1_U2900) );
  OAI21_X1 U17196 ( .B1(n13784), .B2(n13762), .A(n15359), .ZN(n18882) );
  INV_X1 U17197 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19013) );
  OAI222_X1 U17198 ( .A1(n18882), .A2(n18982), .B1(n14964), .B2(n19002), .C1(
        n19013), .C2(n18973), .ZN(P2_U2908) );
  INV_X1 U17199 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13986) );
  INV_X1 U17200 ( .A(n13771), .ZN(n13788) );
  INV_X1 U17201 ( .A(n13785), .ZN(n13786) );
  OAI211_X1 U17202 ( .C1(n13788), .C2(n13787), .A(n13786), .B(n14175), .ZN(
        n13793) );
  OR2_X1 U17203 ( .A1(n13789), .A2(n13767), .ZN(n13791) );
  AND2_X1 U17204 ( .A1(n13791), .A2(n13790), .ZN(n16201) );
  NAND2_X1 U17205 ( .A1(n14915), .A2(n16201), .ZN(n13792) );
  OAI211_X1 U17206 ( .C1(n14915), .C2(n13986), .A(n13793), .B(n13792), .ZN(
        P2_U2879) );
  OR2_X1 U17207 ( .A1(n13796), .A2(n13795), .ZN(n13797) );
  AND2_X1 U17208 ( .A1(n13794), .A2(n13797), .ZN(n19862) );
  INV_X1 U17209 ( .A(n19862), .ZN(n13852) );
  OAI222_X1 U17210 ( .A1(n13852), .A2(n14543), .B1(n14542), .B2(n20029), .C1(
        n14539), .C2(n19926), .ZN(P1_U2899) );
  OAI211_X1 U17211 ( .C1(n13785), .C2(n13799), .A(n13798), .B(n14175), .ZN(
        n13805) );
  NAND2_X1 U17212 ( .A1(n13800), .A2(n13790), .ZN(n13803) );
  INV_X1 U17213 ( .A(n13801), .ZN(n13802) );
  AND2_X1 U17214 ( .A1(n13803), .A2(n13802), .ZN(n18901) );
  NAND2_X1 U17215 ( .A1(n14915), .A2(n18901), .ZN(n13804) );
  OAI211_X1 U17216 ( .C1(n14915), .C2(n13806), .A(n13805), .B(n13804), .ZN(
        P2_U2878) );
  NOR2_X1 U17217 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15944), .ZN(n13831) );
  MUX2_X1 U17218 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13807), .S(
        n15548), .Z(n15552) );
  AOI22_X1 U17219 ( .A1(n13831), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15552), .B2(n15944), .ZN(n13823) );
  AOI21_X1 U17220 ( .B1(n15541), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11330), .ZN(n13809) );
  NOR2_X1 U17221 ( .A1(n13810), .A2(n13809), .ZN(n14820) );
  MUX2_X1 U17222 ( .A(n13811), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15541), .Z(n13812) );
  XNOR2_X1 U17223 ( .A(n13813), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13814) );
  NOR2_X1 U17224 ( .A1(n15544), .A2(n13814), .ZN(n13815) );
  AOI21_X1 U17225 ( .B1(n13817), .B2(n13816), .A(n13815), .ZN(n13818) );
  OAI21_X1 U17226 ( .B1(n13819), .B2(n14820), .A(n13818), .ZN(n13820) );
  AOI21_X1 U17227 ( .B1(n20314), .B2(n15546), .A(n13820), .ZN(n14821) );
  MUX2_X1 U17228 ( .A(n11330), .B(n14821), .S(n15548), .Z(n15553) );
  INV_X1 U17229 ( .A(n15553), .ZN(n13821) );
  AOI22_X1 U17230 ( .A1(n13821), .A2(n15944), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13831), .ZN(n13822) );
  OR2_X1 U17231 ( .A1(n13823), .A2(n13822), .ZN(n15562) );
  NOR2_X1 U17232 ( .A1(n15562), .A2(n13824), .ZN(n13834) );
  INV_X1 U17233 ( .A(n20157), .ZN(n20481) );
  NOR2_X1 U17234 ( .A1(n13825), .A2(n20481), .ZN(n13826) );
  XNOR2_X1 U17235 ( .A(n13826), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19876) );
  INV_X1 U17236 ( .A(n19876), .ZN(n15936) );
  INV_X1 U17237 ( .A(n13233), .ZN(n15935) );
  AOI21_X1 U17238 ( .B1(n15936), .B2(n15935), .A(n13829), .ZN(n13827) );
  AOI211_X1 U17239 ( .C1(n13829), .C2(n13828), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n13827), .ZN(n13830) );
  AOI21_X1 U17240 ( .B1(n13831), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13830), .ZN(n15561) );
  INV_X1 U17241 ( .A(n15561), .ZN(n13832) );
  NOR3_X1 U17242 ( .A1(n13834), .A2(n13832), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n13833) );
  NOR2_X1 U17243 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20801) );
  OAI21_X1 U17244 ( .B1(n13833), .B2(n15945), .A(n20165), .ZN(n19992) );
  INV_X1 U17245 ( .A(n13834), .ZN(n13836) );
  NAND3_X1 U17246 ( .A1(n13836), .A2(n15561), .A3(n13835), .ZN(n15576) );
  INV_X1 U17247 ( .A(n15576), .ZN(n13838) );
  INV_X1 U17248 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20323) );
  AND2_X1 U17249 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20323), .ZN(n14816) );
  OAI22_X1 U17250 ( .A1(n12563), .A2(n20567), .B1(n13963), .B2(n14816), .ZN(
        n13837) );
  OAI21_X1 U17251 ( .B1(n13838), .B2(n13837), .A(n19992), .ZN(n13839) );
  OAI21_X1 U17252 ( .B1(n19992), .B2(n20521), .A(n13839), .ZN(P1_U3478) );
  NOR2_X1 U17253 ( .A1(n13583), .A2(n14816), .ZN(n13845) );
  NAND2_X1 U17254 ( .A1(n13840), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14812) );
  NOR2_X1 U17255 ( .A1(n14812), .A2(n20567), .ZN(n13843) );
  MUX2_X1 U17256 ( .A(n20621), .B(n13843), .S(n13842), .Z(n13844) );
  OAI21_X1 U17257 ( .B1(n13845), .B2(n13844), .A(n19992), .ZN(n13846) );
  OAI21_X1 U17258 ( .B1(n19992), .B2(n20394), .A(n13846), .ZN(P1_U3476) );
  OAI21_X1 U17259 ( .B1(n13849), .B2(n13848), .A(n13847), .ZN(n18868) );
  INV_X1 U17260 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19009) );
  OAI222_X1 U17261 ( .A1(n18868), .A2(n18982), .B1(n14948), .B2(n19002), .C1(
        n19009), .C2(n18973), .ZN(P2_U2906) );
  NOR2_X1 U17262 ( .A1(n13940), .A2(n13850), .ZN(n13851) );
  OR2_X1 U17263 ( .A1(n15914), .A2(n13851), .ZN(n19854) );
  INV_X1 U17264 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13853) );
  OAI222_X1 U17265 ( .A1(n19854), .A2(n14472), .B1(n13853), .B2(n19904), .C1(
        n14470), .C2(n13852), .ZN(P1_U2867) );
  OAI211_X1 U17266 ( .C1(n10219), .C2(n9917), .A(n14175), .B(n13854), .ZN(
        n13858) );
  OAI21_X1 U17267 ( .B1(n13856), .B2(n13801), .A(n13855), .ZN(n14001) );
  INV_X1 U17268 ( .A(n14001), .ZN(n16187) );
  NAND2_X1 U17269 ( .A1(n14915), .A2(n16187), .ZN(n13857) );
  OAI211_X1 U17270 ( .C1(n14915), .C2(n13997), .A(n13858), .B(n13857), .ZN(
        P2_U2877) );
  OAI222_X1 U17271 ( .A1(n13967), .A2(n14472), .B1(n14464), .B2(n13859), .C1(
        n13961), .C2(n14470), .ZN(P1_U2872) );
  NOR2_X1 U17272 ( .A1(n13861), .A2(n13862), .ZN(n13863) );
  OR2_X1 U17273 ( .A1(n13860), .A2(n13863), .ZN(n19823) );
  AOI22_X1 U17274 ( .A1(n14534), .A2(n14494), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14532), .ZN(n13864) );
  OAI21_X1 U17275 ( .B1(n19823), .B2(n14543), .A(n13864), .ZN(P1_U2895) );
  XOR2_X1 U17276 ( .A(n13794), .B(n13865), .Z(n19901) );
  INV_X1 U17277 ( .A(n19901), .ZN(n13866) );
  OAI222_X1 U17278 ( .A1(n14539), .A2(n13868), .B1(n14542), .B2(n13867), .C1(
        n14543), .C2(n13866), .ZN(P1_U2898) );
  INV_X1 U17279 ( .A(n20314), .ZN(n14817) );
  AND2_X1 U17280 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n19998), .ZN(n13870) );
  NAND2_X1 U17281 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20801), .ZN(n15573) );
  INV_X1 U17282 ( .A(n15573), .ZN(n13869) );
  AOI22_X1 U17283 ( .A1(n9602), .A2(n13870), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n13869), .ZN(n13871) );
  NAND2_X1 U17284 ( .A1(n19957), .A2(n13871), .ZN(n13872) );
  NAND2_X1 U17285 ( .A1(n14417), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13883) );
  INV_X1 U17286 ( .A(n13883), .ZN(n13876) );
  NAND2_X1 U17287 ( .A1(n13876), .A2(n13873), .ZN(n19887) );
  NOR2_X1 U17288 ( .A1(n13886), .A2(n15944), .ZN(n13874) );
  NAND2_X1 U17289 ( .A1(n13876), .A2(n13875), .ZN(n13877) );
  NAND2_X1 U17290 ( .A1(n14414), .A2(n13877), .ZN(n19889) );
  NAND2_X1 U17291 ( .A1(n13878), .A2(n19889), .ZN(n13900) );
  INV_X1 U17292 ( .A(n13939), .ZN(n13880) );
  AOI21_X1 U17293 ( .B1(n13879), .B2(n13881), .A(n13880), .ZN(n19968) );
  NAND2_X1 U17294 ( .A1(n11136), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13889) );
  AND2_X1 U17295 ( .A1(n20797), .A2(n20359), .ZN(n13884) );
  NOR2_X1 U17296 ( .A1(n13889), .A2(n13884), .ZN(n13885) );
  AND2_X1 U17297 ( .A1(n13886), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13887) );
  AND2_X2 U17298 ( .A1(n14417), .A2(n13887), .ZN(n19883) );
  INV_X1 U17299 ( .A(n19883), .ZN(n15712) );
  OR2_X1 U17300 ( .A1(n13888), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15567) );
  AND2_X1 U17301 ( .A1(n15567), .A2(n13889), .ZN(n13890) );
  NAND2_X1 U17302 ( .A1(n13892), .A2(n13890), .ZN(n19833) );
  NAND2_X1 U17303 ( .A1(n19879), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n13895) );
  INV_X1 U17304 ( .A(n15567), .ZN(n13891) );
  OAI221_X1 U17305 ( .B1(n19877), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n19877), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n14417), .ZN(n13893) );
  AOI22_X1 U17306 ( .A1(n19884), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13893), .ZN(n13894) );
  OAI211_X1 U17307 ( .C1(n15712), .C2(n13896), .A(n13895), .B(n13894), .ZN(
        n13898) );
  INV_X1 U17308 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20709) );
  AND4_X1 U17309 ( .A1(n15642), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n20709), .A4(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13897) );
  AOI211_X1 U17310 ( .C1(n19968), .C2(n19860), .A(n13898), .B(n13897), .ZN(
        n13899) );
  OAI211_X1 U17311 ( .C1(n14817), .C2(n19887), .A(n13900), .B(n13899), .ZN(
        P1_U2837) );
  XNOR2_X1 U17312 ( .A(n13902), .B(n13901), .ZN(n14804) );
  AOI22_X1 U17313 ( .A1(n19899), .A2(n14804), .B1(n14468), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13903) );
  OAI21_X1 U17314 ( .B1(n14415), .B2(n14470), .A(n13903), .ZN(P1_U2871) );
  INV_X1 U17315 ( .A(n13976), .ZN(n13904) );
  AOI21_X1 U17316 ( .B1(n13905), .B2(n14406), .A(n13904), .ZN(n19820) );
  AOI22_X1 U17317 ( .A1(n19820), .A2(n19899), .B1(n14468), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n13906) );
  OAI21_X1 U17318 ( .B1(n19823), .B2(n14470), .A(n13906), .ZN(P1_U2863) );
  AOI22_X1 U17319 ( .A1(n19968), .A2(n19899), .B1(n14468), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13907) );
  OAI21_X1 U17320 ( .B1(n13908), .B2(n14470), .A(n13907), .ZN(P1_U2869) );
  NAND2_X1 U17321 ( .A1(n13909), .A2(n13855), .ZN(n13911) );
  AND2_X1 U17322 ( .A1(n13911), .A2(n9742), .ZN(n18889) );
  INV_X1 U17323 ( .A(n18889), .ZN(n13918) );
  INV_X1 U17324 ( .A(n13854), .ZN(n13915) );
  INV_X1 U17325 ( .A(n13912), .ZN(n13914) );
  OAI211_X1 U17326 ( .C1(n13915), .C2(n13914), .A(n14175), .B(n9857), .ZN(
        n13917) );
  NAND2_X1 U17327 ( .A1(n14932), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13916) );
  OAI211_X1 U17328 ( .C1(n13918), .C2(n14932), .A(n13917), .B(n13916), .ZN(
        P2_U2876) );
  NAND2_X1 U17329 ( .A1(n14070), .A2(n13919), .ZN(n13920) );
  XNOR2_X1 U17330 ( .A(n16114), .B(n13920), .ZN(n13931) );
  NOR2_X1 U17331 ( .A1(n19730), .A2(n18955), .ZN(n13930) );
  XNOR2_X1 U17332 ( .A(n13921), .B(n13922), .ZN(n19728) );
  INV_X1 U17333 ( .A(n13617), .ZN(n16232) );
  NAND2_X1 U17334 ( .A1(n18927), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13923) );
  OAI21_X1 U17335 ( .B1(n18924), .B2(n13924), .A(n13923), .ZN(n13925) );
  AOI21_X1 U17336 ( .B1(n16232), .B2(n18932), .A(n13925), .ZN(n13928) );
  OAI22_X1 U17337 ( .A1(n16125), .A2(n18922), .B1(n12910), .B2(n18921), .ZN(
        n13926) );
  INV_X1 U17338 ( .A(n13926), .ZN(n13927) );
  OAI211_X1 U17339 ( .C1(n19728), .C2(n18937), .A(n13928), .B(n13927), .ZN(
        n13929) );
  AOI211_X1 U17340 ( .C1(n13931), .C2(n18933), .A(n13930), .B(n13929), .ZN(
        n13932) );
  INV_X1 U17341 ( .A(n13932), .ZN(P2_U2852) );
  OR2_X1 U17342 ( .A1(n13934), .A2(n13933), .ZN(n13935) );
  NAND2_X1 U17343 ( .A1(n13879), .A2(n13935), .ZN(n19984) );
  INV_X1 U17344 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13937) );
  OAI222_X1 U17345 ( .A1(n19984), .A2(n14472), .B1(n14464), .B2(n13937), .C1(
        n14470), .C2(n13936), .ZN(P1_U2870) );
  AND2_X1 U17346 ( .A1(n13939), .A2(n13938), .ZN(n13941) );
  OR2_X1 U17347 ( .A1(n13941), .A2(n13940), .ZN(n19958) );
  OAI22_X1 U17348 ( .A1(n19958), .A2(n14472), .B1(n13942), .B2(n19904), .ZN(
        n13943) );
  AOI21_X1 U17349 ( .B1(n19946), .B2(n19900), .A(n13943), .ZN(n13944) );
  INV_X1 U17350 ( .A(n13944), .ZN(P1_U2868) );
  NOR2_X1 U17351 ( .A1(n18939), .A2(n19638), .ZN(n18888) );
  INV_X1 U17352 ( .A(n18888), .ZN(n13955) );
  INV_X1 U17353 ( .A(n14057), .ZN(n14071) );
  AOI22_X1 U17354 ( .A1(n18958), .A2(n18999), .B1(P2_REIP_REG_0__SCAN_IN), 
        .B2(n9691), .ZN(n13945) );
  OAI21_X1 U17355 ( .B1(n18924), .B2(n13946), .A(n13945), .ZN(n13947) );
  AOI21_X1 U17356 ( .B1(n15402), .B2(n18932), .A(n13947), .ZN(n13948) );
  OAI21_X1 U17357 ( .B1(n18952), .B2(n12146), .A(n13948), .ZN(n13952) );
  NOR2_X1 U17358 ( .A1(n14070), .A2(n19638), .ZN(n18891) );
  INV_X1 U17359 ( .A(n18891), .ZN(n18854) );
  AOI21_X1 U17360 ( .B1(n18922), .B2(n18854), .A(n13950), .ZN(n13951) );
  AOI211_X1 U17361 ( .C1(n13953), .C2(n19507), .A(n13952), .B(n13951), .ZN(
        n13954) );
  OAI21_X1 U17362 ( .B1(n13955), .B2(n14071), .A(n13954), .ZN(P2_U2855) );
  OR2_X1 U17363 ( .A1(n13957), .A2(n13956), .ZN(n13959) );
  NAND2_X1 U17364 ( .A1(n13959), .A2(n14156), .ZN(n18841) );
  INV_X1 U17365 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19005) );
  OAI222_X1 U17366 ( .A1(n18841), .A2(n18982), .B1(n18973), .B2(n19005), .C1(
        n13960), .C2(n19002), .ZN(P2_U2904) );
  INV_X1 U17367 ( .A(n13961), .ZN(n13969) );
  OAI21_X1 U17368 ( .B1(n19884), .B2(n19883), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13962) );
  OAI21_X1 U17369 ( .B1(n19887), .B2(n13963), .A(n13962), .ZN(n13964) );
  AOI21_X1 U17370 ( .B1(P1_EBX_REG_0__SCAN_IN), .B2(n19879), .A(n13964), .ZN(
        n13966) );
  NAND2_X1 U17371 ( .A1(n19877), .A2(n14417), .ZN(n14376) );
  NAND2_X1 U17372 ( .A1(n14376), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13965) );
  OAI211_X1 U17373 ( .C1(n13967), .C2(n19893), .A(n13966), .B(n13965), .ZN(
        n13968) );
  AOI21_X1 U17374 ( .B1(n13969), .B2(n19889), .A(n13968), .ZN(n13970) );
  INV_X1 U17375 ( .A(n13970), .ZN(P1_U2840) );
  INV_X1 U17376 ( .A(n13971), .ZN(n13974) );
  INV_X1 U17377 ( .A(n13860), .ZN(n13973) );
  AOI21_X1 U17378 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n14649) );
  AND2_X1 U17379 ( .A1(n13976), .A2(n13975), .ZN(n13977) );
  OR2_X1 U17380 ( .A1(n13977), .A2(n15709), .ZN(n15875) );
  OAI22_X1 U17381 ( .A1(n15875), .A2(n14472), .B1(n14049), .B2(n19904), .ZN(
        n13978) );
  AOI21_X1 U17382 ( .B1(n14649), .B2(n19900), .A(n13978), .ZN(n13979) );
  INV_X1 U17383 ( .A(n13979), .ZN(P1_U2862) );
  NOR2_X1 U17384 ( .A1(n18939), .A2(n13980), .ZN(n13981) );
  XNOR2_X1 U17385 ( .A(n13981), .B(n16106), .ZN(n13982) );
  NAND2_X1 U17386 ( .A1(n13982), .A2(n18933), .ZN(n13991) );
  INV_X1 U17387 ( .A(n13983), .ZN(n13989) );
  AOI22_X1 U17388 ( .A1(n18958), .A2(n16200), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18947), .ZN(n13985) );
  NAND2_X1 U17389 ( .A1(n18932), .A2(n16201), .ZN(n13984) );
  OAI211_X1 U17390 ( .C1(n18952), .C2(n13986), .A(n13985), .B(n13984), .ZN(
        n13988) );
  OAI21_X1 U17391 ( .B1(n12929), .B2(n18921), .A(n18920), .ZN(n13987) );
  AOI211_X1 U17392 ( .C1(n13079), .C2(n13989), .A(n13988), .B(n13987), .ZN(
        n13990) );
  NAND2_X1 U17393 ( .A1(n13991), .A2(n13990), .ZN(P2_U2847) );
  NOR2_X1 U17394 ( .A1(n18939), .A2(n13992), .ZN(n13993) );
  XNOR2_X1 U17395 ( .A(n13993), .B(n16086), .ZN(n14003) );
  INV_X1 U17396 ( .A(n13994), .ZN(n13995) );
  AOI22_X1 U17397 ( .A1(n13995), .A2(n13079), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18947), .ZN(n13996) );
  OAI21_X1 U17398 ( .B1(n18952), .B2(n13997), .A(n13996), .ZN(n13998) );
  AOI211_X1 U17399 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n9691), .A(n13998), .B(
        n19040), .ZN(n14000) );
  NAND2_X1 U17400 ( .A1(n18958), .A2(n16186), .ZN(n13999) );
  OAI211_X1 U17401 ( .C1(n18954), .C2(n14001), .A(n14000), .B(n13999), .ZN(
        n14002) );
  AOI21_X1 U17402 ( .B1(n14003), .B2(n18933), .A(n14002), .ZN(n14004) );
  INV_X1 U17403 ( .A(n14004), .ZN(P2_U2845) );
  INV_X1 U17404 ( .A(n14649), .ZN(n14054) );
  AOI22_X1 U17405 ( .A1(n14534), .A2(n14487), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14532), .ZN(n14005) );
  OAI21_X1 U17406 ( .B1(n14054), .B2(n14543), .A(n14005), .ZN(P1_U2894) );
  NOR2_X1 U17407 ( .A1(n18939), .A2(n14006), .ZN(n14007) );
  XNOR2_X1 U17408 ( .A(n14007), .B(n14199), .ZN(n14008) );
  NAND2_X1 U17409 ( .A1(n14008), .A2(n18933), .ZN(n14016) );
  OAI21_X1 U17410 ( .B1(n19666), .B2(n18921), .A(n18920), .ZN(n14014) );
  INV_X1 U17411 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14009) );
  OAI22_X1 U17412 ( .A1(n18937), .A2(n14195), .B1(n14009), .B2(n18922), .ZN(
        n14010) );
  AOI21_X1 U17413 ( .B1(P2_EBX_REG_6__SCAN_IN), .B2(n18927), .A(n14010), .ZN(
        n14011) );
  OAI21_X1 U17414 ( .B1(n14012), .B2(n18924), .A(n14011), .ZN(n14013) );
  NOR2_X1 U17415 ( .A1(n14014), .A2(n14013), .ZN(n14015) );
  OAI211_X1 U17416 ( .C1(n14202), .C2(n18954), .A(n14016), .B(n14015), .ZN(
        P2_U2849) );
  NOR2_X1 U17417 ( .A1(n18939), .A2(n14055), .ZN(n14018) );
  XNOR2_X1 U17418 ( .A(n14018), .B(n14017), .ZN(n14019) );
  NAND2_X1 U17419 ( .A1(n14019), .A2(n18933), .ZN(n14029) );
  INV_X1 U17420 ( .A(n14020), .ZN(n14021) );
  AOI22_X1 U17421 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n18927), .B1(n13079), .B2(
        n14021), .ZN(n14022) );
  OAI21_X1 U17422 ( .B1(n14023), .B2(n18954), .A(n14022), .ZN(n14026) );
  OAI22_X1 U17423 ( .A1(n14024), .A2(n18922), .B1(n19661), .B2(n18921), .ZN(
        n14025) );
  AOI211_X1 U17424 ( .C1(n18958), .C2(n14027), .A(n14026), .B(n14025), .ZN(
        n14028) );
  OAI211_X1 U17425 ( .C1(n19738), .C2(n18955), .A(n14029), .B(n14028), .ZN(
        P2_U2853) );
  INV_X1 U17426 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n14036) );
  OAI211_X1 U17427 ( .C1(n13913), .C2(n9913), .A(n9855), .B(n14175), .ZN(
        n14035) );
  NOR2_X1 U17428 ( .A1(n14032), .A2(n13910), .ZN(n14033) );
  OR2_X1 U17429 ( .A1(n14031), .A2(n14033), .ZN(n18874) );
  INV_X1 U17430 ( .A(n18874), .ZN(n16056) );
  NAND2_X1 U17431 ( .A1(n14915), .A2(n16056), .ZN(n14034) );
  OAI211_X1 U17432 ( .C1(n14915), .C2(n14036), .A(n14035), .B(n14034), .ZN(
        P2_U2875) );
  NOR2_X1 U17433 ( .A1(n14031), .A2(n14037), .ZN(n14038) );
  OR2_X1 U17434 ( .A1(n14107), .A2(n14038), .ZN(n18857) );
  OAI211_X1 U17435 ( .C1(n14030), .C2(n14040), .A(n14039), .B(n14175), .ZN(
        n14042) );
  NAND2_X1 U17436 ( .A1(n14932), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n14041) );
  OAI211_X1 U17437 ( .C1(n18857), .C2(n14932), .A(n14042), .B(n14041), .ZN(
        P2_U2874) );
  INV_X1 U17438 ( .A(n14376), .ZN(n19838) );
  INV_X1 U17439 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20720) );
  INV_X1 U17440 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20717) );
  NAND3_X1 U17441 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14408) );
  NOR2_X1 U17442 ( .A1(n20717), .A2(n14408), .ZN(n19821) );
  NAND2_X1 U17443 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19821), .ZN(n14050) );
  NOR2_X1 U17444 ( .A1(n20720), .A2(n14050), .ZN(n14253) );
  INV_X1 U17445 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20711) );
  NAND3_X1 U17446 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19866) );
  NOR2_X1 U17447 ( .A1(n20711), .A2(n19866), .ZN(n14254) );
  NAND2_X1 U17448 ( .A1(n14417), .A2(n14254), .ZN(n14043) );
  NAND2_X1 U17449 ( .A1(n14043), .A2(n14376), .ZN(n19871) );
  OAI21_X1 U17450 ( .B1(n19838), .B2(n14253), .A(n19871), .ZN(n15715) );
  NAND2_X1 U17451 ( .A1(n14417), .A2(n14044), .ZN(n19839) );
  NOR2_X1 U17452 ( .A1(n19893), .A2(n15875), .ZN(n14045) );
  NOR2_X1 U17453 ( .A1(n19868), .A2(n14045), .ZN(n14048) );
  INV_X1 U17454 ( .A(n14647), .ZN(n14046) );
  AOI22_X1 U17455 ( .A1(n14046), .A2(n19883), .B1(n19884), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14047) );
  OAI211_X1 U17456 ( .C1(n19833), .C2(n14049), .A(n14048), .B(n14047), .ZN(
        n14052) );
  NOR3_X1 U17457 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14050), .A3(n19857), 
        .ZN(n14051) );
  AOI211_X1 U17458 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n15715), .A(n14052), 
        .B(n14051), .ZN(n14053) );
  OAI21_X1 U17459 ( .B1(n14054), .B2(n14414), .A(n14053), .ZN(P1_U2830) );
  AOI211_X1 U17460 ( .C1(n14057), .C2(n14056), .A(n18939), .B(n14055), .ZN(
        n14069) );
  INV_X1 U17461 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15173) );
  AOI22_X1 U17462 ( .A1(n14069), .A2(n18933), .B1(n18891), .B2(n15173), .ZN(
        n14064) );
  NAND2_X1 U17463 ( .A1(n18927), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U17464 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n9691), .ZN(n14058) );
  OAI211_X1 U17465 ( .C1(n18924), .C2(n15171), .A(n14059), .B(n14058), .ZN(
        n14062) );
  NOR2_X1 U17466 ( .A1(n14060), .A2(n18954), .ZN(n14061) );
  AOI211_X1 U17467 ( .C1(n18958), .C2(n19749), .A(n14062), .B(n14061), .ZN(
        n14063) );
  OAI211_X1 U17468 ( .C1(n19744), .C2(n18955), .A(n14064), .B(n14063), .ZN(
        P2_U2854) );
  NOR2_X1 U17469 ( .A1(n14065), .A2(n14066), .ZN(n14067) );
  OR2_X1 U17470 ( .A1(n9641), .A2(n14067), .ZN(n14626) );
  AOI22_X1 U17471 ( .A1(n14534), .A2(n14473), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14532), .ZN(n14068) );
  OAI21_X1 U17472 ( .B1(n14626), .B2(n14543), .A(n14068), .ZN(P1_U2890) );
  AOI21_X1 U17473 ( .B1(n18939), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n14069), .ZN(n19716) );
  AOI22_X1 U17474 ( .A1(n18939), .A2(n13308), .B1(n14071), .B2(n14070), .ZN(
        n15403) );
  NAND2_X1 U17475 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15403), .ZN(n19717) );
  INV_X1 U17476 ( .A(n19717), .ZN(n14080) );
  INV_X1 U17477 ( .A(n14072), .ZN(n14073) );
  OR2_X1 U17478 ( .A1(n14073), .A2(n10552), .ZN(n15400) );
  OAI21_X1 U17479 ( .B1(n14075), .B2(n14074), .A(n15400), .ZN(n14077) );
  NAND2_X1 U17480 ( .A1(n13210), .A2(n9854), .ZN(n14076) );
  NAND2_X1 U17481 ( .A1(n14077), .A2(n14076), .ZN(n14078) );
  AOI21_X1 U17482 ( .B1(n15393), .B2(n16243), .A(n14078), .ZN(n16248) );
  OAI22_X1 U17483 ( .A1(n19744), .A2(n19719), .B1(n16248), .B2(n19726), .ZN(
        n14079) );
  AOI21_X1 U17484 ( .B1(n19716), .B2(n14080), .A(n14079), .ZN(n14082) );
  NAND2_X1 U17485 ( .A1(n19720), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14081) );
  OAI21_X1 U17486 ( .B1(n14082), .B2(n19720), .A(n14081), .ZN(P2_U3600) );
  XNOR2_X1 U17487 ( .A(n14083), .B(n14084), .ZN(n16110) );
  INV_X1 U17488 ( .A(n14085), .ZN(n14089) );
  NAND2_X1 U17489 ( .A1(n14086), .A2(n14085), .ZN(n14087) );
  NAND2_X1 U17490 ( .A1(n9682), .A2(n14087), .ZN(n14088) );
  OAI21_X1 U17491 ( .B1(n14090), .B2(n14089), .A(n14088), .ZN(n16107) );
  INV_X1 U17492 ( .A(n15273), .ZN(n14091) );
  OR2_X1 U17493 ( .A1(n16214), .A2(n14091), .ZN(n19060) );
  INV_X1 U17494 ( .A(n19060), .ZN(n14096) );
  NOR2_X1 U17495 ( .A1(n12919), .A2(n18920), .ZN(n14095) );
  INV_X1 U17496 ( .A(n19055), .ZN(n14092) );
  AOI211_X1 U17497 ( .C1(n14093), .C2(n19059), .A(n14190), .B(n14092), .ZN(
        n14094) );
  AOI211_X1 U17498 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n14096), .A(
        n14095), .B(n14094), .ZN(n14101) );
  XNOR2_X1 U17499 ( .A(n14097), .B(n18943), .ZN(n18981) );
  OAI22_X1 U17500 ( .A1(n14098), .A2(n15384), .B1(n18981), .B2(n19058), .ZN(
        n14099) );
  INV_X1 U17501 ( .A(n14099), .ZN(n14100) );
  OAI211_X1 U17502 ( .C1(n16107), .C2(n16207), .A(n14101), .B(n14100), .ZN(
        n14102) );
  INV_X1 U17503 ( .A(n14102), .ZN(n14103) );
  OAI21_X1 U17504 ( .B1(n16191), .B2(n16110), .A(n14103), .ZN(P2_U3041) );
  INV_X1 U17505 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n18845) );
  INV_X1 U17506 ( .A(n14039), .ZN(n14106) );
  OAI211_X1 U17507 ( .C1(n14106), .C2(n14105), .A(n14175), .B(n14174), .ZN(
        n14113) );
  INV_X1 U17508 ( .A(n14107), .ZN(n14110) );
  INV_X1 U17509 ( .A(n14108), .ZN(n14109) );
  NAND2_X1 U17510 ( .A1(n14110), .A2(n14109), .ZN(n14111) );
  AND2_X1 U17511 ( .A1(n14171), .A2(n14111), .ZN(n18850) );
  NAND2_X1 U17512 ( .A1(n14915), .A2(n18850), .ZN(n14112) );
  OAI211_X1 U17513 ( .C1(n14915), .C2(n18845), .A(n14113), .B(n14112), .ZN(
        P2_U2873) );
  AND2_X1 U17514 ( .A1(n14125), .A2(n14114), .ZN(n14115) );
  OR2_X1 U17515 ( .A1(n14115), .A2(n15682), .ZN(n15847) );
  INV_X1 U17516 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14116) );
  OAI222_X1 U17517 ( .A1(n15847), .A2(n14472), .B1(n14464), .B2(n14116), .C1(
        n14470), .C2(n14626), .ZN(P1_U2858) );
  OR2_X1 U17518 ( .A1(n13972), .A2(n14117), .ZN(n14118) );
  AND2_X1 U17519 ( .A1(n14118), .A2(n14119), .ZN(n14138) );
  INV_X1 U17520 ( .A(n14119), .ZN(n14120) );
  AOI21_X1 U17521 ( .B1(n14138), .B2(n14139), .A(n14120), .ZN(n14182) );
  INV_X1 U17522 ( .A(n14121), .ZN(n14181) );
  NOR2_X1 U17523 ( .A1(n14182), .A2(n14181), .ZN(n14180) );
  OAI21_X1 U17524 ( .B1(n14180), .B2(n14122), .A(n9871), .ZN(n14641) );
  INV_X1 U17525 ( .A(n14793), .ZN(n14124) );
  NOR2_X1 U17526 ( .A1(n14123), .A2(n14124), .ZN(n14127) );
  OAI21_X1 U17527 ( .B1(n14127), .B2(n14126), .A(n14125), .ZN(n14169) );
  INV_X1 U17528 ( .A(n14169), .ZN(n15859) );
  AOI22_X1 U17529 ( .A1(n15859), .A2(n19860), .B1(n19879), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14128) );
  OAI211_X1 U17530 ( .C1(n19855), .C2(n14129), .A(n14128), .B(n19839), .ZN(
        n14135) );
  NAND2_X1 U17531 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14131) );
  INV_X1 U17532 ( .A(n14253), .ZN(n14130) );
  INV_X1 U17533 ( .A(n15701), .ZN(n15718) );
  NOR2_X1 U17534 ( .A1(n14131), .A2(n15718), .ZN(n14133) );
  AOI21_X1 U17535 ( .B1(n15642), .B2(n14131), .A(n15715), .ZN(n15707) );
  INV_X1 U17536 ( .A(n15707), .ZN(n14132) );
  MUX2_X1 U17537 ( .A(n14133), .B(n14132), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14134) );
  AOI211_X1 U17538 ( .C1(n14638), .C2(n19883), .A(n14135), .B(n14134), .ZN(
        n14136) );
  OAI21_X1 U17539 ( .B1(n14641), .B2(n14414), .A(n14136), .ZN(P1_U2827) );
  AOI22_X1 U17540 ( .A1(n14534), .A2(n14476), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14532), .ZN(n14137) );
  OAI21_X1 U17541 ( .B1(n14641), .B2(n14543), .A(n14137), .ZN(P1_U2891) );
  XOR2_X1 U17542 ( .A(n14139), .B(n14138), .Z(n15789) );
  INV_X1 U17543 ( .A(n15789), .ZN(n14141) );
  AOI22_X1 U17544 ( .A1(n14534), .A2(n14484), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14532), .ZN(n14140) );
  OAI21_X1 U17545 ( .B1(n14141), .B2(n14543), .A(n14140), .ZN(P1_U2893) );
  OAI21_X1 U17546 ( .B1(n9641), .B2(n14143), .A(n14142), .ZN(n15680) );
  OAI222_X1 U17547 ( .A1(n15680), .A2(n14543), .B1(n14542), .B2(n14144), .C1(
        n14539), .C2(n20885), .ZN(P1_U2889) );
  NAND2_X1 U17548 ( .A1(n9681), .A2(n14146), .ZN(n14147) );
  XNOR2_X1 U17549 ( .A(n14145), .B(n14147), .ZN(n15883) );
  NAND2_X1 U17550 ( .A1(n15883), .A2(n19948), .ZN(n14150) );
  NAND2_X1 U17551 ( .A1(n19940), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15880) );
  OAI21_X1 U17552 ( .B1(n14636), .B2(n11419), .A(n15880), .ZN(n14148) );
  AOI21_X1 U17553 ( .B1(n15781), .B2(n19819), .A(n14148), .ZN(n14149) );
  OAI211_X1 U17554 ( .C1(n19995), .C2(n19823), .A(n14150), .B(n14149), .ZN(
        P1_U2990) );
  INV_X1 U17555 ( .A(n14151), .ZN(n14167) );
  NOR2_X1 U17556 ( .A1(n18939), .A2(n14152), .ZN(n14153) );
  XNOR2_X1 U17557 ( .A(n14153), .B(n16040), .ZN(n14154) );
  NAND2_X1 U17558 ( .A1(n14154), .A2(n18933), .ZN(n14166) );
  AOI21_X1 U17559 ( .B1(n14157), .B2(n14156), .A(n14155), .ZN(n15320) );
  AOI22_X1 U17560 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18947), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n18927), .ZN(n14158) );
  OAI211_X1 U17561 ( .C1(n14159), .C2(n18921), .A(n18920), .B(n14158), .ZN(
        n14164) );
  OAI21_X1 U17562 ( .B1(n14160), .B2(n14162), .A(n14161), .ZN(n16033) );
  NOR2_X1 U17563 ( .A1(n16033), .A2(n18954), .ZN(n14163) );
  AOI211_X1 U17564 ( .C1(n15320), .C2(n18958), .A(n14164), .B(n14163), .ZN(
        n14165) );
  OAI211_X1 U17565 ( .C1(n18924), .C2(n14167), .A(n14166), .B(n14165), .ZN(
        P2_U2839) );
  INV_X1 U17566 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14168) );
  OAI222_X1 U17567 ( .A1(n14169), .A2(n14472), .B1(n14168), .B2(n19904), .C1(
        n14470), .C2(n14641), .ZN(P1_U2859) );
  AND2_X1 U17568 ( .A1(n14171), .A2(n14170), .ZN(n14172) );
  OR2_X1 U17569 ( .A1(n14160), .A2(n14172), .ZN(n15336) );
  INV_X1 U17570 ( .A(n14218), .ZN(n14176) );
  OAI211_X1 U17571 ( .C1(n14104), .C2(n14177), .A(n14176), .B(n14175), .ZN(
        n14179) );
  NAND2_X1 U17572 ( .A1(n14932), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14178) );
  OAI211_X1 U17573 ( .C1(n15336), .C2(n14932), .A(n14179), .B(n14178), .ZN(
        P2_U2872) );
  AOI21_X1 U17574 ( .B1(n14182), .B2(n14181), .A(n14180), .ZN(n15779) );
  INV_X1 U17575 ( .A(n15779), .ZN(n14185) );
  OAI222_X1 U17576 ( .A1(n14185), .A2(n14543), .B1(n14542), .B2(n14184), .C1(
        n14183), .C2(n14539), .ZN(P1_U2892) );
  XNOR2_X1 U17577 ( .A(n14186), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14206) );
  XOR2_X1 U17578 ( .A(n14187), .B(n14189), .Z(n14204) );
  NAND2_X1 U17579 ( .A1(n14190), .A2(n19055), .ZN(n14194) );
  NAND2_X1 U17580 ( .A1(n15273), .A2(n14191), .ZN(n16196) );
  NAND2_X1 U17581 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19040), .ZN(n14192) );
  OAI221_X1 U17582 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14194), .C1(
        n14193), .C2(n16196), .A(n14192), .ZN(n14197) );
  OAI22_X1 U17583 ( .A1(n14202), .A2(n15384), .B1(n19058), .B2(n14195), .ZN(
        n14196) );
  AOI211_X1 U17584 ( .C1(n14204), .C2(n19064), .A(n14197), .B(n14196), .ZN(
        n14198) );
  OAI21_X1 U17585 ( .B1(n14206), .B2(n16207), .A(n14198), .ZN(P2_U3040) );
  OAI22_X1 U17586 ( .A1(n19666), .A2(n18920), .B1(n19052), .B2(n14199), .ZN(
        n14200) );
  AOI21_X1 U17587 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19041), .A(
        n14200), .ZN(n14201) );
  OAI21_X1 U17588 ( .B1(n14202), .B2(n16034), .A(n14201), .ZN(n14203) );
  AOI21_X1 U17589 ( .B1(n14204), .B2(n19046), .A(n14203), .ZN(n14205) );
  OAI21_X1 U17590 ( .B1(n14206), .B2(n16108), .A(n14205), .ZN(P2_U3008) );
  XOR2_X1 U17591 ( .A(n14207), .B(n14142), .Z(n15767) );
  INV_X1 U17592 ( .A(n15767), .ZN(n14215) );
  OAI21_X1 U17593 ( .B1(n15684), .B2(n14208), .A(n14391), .ZN(n15673) );
  INV_X1 U17594 ( .A(n15673), .ZN(n14778) );
  AOI22_X1 U17595 ( .A1(n14778), .A2(n19899), .B1(n14468), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14209) );
  OAI21_X1 U17596 ( .B1(n14215), .B2(n14470), .A(n14209), .ZN(P1_U2856) );
  AOI22_X1 U17597 ( .A1(n14526), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14532), .ZN(n14214) );
  NOR3_X1 U17598 ( .A1(n14532), .A2(n14210), .A3(n11135), .ZN(n14211) );
  INV_X1 U17599 ( .A(n20005), .ZN(n14212) );
  AOI22_X1 U17600 ( .A1(n14528), .A2(n14212), .B1(n14527), .B2(DATAI_16_), 
        .ZN(n14213) );
  OAI211_X1 U17601 ( .C1(n14215), .C2(n14543), .A(n14214), .B(n14213), .ZN(
        P1_U2888) );
  INV_X1 U17602 ( .A(n14938), .ZN(n14216) );
  OAI21_X1 U17603 ( .B1(n14218), .B2(n14217), .A(n14216), .ZN(n14225) );
  MUX2_X1 U17604 ( .A(n16033), .B(n12350), .S(n14932), .Z(n14219) );
  OAI21_X1 U17605 ( .B1(n14225), .B2(n14942), .A(n14219), .ZN(P2_U2871) );
  OAI22_X1 U17606 ( .A1(n19081), .A2(n16003), .B1(n18973), .B2(n14220), .ZN(
        n14223) );
  AOI22_X1 U17607 ( .A1(n18963), .A2(BUF2_REG_16__SCAN_IN), .B1(n18962), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14221) );
  INV_X1 U17608 ( .A(n14221), .ZN(n14222) );
  AOI211_X1 U17609 ( .C1(n18996), .C2(n15320), .A(n14223), .B(n14222), .ZN(
        n14224) );
  OAI21_X1 U17610 ( .B1(n14225), .B2(n18978), .A(n14224), .ZN(P2_U2903) );
  INV_X2 U17611 ( .A(n18532), .ZN(n18563) );
  OAI21_X1 U17612 ( .B1(n18562), .B2(n18711), .A(n18545), .ZN(n14226) );
  NAND2_X1 U17613 ( .A1(n18563), .A2(n14226), .ZN(n18544) );
  NOR2_X1 U17614 ( .A1(n18708), .A2(n18544), .ZN(n14233) );
  INV_X1 U17615 ( .A(n18759), .ZN(n18750) );
  NOR2_X1 U17616 ( .A1(n18535), .A2(n18750), .ZN(n14230) );
  INV_X1 U17617 ( .A(n14227), .ZN(n14228) );
  NAND2_X1 U17618 ( .A1(n17332), .A2(n10902), .ZN(n18597) );
  INV_X1 U17619 ( .A(n18748), .ZN(n18619) );
  AOI21_X1 U17620 ( .B1(n14230), .B2(n17292), .A(n14229), .ZN(n14231) );
  OAI211_X1 U17621 ( .C1(n15487), .C2(n15488), .A(n14231), .B(n15610), .ZN(
        n18580) );
  INV_X1 U17622 ( .A(n18580), .ZN(n18569) );
  NAND2_X1 U17623 ( .A1(n18753), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18102) );
  INV_X1 U17624 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18096) );
  NAND3_X1 U17625 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n18702)
         );
  OR2_X1 U17626 ( .A1(n18096), .A2(n18702), .ZN(n14232) );
  OAI211_X1 U17627 ( .C1(n18603), .C2(n18569), .A(n18102), .B(n14232), .ZN(
        n18731) );
  INV_X1 U17628 ( .A(n18731), .ZN(n18734) );
  MUX2_X1 U17629 ( .A(n14233), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18734), .Z(P3_U3284) );
  OAI211_X1 U17630 ( .C1(n18711), .C2(n18562), .A(n16957), .B(n18545), .ZN(
        n18095) );
  NOR2_X1 U17631 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18095), .ZN(n14234) );
  INV_X1 U17632 ( .A(n18385), .ZN(n18200) );
  OAI21_X1 U17633 ( .B1(n14234), .B2(n18702), .A(n18200), .ZN(n18101) );
  INV_X1 U17634 ( .A(n18101), .ZN(n14235) );
  INV_X1 U17635 ( .A(n17721), .ZN(n17659) );
  NOR2_X1 U17636 ( .A1(n17659), .A2(n18756), .ZN(n15511) );
  AOI21_X1 U17637 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n15511), .ZN(n15512) );
  NOR2_X1 U17638 ( .A1(n14235), .A2(n15512), .ZN(n14237) );
  NOR2_X1 U17639 ( .A1(n18704), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18138) );
  OR2_X1 U17640 ( .A1(n18138), .A2(n14235), .ZN(n15510) );
  OR2_X1 U17641 ( .A1(n18441), .A2(n15510), .ZN(n14236) );
  MUX2_X1 U17642 ( .A(n14237), .B(n14236), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NAND2_X1 U17643 ( .A1(n14239), .A2(n14238), .ZN(n14242) );
  NOR2_X1 U17644 ( .A1(n14240), .A2(n9646), .ZN(n14241) );
  XOR2_X1 U17645 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14243), .Z(
        n15054) );
  NOR2_X1 U17646 ( .A1(n15204), .A2(n14244), .ZN(n14246) );
  OAI21_X1 U17647 ( .B1(n14246), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14245), .ZN(n14249) );
  AND2_X1 U17648 ( .A1(n19040), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15049) );
  OAI211_X1 U17649 ( .C1(n15052), .C2(n15384), .A(n14249), .B(n14248), .ZN(
        n14250) );
  OAI21_X1 U17650 ( .B1(n15056), .B2(n16191), .A(n14251), .ZN(P2_U3016) );
  NAND2_X1 U17651 ( .A1(n14252), .A2(n19847), .ZN(n14266) );
  AND2_X1 U17652 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14261) );
  INV_X1 U17653 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20741) );
  INV_X1 U17654 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20734) );
  NAND4_X1 U17655 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14375) );
  NAND3_X1 U17656 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14379) );
  NOR3_X1 U17657 ( .A1(n20734), .A2(n14375), .A3(n14379), .ZN(n15660) );
  NAND4_X1 U17658 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n14254), .A3(n14253), 
        .A4(n15660), .ZN(n14368) );
  NAND3_X1 U17659 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14369) );
  NOR3_X1 U17660 ( .A1(n20741), .A2(n14368), .A3(n14369), .ZN(n14353) );
  NAND2_X1 U17661 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14353), .ZN(n15616) );
  NAND2_X1 U17662 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14255) );
  NOR2_X1 U17663 ( .A1(n15616), .A2(n14255), .ZN(n14323) );
  AND2_X1 U17664 ( .A1(n14323), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14256) );
  NAND2_X1 U17665 ( .A1(n14417), .A2(n14256), .ZN(n14314) );
  INV_X1 U17666 ( .A(n14314), .ZN(n14257) );
  NAND2_X1 U17667 ( .A1(n14257), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14259) );
  NAND2_X1 U17668 ( .A1(n14376), .A2(n14259), .ZN(n14313) );
  OAI21_X1 U17669 ( .B1(n19838), .B2(n14261), .A(n14313), .ZN(n14288) );
  INV_X1 U17670 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14428) );
  OAI22_X1 U17671 ( .A1(n19833), .A2(n14428), .B1(n14258), .B2(n19855), .ZN(
        n14264) );
  INV_X1 U17672 ( .A(n14259), .ZN(n14260) );
  NAND2_X1 U17673 ( .A1(n15642), .A2(n14260), .ZN(n14300) );
  INV_X1 U17674 ( .A(n14261), .ZN(n14262) );
  NOR3_X1 U17675 ( .A1(n14300), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14262), 
        .ZN(n14263) );
  AOI211_X1 U17676 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14288), .A(n14264), 
        .B(n14263), .ZN(n14265) );
  OAI211_X1 U17677 ( .C1(n14429), .C2(n19893), .A(n14266), .B(n14265), .ZN(
        P1_U2809) );
  NOR2_X1 U17678 ( .A1(n14267), .A2(n19052), .ZN(n14270) );
  AOI21_X1 U17679 ( .B1(n19041), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14268), .ZN(n14269) );
  OAI21_X1 U17680 ( .B1(n14273), .B2(n16109), .A(n14272), .ZN(P2_U2983) );
  INV_X1 U17681 ( .A(n14274), .ZN(n14283) );
  NAND2_X1 U17682 ( .A1(n14275), .A2(n18888), .ZN(n14282) );
  AOI22_X1 U17683 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n9691), .ZN(n14276) );
  OAI21_X1 U17684 ( .B1(n14278), .B2(n14277), .A(n14276), .ZN(n14280) );
  NOR2_X1 U17685 ( .A1(n14865), .A2(n18954), .ZN(n14279) );
  OAI211_X1 U17686 ( .C1(n18924), .C2(n14283), .A(n14282), .B(n14281), .ZN(
        P2_U2824) );
  NOR2_X1 U17687 ( .A1(n15052), .A2(n13608), .ZN(n14284) );
  AOI21_X1 U17688 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n13608), .A(n14284), .ZN(
        n14285) );
  OAI21_X1 U17689 ( .B1(n14286), .B2(n14942), .A(n14285), .ZN(P2_U2857) );
  NOR2_X1 U17690 ( .A1(n14300), .A2(n20753), .ZN(n14289) );
  OAI21_X1 U17691 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14289), .A(n14288), 
        .ZN(n14291) );
  AOI22_X1 U17692 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19884), .B1(
        n19883), .B2(n14547), .ZN(n14290) );
  OAI211_X1 U17693 ( .C1(n19833), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        n14293) );
  AOI21_X1 U17694 ( .B1(n14661), .B2(n19860), .A(n14293), .ZN(n14294) );
  OAI21_X1 U17695 ( .B1(n14553), .B2(n14414), .A(n14294), .ZN(P1_U2810) );
  INV_X1 U17696 ( .A(n14295), .ZN(n14479) );
  INV_X1 U17697 ( .A(n14313), .ZN(n14305) );
  OAI22_X1 U17698 ( .A1(n14297), .A2(n19855), .B1(n15712), .B2(n14296), .ZN(
        n14298) );
  AOI21_X1 U17699 ( .B1(n19879), .B2(P1_EBX_REG_29__SCAN_IN), .A(n14298), .ZN(
        n14299) );
  OAI21_X1 U17700 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14300), .A(n14299), 
        .ZN(n14304) );
  OAI21_X1 U17701 ( .B1(n14309), .B2(n14302), .A(n14301), .ZN(n14666) );
  NOR2_X1 U17702 ( .A1(n14666), .A2(n19893), .ZN(n14303) );
  AOI211_X1 U17703 ( .C1(n14305), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14304), 
        .B(n14303), .ZN(n14306) );
  OAI21_X1 U17704 ( .B1(n14479), .B2(n14414), .A(n14306), .ZN(P1_U2811) );
  NOR2_X1 U17705 ( .A1(n14328), .A2(n14307), .ZN(n14308) );
  OR2_X1 U17706 ( .A1(n14309), .A2(n14308), .ZN(n14683) );
  AOI21_X1 U17707 ( .B1(n14311), .B2(n14321), .A(n12778), .ZN(n14570) );
  NAND2_X1 U17708 ( .A1(n14570), .A2(n19847), .ZN(n14319) );
  INV_X1 U17709 ( .A(n14566), .ZN(n14312) );
  OAI22_X1 U17710 ( .A1(n14568), .A2(n19855), .B1(n15712), .B2(n14312), .ZN(
        n14317) );
  INV_X1 U17711 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14315) );
  AOI21_X1 U17712 ( .B1(n14315), .B2(n14314), .A(n14313), .ZN(n14316) );
  AOI211_X1 U17713 ( .C1(n19879), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14317), .B(
        n14316), .ZN(n14318) );
  OAI211_X1 U17714 ( .C1(n19893), .C2(n14683), .A(n14319), .B(n14318), .ZN(
        P1_U2812) );
  AOI21_X1 U17715 ( .B1(n14323), .B2(n14417), .A(n19838), .ZN(n14338) );
  INV_X1 U17716 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14432) );
  INV_X1 U17717 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20750) );
  NAND3_X1 U17718 ( .A1(n15642), .A2(n14323), .A3(n20750), .ZN(n14325) );
  AOI22_X1 U17719 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19884), .B1(
        n19883), .B2(n14580), .ZN(n14324) );
  OAI211_X1 U17720 ( .C1(n14432), .C2(n19833), .A(n14325), .B(n14324), .ZN(
        n14330) );
  NOR2_X1 U17721 ( .A1(n14336), .A2(n14326), .ZN(n14327) );
  OR2_X1 U17722 ( .A1(n14328), .A2(n14327), .ZN(n14691) );
  NOR2_X1 U17723 ( .A1(n14691), .A2(n19893), .ZN(n14329) );
  AOI211_X1 U17724 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14338), .A(n14330), 
        .B(n14329), .ZN(n14331) );
  OAI21_X1 U17725 ( .B1(n14577), .B2(n14414), .A(n14331), .ZN(P1_U2813) );
  INV_X1 U17726 ( .A(n14332), .ZN(n14333) );
  AOI21_X1 U17727 ( .B1(n14334), .B2(n14333), .A(n14320), .ZN(n14583) );
  INV_X1 U17728 ( .A(n14583), .ZN(n14490) );
  AND2_X1 U17729 ( .A1(n15625), .A2(n14335), .ZN(n14337) );
  OR2_X1 U17730 ( .A1(n14337), .A2(n14336), .ZN(n14701) );
  INV_X1 U17731 ( .A(n14701), .ZN(n14344) );
  INV_X1 U17732 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14342) );
  INV_X1 U17733 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20745) );
  NOR3_X1 U17734 ( .A1(n19877), .A2(n15616), .A3(n20745), .ZN(n14339) );
  OAI21_X1 U17735 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n14339), .A(n14338), 
        .ZN(n14341) );
  AOI22_X1 U17736 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19884), .B1(
        n19883), .B2(n14586), .ZN(n14340) );
  OAI211_X1 U17737 ( .C1(n19833), .C2(n14342), .A(n14341), .B(n14340), .ZN(
        n14343) );
  AOI21_X1 U17738 ( .B1(n14344), .B2(n19860), .A(n14343), .ZN(n14345) );
  OAI21_X1 U17739 ( .B1(n14490), .B2(n14414), .A(n14345), .ZN(P1_U2814) );
  OAI21_X1 U17740 ( .B1(n14362), .B2(n14346), .A(n15623), .ZN(n14711) );
  OR2_X1 U17741 ( .A1(n14348), .A2(n14349), .ZN(n14350) );
  AND2_X1 U17742 ( .A1(n14347), .A2(n14350), .ZN(n14597) );
  NAND2_X1 U17743 ( .A1(n14597), .A2(n19847), .ZN(n14357) );
  OAI21_X1 U17744 ( .B1(n14353), .B2(n19877), .A(n14417), .ZN(n15615) );
  AOI22_X1 U17745 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19884), .B1(
        n19883), .B2(n14594), .ZN(n14351) );
  OAI21_X1 U17746 ( .B1(n19833), .B2(n14352), .A(n14351), .ZN(n14355) );
  INV_X1 U17747 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20743) );
  AND3_X1 U17748 ( .A1(n20743), .A2(n15642), .A3(n14353), .ZN(n14354) );
  AOI211_X1 U17749 ( .C1(n15615), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14355), 
        .B(n14354), .ZN(n14356) );
  OAI211_X1 U17750 ( .C1(n19893), .C2(n14711), .A(n14357), .B(n14356), .ZN(
        P1_U2816) );
  AND2_X1 U17751 ( .A1(n14358), .A2(n14359), .ZN(n14360) );
  NOR2_X1 U17752 ( .A1(n14348), .A2(n14360), .ZN(n15741) );
  INV_X1 U17753 ( .A(n15741), .ZN(n14503) );
  AND2_X1 U17754 ( .A1(n14440), .A2(n14361), .ZN(n14363) );
  OR2_X1 U17755 ( .A1(n14363), .A2(n14362), .ZN(n15822) );
  INV_X1 U17756 ( .A(n15822), .ZN(n14367) );
  INV_X1 U17757 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14435) );
  INV_X1 U17758 ( .A(n15744), .ZN(n14364) );
  AOI22_X1 U17759 ( .A1(n14364), .A2(n19883), .B1(n19884), .B2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14365) );
  OAI21_X1 U17760 ( .B1(n19833), .B2(n14435), .A(n14365), .ZN(n14366) );
  AOI21_X1 U17761 ( .B1(n14367), .B2(n19860), .A(n14366), .ZN(n14372) );
  INV_X1 U17762 ( .A(n14368), .ZN(n15635) );
  NAND2_X1 U17763 ( .A1(n15642), .A2(n15635), .ZN(n15653) );
  OAI21_X1 U17764 ( .B1(n14369), .B2(n15653), .A(n20741), .ZN(n14370) );
  NAND2_X1 U17765 ( .A1(n15615), .A2(n14370), .ZN(n14371) );
  OAI211_X1 U17766 ( .C1(n14503), .C2(n14414), .A(n14372), .B(n14371), .ZN(
        P1_U2817) );
  XOR2_X1 U17767 ( .A(n14374), .B(n14373), .Z(n14615) );
  INV_X1 U17768 ( .A(n14615), .ZN(n14525) );
  INV_X1 U17769 ( .A(n14379), .ZN(n14377) );
  AOI21_X1 U17770 ( .B1(n14376), .B2(n14375), .A(n15715), .ZN(n15700) );
  OAI21_X1 U17771 ( .B1(n14377), .B2(n19877), .A(n15700), .ZN(n15667) );
  NAND3_X1 U17772 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14378) );
  NOR2_X1 U17773 ( .A1(n14378), .A2(n15718), .ZN(n15691) );
  NAND2_X1 U17774 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15691), .ZN(n15675) );
  NOR3_X1 U17775 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14379), .A3(n15675), 
        .ZN(n15668) );
  AND2_X1 U17776 ( .A1(n9643), .A2(n14380), .ZN(n14381) );
  OR2_X1 U17777 ( .A1(n14381), .A2(n14459), .ZN(n15827) );
  AOI21_X1 U17778 ( .B1(n19884), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19868), .ZN(n14383) );
  AOI22_X1 U17779 ( .A1(n14611), .A2(n19883), .B1(n19879), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n14382) );
  OAI211_X1 U17780 ( .C1(n19893), .C2(n15827), .A(n14383), .B(n14382), .ZN(
        n14384) );
  AOI211_X1 U17781 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15667), .A(n15668), 
        .B(n14384), .ZN(n14385) );
  OAI21_X1 U17782 ( .B1(n14525), .B2(n14414), .A(n14385), .ZN(P1_U2822) );
  INV_X1 U17783 ( .A(n14386), .ZN(n14388) );
  INV_X1 U17784 ( .A(n14373), .ZN(n14387) );
  AOI21_X1 U17785 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(n15761) );
  INV_X1 U17786 ( .A(n15761), .ZN(n14531) );
  NAND2_X1 U17787 ( .A1(n14391), .A2(n14390), .ZN(n14392) );
  AND2_X1 U17788 ( .A1(n9643), .A2(n14392), .ZN(n14756) );
  INV_X1 U17789 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14395) );
  NAND2_X1 U17790 ( .A1(n15760), .A2(n19883), .ZN(n14394) );
  AOI21_X1 U17791 ( .B1(n19884), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n19868), .ZN(n14393) );
  OAI211_X1 U17792 ( .C1(n14395), .C2(n19833), .A(n14394), .B(n14393), .ZN(
        n14396) );
  AOI21_X1 U17793 ( .B1(n14756), .B2(n19860), .A(n14396), .ZN(n14400) );
  NAND2_X1 U17794 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14397) );
  INV_X1 U17795 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20732) );
  OAI21_X1 U17796 ( .B1(n14397), .B2(n15675), .A(n20732), .ZN(n14398) );
  NAND2_X1 U17797 ( .A1(n15667), .A2(n14398), .ZN(n14399) );
  OAI211_X1 U17798 ( .C1(n14531), .C2(n14414), .A(n14400), .B(n14399), .ZN(
        P1_U2823) );
  OR2_X1 U17799 ( .A1(n14401), .A2(n14402), .ZN(n14538) );
  AOI21_X1 U17800 ( .B1(n14403), .B2(n14538), .A(n13861), .ZN(n14657) );
  INV_X1 U17801 ( .A(n14657), .ZN(n14536) );
  OAI21_X1 U17802 ( .B1(n19838), .B2(n19821), .A(n19871), .ZN(n19824) );
  NAND2_X1 U17803 ( .A1(n15906), .A2(n14404), .ZN(n14405) );
  NAND2_X1 U17804 ( .A1(n14406), .A2(n14405), .ZN(n15898) );
  INV_X1 U17805 ( .A(n14655), .ZN(n14407) );
  AOI22_X1 U17806 ( .A1(n19879), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n14407), .B2(
        n19883), .ZN(n14411) );
  NOR3_X1 U17807 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14408), .A3(n19857), .ZN(
        n14409) );
  AOI211_X1 U17808 ( .C1(n19884), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19868), .B(n14409), .ZN(n14410) );
  OAI211_X1 U17809 ( .C1(n19893), .C2(n15898), .A(n14411), .B(n14410), .ZN(
        n14412) );
  AOI21_X1 U17810 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n19824), .A(n14412), .ZN(
        n14413) );
  OAI21_X1 U17811 ( .B1(n14536), .B2(n14414), .A(n14413), .ZN(P1_U2832) );
  INV_X1 U17812 ( .A(n14415), .ZN(n14416) );
  NAND2_X1 U17813 ( .A1(n14416), .A2(n19889), .ZN(n14427) );
  NOR2_X1 U17814 ( .A1(n19877), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19881) );
  INV_X1 U17815 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14421) );
  INV_X1 U17816 ( .A(n14417), .ZN(n19880) );
  AOI22_X1 U17817 ( .A1(n19883), .A2(n14418), .B1(n19880), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14420) );
  NAND2_X1 U17818 ( .A1(n19884), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14419) );
  OAI211_X1 U17819 ( .C1(n19833), .C2(n14421), .A(n14420), .B(n14419), .ZN(
        n14422) );
  NOR2_X1 U17820 ( .A1(n19881), .A2(n14422), .ZN(n14426) );
  OR2_X1 U17821 ( .A1(n20315), .A2(n19887), .ZN(n14425) );
  NAND2_X1 U17822 ( .A1(n19860), .A2(n14804), .ZN(n14424) );
  NAND4_X1 U17823 ( .A1(n14427), .A2(n14426), .A3(n14425), .A4(n14424), .ZN(
        P1_U2839) );
  OAI22_X1 U17824 ( .A1(n14429), .A2(n14472), .B1(n14428), .B2(n14464), .ZN(
        P1_U2841) );
  OAI222_X1 U17825 ( .A1(n14430), .A2(n19904), .B1(n14472), .B2(n14666), .C1(
        n14479), .C2(n14470), .ZN(P1_U2843) );
  INV_X1 U17826 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14431) );
  INV_X1 U17827 ( .A(n14570), .ZN(n14483) );
  OAI222_X1 U17828 ( .A1(n14431), .A2(n19904), .B1(n14472), .B2(n14683), .C1(
        n14483), .C2(n14470), .ZN(P1_U2844) );
  OAI222_X1 U17829 ( .A1(n14432), .A2(n19904), .B1(n14472), .B2(n14691), .C1(
        n14577), .C2(n14470), .ZN(P1_U2845) );
  OAI222_X1 U17830 ( .A1(n14470), .A2(n14490), .B1(n14464), .B2(n14342), .C1(
        n14701), .C2(n14472), .ZN(P1_U2846) );
  INV_X1 U17831 ( .A(n14597), .ZN(n14500) );
  INV_X1 U17832 ( .A(n14711), .ZN(n14433) );
  AOI22_X1 U17833 ( .A1(n14433), .A2(n19899), .B1(n14468), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14434) );
  OAI21_X1 U17834 ( .B1(n14500), .B2(n14470), .A(n14434), .ZN(P1_U2848) );
  OAI222_X1 U17835 ( .A1(n14435), .A2(n19904), .B1(n14470), .B2(n14503), .C1(
        n14472), .C2(n15822), .ZN(P1_U2849) );
  INV_X1 U17836 ( .A(n14358), .ZN(n14436) );
  AOI21_X1 U17837 ( .B1(n14437), .B2(n9639), .A(n14436), .ZN(n15637) );
  NAND2_X1 U17838 ( .A1(n14449), .A2(n14438), .ZN(n14439) );
  NAND2_X1 U17839 ( .A1(n14440), .A2(n14439), .ZN(n15640) );
  OAI22_X1 U17840 ( .A1(n15640), .A2(n14472), .B1(n15631), .B2(n14464), .ZN(
        n14441) );
  AOI21_X1 U17841 ( .B1(n15637), .B2(n19900), .A(n14441), .ZN(n14442) );
  INV_X1 U17842 ( .A(n14442), .ZN(P1_U2850) );
  NAND2_X1 U17843 ( .A1(n14443), .A2(n14444), .ZN(n14445) );
  AND2_X1 U17844 ( .A1(n9639), .A2(n14445), .ZN(n15745) );
  INV_X1 U17845 ( .A(n15745), .ZN(n14510) );
  NAND2_X1 U17846 ( .A1(n14446), .A2(n14447), .ZN(n14448) );
  AND2_X1 U17847 ( .A1(n14449), .A2(n14448), .ZN(n15649) );
  AOI22_X1 U17848 ( .A1(n15649), .A2(n19899), .B1(n14468), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n14450) );
  OAI21_X1 U17849 ( .B1(n14510), .B2(n14470), .A(n14450), .ZN(P1_U2851) );
  OR2_X1 U17850 ( .A1(n14461), .A2(n14451), .ZN(n14452) );
  NAND2_X1 U17851 ( .A1(n14446), .A2(n14452), .ZN(n15659) );
  INV_X1 U17852 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15655) );
  XOR2_X1 U17853 ( .A(n14454), .B(n14453), .Z(n15751) );
  INV_X1 U17854 ( .A(n15751), .ZN(n14515) );
  OAI222_X1 U17855 ( .A1(n15659), .A2(n14472), .B1(n15655), .B2(n19904), .C1(
        n14515), .C2(n14470), .ZN(P1_U2852) );
  NOR2_X1 U17856 ( .A1(n14455), .A2(n14456), .ZN(n14457) );
  NOR2_X1 U17857 ( .A1(n14457), .A2(n14453), .ZN(n15755) );
  NOR2_X1 U17858 ( .A1(n14459), .A2(n14458), .ZN(n14460) );
  OR2_X1 U17859 ( .A1(n14461), .A2(n14460), .ZN(n15671) );
  INV_X1 U17860 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n20829) );
  OAI22_X1 U17861 ( .A1(n15671), .A2(n14472), .B1(n20829), .B2(n14464), .ZN(
        n14462) );
  AOI21_X1 U17862 ( .B1(n15755), .B2(n19900), .A(n14462), .ZN(n14463) );
  INV_X1 U17863 ( .A(n14463), .ZN(P1_U2853) );
  OAI22_X1 U17864 ( .A1(n15827), .A2(n14472), .B1(n14465), .B2(n14464), .ZN(
        n14466) );
  AOI21_X1 U17865 ( .B1(n14615), .B2(n19900), .A(n14466), .ZN(n14467) );
  INV_X1 U17866 ( .A(n14467), .ZN(P1_U2854) );
  AOI22_X1 U17867 ( .A1(n14756), .A2(n19899), .B1(n14468), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14469) );
  OAI21_X1 U17868 ( .B1(n14531), .B2(n14470), .A(n14469), .ZN(P1_U2855) );
  INV_X1 U17869 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14471) );
  OAI222_X1 U17870 ( .A1(n15898), .A2(n14472), .B1(n19904), .B2(n14471), .C1(
        n14470), .C2(n14536), .ZN(P1_U2864) );
  AOI22_X1 U17871 ( .A1(n14526), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14532), .ZN(n14475) );
  AOI22_X1 U17872 ( .A1(n14528), .A2(n14473), .B1(n14527), .B2(DATAI_30_), 
        .ZN(n14474) );
  OAI211_X1 U17873 ( .C1(n14553), .C2(n14543), .A(n14475), .B(n14474), .ZN(
        P1_U2874) );
  AOI22_X1 U17874 ( .A1(n14526), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14532), .ZN(n14478) );
  AOI22_X1 U17875 ( .A1(n14528), .A2(n14476), .B1(n14527), .B2(DATAI_29_), 
        .ZN(n14477) );
  OAI211_X1 U17876 ( .C1(n14479), .C2(n14543), .A(n14478), .B(n14477), .ZN(
        P1_U2875) );
  AOI22_X1 U17877 ( .A1(n14526), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14532), .ZN(n14482) );
  AOI22_X1 U17878 ( .A1(n14528), .A2(n14480), .B1(n14527), .B2(DATAI_28_), 
        .ZN(n14481) );
  OAI211_X1 U17879 ( .C1(n14483), .C2(n14543), .A(n14482), .B(n14481), .ZN(
        P1_U2876) );
  AOI22_X1 U17880 ( .A1(n14526), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14532), .ZN(n14486) );
  AOI22_X1 U17881 ( .A1(n14528), .A2(n14484), .B1(n14527), .B2(DATAI_27_), 
        .ZN(n14485) );
  OAI211_X1 U17882 ( .C1(n14577), .C2(n14543), .A(n14486), .B(n14485), .ZN(
        P1_U2877) );
  AOI22_X1 U17883 ( .A1(n14526), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14532), .ZN(n14489) );
  AOI22_X1 U17884 ( .A1(n14528), .A2(n14487), .B1(n14527), .B2(DATAI_26_), 
        .ZN(n14488) );
  OAI211_X1 U17885 ( .C1(n14490), .C2(n14543), .A(n14489), .B(n14488), .ZN(
        P1_U2878) );
  AOI21_X1 U17886 ( .B1(n14491), .B2(n14347), .A(n14332), .ZN(n15732) );
  INV_X1 U17887 ( .A(n15732), .ZN(n14497) );
  INV_X1 U17888 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16349) );
  OAI22_X1 U17889 ( .A1(n14518), .A2(n16349), .B1(n14492), .B2(n14539), .ZN(
        n14493) );
  INV_X1 U17890 ( .A(n14493), .ZN(n14496) );
  AOI22_X1 U17891 ( .A1(n14528), .A2(n14494), .B1(n14527), .B2(DATAI_25_), 
        .ZN(n14495) );
  OAI211_X1 U17892 ( .C1(n14497), .C2(n14543), .A(n14496), .B(n14495), .ZN(
        P1_U2879) );
  AOI22_X1 U17893 ( .A1(n14526), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14532), .ZN(n14499) );
  AOI22_X1 U17894 ( .A1(n14528), .A2(n14533), .B1(n14527), .B2(DATAI_24_), 
        .ZN(n14498) );
  OAI211_X1 U17895 ( .C1(n14500), .C2(n14543), .A(n14499), .B(n14498), .ZN(
        P1_U2880) );
  AOI22_X1 U17896 ( .A1(n14526), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14532), .ZN(n14502) );
  AOI22_X1 U17897 ( .A1(n14528), .A2(n20042), .B1(n14527), .B2(DATAI_23_), 
        .ZN(n14501) );
  OAI211_X1 U17898 ( .C1(n14503), .C2(n14543), .A(n14502), .B(n14501), .ZN(
        P1_U2881) );
  INV_X1 U17899 ( .A(n15637), .ZN(n14506) );
  AOI22_X1 U17900 ( .A1(n14526), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14532), .ZN(n14505) );
  AOI22_X1 U17901 ( .A1(n14528), .A2(n20033), .B1(n14527), .B2(DATAI_22_), 
        .ZN(n14504) );
  OAI211_X1 U17902 ( .C1(n14506), .C2(n14543), .A(n14505), .B(n14504), .ZN(
        P1_U2882) );
  AOI22_X1 U17903 ( .A1(n14526), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14532), .ZN(n14509) );
  INV_X1 U17904 ( .A(n20029), .ZN(n14507) );
  AOI22_X1 U17905 ( .A1(n14528), .A2(n14507), .B1(n14527), .B2(DATAI_21_), 
        .ZN(n14508) );
  OAI211_X1 U17906 ( .C1(n14510), .C2(n14543), .A(n14509), .B(n14508), .ZN(
        P1_U2883) );
  INV_X1 U17907 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19101) );
  OAI22_X1 U17908 ( .A1(n14518), .A2(n19101), .B1(n13648), .B2(n14539), .ZN(
        n14513) );
  INV_X1 U17909 ( .A(n14528), .ZN(n14511) );
  NOR2_X1 U17910 ( .A1(n14511), .A2(n20025), .ZN(n14512) );
  AOI211_X1 U17911 ( .C1(n14527), .C2(DATAI_20_), .A(n14513), .B(n14512), .ZN(
        n14514) );
  OAI21_X1 U17912 ( .B1(n14515), .B2(n14543), .A(n14514), .ZN(P1_U2884) );
  INV_X1 U17913 ( .A(n15755), .ZN(n14522) );
  INV_X1 U17914 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14517) );
  OAI22_X1 U17915 ( .A1(n14518), .A2(n14517), .B1(n14516), .B2(n14539), .ZN(
        n14519) );
  INV_X1 U17916 ( .A(n14519), .ZN(n14521) );
  AOI22_X1 U17917 ( .A1(n14528), .A2(n20021), .B1(n14527), .B2(DATAI_19_), 
        .ZN(n14520) );
  OAI211_X1 U17918 ( .C1(n14522), .C2(n14543), .A(n14521), .B(n14520), .ZN(
        P1_U2885) );
  AOI22_X1 U17919 ( .A1(n14526), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14532), .ZN(n14524) );
  AOI22_X1 U17920 ( .A1(n14528), .A2(n20017), .B1(n14527), .B2(DATAI_18_), 
        .ZN(n14523) );
  OAI211_X1 U17921 ( .C1(n14525), .C2(n14543), .A(n14524), .B(n14523), .ZN(
        P1_U2886) );
  AOI22_X1 U17922 ( .A1(n14526), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14532), .ZN(n14530) );
  AOI22_X1 U17923 ( .A1(n14528), .A2(n20013), .B1(n14527), .B2(DATAI_17_), 
        .ZN(n14529) );
  OAI211_X1 U17924 ( .C1(n14531), .C2(n14543), .A(n14530), .B(n14529), .ZN(
        P1_U2887) );
  AOI22_X1 U17925 ( .A1(n14534), .A2(n14533), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14532), .ZN(n14535) );
  OAI21_X1 U17926 ( .B1(n14536), .B2(n14543), .A(n14535), .ZN(P1_U2896) );
  NAND2_X1 U17927 ( .A1(n14401), .A2(n14402), .ZN(n14537) );
  AND2_X1 U17928 ( .A1(n14538), .A2(n14537), .ZN(n19895) );
  INV_X1 U17929 ( .A(n19895), .ZN(n14544) );
  OAI222_X1 U17930 ( .A1(n14544), .A2(n14543), .B1(n14542), .B2(n14541), .C1(
        n14540), .C2(n14539), .ZN(P1_U2897) );
  INV_X1 U17931 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20757) );
  NOR2_X1 U17932 ( .A1(n19957), .A2(n20757), .ZN(n14660) );
  NOR2_X1 U17933 ( .A1(n14636), .A2(n14545), .ZN(n14546) );
  AOI211_X1 U17934 ( .C1(n15781), .C2(n14547), .A(n14660), .B(n14546), .ZN(
        n14552) );
  NAND2_X1 U17935 ( .A1(n14659), .A2(n19948), .ZN(n14551) );
  OAI211_X1 U17936 ( .C1(n14553), .C2(n19995), .A(n14552), .B(n14551), .ZN(
        P1_U2969) );
  NAND2_X1 U17937 ( .A1(n14591), .A2(n14556), .ZN(n14573) );
  NAND2_X1 U17938 ( .A1(n15740), .A2(n14573), .ZN(n14562) );
  NOR2_X1 U17939 ( .A1(n14557), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14558) );
  NAND2_X1 U17940 ( .A1(n15772), .A2(n14696), .ZN(n14559) );
  NAND2_X1 U17941 ( .A1(n14574), .A2(n14563), .ZN(n14565) );
  XNOR2_X1 U17942 ( .A(n14565), .B(n14564), .ZN(n14686) );
  NAND2_X1 U17943 ( .A1(n15781), .A2(n14566), .ZN(n14567) );
  NAND2_X1 U17944 ( .A1(n19940), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14682) );
  OAI211_X1 U17945 ( .C1(n14636), .C2(n14568), .A(n14567), .B(n14682), .ZN(
        n14569) );
  AOI21_X1 U17946 ( .B1(n14570), .B2(n19947), .A(n14569), .ZN(n14571) );
  OAI21_X1 U17947 ( .B1(n19803), .B2(n14686), .A(n14571), .ZN(P1_U2971) );
  AOI21_X1 U17948 ( .B1(n15772), .B2(n14573), .A(n14572), .ZN(n14582) );
  NAND2_X1 U17949 ( .A1(n14582), .A2(n14574), .ZN(n14575) );
  XNOR2_X1 U17950 ( .A(n14575), .B(n14687), .ZN(n14695) );
  NAND2_X1 U17951 ( .A1(n19940), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14690) );
  OAI21_X1 U17952 ( .B1(n14636), .B2(n14576), .A(n14690), .ZN(n14579) );
  NOR2_X1 U17953 ( .A1(n14577), .A2(n19995), .ZN(n14578) );
  OAI21_X1 U17954 ( .B1(n19803), .B2(n14695), .A(n14581), .ZN(P1_U2972) );
  XNOR2_X1 U17955 ( .A(n14582), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14704) );
  NAND2_X1 U17956 ( .A1(n14583), .A2(n19947), .ZN(n14588) );
  INV_X1 U17957 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20747) );
  NOR2_X1 U17958 ( .A1(n19957), .A2(n20747), .ZN(n14698) );
  INV_X1 U17959 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14584) );
  NOR2_X1 U17960 ( .A1(n14636), .A2(n14584), .ZN(n14585) );
  AOI211_X1 U17961 ( .C1(n15781), .C2(n14586), .A(n14698), .B(n14585), .ZN(
        n14587) );
  OAI211_X1 U17962 ( .C1(n14704), .C2(n19803), .A(n14588), .B(n14587), .ZN(
        P1_U2973) );
  INV_X1 U17963 ( .A(n14589), .ZN(n14590) );
  NOR2_X1 U17964 ( .A1(n14590), .A2(n15739), .ZN(n15730) );
  NOR2_X1 U17965 ( .A1(n15730), .A2(n14591), .ZN(n14592) );
  MUX2_X1 U17966 ( .A(n15730), .B(n14592), .S(n9588), .Z(n14593) );
  XNOR2_X1 U17967 ( .A(n14593), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14716) );
  NAND2_X1 U17968 ( .A1(n15781), .A2(n14594), .ZN(n14595) );
  NAND2_X1 U17969 ( .A1(n19940), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14710) );
  OAI211_X1 U17970 ( .C1(n14636), .C2(n11668), .A(n14595), .B(n14710), .ZN(
        n14596) );
  AOI21_X1 U17971 ( .B1(n14597), .B2(n19947), .A(n14596), .ZN(n14598) );
  OAI21_X1 U17972 ( .B1(n14716), .B2(n19803), .A(n14598), .ZN(P1_U2975) );
  NAND2_X1 U17973 ( .A1(n14601), .A2(n14600), .ZN(n14603) );
  XNOR2_X1 U17974 ( .A(n14603), .B(n14602), .ZN(n14722) );
  INV_X1 U17975 ( .A(n15634), .ZN(n14605) );
  NAND2_X1 U17976 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14604) );
  NAND2_X1 U17977 ( .A1(n19940), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14718) );
  OAI211_X1 U17978 ( .C1(n19953), .C2(n14605), .A(n14604), .B(n14718), .ZN(
        n14606) );
  AOI21_X1 U17979 ( .B1(n15637), .B2(n19947), .A(n14606), .ZN(n14607) );
  OAI21_X1 U17980 ( .B1(n19803), .B2(n14722), .A(n14607), .ZN(P1_U2977) );
  OAI21_X1 U17981 ( .B1(n14610), .B2(n14609), .A(n14741), .ZN(n15828) );
  INV_X1 U17982 ( .A(n14611), .ZN(n14613) );
  AOI22_X1 U17983 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14612) );
  OAI21_X1 U17984 ( .B1(n14613), .B2(n19953), .A(n14612), .ZN(n14614) );
  AOI21_X1 U17985 ( .B1(n14615), .B2(n19947), .A(n14614), .ZN(n14616) );
  OAI21_X1 U17986 ( .B1(n15828), .B2(n19803), .A(n14616), .ZN(P1_U2981) );
  AOI22_X1 U17987 ( .A1(n15785), .A2(n15852), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15772), .ZN(n14625) );
  INV_X1 U17988 ( .A(n14618), .ZN(n14619) );
  NAND2_X1 U17989 ( .A1(n15785), .A2(n14619), .ZN(n14620) );
  INV_X1 U17990 ( .A(n14621), .ZN(n14623) );
  OAI21_X1 U17991 ( .B1(n14765), .B2(n14623), .A(n14622), .ZN(n14624) );
  XOR2_X1 U17992 ( .A(n14625), .B(n14624), .Z(n15844) );
  INV_X1 U17993 ( .A(n14626), .ZN(n15696) );
  AOI22_X1 U17994 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14627) );
  OAI21_X1 U17995 ( .B1(n19953), .B2(n15692), .A(n14627), .ZN(n14628) );
  AOI21_X1 U17996 ( .B1(n15696), .B2(n19947), .A(n14628), .ZN(n14629) );
  OAI21_X1 U17997 ( .B1(n15844), .B2(n19803), .A(n14629), .ZN(P1_U2985) );
  OAI22_X1 U17998 ( .A1(n14617), .A2(n14631), .B1(n14630), .B2(n15772), .ZN(
        n14782) );
  INV_X1 U17999 ( .A(n14633), .ZN(n14632) );
  OAI21_X1 U18000 ( .B1(n14791), .B2(n15772), .A(n14632), .ZN(n14781) );
  NOR2_X1 U18001 ( .A1(n14782), .A2(n14781), .ZN(n14780) );
  NOR2_X1 U18002 ( .A1(n14780), .A2(n14633), .ZN(n14635) );
  XNOR2_X1 U18003 ( .A(n14635), .B(n14634), .ZN(n15861) );
  NAND2_X1 U18004 ( .A1(n15861), .A2(n19948), .ZN(n14640) );
  NAND2_X1 U18005 ( .A1(n19940), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15857) );
  OAI21_X1 U18006 ( .B1(n14636), .B2(n14129), .A(n15857), .ZN(n14637) );
  AOI21_X1 U18007 ( .B1(n15781), .B2(n14638), .A(n14637), .ZN(n14639) );
  OAI211_X1 U18008 ( .C1(n19995), .C2(n14641), .A(n14640), .B(n14639), .ZN(
        P1_U2986) );
  AND2_X1 U18009 ( .A1(n14642), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14644) );
  XNOR2_X1 U18010 ( .A(n14617), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14643) );
  MUX2_X1 U18011 ( .A(n14644), .B(n14643), .S(n15772), .Z(n14645) );
  NOR3_X1 U18012 ( .A1(n14642), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15772), .ZN(n15786) );
  NOR2_X1 U18013 ( .A1(n14645), .A2(n15786), .ZN(n15874) );
  AOI22_X1 U18014 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14646) );
  OAI21_X1 U18015 ( .B1(n19953), .B2(n14647), .A(n14646), .ZN(n14648) );
  AOI21_X1 U18016 ( .B1(n14649), .B2(n19947), .A(n14648), .ZN(n14650) );
  OAI21_X1 U18017 ( .B1(n15874), .B2(n19803), .A(n14650), .ZN(P1_U2989) );
  XNOR2_X1 U18018 ( .A(n14652), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14653) );
  XNOR2_X1 U18019 ( .A(n14651), .B(n14653), .ZN(n15897) );
  AOI22_X1 U18020 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14654) );
  OAI21_X1 U18021 ( .B1(n19953), .B2(n14655), .A(n14654), .ZN(n14656) );
  AOI21_X1 U18022 ( .B1(n14657), .B2(n19947), .A(n14656), .ZN(n14658) );
  OAI21_X1 U18023 ( .B1(n15897), .B2(n19803), .A(n14658), .ZN(P1_U2991) );
  AOI21_X1 U18024 ( .B1(n14661), .B2(n19967), .A(n14660), .ZN(n14665) );
  OAI21_X1 U18025 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14663), .A(
        n14662), .ZN(n14664) );
  INV_X1 U18026 ( .A(n14666), .ZN(n14675) );
  AOI21_X1 U18027 ( .B1(n14680), .B2(n14668), .A(n14667), .ZN(n14672) );
  INV_X1 U18028 ( .A(n14669), .ZN(n14688) );
  AOI21_X1 U18029 ( .B1(n14688), .B2(n14670), .A(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14671) );
  NOR2_X1 U18030 ( .A1(n14672), .A2(n14671), .ZN(n14673) );
  AOI211_X1 U18031 ( .C1(n19967), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14676) );
  OAI21_X1 U18032 ( .B1(n14677), .B2(n19977), .A(n14676), .ZN(P1_U3002) );
  INV_X1 U18033 ( .A(n14678), .ZN(n14693) );
  NAND3_X1 U18034 ( .A1(n14688), .A2(n14680), .A3(n14679), .ZN(n14681) );
  OAI211_X1 U18035 ( .C1(n14683), .C2(n19983), .A(n14682), .B(n14681), .ZN(
        n14684) );
  AOI21_X1 U18036 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14693), .A(
        n14684), .ZN(n14685) );
  OAI21_X1 U18037 ( .B1(n14686), .B2(n19977), .A(n14685), .ZN(P1_U3003) );
  NAND2_X1 U18038 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  OAI211_X1 U18039 ( .C1(n14691), .C2(n19983), .A(n14690), .B(n14689), .ZN(
        n14692) );
  AOI21_X1 U18040 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14693), .A(
        n14692), .ZN(n14694) );
  OAI21_X1 U18041 ( .B1(n14695), .B2(n19977), .A(n14694), .ZN(P1_U3004) );
  AOI22_X1 U18042 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15815), .B1(
        n14697), .B2(n14696), .ZN(n14700) );
  INV_X1 U18043 ( .A(n14698), .ZN(n14699) );
  OAI211_X1 U18044 ( .C1(n14701), .C2(n19983), .A(n14700), .B(n14699), .ZN(
        n14702) );
  INV_X1 U18045 ( .A(n14702), .ZN(n14703) );
  OAI21_X1 U18046 ( .B1(n14704), .B2(n19977), .A(n14703), .ZN(P1_U3005) );
  INV_X1 U18047 ( .A(n14705), .ZN(n14709) );
  NAND3_X1 U18048 ( .A1(n14707), .A2(n14706), .A3(n15739), .ZN(n15820) );
  OAI211_X1 U18049 ( .C1(n14709), .C2(n15820), .A(n14708), .B(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14714) );
  OAI21_X1 U18050 ( .B1(n15739), .B2(n15810), .A(n12646), .ZN(n14713) );
  OAI21_X1 U18051 ( .B1(n14711), .B2(n19983), .A(n14710), .ZN(n14712) );
  AOI21_X1 U18052 ( .B1(n14714), .B2(n14713), .A(n14712), .ZN(n14715) );
  OAI21_X1 U18053 ( .B1(n14716), .B2(n19977), .A(n14715), .ZN(P1_U3007) );
  NOR2_X1 U18054 ( .A1(n14733), .A2(n14732), .ZN(n14717) );
  OAI21_X1 U18055 ( .B1(n14717), .B2(n14772), .A(n14735), .ZN(n15578) );
  OAI21_X1 U18056 ( .B1(n15640), .B2(n19983), .A(n14718), .ZN(n14720) );
  NAND3_X1 U18057 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n14740), .ZN(n15585) );
  AOI221_X1 U18058 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C1(n12639), .C2(n14602), .A(
        n15585), .ZN(n14719) );
  AOI211_X1 U18059 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15578), .A(
        n14720), .B(n14719), .ZN(n14721) );
  OAI21_X1 U18060 ( .B1(n14722), .B2(n19977), .A(n14721), .ZN(P1_U3009) );
  NAND2_X1 U18061 ( .A1(n14723), .A2(n15785), .ZN(n14725) );
  NAND2_X1 U18062 ( .A1(n15772), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14724) );
  OR2_X1 U18063 ( .A1(n14741), .A2(n14724), .ZN(n15579) );
  NOR2_X1 U18064 ( .A1(n14726), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15581) );
  AOI21_X1 U18065 ( .B1(n14726), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15581), .ZN(n15754) );
  INV_X1 U18066 ( .A(n15659), .ZN(n14738) );
  INV_X1 U18067 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14728) );
  NAND2_X1 U18068 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n14740), .ZN(
        n14727) );
  OAI22_X1 U18069 ( .A1(n19957), .A2(n14728), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14727), .ZN(n14737) );
  NAND2_X1 U18070 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15855), .ZN(
        n14730) );
  OAI22_X1 U18071 ( .A1(n14731), .A2(n14730), .B1(n19981), .B2(n14729), .ZN(
        n15854) );
  OAI21_X1 U18072 ( .B1(n15856), .B2(n15854), .A(n14732), .ZN(n14734) );
  AOI21_X1 U18073 ( .B1(n14735), .B2(n14734), .A(n14733), .ZN(n14736) );
  AOI211_X1 U18074 ( .C1(n19967), .C2(n14738), .A(n14737), .B(n14736), .ZN(
        n14739) );
  OAI21_X1 U18075 ( .B1(n15754), .B2(n19977), .A(n14739), .ZN(P1_U3011) );
  INV_X1 U18076 ( .A(n14740), .ZN(n14749) );
  NAND2_X1 U18077 ( .A1(n9588), .A2(n15831), .ZN(n14742) );
  MUX2_X1 U18078 ( .A(n15785), .B(n14742), .S(n14741), .Z(n14743) );
  XNOR2_X1 U18079 ( .A(n14743), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15756) );
  NAND2_X1 U18080 ( .A1(n15756), .A2(n19970), .ZN(n14748) );
  INV_X1 U18081 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14744) );
  OAI22_X1 U18082 ( .A1(n15671), .A2(n19983), .B1(n19957), .B2(n14744), .ZN(
        n14745) );
  AOI21_X1 U18083 ( .B1(n14746), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14745), .ZN(n14747) );
  OAI211_X1 U18084 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n14749), .A(
        n14748), .B(n14747), .ZN(P1_U3012) );
  AND2_X1 U18085 ( .A1(n14765), .A2(n14750), .ZN(n14752) );
  NOR2_X1 U18086 ( .A1(n14752), .A2(n14751), .ZN(n14754) );
  NOR2_X1 U18087 ( .A1(n15772), .A2(n14754), .ZN(n14753) );
  AOI22_X1 U18088 ( .A1(n15772), .A2(n14754), .B1(n11919), .B2(n14753), .ZN(
        n14755) );
  XNOR2_X1 U18089 ( .A(n14757), .B(n14755), .ZN(n15764) );
  AOI22_X1 U18090 ( .A1(n14756), .A2(n19967), .B1(n19940), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14761) );
  OAI21_X1 U18091 ( .B1(n15821), .B2(n14758), .A(n14757), .ZN(n14759) );
  OAI21_X1 U18092 ( .B1(n14772), .B2(n15832), .A(n15853), .ZN(n15830) );
  NAND2_X1 U18093 ( .A1(n14759), .A2(n15830), .ZN(n14760) );
  OAI211_X1 U18094 ( .C1(n15764), .C2(n19977), .A(n14761), .B(n14760), .ZN(
        P1_U3014) );
  NOR2_X1 U18095 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14774) );
  INV_X1 U18096 ( .A(n14762), .ZN(n14763) );
  OAI21_X1 U18097 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n15774) );
  NOR2_X1 U18098 ( .A1(n15771), .A2(n15774), .ZN(n14769) );
  NOR2_X1 U18099 ( .A1(n14774), .A2(n14769), .ZN(n14771) );
  INV_X1 U18100 ( .A(n14766), .ZN(n14770) );
  INV_X1 U18101 ( .A(n14767), .ZN(n14768) );
  OAI22_X1 U18102 ( .A1(n14771), .A2(n14770), .B1(n14769), .B2(n14768), .ZN(
        n15770) );
  INV_X1 U18103 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14773) );
  INV_X1 U18104 ( .A(n14772), .ZN(n15896) );
  AOI21_X1 U18105 ( .B1(n15852), .B2(n15896), .A(n15860), .ZN(n15843) );
  OAI22_X1 U18106 ( .A1(n19957), .A2(n14773), .B1(n11919), .B2(n15843), .ZN(
        n14777) );
  INV_X1 U18107 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15842) );
  NOR2_X1 U18108 ( .A1(n15842), .A2(n11919), .ZN(n14775) );
  NOR4_X1 U18109 ( .A1(n15821), .A2(n14775), .A3(n14774), .A4(n15852), .ZN(
        n14776) );
  AOI211_X1 U18110 ( .C1(n19967), .C2(n14778), .A(n14777), .B(n14776), .ZN(
        n14779) );
  OAI21_X1 U18111 ( .B1(n15770), .B2(n19977), .A(n14779), .ZN(P1_U3015) );
  AOI21_X1 U18112 ( .B1(n14782), .B2(n14781), .A(n14780), .ZN(n15784) );
  INV_X1 U18113 ( .A(n15888), .ZN(n15893) );
  AOI21_X1 U18114 ( .B1(n15871), .B2(n14788), .A(n15893), .ZN(n14786) );
  AND2_X1 U18115 ( .A1(n14783), .A2(n15872), .ZN(n14792) );
  INV_X1 U18116 ( .A(n15887), .ZN(n14784) );
  OAI21_X1 U18117 ( .B1(n19981), .B2(n14792), .A(n14784), .ZN(n14785) );
  OR2_X1 U18118 ( .A1(n14786), .A2(n14785), .ZN(n15866) );
  INV_X1 U18119 ( .A(n15866), .ZN(n14789) );
  INV_X1 U18120 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14787) );
  NAND2_X1 U18121 ( .A1(n14788), .A2(n14787), .ZN(n15870) );
  AOI221_X1 U18122 ( .B1(n14790), .B2(n14789), .C1(n15870), .C2(n14789), .A(
        n14791), .ZN(n14797) );
  INV_X1 U18123 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20723) );
  NOR2_X1 U18124 ( .A1(n15889), .A2(n14790), .ZN(n19976) );
  NAND2_X1 U18125 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19976), .ZN(
        n15895) );
  NAND2_X1 U18126 ( .A1(n19981), .A2(n15895), .ZN(n15922) );
  NAND3_X1 U18127 ( .A1(n14792), .A2(n14791), .A3(n15922), .ZN(n14795) );
  XNOR2_X1 U18128 ( .A(n14123), .B(n14793), .ZN(n15723) );
  NAND2_X1 U18129 ( .A1(n15723), .A2(n19967), .ZN(n14794) );
  OAI211_X1 U18130 ( .C1(n20723), .C2(n19957), .A(n14795), .B(n14794), .ZN(
        n14796) );
  NOR2_X1 U18131 ( .A1(n14797), .A2(n14796), .ZN(n14798) );
  OAI21_X1 U18132 ( .B1(n15784), .B2(n19977), .A(n14798), .ZN(P1_U3019) );
  NAND3_X1 U18133 ( .A1(n15889), .A2(n15896), .A3(n14799), .ZN(n14808) );
  AOI21_X1 U18134 ( .B1(n14801), .B2(n14800), .A(n15889), .ZN(n14803) );
  NOR2_X1 U18135 ( .A1(n19957), .A2(n13525), .ZN(n14802) );
  AOI211_X1 U18136 ( .C1(n19967), .C2(n14804), .A(n14803), .B(n14802), .ZN(
        n14807) );
  NAND3_X1 U18137 ( .A1(n14805), .A2(n19970), .A3(n13528), .ZN(n14806) );
  NAND3_X1 U18138 ( .A1(n14808), .A2(n14807), .A3(n14806), .ZN(P1_U3030) );
  XNOR2_X1 U18139 ( .A(n13840), .B(P1_STATEBS16_REG_SCAN_IN), .ZN(n14809) );
  OAI22_X1 U18140 ( .A1(n14809), .A2(n20567), .B1(n20315), .B2(n14816), .ZN(
        n14810) );
  MUX2_X1 U18141 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14810), .S(
        n19992), .Z(P1_U3477) );
  INV_X1 U18142 ( .A(n14814), .ZN(n14811) );
  OAI22_X1 U18143 ( .A1(n14812), .A2(n20283), .B1(n12577), .B2(
        P1_STATEBS16_REG_SCAN_IN), .ZN(n14813) );
  OAI21_X1 U18144 ( .B1(n14813), .B2(n20446), .A(n20625), .ZN(n14815) );
  OR2_X1 U18145 ( .A1(n13842), .A2(n14814), .ZN(n20622) );
  NOR2_X1 U18146 ( .A1(n20622), .A2(n13840), .ZN(n20529) );
  NAND3_X1 U18147 ( .A1(n20529), .A2(n20625), .A3(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20520) );
  OAI211_X1 U18148 ( .C1(n14817), .C2(n14816), .A(n14815), .B(n20520), .ZN(
        n14818) );
  MUX2_X1 U18149 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n14818), .S(
        n19992), .Z(P1_U3475) );
  INV_X1 U18150 ( .A(n15934), .ZN(n20772) );
  OAI22_X1 U18151 ( .A1(n14821), .A2(n20772), .B1(n14820), .B2(n14819), .ZN(
        n14822) );
  MUX2_X1 U18152 ( .A(n14822), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20781), .Z(P1_U3469) );
  INV_X1 U18153 ( .A(n14823), .ZN(n14835) );
  AOI211_X1 U18154 ( .C1(n14826), .C2(n14824), .A(n14825), .B(n19638), .ZN(
        n14827) );
  INV_X1 U18155 ( .A(n14827), .ZN(n14834) );
  NAND2_X1 U18156 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18927), .ZN(n14831) );
  AOI22_X1 U18157 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n9691), .ZN(n14830) );
  OAI211_X1 U18158 ( .C1(n18937), .C2(n15198), .A(n14831), .B(n14830), .ZN(
        n14832) );
  AOI21_X1 U18159 ( .B1(n15201), .B2(n18932), .A(n14832), .ZN(n14833) );
  OAI211_X1 U18160 ( .C1(n18924), .C2(n14835), .A(n14834), .B(n14833), .ZN(
        P2_U2827) );
  AOI211_X1 U18161 ( .C1(n15113), .C2(n14850), .A(n14836), .B(n19638), .ZN(
        n14838) );
  OAI22_X1 U18162 ( .A1(n20815), .A2(n18922), .B1(n19686), .B2(n18921), .ZN(
        n14837) );
  AOI211_X1 U18163 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n18927), .A(n14838), .B(
        n14837), .ZN(n14847) );
  NOR2_X1 U18164 ( .A1(n14840), .A2(n14841), .ZN(n14842) );
  OR2_X1 U18165 ( .A1(n14839), .A2(n14842), .ZN(n15110) );
  OAI21_X1 U18166 ( .B1(n14843), .B2(n14844), .A(n15004), .ZN(n15013) );
  OAI22_X1 U18167 ( .A1(n15110), .A2(n18954), .B1(n15013), .B2(n18937), .ZN(
        n14845) );
  INV_X1 U18168 ( .A(n14845), .ZN(n14846) );
  OAI211_X1 U18169 ( .C1(n14848), .C2(n18924), .A(n14847), .B(n14846), .ZN(
        P2_U2834) );
  INV_X1 U18170 ( .A(n15128), .ZN(n14849) );
  AOI22_X1 U18171 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n18927), .B1(n14849), 
        .B2(n18891), .ZN(n14864) );
  OAI211_X1 U18172 ( .C1(n14851), .C2(n15128), .A(n18933), .B(n14850), .ZN(
        n14863) );
  AND2_X1 U18173 ( .A1(n14853), .A2(n14852), .ZN(n14854) );
  OR2_X1 U18174 ( .A1(n14854), .A2(n14840), .ZN(n15282) );
  AOI22_X1 U18175 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n9691), .ZN(n14859) );
  NOR2_X1 U18176 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  NOR2_X1 U18177 ( .A1(n14843), .A2(n14857), .ZN(n15279) );
  NAND2_X1 U18178 ( .A1(n18958), .A2(n15279), .ZN(n14858) );
  OAI211_X1 U18179 ( .C1(n18954), .C2(n15282), .A(n14859), .B(n14858), .ZN(
        n14860) );
  AOI21_X1 U18180 ( .B1(n14861), .B2(n13079), .A(n14860), .ZN(n14862) );
  NAND3_X1 U18181 ( .A1(n14864), .A2(n14863), .A3(n14862), .ZN(P2_U2835) );
  INV_X1 U18182 ( .A(n14865), .ZN(n14866) );
  NAND2_X1 U18183 ( .A1(n14866), .A2(n14915), .ZN(n14867) );
  OAI21_X1 U18184 ( .B1(n14915), .B2(n14277), .A(n14867), .ZN(P2_U2856) );
  XNOR2_X1 U18185 ( .A(n14868), .B(n14869), .ZN(n14952) );
  NOR2_X1 U18186 ( .A1(n15947), .A2(n13608), .ZN(n14870) );
  AOI21_X1 U18187 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n13608), .A(n14870), .ZN(
        n14871) );
  OAI21_X1 U18188 ( .B1(n14952), .B2(n14942), .A(n14871), .ZN(P2_U2858) );
  NOR2_X1 U18189 ( .A1(n14873), .A2(n14872), .ZN(n14874) );
  XOR2_X1 U18190 ( .A(n14875), .B(n14874), .Z(n14958) );
  NAND2_X1 U18191 ( .A1(n13608), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14877) );
  NAND2_X1 U18192 ( .A1(n15201), .A2(n14915), .ZN(n14876) );
  OAI211_X1 U18193 ( .C1(n14958), .C2(n14942), .A(n14877), .B(n14876), .ZN(
        P2_U2859) );
  XNOR2_X1 U18194 ( .A(n14878), .B(n14879), .ZN(n14977) );
  OR2_X1 U18195 ( .A1(n14880), .A2(n14881), .ZN(n14882) );
  AND2_X1 U18196 ( .A1(n9660), .A2(n14882), .ZN(n15072) );
  NOR2_X1 U18197 ( .A1(n14932), .A2(n15977), .ZN(n14883) );
  AOI21_X1 U18198 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14932), .A(n14883), .ZN(
        n14884) );
  OAI21_X1 U18199 ( .B1(n14977), .B2(n14942), .A(n14884), .ZN(P2_U2861) );
  OAI21_X1 U18200 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n14986) );
  AND2_X1 U18201 ( .A1(n13275), .A2(n14888), .ZN(n14889) );
  OR2_X1 U18202 ( .A1(n14880), .A2(n14889), .ZN(n15983) );
  NOR2_X1 U18203 ( .A1(n14932), .A2(n15983), .ZN(n14890) );
  AOI21_X1 U18204 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n14932), .A(n14890), .ZN(
        n14891) );
  OAI21_X1 U18205 ( .B1(n14986), .B2(n14942), .A(n14891), .ZN(P2_U2862) );
  AOI21_X1 U18206 ( .B1(n13146), .B2(n14893), .A(n14892), .ZN(n14895) );
  XOR2_X1 U18207 ( .A(n14895), .B(n14894), .Z(n14993) );
  NAND2_X1 U18208 ( .A1(n14932), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n14897) );
  NAND2_X1 U18209 ( .A1(n14915), .A2(n16014), .ZN(n14896) );
  OAI211_X1 U18210 ( .C1(n14993), .C2(n14942), .A(n14897), .B(n14896), .ZN(
        P2_U2863) );
  OAI21_X1 U18211 ( .B1(n14900), .B2(n14899), .A(n14898), .ZN(n15003) );
  AOI21_X1 U18212 ( .B1(n14901), .B2(n14907), .A(n13276), .ZN(n16144) );
  INV_X1 U18213 ( .A(n16144), .ZN(n15096) );
  NOR2_X1 U18214 ( .A1(n14932), .A2(n15096), .ZN(n14902) );
  AOI21_X1 U18215 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n14932), .A(n14902), .ZN(
        n14903) );
  OAI21_X1 U18216 ( .B1(n15003), .B2(n14942), .A(n14903), .ZN(P2_U2864) );
  AND2_X1 U18217 ( .A1(n14935), .A2(n14904), .ZN(n14912) );
  OAI21_X1 U18218 ( .B1(n14912), .B2(n14905), .A(n10439), .ZN(n15012) );
  OR2_X1 U18219 ( .A1(n14839), .A2(n14906), .ZN(n14908) );
  AND2_X1 U18220 ( .A1(n14908), .A2(n14907), .ZN(n16023) );
  INV_X1 U18221 ( .A(n16023), .ZN(n15252) );
  NOR2_X1 U18222 ( .A1(n15252), .A2(n13608), .ZN(n14909) );
  AOI21_X1 U18223 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n14932), .A(n14909), .ZN(
        n14910) );
  OAI21_X1 U18224 ( .B1(n15012), .B2(n14942), .A(n14910), .ZN(P2_U2865) );
  AND2_X1 U18225 ( .A1(n14935), .A2(n14911), .ZN(n14918) );
  INV_X1 U18226 ( .A(n14912), .ZN(n14913) );
  OAI21_X1 U18227 ( .B1(n14918), .B2(n14914), .A(n14913), .ZN(n15020) );
  NAND2_X1 U18228 ( .A1(n13608), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14917) );
  INV_X1 U18229 ( .A(n15110), .ZN(n15262) );
  NAND2_X1 U18230 ( .A1(n15262), .A2(n14915), .ZN(n14916) );
  OAI211_X1 U18231 ( .C1(n15020), .C2(n14942), .A(n14917), .B(n14916), .ZN(
        P2_U2866) );
  NAND2_X1 U18232 ( .A1(n14935), .A2(n14930), .ZN(n14929) );
  AOI21_X1 U18233 ( .B1(n14919), .B2(n14925), .A(n14918), .ZN(n14920) );
  INV_X1 U18234 ( .A(n14920), .ZN(n15026) );
  MUX2_X1 U18235 ( .A(n15282), .B(n14921), .S(n13608), .Z(n14922) );
  OAI21_X1 U18236 ( .B1(n15026), .B2(n14942), .A(n14922), .ZN(P2_U2867) );
  NAND2_X1 U18237 ( .A1(n14929), .A2(n14923), .ZN(n14924) );
  INV_X1 U18238 ( .A(n16009), .ZN(n14928) );
  MUX2_X1 U18239 ( .A(n14926), .B(n12334), .S(n13608), .Z(n14927) );
  OAI21_X1 U18240 ( .B1(n14928), .B2(n14942), .A(n14927), .ZN(P2_U2868) );
  OAI21_X1 U18241 ( .B1(n14935), .B2(n14930), .A(n14929), .ZN(n15035) );
  INV_X1 U18242 ( .A(n14931), .ZN(n18813) );
  NOR2_X1 U18243 ( .A1(n14932), .A2(n18813), .ZN(n14933) );
  AOI21_X1 U18244 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n14932), .A(n14933), .ZN(
        n14934) );
  OAI21_X1 U18245 ( .B1(n15035), .B2(n14942), .A(n14934), .ZN(P2_U2869) );
  INV_X1 U18246 ( .A(n14935), .ZN(n14936) );
  OAI21_X1 U18247 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n15047) );
  AOI21_X1 U18248 ( .B1(n14939), .B2(n14161), .A(n12525), .ZN(n18825) );
  INV_X1 U18249 ( .A(n18825), .ZN(n14940) );
  INV_X1 U18250 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n18818) );
  MUX2_X1 U18251 ( .A(n14940), .B(n18818), .S(n13608), .Z(n14941) );
  OAI21_X1 U18252 ( .B1(n15047), .B2(n14942), .A(n14941), .ZN(P2_U2870) );
  OR2_X1 U18253 ( .A1(n14944), .A2(n14943), .ZN(n14945) );
  NAND2_X1 U18254 ( .A1(n14946), .A2(n14945), .ZN(n15185) );
  INV_X1 U18255 ( .A(n15185), .ZN(n15948) );
  OAI22_X1 U18256 ( .A1(n14948), .A2(n16003), .B1(n18973), .B2(n14947), .ZN(
        n14949) );
  AOI21_X1 U18257 ( .B1(n18996), .B2(n15948), .A(n14949), .ZN(n14951) );
  AOI22_X1 U18258 ( .A1(n18963), .A2(BUF2_REG_29__SCAN_IN), .B1(n18962), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14950) );
  OAI211_X1 U18259 ( .C1(n14952), .C2(n18978), .A(n14951), .B(n14950), .ZN(
        P2_U2890) );
  INV_X1 U18260 ( .A(n15198), .ZN(n14955) );
  OAI22_X1 U18261 ( .A1(n14953), .A2(n16003), .B1(n18973), .B2(n13432), .ZN(
        n14954) );
  AOI21_X1 U18262 ( .B1(n18996), .B2(n14955), .A(n14954), .ZN(n14957) );
  AOI22_X1 U18263 ( .A1(n18963), .A2(BUF2_REG_28__SCAN_IN), .B1(n18962), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14956) );
  OAI211_X1 U18264 ( .C1(n14958), .C2(n18978), .A(n14957), .B(n14956), .ZN(
        P2_U2891) );
  INV_X1 U18265 ( .A(n14959), .ZN(n14968) );
  NOR2_X1 U18266 ( .A1(n14970), .A2(n14961), .ZN(n14962) );
  OR2_X1 U18267 ( .A1(n14828), .A2(n14962), .ZN(n15211) );
  INV_X1 U18268 ( .A(n15211), .ZN(n15958) );
  OAI22_X1 U18269 ( .A1(n14964), .A2(n16003), .B1(n18973), .B2(n14963), .ZN(
        n14965) );
  AOI21_X1 U18270 ( .B1(n18996), .B2(n15958), .A(n14965), .ZN(n14967) );
  AOI22_X1 U18271 ( .A1(n18963), .A2(BUF2_REG_27__SCAN_IN), .B1(n18962), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14966) );
  OAI211_X1 U18272 ( .C1(n14968), .C2(n18978), .A(n14967), .B(n14966), .ZN(
        P2_U2892) );
  AOI21_X1 U18273 ( .B1(n14971), .B2(n14969), .A(n14970), .ZN(n15980) );
  OAI22_X1 U18274 ( .A1(n14973), .A2(n16003), .B1(n18973), .B2(n14972), .ZN(
        n14974) );
  AOI21_X1 U18275 ( .B1(n18996), .B2(n15980), .A(n14974), .ZN(n14976) );
  AOI22_X1 U18276 ( .A1(n18963), .A2(BUF2_REG_26__SCAN_IN), .B1(n18962), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14975) );
  OAI211_X1 U18277 ( .C1(n14977), .C2(n18978), .A(n14976), .B(n14975), .ZN(
        P2_U2893) );
  OAI21_X1 U18278 ( .B1(n14979), .B2(n14978), .A(n14969), .ZN(n16126) );
  INV_X1 U18279 ( .A(n16126), .ZN(n15984) );
  NAND2_X1 U18280 ( .A1(n18995), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n14980) );
  OAI21_X1 U18281 ( .B1(n16003), .B2(n14981), .A(n14980), .ZN(n14984) );
  INV_X1 U18282 ( .A(n18963), .ZN(n15042) );
  INV_X1 U18283 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n14982) );
  INV_X1 U18284 ( .A(n18962), .ZN(n15040) );
  OAI22_X1 U18285 ( .A1(n15042), .A2(n14982), .B1(n15040), .B2(n16349), .ZN(
        n14983) );
  AOI211_X1 U18286 ( .C1(n18996), .C2(n15984), .A(n14984), .B(n14983), .ZN(
        n14985) );
  OAI21_X1 U18287 ( .B1(n14986), .B2(n18978), .A(n14985), .ZN(P2_U2894) );
  INV_X1 U18288 ( .A(n15235), .ZN(n14990) );
  OAI22_X1 U18289 ( .A1(n14988), .A2(n16003), .B1(n18973), .B2(n14987), .ZN(
        n14989) );
  AOI21_X1 U18290 ( .B1(n18996), .B2(n14990), .A(n14989), .ZN(n14992) );
  AOI22_X1 U18291 ( .A1(n18963), .A2(BUF2_REG_24__SCAN_IN), .B1(n18962), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14991) );
  OAI211_X1 U18292 ( .C1(n14993), .C2(n18978), .A(n14992), .B(n14991), .ZN(
        P2_U2895) );
  OAI21_X1 U18293 ( .B1(n14996), .B2(n14994), .A(n14995), .ZN(n16137) );
  INV_X1 U18294 ( .A(n16137), .ZN(n15994) );
  NAND2_X1 U18295 ( .A1(n18995), .A2(P2_EAX_REG_23__SCAN_IN), .ZN(n14997) );
  OAI21_X1 U18296 ( .B1(n16003), .B2(n19120), .A(n14997), .ZN(n15001) );
  INV_X1 U18297 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n14999) );
  INV_X1 U18298 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14998) );
  OAI22_X1 U18299 ( .A1(n15042), .A2(n14999), .B1(n15040), .B2(n14998), .ZN(
        n15000) );
  AOI211_X1 U18300 ( .C1(n18996), .C2(n15994), .A(n15001), .B(n15000), .ZN(
        n15002) );
  OAI21_X1 U18301 ( .B1(n15003), .B2(n18978), .A(n15002), .ZN(P2_U2896) );
  AOI21_X1 U18302 ( .B1(n15005), .B2(n15004), .A(n14994), .ZN(n15530) );
  OAI22_X1 U18303 ( .A1(n19109), .A2(n16003), .B1(n18973), .B2(n15006), .ZN(
        n15010) );
  INV_X1 U18304 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n15008) );
  INV_X1 U18305 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n15007) );
  OAI22_X1 U18306 ( .A1(n15042), .A2(n15008), .B1(n15040), .B2(n15007), .ZN(
        n15009) );
  AOI211_X1 U18307 ( .C1(n18996), .C2(n15530), .A(n15010), .B(n15009), .ZN(
        n15011) );
  OAI21_X1 U18308 ( .B1(n15012), .B2(n18978), .A(n15011), .ZN(P2_U2897) );
  INV_X1 U18309 ( .A(n15013), .ZN(n15261) );
  NAND2_X1 U18310 ( .A1(n18995), .A2(P2_EAX_REG_21__SCAN_IN), .ZN(n15014) );
  OAI21_X1 U18311 ( .B1(n16003), .B2(n19106), .A(n15014), .ZN(n15018) );
  INV_X1 U18312 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15016) );
  INV_X1 U18313 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15015) );
  OAI22_X1 U18314 ( .A1(n15042), .A2(n15016), .B1(n15040), .B2(n15015), .ZN(
        n15017) );
  AOI211_X1 U18315 ( .C1(n18996), .C2(n15261), .A(n15018), .B(n15017), .ZN(
        n15019) );
  OAI21_X1 U18316 ( .B1(n15020), .B2(n18978), .A(n15019), .ZN(P2_U2898) );
  OAI22_X1 U18317 ( .A1(n19103), .A2(n16003), .B1(n18973), .B2(n15021), .ZN(
        n15024) );
  INV_X1 U18318 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n15022) );
  OAI22_X1 U18319 ( .A1(n15042), .A2(n15022), .B1(n15040), .B2(n19101), .ZN(
        n15023) );
  AOI211_X1 U18320 ( .C1(n18996), .C2(n15279), .A(n15024), .B(n15023), .ZN(
        n15025) );
  OAI21_X1 U18321 ( .B1(n15026), .B2(n18978), .A(n15025), .ZN(P2_U2899) );
  XNOR2_X1 U18322 ( .A(n15028), .B(n15036), .ZN(n18812) );
  INV_X1 U18323 ( .A(n18812), .ZN(n15033) );
  OAI22_X1 U18324 ( .A1(n19094), .A2(n16003), .B1(n18973), .B2(n15029), .ZN(
        n15032) );
  AOI22_X1 U18325 ( .A1(n18963), .A2(BUF2_REG_18__SCAN_IN), .B1(n18962), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15030) );
  INV_X1 U18326 ( .A(n15030), .ZN(n15031) );
  AOI211_X1 U18327 ( .C1(n18996), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        n15034) );
  OAI21_X1 U18328 ( .B1(n15035), .B2(n18978), .A(n15034), .ZN(P2_U2901) );
  OAI21_X1 U18329 ( .B1(n15037), .B2(n14155), .A(n15036), .ZN(n18829) );
  INV_X1 U18330 ( .A(n18829), .ZN(n15045) );
  NAND2_X1 U18331 ( .A1(n18995), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n15038) );
  OAI21_X1 U18332 ( .B1(n16003), .B2(n19089), .A(n15038), .ZN(n15044) );
  INV_X1 U18333 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15041) );
  INV_X1 U18334 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n15039) );
  OAI22_X1 U18335 ( .A1(n15042), .A2(n15041), .B1(n15040), .B2(n15039), .ZN(
        n15043) );
  AOI211_X1 U18336 ( .C1(n18996), .C2(n15045), .A(n15044), .B(n15043), .ZN(
        n15046) );
  OAI21_X1 U18337 ( .B1(n15047), .B2(n18978), .A(n15046), .ZN(P2_U2902) );
  NAND2_X1 U18338 ( .A1(n15048), .A2(n16115), .ZN(n15051) );
  AOI21_X1 U18339 ( .B1(n19041), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15049), .ZN(n15050) );
  OAI211_X1 U18340 ( .C1(n15052), .C2(n16034), .A(n15051), .B(n15050), .ZN(
        n15053) );
  AOI21_X1 U18341 ( .B1(n15054), .B2(n19048), .A(n15053), .ZN(n15055) );
  OAI21_X1 U18342 ( .B1(n15056), .B2(n16109), .A(n15055), .ZN(P2_U2984) );
  XNOR2_X1 U18343 ( .A(n15057), .B(n15062), .ZN(n15218) );
  NAND2_X1 U18344 ( .A1(n15959), .A2(n19047), .ZN(n15058) );
  NAND2_X1 U18345 ( .A1(n19040), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15209) );
  OAI211_X1 U18346 ( .C1(n16124), .C2(n15059), .A(n15058), .B(n15209), .ZN(
        n15060) );
  AOI21_X1 U18347 ( .B1(n15962), .B2(n16115), .A(n15060), .ZN(n15065) );
  NAND2_X1 U18348 ( .A1(n15063), .A2(n15062), .ZN(n15215) );
  NAND3_X1 U18349 ( .A1(n12511), .A2(n19048), .A3(n15215), .ZN(n15064) );
  OAI211_X1 U18350 ( .C1(n15218), .C2(n16109), .A(n15065), .B(n15064), .ZN(
        P2_U2987) );
  OAI21_X1 U18351 ( .B1(n15066), .B2(n15081), .A(n15082), .ZN(n15067) );
  XOR2_X1 U18352 ( .A(n15068), .B(n15067), .Z(n15228) );
  AOI21_X1 U18353 ( .B1(n15069), .B2(n9630), .A(n15061), .ZN(n15226) );
  INV_X1 U18354 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15070) );
  NAND2_X1 U18355 ( .A1(n19040), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15219) );
  OAI21_X1 U18356 ( .B1(n16124), .B2(n15070), .A(n15219), .ZN(n15071) );
  AOI21_X1 U18357 ( .B1(n19047), .B2(n15072), .A(n15071), .ZN(n15073) );
  OAI21_X1 U18358 ( .B1(n15074), .B2(n19052), .A(n15073), .ZN(n15075) );
  AOI21_X1 U18359 ( .B1(n15226), .B2(n19048), .A(n15075), .ZN(n15076) );
  OAI21_X1 U18360 ( .B1(n15228), .B2(n16109), .A(n15076), .ZN(P2_U2988) );
  OAI21_X1 U18361 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15077), .A(
        n9630), .ZN(n16135) );
  OAI22_X1 U18362 ( .A1(n16124), .A2(n15078), .B1(n19691), .B2(n18920), .ZN(
        n15080) );
  NOR2_X1 U18363 ( .A1(n16034), .A2(n15983), .ZN(n15079) );
  AOI211_X1 U18364 ( .C1(n16115), .C2(n15987), .A(n15080), .B(n15079), .ZN(
        n15085) );
  NAND2_X1 U18365 ( .A1(n9893), .A2(n15082), .ZN(n15083) );
  XOR2_X1 U18366 ( .A(n15083), .B(n15066), .Z(n16132) );
  NAND2_X1 U18367 ( .A1(n16132), .A2(n19046), .ZN(n15084) );
  OAI211_X1 U18368 ( .C1(n16135), .C2(n16108), .A(n15085), .B(n15084), .ZN(
        P2_U2989) );
  NAND2_X1 U18369 ( .A1(n15086), .A2(n15255), .ZN(n15087) );
  NAND2_X1 U18370 ( .A1(n15087), .A2(n15256), .ZN(n15092) );
  AND2_X1 U18371 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  OAI21_X1 U18372 ( .B1(n15092), .B2(n15091), .A(n15090), .ZN(n16143) );
  NAND2_X1 U18373 ( .A1(n15123), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15244) );
  NOR2_X1 U18374 ( .A1(n15243), .A2(n15244), .ZN(n15245) );
  OAI21_X1 U18375 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15245), .A(
        n15094), .ZN(n16148) );
  OR2_X1 U18376 ( .A1(n16148), .A2(n16108), .ZN(n15100) );
  OAI22_X1 U18377 ( .A1(n16124), .A2(n15095), .B1(n19688), .B2(n18920), .ZN(
        n15098) );
  NOR2_X1 U18378 ( .A1(n16034), .A2(n15096), .ZN(n15097) );
  AOI211_X1 U18379 ( .C1(n15997), .C2(n16115), .A(n15098), .B(n15097), .ZN(
        n15099) );
  OAI211_X1 U18380 ( .C1(n16109), .C2(n16143), .A(n15100), .B(n15099), .ZN(
        P2_U2991) );
  NAND2_X1 U18381 ( .A1(n15102), .A2(n15101), .ZN(n15116) );
  INV_X1 U18382 ( .A(n15117), .ZN(n15103) );
  AOI21_X1 U18383 ( .B1(n15116), .B2(n15104), .A(n15103), .ZN(n15108) );
  NAND2_X1 U18384 ( .A1(n15106), .A2(n15105), .ZN(n15107) );
  XNOR2_X1 U18385 ( .A(n15108), .B(n15107), .ZN(n15271) );
  NAND2_X1 U18386 ( .A1(n19040), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15265) );
  NAND2_X1 U18387 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15109) );
  OAI211_X1 U18388 ( .C1(n16034), .C2(n15110), .A(n15265), .B(n15109), .ZN(
        n15112) );
  OAI21_X1 U18389 ( .B1(n15123), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15244), .ZN(n15267) );
  NOR2_X1 U18390 ( .A1(n15267), .A2(n16108), .ZN(n15111) );
  AOI211_X1 U18391 ( .C1(n16115), .C2(n15113), .A(n15112), .B(n15111), .ZN(
        n15114) );
  OAI21_X1 U18392 ( .B1(n15271), .B2(n16109), .A(n15114), .ZN(P2_U2993) );
  NAND2_X1 U18393 ( .A1(n15116), .A2(n15115), .ZN(n15120) );
  NAND2_X1 U18394 ( .A1(n15118), .A2(n15117), .ZN(n15119) );
  XNOR2_X1 U18395 ( .A(n15120), .B(n15119), .ZN(n15291) );
  AOI21_X1 U18396 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15121), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15122) );
  INV_X1 U18397 ( .A(n15282), .ZN(n15126) );
  INV_X1 U18398 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15124) );
  NAND2_X1 U18399 ( .A1(n19040), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15280) );
  OAI21_X1 U18400 ( .B1(n16124), .B2(n15124), .A(n15280), .ZN(n15125) );
  AOI21_X1 U18401 ( .B1(n19047), .B2(n15126), .A(n15125), .ZN(n15127) );
  OAI21_X1 U18402 ( .B1(n15128), .B2(n19052), .A(n15127), .ZN(n15129) );
  AOI21_X1 U18403 ( .B1(n15289), .B2(n19048), .A(n15129), .ZN(n15130) );
  OAI21_X1 U18404 ( .B1(n16109), .B2(n15291), .A(n15130), .ZN(P2_U2994) );
  XNOR2_X1 U18405 ( .A(n15132), .B(n15131), .ZN(n15308) );
  INV_X1 U18406 ( .A(n15308), .ZN(n15143) );
  NOR2_X1 U18407 ( .A1(n19680), .A2(n18920), .ZN(n15137) );
  INV_X1 U18408 ( .A(n16031), .ZN(n15303) );
  INV_X1 U18409 ( .A(n15133), .ZN(n15134) );
  AOI211_X1 U18410 ( .C1(n15135), .C2(n15303), .A(n15134), .B(n16108), .ZN(
        n15136) );
  AOI211_X1 U18411 ( .C1(n18825), .C2(n19047), .A(n15137), .B(n15136), .ZN(
        n15142) );
  INV_X1 U18412 ( .A(n15138), .ZN(n18824) );
  OAI22_X1 U18413 ( .A1(n16124), .A2(n15139), .B1(n19052), .B2(n18824), .ZN(
        n15140) );
  INV_X1 U18414 ( .A(n15140), .ZN(n15141) );
  OAI211_X1 U18415 ( .C1(n15143), .C2(n16109), .A(n15142), .B(n15141), .ZN(
        P2_U2997) );
  NAND2_X1 U18416 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15355), .ZN(
        n15354) );
  NAND2_X1 U18417 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16158) );
  INV_X1 U18418 ( .A(n15355), .ZN(n16060) );
  NOR2_X1 U18419 ( .A1(n16158), .A2(n16060), .ZN(n16047) );
  AOI21_X1 U18420 ( .B1(n12377), .B2(n15354), .A(n16047), .ZN(n15145) );
  INV_X1 U18421 ( .A(n15145), .ZN(n15353) );
  NAND2_X1 U18422 ( .A1(n15148), .A2(n15147), .ZN(n15149) );
  XNOR2_X1 U18423 ( .A(n15146), .B(n15149), .ZN(n15351) );
  INV_X1 U18424 ( .A(n15150), .ZN(n18864) );
  OAI22_X1 U18425 ( .A1(n16124), .A2(n15151), .B1(n19052), .B2(n18864), .ZN(
        n15154) );
  OAI22_X1 U18426 ( .A1(n16034), .A2(n18857), .B1(n18920), .B2(n15152), .ZN(
        n15153) );
  AOI211_X1 U18427 ( .C1(n15351), .C2(n19046), .A(n15154), .B(n15153), .ZN(
        n15155) );
  OAI21_X1 U18428 ( .B1(n15353), .B2(n16108), .A(n15155), .ZN(P2_U3001) );
  INV_X1 U18429 ( .A(n15156), .ZN(n15157) );
  AOI21_X1 U18430 ( .B1(n15159), .B2(n15158), .A(n15157), .ZN(n15160) );
  INV_X1 U18431 ( .A(n16095), .ZN(n15162) );
  NAND2_X1 U18432 ( .A1(n15162), .A2(n16096), .ZN(n15163) );
  XNOR2_X1 U18433 ( .A(n15161), .B(n15163), .ZN(n15387) );
  OAI22_X1 U18434 ( .A1(n16124), .A2(n15164), .B1(n19668), .B2(n18920), .ZN(
        n15167) );
  INV_X1 U18435 ( .A(n18908), .ZN(n15165) );
  OAI22_X1 U18436 ( .A1(n19052), .A2(n15165), .B1(n16034), .B2(n18913), .ZN(
        n15166) );
  AOI211_X1 U18437 ( .C1(n15387), .C2(n19046), .A(n15167), .B(n15166), .ZN(
        n15168) );
  OAI21_X1 U18438 ( .B1(n9930), .B2(n16108), .A(n15168), .ZN(P2_U3007) );
  OAI21_X1 U18439 ( .B1(n15171), .B2(n15170), .A(n15169), .ZN(n15172) );
  XNOR2_X1 U18440 ( .A(n15172), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15395) );
  AOI22_X1 U18441 ( .A1(n16115), .A2(n15173), .B1(n19046), .B2(n15395), .ZN(
        n15180) );
  AOI21_X1 U18442 ( .B1(n15176), .B2(n15175), .A(n15174), .ZN(n15391) );
  AND2_X1 U18443 ( .A1(n19040), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15392) );
  AOI21_X1 U18444 ( .B1(n19048), .B2(n15391), .A(n15392), .ZN(n15179) );
  OR2_X1 U18445 ( .A1(n16124), .A2(n15173), .ZN(n15178) );
  NAND2_X1 U18446 ( .A1(n19047), .A2(n15393), .ZN(n15177) );
  NAND4_X1 U18447 ( .A1(n15180), .A2(n15179), .A3(n15178), .A4(n15177), .ZN(
        P2_U3013) );
  INV_X1 U18448 ( .A(n15182), .ZN(n15181) );
  NAND2_X1 U18449 ( .A1(n15181), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15190) );
  OAI21_X1 U18450 ( .B1(n15195), .B2(n15182), .A(n15196), .ZN(n15183) );
  NAND2_X1 U18451 ( .A1(n15183), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15189) );
  OAI21_X1 U18452 ( .B1(n15384), .B2(n15947), .A(n15184), .ZN(n15187) );
  NOR2_X1 U18453 ( .A1(n19058), .A2(n15185), .ZN(n15186) );
  NOR2_X1 U18454 ( .A1(n15187), .A2(n15186), .ZN(n15188) );
  OAI211_X1 U18455 ( .C1(n15204), .C2(n15190), .A(n15189), .B(n15188), .ZN(
        n15191) );
  AOI21_X1 U18456 ( .B1(n15192), .B2(n19063), .A(n15191), .ZN(n15193) );
  OAI21_X1 U18457 ( .B1(n15194), .B2(n16191), .A(n15193), .ZN(P2_U3017) );
  NOR2_X1 U18458 ( .A1(n15195), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15212) );
  INV_X1 U18459 ( .A(n15196), .ZN(n15214) );
  OAI21_X1 U18460 ( .B1(n15212), .B2(n15214), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15203) );
  INV_X1 U18461 ( .A(n15197), .ZN(n15200) );
  AOI211_X1 U18462 ( .C1(n15201), .C2(n19053), .A(n15200), .B(n15199), .ZN(
        n15202) );
  OAI211_X1 U18463 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15204), .A(
        n15203), .B(n15202), .ZN(n15205) );
  AOI21_X1 U18464 ( .B1(n15206), .B2(n19063), .A(n15205), .ZN(n15207) );
  OAI21_X1 U18465 ( .B1(n15208), .B2(n16191), .A(n15207), .ZN(P2_U3018) );
  NAND2_X1 U18466 ( .A1(n19053), .A2(n15959), .ZN(n15210) );
  OAI211_X1 U18467 ( .C1(n19058), .C2(n15211), .A(n15210), .B(n15209), .ZN(
        n15213) );
  AOI211_X1 U18468 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15214), .A(
        n15213), .B(n15212), .ZN(n15217) );
  NAND3_X1 U18469 ( .A1(n12511), .A2(n19063), .A3(n15215), .ZN(n15216) );
  OAI211_X1 U18470 ( .C1(n15218), .C2(n16191), .A(n15217), .B(n15216), .ZN(
        P2_U3019) );
  INV_X1 U18471 ( .A(n16130), .ZN(n15224) );
  XNOR2_X1 U18472 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15223) );
  NAND2_X1 U18473 ( .A1(n16199), .A2(n15980), .ZN(n15220) );
  OAI211_X1 U18474 ( .C1(n15977), .C2(n15384), .A(n15220), .B(n15219), .ZN(
        n15221) );
  AOI21_X1 U18475 ( .B1(n16128), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15221), .ZN(n15222) );
  OAI21_X1 U18476 ( .B1(n15224), .B2(n15223), .A(n15222), .ZN(n15225) );
  AOI21_X1 U18477 ( .B1(n15226), .B2(n19063), .A(n15225), .ZN(n15227) );
  OAI21_X1 U18478 ( .B1(n15228), .B2(n16191), .A(n15227), .ZN(P2_U3020) );
  INV_X1 U18479 ( .A(n15230), .ZN(n15232) );
  NOR2_X1 U18480 ( .A1(n15232), .A2(n15231), .ZN(n15233) );
  XNOR2_X1 U18481 ( .A(n9612), .B(n15233), .ZN(n16017) );
  AOI21_X1 U18482 ( .B1(n13196), .B2(n15094), .A(n15077), .ZN(n16013) );
  NAND2_X1 U18483 ( .A1(n15234), .A2(n13196), .ZN(n15239) );
  NOR2_X1 U18484 ( .A1(n12978), .A2(n18920), .ZN(n15237) );
  NOR2_X1 U18485 ( .A1(n19058), .A2(n15235), .ZN(n15236) );
  AOI211_X1 U18486 ( .C1(n16014), .C2(n19053), .A(n15237), .B(n15236), .ZN(
        n15238) );
  OAI211_X1 U18487 ( .C1(n15240), .C2(n13196), .A(n15239), .B(n15238), .ZN(
        n15241) );
  AOI21_X1 U18488 ( .B1(n16013), .B2(n19063), .A(n15241), .ZN(n15242) );
  OAI21_X1 U18489 ( .B1(n16017), .B2(n16191), .A(n15242), .ZN(P2_U3022) );
  NAND2_X1 U18490 ( .A1(n15244), .A2(n15243), .ZN(n15247) );
  INV_X1 U18491 ( .A(n15245), .ZN(n15246) );
  NAND2_X1 U18492 ( .A1(n15247), .A2(n15246), .ZN(n16026) );
  NAND2_X1 U18493 ( .A1(n15390), .A2(n15248), .ZN(n15249) );
  NAND2_X1 U18494 ( .A1(n15374), .A2(n15249), .ZN(n16142) );
  NAND2_X1 U18495 ( .A1(n16199), .A2(n15530), .ZN(n15251) );
  NAND2_X1 U18496 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19040), .ZN(n15250) );
  OAI211_X1 U18497 ( .C1(n15252), .C2(n15384), .A(n15251), .B(n15250), .ZN(
        n15254) );
  NOR2_X1 U18498 ( .A1(n16139), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15253) );
  AOI211_X1 U18499 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n16142), .A(
        n15254), .B(n15253), .ZN(n15259) );
  NAND2_X1 U18500 ( .A1(n15256), .A2(n15255), .ZN(n15257) );
  XNOR2_X1 U18501 ( .A(n15086), .B(n15257), .ZN(n16022) );
  NAND2_X1 U18502 ( .A1(n16022), .A2(n19064), .ZN(n15258) );
  OAI211_X1 U18503 ( .C1(n16026), .C2(n16207), .A(n15259), .B(n15258), .ZN(
        P2_U3024) );
  NAND3_X1 U18504 ( .A1(n15260), .A2(n16172), .A3(n12364), .ZN(n15266) );
  NAND2_X1 U18505 ( .A1(n16199), .A2(n15261), .ZN(n15264) );
  NAND2_X1 U18506 ( .A1(n19053), .A2(n15262), .ZN(n15263) );
  NAND4_X1 U18507 ( .A1(n15266), .A2(n15265), .A3(n15264), .A4(n15263), .ZN(
        n15269) );
  NOR2_X1 U18508 ( .A1(n15267), .A2(n16207), .ZN(n15268) );
  AOI211_X1 U18509 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n16142), .A(
        n15269), .B(n15268), .ZN(n15270) );
  OAI21_X1 U18510 ( .B1(n15271), .B2(n16191), .A(n15270), .ZN(P2_U3025) );
  INV_X1 U18511 ( .A(n15272), .ZN(n16173) );
  OAI21_X1 U18512 ( .B1(n15274), .B2(n12315), .A(n15273), .ZN(n16182) );
  OAI21_X1 U18513 ( .B1(n16173), .B2(n15277), .A(n16182), .ZN(n16160) );
  NAND3_X1 U18514 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15275) );
  AND2_X1 U18515 ( .A1(n15390), .A2(n15275), .ZN(n15276) );
  NOR2_X1 U18516 ( .A1(n16160), .A2(n15276), .ZN(n15332) );
  OAI21_X1 U18517 ( .B1(n15294), .B2(n15277), .A(n15332), .ZN(n15296) );
  AND2_X1 U18518 ( .A1(n15390), .A2(n20842), .ZN(n15278) );
  NOR2_X1 U18519 ( .A1(n15296), .A2(n15278), .ZN(n16150) );
  NAND4_X1 U18520 ( .A1(n15293), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15294), .A4(n16172), .ZN(n16152) );
  INV_X1 U18521 ( .A(n16152), .ZN(n15285) );
  XNOR2_X1 U18522 ( .A(n15287), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15284) );
  NAND2_X1 U18523 ( .A1(n16199), .A2(n15279), .ZN(n15281) );
  OAI211_X1 U18524 ( .C1(n15282), .C2(n15384), .A(n15281), .B(n15280), .ZN(
        n15283) );
  AOI21_X1 U18525 ( .B1(n15285), .B2(n15284), .A(n15283), .ZN(n15286) );
  OAI21_X1 U18526 ( .B1(n16150), .B2(n15287), .A(n15286), .ZN(n15288) );
  AOI21_X1 U18527 ( .B1(n15289), .B2(n19063), .A(n15288), .ZN(n15290) );
  OAI21_X1 U18528 ( .B1(n16191), .B2(n15291), .A(n15290), .ZN(P2_U3026) );
  INV_X1 U18529 ( .A(n15292), .ZN(n15302) );
  NAND2_X1 U18530 ( .A1(n15293), .A2(n16172), .ZN(n15309) );
  INV_X1 U18531 ( .A(n15309), .ZN(n15335) );
  AND2_X1 U18532 ( .A1(n15294), .A2(n15335), .ZN(n15297) );
  NOR2_X1 U18533 ( .A1(n12964), .A2(n18920), .ZN(n15295) );
  AOI221_X1 U18534 ( .B1(n15297), .B2(n20842), .C1(n15296), .C2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(n15295), .ZN(n15301) );
  OAI22_X1 U18535 ( .A1(n19058), .A2(n18812), .B1(n15384), .B2(n18813), .ZN(
        n15298) );
  AOI21_X1 U18536 ( .B1(n19063), .B2(n15299), .A(n15298), .ZN(n15300) );
  OAI211_X1 U18537 ( .C1(n15302), .C2(n16191), .A(n15301), .B(n15300), .ZN(
        P2_U3028) );
  OAI21_X1 U18538 ( .B1(n15304), .B2(n19063), .A(n15303), .ZN(n15305) );
  OAI211_X1 U18539 ( .C1(n15306), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15332), .B(n15305), .ZN(n15323) );
  AOI21_X1 U18540 ( .B1(n15307), .B2(n15390), .A(n15323), .ZN(n15315) );
  NAND2_X1 U18541 ( .A1(n15308), .A2(n19064), .ZN(n15314) );
  OAI22_X1 U18542 ( .A1(n12373), .A2(n15309), .B1(n16207), .B2(n16032), .ZN(
        n15319) );
  NAND3_X1 U18543 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15135), .A3(
        n15319), .ZN(n15310) );
  OAI21_X1 U18544 ( .B1(n18920), .B2(n19680), .A(n15310), .ZN(n15312) );
  NOR2_X1 U18545 ( .A1(n19058), .A2(n18829), .ZN(n15311) );
  AOI211_X1 U18546 ( .C1(n19053), .C2(n18825), .A(n15312), .B(n15311), .ZN(
        n15313) );
  OAI211_X1 U18547 ( .C1(n15135), .C2(n15315), .A(n15314), .B(n15313), .ZN(
        P2_U3029) );
  OAI21_X1 U18548 ( .B1(n15318), .B2(n15317), .A(n15316), .ZN(n16035) );
  NAND2_X1 U18549 ( .A1(n15319), .A2(n15307), .ZN(n15325) );
  AOI22_X1 U18550 ( .A1(n16199), .A2(n15320), .B1(n19040), .B2(
        P2_REIP_REG_16__SCAN_IN), .ZN(n15321) );
  OAI21_X1 U18551 ( .B1(n15384), .B2(n16033), .A(n15321), .ZN(n15322) );
  AOI21_X1 U18552 ( .B1(n15323), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15322), .ZN(n15324) );
  OAI211_X1 U18553 ( .C1(n16191), .C2(n16035), .A(n15325), .B(n15324), .ZN(
        P2_U3030) );
  NAND2_X1 U18554 ( .A1(n15327), .A2(n15326), .ZN(n15330) );
  NAND2_X1 U18555 ( .A1(n15328), .A2(n16048), .ZN(n15329) );
  XOR2_X1 U18556 ( .A(n15330), .B(n15329), .Z(n16041) );
  OAI21_X1 U18557 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15331), .A(
        n16032), .ZN(n16042) );
  INV_X1 U18558 ( .A(n16042), .ZN(n15340) );
  INV_X1 U18559 ( .A(n15332), .ZN(n15334) );
  NOR2_X1 U18560 ( .A1(n12959), .A2(n18920), .ZN(n15333) );
  AOI221_X1 U18561 ( .B1(n15335), .B2(n12373), .C1(n15334), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n15333), .ZN(n15338) );
  INV_X1 U18562 ( .A(n15336), .ZN(n18837) );
  NAND2_X1 U18563 ( .A1(n19053), .A2(n18837), .ZN(n15337) );
  OAI211_X1 U18564 ( .C1(n19058), .C2(n18841), .A(n15338), .B(n15337), .ZN(
        n15339) );
  AOI21_X1 U18565 ( .B1(n15340), .B2(n19063), .A(n15339), .ZN(n15341) );
  OAI21_X1 U18566 ( .B1(n16041), .B2(n16191), .A(n15341), .ZN(P2_U3031) );
  NAND2_X1 U18567 ( .A1(n15342), .A2(n16172), .ZN(n16159) );
  NOR2_X1 U18568 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16159), .ZN(
        n15358) );
  NOR2_X1 U18569 ( .A1(n15358), .A2(n16160), .ZN(n15349) );
  INV_X1 U18570 ( .A(n18857), .ZN(n15345) );
  NOR2_X1 U18571 ( .A1(n15152), .A2(n18920), .ZN(n15344) );
  NOR2_X1 U18572 ( .A1(n19058), .A2(n18868), .ZN(n15343) );
  AOI211_X1 U18573 ( .C1(n15345), .C2(n19053), .A(n15344), .B(n15343), .ZN(
        n15348) );
  NOR2_X1 U18574 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16159), .ZN(
        n15346) );
  NAND2_X1 U18575 ( .A1(n15346), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15347) );
  OAI211_X1 U18576 ( .C1(n15349), .C2(n12377), .A(n15348), .B(n15347), .ZN(
        n15350) );
  AOI21_X1 U18577 ( .B1(n15351), .B2(n19064), .A(n15350), .ZN(n15352) );
  OAI21_X1 U18578 ( .B1(n15353), .B2(n16207), .A(n15352), .ZN(P2_U3033) );
  OAI21_X1 U18579 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15355), .A(
        n15354), .ZN(n15356) );
  INV_X1 U18580 ( .A(n15356), .ZN(n16055) );
  NAND2_X1 U18581 ( .A1(n16055), .A2(n19063), .ZN(n15368) );
  NOR2_X1 U18582 ( .A1(n12945), .A2(n18920), .ZN(n15357) );
  AOI211_X1 U18583 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16160), .A(
        n15358), .B(n15357), .ZN(n15367) );
  XNOR2_X1 U18584 ( .A(n15360), .B(n15359), .ZN(n18972) );
  OAI22_X1 U18585 ( .A1(n19058), .A2(n18972), .B1(n15384), .B2(n18874), .ZN(
        n15361) );
  INV_X1 U18586 ( .A(n15361), .ZN(n15366) );
  XNOR2_X1 U18587 ( .A(n15363), .B(n12325), .ZN(n15364) );
  XNOR2_X1 U18588 ( .A(n15362), .B(n15364), .ZN(n16057) );
  NAND2_X1 U18589 ( .A1(n16057), .A2(n19064), .ZN(n15365) );
  NAND4_X1 U18590 ( .A1(n15368), .A2(n15367), .A3(n15366), .A4(n15365), .ZN(
        P2_U3034) );
  OAI21_X1 U18591 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15144), .A(
        n16082), .ZN(n16088) );
  NAND2_X1 U18592 ( .A1(n16061), .A2(n15369), .ZN(n15373) );
  INV_X1 U18593 ( .A(n15370), .ZN(n16075) );
  OR2_X1 U18594 ( .A1(n16075), .A2(n15371), .ZN(n15372) );
  XNOR2_X1 U18595 ( .A(n15373), .B(n15372), .ZN(n16087) );
  INV_X1 U18596 ( .A(n15374), .ZN(n15376) );
  NOR2_X1 U18597 ( .A1(n12936), .A2(n18920), .ZN(n15375) );
  AOI221_X1 U18598 ( .B1(n15376), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n16172), .C2(n12315), .A(n15375), .ZN(n15380) );
  INV_X1 U18599 ( .A(n18901), .ZN(n15377) );
  OAI22_X1 U18600 ( .A1(n19058), .A2(n18905), .B1(n15384), .B2(n15377), .ZN(
        n15378) );
  INV_X1 U18601 ( .A(n15378), .ZN(n15379) );
  OAI211_X1 U18602 ( .C1(n16087), .C2(n16191), .A(n15380), .B(n15379), .ZN(
        n15381) );
  INV_X1 U18603 ( .A(n15381), .ZN(n15382) );
  OAI21_X1 U18604 ( .B1(n16088), .B2(n16207), .A(n15382), .ZN(P2_U3037) );
  NAND2_X1 U18605 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19040), .ZN(n15383) );
  OAI221_X1 U18606 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16195), .C1(
        n12304), .C2(n16196), .A(n15383), .ZN(n15386) );
  OAI22_X1 U18607 ( .A1(n19058), .A2(n18914), .B1(n15384), .B2(n18913), .ZN(
        n15385) );
  AOI211_X1 U18608 ( .C1(n15387), .C2(n19064), .A(n15386), .B(n15385), .ZN(
        n15388) );
  OAI21_X1 U18609 ( .B1(n9930), .B2(n16207), .A(n15388), .ZN(P2_U3039) );
  OAI211_X1 U18610 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15390), .B(n15389), .ZN(n15399) );
  AOI22_X1 U18611 ( .A1(n19063), .A2(n15391), .B1(n16199), .B2(n19749), .ZN(
        n15398) );
  AOI21_X1 U18612 ( .B1(n19053), .B2(n15393), .A(n15392), .ZN(n15397) );
  AOI22_X1 U18613 ( .A1(n19064), .A2(n15395), .B1(n15394), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15396) );
  NAND4_X1 U18614 ( .A1(n15399), .A2(n15398), .A3(n15397), .A4(n15396), .ZN(
        P2_U3045) );
  MUX2_X1 U18615 ( .A(n15400), .B(n13210), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15401) );
  AOI21_X1 U18616 ( .B1(n15402), .B2(n16243), .A(n15401), .ZN(n16246) );
  OAI222_X1 U18617 ( .A1(n19719), .A2(n10139), .B1(n19726), .B2(n16246), .C1(
        n15404), .C2(n15403), .ZN(n15405) );
  MUX2_X1 U18618 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15405), .S(
        n19714), .Z(P2_U3601) );
  OAI22_X1 U18619 ( .A1(n17061), .A2(n17021), .B1(n9644), .B2(n17013), .ZN(
        n15415) );
  AOI22_X1 U18620 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U18621 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15412) );
  OAI22_X1 U18622 ( .A1(n16957), .A2(n17010), .B1(n9598), .B2(n16905), .ZN(
        n15410) );
  AOI22_X1 U18623 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U18624 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U18625 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15406) );
  NAND3_X1 U18626 ( .A1(n15408), .A2(n15407), .A3(n15406), .ZN(n15409) );
  AOI211_X1 U18627 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15410), .B(n15409), .ZN(n15411) );
  NAND3_X1 U18628 ( .A1(n15413), .A2(n15412), .A3(n15411), .ZN(n15414) );
  AOI211_X1 U18629 ( .C1(n17030), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n15415), .B(n15414), .ZN(n16844) );
  AOI22_X1 U18630 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15416) );
  OAI21_X1 U18631 ( .B1(n10714), .B2(n17046), .A(n15416), .ZN(n15426) );
  AOI22_X1 U18632 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16828), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15424) );
  OAI22_X1 U18633 ( .A1(n10692), .A2(n17044), .B1(n17011), .B2(n15417), .ZN(
        n15422) );
  AOI22_X1 U18634 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15420) );
  AOI22_X1 U18635 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U18636 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15418) );
  NAND3_X1 U18637 ( .A1(n15420), .A2(n15419), .A3(n15418), .ZN(n15421) );
  AOI211_X1 U18638 ( .C1(n9595), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n15422), .B(n15421), .ZN(n15423) );
  OAI211_X1 U18639 ( .C1(n16957), .C2(n16935), .A(n15424), .B(n15423), .ZN(
        n15425) );
  AOI211_X1 U18640 ( .C1(n9591), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15426), .B(n15425), .ZN(n16857) );
  AOI22_X1 U18641 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15427) );
  OAI21_X1 U18642 ( .B1(n15507), .B2(n17100), .A(n15427), .ZN(n15437) );
  AOI22_X1 U18643 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10657), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15435) );
  AOI22_X1 U18644 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15428) );
  OAI21_X1 U18645 ( .B1(n10692), .B2(n17086), .A(n15428), .ZN(n15433) );
  AOI22_X1 U18646 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U18647 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15429) );
  OAI211_X1 U18648 ( .C1(n16821), .C2(n15431), .A(n15430), .B(n15429), .ZN(
        n15432) );
  AOI211_X1 U18649 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n15433), .B(n15432), .ZN(n15434) );
  OAI211_X1 U18650 ( .C1(n17061), .C2(n17084), .A(n15435), .B(n15434), .ZN(
        n15436) );
  AOI211_X1 U18651 ( .C1(n9592), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n15437), .B(n15436), .ZN(n16867) );
  AOI22_X1 U18652 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15438) );
  OAI21_X1 U18653 ( .B1(n17087), .B2(n20927), .A(n15438), .ZN(n15447) );
  INV_X1 U18654 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U18655 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15445) );
  OAI22_X1 U18656 ( .A1(n9586), .A2(n16987), .B1(n16957), .B2(n16982), .ZN(
        n15443) );
  AOI22_X1 U18657 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15441) );
  AOI22_X1 U18658 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15440) );
  AOI22_X1 U18659 ( .A1(n16828), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15439) );
  NAND3_X1 U18660 ( .A1(n15441), .A2(n15440), .A3(n15439), .ZN(n15442) );
  AOI211_X1 U18661 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n15443), .B(n15442), .ZN(n15444) );
  OAI211_X1 U18662 ( .C1(n9598), .C2(n16977), .A(n15445), .B(n15444), .ZN(
        n15446) );
  AOI211_X1 U18663 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n15447), .B(n15446), .ZN(n16868) );
  NOR2_X1 U18664 ( .A1(n16867), .A2(n16868), .ZN(n16866) );
  AOI22_X1 U18665 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15458) );
  AOI22_X1 U18666 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U18667 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16828), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15456) );
  OAI22_X1 U18668 ( .A1(n10692), .A2(n15448), .B1(n16821), .B2(n17073), .ZN(
        n15454) );
  AOI22_X1 U18669 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U18670 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U18671 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10721), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15450) );
  NAND2_X1 U18672 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n15449) );
  NAND4_X1 U18673 ( .A1(n15452), .A2(n15451), .A3(n15450), .A4(n15449), .ZN(
        n15453) );
  AOI211_X1 U18674 ( .C1(n17082), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n15454), .B(n15453), .ZN(n15455) );
  NAND4_X1 U18675 ( .A1(n15458), .A2(n15457), .A3(n15456), .A4(n15455), .ZN(
        n16862) );
  NAND2_X1 U18676 ( .A1(n16866), .A2(n16862), .ZN(n16861) );
  NOR2_X1 U18677 ( .A1(n16857), .A2(n16861), .ZN(n16856) );
  AOI22_X1 U18678 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U18679 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15469) );
  AOI22_X1 U18680 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15468) );
  OAI22_X1 U18681 ( .A1(n10692), .A2(n15460), .B1(n10732), .B2(n15459), .ZN(
        n15466) );
  AOI22_X1 U18682 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15464) );
  AOI22_X1 U18683 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15463) );
  AOI22_X1 U18684 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U18685 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n15461) );
  NAND4_X1 U18686 ( .A1(n15464), .A2(n15463), .A3(n15462), .A4(n15461), .ZN(
        n15465) );
  AOI211_X1 U18687 ( .C1(n9599), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n15466), .B(n15465), .ZN(n15467) );
  NAND4_X1 U18688 ( .A1(n15470), .A2(n15469), .A3(n15468), .A4(n15467), .ZN(
        n16849) );
  NAND2_X1 U18689 ( .A1(n16856), .A2(n16849), .ZN(n16848) );
  NOR2_X1 U18690 ( .A1(n16844), .A2(n16848), .ZN(n16843) );
  AOI22_X1 U18691 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U18692 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15482) );
  AOI22_X1 U18693 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16828), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15481) );
  OAI22_X1 U18694 ( .A1(n15507), .A2(n16889), .B1(n17061), .B2(n15472), .ZN(
        n15479) );
  AOI22_X1 U18695 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U18696 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U18697 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U18698 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n15474) );
  NAND4_X1 U18699 ( .A1(n15477), .A2(n15476), .A3(n15475), .A4(n15474), .ZN(
        n15478) );
  AOI211_X1 U18700 ( .C1(n10657), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n15479), .B(n15478), .ZN(n15480) );
  NAND4_X1 U18701 ( .A1(n15483), .A2(n15482), .A3(n15481), .A4(n15480), .ZN(
        n15484) );
  NAND2_X1 U18702 ( .A1(n16843), .A2(n15484), .ZN(n16838) );
  OAI21_X1 U18703 ( .B1(n16843), .B2(n15484), .A(n16838), .ZN(n17158) );
  NAND2_X1 U18704 ( .A1(n18134), .A2(n18119), .ZN(n15485) );
  OAI22_X1 U18705 ( .A1(n15488), .A2(n15487), .B1(n15486), .B2(n15485), .ZN(
        n15608) );
  NAND4_X1 U18706 ( .A1(n18757), .A2(n18749), .A3(n10901), .A4(n15608), .ZN(
        n17134) );
  INV_X1 U18707 ( .A(n17134), .ZN(n17131) );
  INV_X1 U18708 ( .A(n18134), .ZN(n17259) );
  AND2_X1 U18709 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16836) );
  NAND2_X1 U18710 ( .A1(n18134), .A2(n17131), .ZN(n17136) );
  INV_X1 U18711 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17116) );
  NAND2_X1 U18712 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16785) );
  INV_X1 U18713 ( .A(n16785), .ZN(n17125) );
  NAND2_X1 U18714 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17125), .ZN(n17115) );
  OR3_X1 U18715 ( .A1(n17116), .A2(n16758), .A3(n17115), .ZN(n17117) );
  INV_X1 U18716 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16704) );
  NOR2_X1 U18717 ( .A1(n17105), .A2(n16704), .ZN(n15493) );
  NAND3_X1 U18718 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n16990) );
  NAND4_X1 U18719 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n15494) );
  NOR4_X1 U18720 ( .A1(n16972), .A2(n16729), .A3(n16990), .A4(n15494), .ZN(
        n15489) );
  NAND4_X1 U18721 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17111), .A3(n15493), 
        .A4(n15489), .ZN(n16973) );
  NAND2_X1 U18722 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16961), .ZN(n16944) );
  NAND2_X1 U18723 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16901), .ZN(n16885) );
  NOR2_X1 U18724 ( .A1(n15490), .A2(n16885), .ZN(n16865) );
  NAND2_X1 U18725 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16871), .ZN(n16851) );
  NAND3_X1 U18726 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16864), .ZN(n16847) );
  NAND2_X1 U18727 ( .A1(n17129), .A2(n16847), .ZN(n16850) );
  OAI21_X1 U18728 ( .B1(n16836), .B2(n17136), .A(n16850), .ZN(n16840) );
  NOR3_X1 U18729 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16846), .A3(n16847), .ZN(
        n15491) );
  AOI21_X1 U18730 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16840), .A(n15491), .ZN(
        n15492) );
  OAI21_X1 U18731 ( .B1(n17158), .B2(n17121), .A(n15492), .ZN(P3_U2675) );
  NAND2_X1 U18732 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17111), .ZN(n17110) );
  INV_X1 U18733 ( .A(n17110), .ZN(n17107) );
  NAND2_X1 U18734 ( .A1(n18134), .A2(n17081), .ZN(n17102) );
  NOR2_X1 U18735 ( .A1(n15494), .A2(n17102), .ZN(n17025) );
  NAND2_X1 U18736 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17025), .ZN(n17024) );
  INV_X1 U18737 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n15495) );
  AND2_X1 U18738 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17081), .ZN(n17079) );
  NAND2_X1 U18739 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17079), .ZN(n17078) );
  INV_X1 U18740 ( .A(n17078), .ZN(n17057) );
  NAND3_X1 U18741 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n17057), .ZN(n17040) );
  OAI21_X1 U18742 ( .B1(n15495), .B2(n17040), .A(n17121), .ZN(n15509) );
  INV_X1 U18743 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U18744 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15505) );
  AOI22_X1 U18745 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U18746 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15496) );
  OAI211_X1 U18747 ( .C1(n10732), .C2(n17113), .A(n15497), .B(n15496), .ZN(
        n15503) );
  AOI22_X1 U18748 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15501) );
  AOI22_X1 U18749 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18750 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15499) );
  NAND2_X1 U18751 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n15498) );
  NAND4_X1 U18752 ( .A1(n15501), .A2(n15500), .A3(n15499), .A4(n15498), .ZN(
        n15502) );
  AOI211_X1 U18753 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15503), .B(n15502), .ZN(n15504) );
  OAI211_X1 U18754 ( .C1(n15507), .C2(n15506), .A(n15505), .B(n15504), .ZN(
        n17234) );
  NAND2_X1 U18755 ( .A1(n17114), .A2(n17234), .ZN(n15508) );
  OAI221_X1 U18756 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17024), .C1(n20860), 
        .C2(n15509), .A(n15508), .ZN(P3_U2690) );
  NAND2_X1 U18757 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18246) );
  AOI221_X1 U18758 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18246), .C1(n15511), 
        .C2(n18246), .A(n15510), .ZN(n18100) );
  NOR2_X1 U18759 ( .A1(n15512), .A2(n18576), .ZN(n15513) );
  OAI21_X1 U18760 ( .B1(n15513), .B2(n18441), .A(n18101), .ZN(n18098) );
  AOI22_X1 U18761 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18100), .B1(
        n18098), .B2(n18411), .ZN(P3_U2865) );
  NAND2_X1 U18762 ( .A1(n15515), .A2(n15514), .ZN(n15516) );
  NOR2_X1 U18763 ( .A1(n18090), .A2(n18539), .ZN(n18089) );
  INV_X1 U18764 ( .A(n16302), .ZN(n16318) );
  NOR3_X1 U18765 ( .A1(n16307), .A2(n18083), .A3(n15517), .ZN(n15518) );
  AOI21_X1 U18766 ( .B1(n18089), .B2(n16318), .A(n15518), .ZN(n15589) );
  INV_X1 U18767 ( .A(n15589), .ZN(n15525) );
  INV_X1 U18768 ( .A(n17811), .ZN(n18004) );
  NAND2_X1 U18769 ( .A1(n18074), .A2(n18004), .ZN(n18076) );
  OAI22_X1 U18770 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18076), .B1(
        n17892), .B2(n15519), .ZN(n15524) );
  NOR2_X1 U18771 ( .A1(n17786), .A2(n15520), .ZN(n16326) );
  INV_X1 U18772 ( .A(n18000), .ZN(n17968) );
  OAI22_X1 U18773 ( .A1(n17968), .A2(n17416), .B1(n18539), .B2(n17772), .ZN(
        n15521) );
  OAI21_X1 U18774 ( .B1(n16326), .B2(n15521), .A(n18074), .ZN(n15594) );
  NOR3_X1 U18775 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15522), .A3(
        n15594), .ZN(n15523) );
  AOI221_X1 U18776 ( .B1(n15525), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), 
        .C1(n15524), .C2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n15523), .ZN(
        n15526) );
  NAND2_X1 U18777 ( .A1(n18050), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16313) );
  OAI211_X1 U18778 ( .C1(n16322), .C2(n17960), .A(n15526), .B(n16313), .ZN(
        P3_U2833) );
  AOI22_X1 U18779 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n9691), .ZN(n15538) );
  INV_X1 U18780 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15527) );
  OAI22_X1 U18781 ( .A1(n15528), .A2(n18924), .B1(n18952), .B2(n15527), .ZN(
        n15529) );
  INV_X1 U18782 ( .A(n15529), .ZN(n15537) );
  AOI22_X1 U18783 ( .A1(n16023), .A2(n18932), .B1(n18958), .B2(n15530), .ZN(
        n15536) );
  AOI21_X1 U18784 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(n15534) );
  NAND2_X1 U18785 ( .A1(n18933), .A2(n15534), .ZN(n15535) );
  NAND4_X1 U18786 ( .A1(n15538), .A2(n15537), .A3(n15536), .A4(n15535), .ZN(
        P2_U2833) );
  NOR3_X1 U18787 ( .A1(n15540), .A2(n15539), .A3(n20521), .ZN(n15550) );
  INV_X1 U18788 ( .A(n20315), .ZN(n20565) );
  INV_X1 U18789 ( .A(n15541), .ZN(n20775) );
  INV_X1 U18790 ( .A(n13824), .ZN(n20776) );
  NAND3_X1 U18791 ( .A1(n15542), .A2(n20775), .A3(n20776), .ZN(n15543) );
  OAI21_X1 U18792 ( .B1(n15544), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15543), .ZN(n15545) );
  AOI21_X1 U18793 ( .B1(n20565), .B2(n15546), .A(n15545), .ZN(n20773) );
  AOI21_X1 U18794 ( .B1(n15550), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n20773), .ZN(n15547) );
  NAND2_X1 U18795 ( .A1(n15548), .A2(n15547), .ZN(n15549) );
  OAI21_X1 U18796 ( .B1(n15550), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15549), .ZN(n15551) );
  AOI222_X1 U18797 ( .A1(n15552), .A2(n20394), .B1(n15552), .B2(n15551), .C1(
        n20394), .C2(n15551), .ZN(n15554) );
  AOI21_X1 U18798 ( .B1(n15554), .B2(n15553), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15556) );
  NOR2_X1 U18799 ( .A1(n15554), .A2(n15553), .ZN(n15555) );
  OAI21_X1 U18800 ( .B1(n15556), .B2(n15555), .A(n19993), .ZN(n15564) );
  OAI21_X1 U18801 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15557), .ZN(n15559) );
  AND4_X1 U18802 ( .A1(n15561), .A2(n15560), .A3(n15559), .A4(n15558), .ZN(
        n15563) );
  NAND3_X1 U18803 ( .A1(n15564), .A2(n15563), .A3(n15562), .ZN(n15569) );
  OAI21_X1 U18804 ( .B1(n15565), .B2(n20797), .A(n20687), .ZN(n15566) );
  OAI21_X1 U18805 ( .B1(n15568), .B2(n15567), .A(n15566), .ZN(n15942) );
  AOI221_X1 U18806 ( .B1(n19998), .B2(n15944), .C1(n15569), .C2(n15944), .A(
        n15942), .ZN(n15571) );
  NOR2_X1 U18807 ( .A1(n15571), .A2(n19998), .ZN(n20690) );
  OAI211_X1 U18808 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20797), .A(n20690), 
        .B(n15573), .ZN(n15943) );
  AOI21_X1 U18809 ( .B1(n15570), .B2(n15569), .A(n15943), .ZN(n15577) );
  INV_X1 U18810 ( .A(n15571), .ZN(n15572) );
  OAI21_X1 U18811 ( .B1(n15574), .B2(n15573), .A(n15572), .ZN(n15575) );
  AOI22_X1 U18812 ( .A1(n15577), .A2(n15576), .B1(n19998), .B2(n15575), .ZN(
        P1_U3161) );
  AOI22_X1 U18813 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15578), .B1(
        n19940), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15584) );
  INV_X1 U18814 ( .A(n15579), .ZN(n15580) );
  AOI22_X1 U18815 ( .A1(n15581), .A2(n9588), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15580), .ZN(n15582) );
  XNOR2_X1 U18816 ( .A(n15582), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15746) );
  AOI22_X1 U18817 ( .A1(n15746), .A2(n19970), .B1(n19967), .B2(n15649), .ZN(
        n15583) );
  OAI211_X1 U18818 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15585), .A(
        n15584), .B(n15583), .ZN(P1_U3010) );
  INV_X1 U18819 ( .A(n18076), .ZN(n15588) );
  AOI22_X1 U18820 ( .A1(n15588), .A2(n15587), .B1(n9600), .B2(n15586), .ZN(
        n16323) );
  AOI21_X1 U18821 ( .B1(n16323), .B2(n15589), .A(n20944), .ZN(n15590) );
  AOI21_X1 U18822 ( .B1(n18009), .B2(n15591), .A(n15590), .ZN(n15593) );
  OAI211_X1 U18823 ( .C1(n15595), .C2(n15594), .A(n15593), .B(n15592), .ZN(
        P3_U2832) );
  INV_X1 U18824 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20704) );
  INV_X1 U18825 ( .A(HOLD), .ZN(n20692) );
  NOR2_X1 U18826 ( .A1(n20704), .A2(n20692), .ZN(n15599) );
  AOI22_X1 U18827 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15598) );
  NAND2_X1 U18828 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20691), .ZN(n15596) );
  OAI211_X1 U18829 ( .C1(n15599), .C2(n15598), .A(n15597), .B(n15596), .ZN(
        P1_U3195) );
  AND2_X1 U18830 ( .A1(n19920), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U18831 ( .A(n15600), .ZN(n19785) );
  NOR2_X1 U18832 ( .A1(n19785), .A2(n19780), .ZN(n19634) );
  NAND2_X1 U18833 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19780), .ZN(n19783) );
  INV_X1 U18834 ( .A(n19783), .ZN(n15601) );
  AOI22_X1 U18835 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19634), .B1(
        P2_STATEBS16_REG_SCAN_IN), .B2(n15601), .ZN(n15602) );
  AOI21_X1 U18836 ( .B1(n15602), .B2(n19784), .A(n15606), .ZN(P2_U3178) );
  NAND2_X1 U18837 ( .A1(n15603), .A2(n19783), .ZN(n19778) );
  NAND2_X1 U18838 ( .A1(n19778), .A2(n15604), .ZN(n15605) );
  AOI221_X1 U18839 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15606), .C1(n19766), .C2(
        n15606), .A(n19576), .ZN(n19758) );
  INV_X1 U18840 ( .A(n19758), .ZN(n19755) );
  NOR2_X1 U18841 ( .A1(n15607), .A2(n19755), .ZN(P2_U3047) );
  NAND3_X1 U18842 ( .A1(n16730), .A2(n17332), .A3(n15608), .ZN(n15609) );
  AND2_X4 U18843 ( .A1(n15611), .A2(n18757), .ZN(n17141) );
  NAND2_X1 U18844 ( .A1(n18134), .A2(n17141), .ZN(n17186) );
  INV_X1 U18845 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17364) );
  NAND2_X1 U18846 ( .A1(n15612), .A2(n17141), .ZN(n17283) );
  AOI22_X1 U18847 ( .A1(n17285), .A2(BUF2_REG_0__SCAN_IN), .B1(n17268), .B2(
        n17758), .ZN(n15614) );
  OAI221_X1 U18848 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17186), .C1(n17364), 
        .C2(n17141), .A(n15614), .ZN(P3_U2735) );
  AOI21_X1 U18849 ( .B1(n15642), .B2(n20743), .A(n15615), .ZN(n15628) );
  INV_X1 U18850 ( .A(n15735), .ZN(n15621) );
  NOR3_X1 U18851 ( .A1(n19877), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n15616), 
        .ZN(n15620) );
  INV_X1 U18852 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15618) );
  INV_X1 U18853 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15617) );
  OAI22_X1 U18854 ( .A1(n19833), .A2(n15618), .B1(n15617), .B2(n19855), .ZN(
        n15619) );
  AOI211_X1 U18855 ( .C1(n15621), .C2(n19883), .A(n15620), .B(n15619), .ZN(
        n15627) );
  NAND2_X1 U18856 ( .A1(n15623), .A2(n15622), .ZN(n15624) );
  AND2_X1 U18857 ( .A1(n15625), .A2(n15624), .ZN(n15814) );
  AOI22_X1 U18858 ( .A1(n15732), .A2(n19847), .B1(n19860), .B2(n15814), .ZN(
        n15626) );
  OAI211_X1 U18859 ( .C1(n15628), .C2(n20745), .A(n15627), .B(n15626), .ZN(
        P1_U2815) );
  NAND2_X1 U18860 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15629) );
  NOR3_X1 U18861 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15629), .A3(n15653), 
        .ZN(n15633) );
  OAI22_X1 U18862 ( .A1(n19833), .A2(n15631), .B1(n15630), .B2(n19855), .ZN(
        n15632) );
  AOI211_X1 U18863 ( .C1(n19883), .C2(n15634), .A(n15633), .B(n15632), .ZN(
        n15639) );
  NAND2_X1 U18864 ( .A1(n15635), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15644) );
  AOI21_X1 U18865 ( .B1(n15642), .B2(n15644), .A(n19880), .ZN(n15652) );
  OAI21_X1 U18866 ( .B1(n19877), .B2(P1_REIP_REG_21__SCAN_IN), .A(n15652), 
        .ZN(n15636) );
  AOI22_X1 U18867 ( .A1(n15637), .A2(n19847), .B1(P1_REIP_REG_22__SCAN_IN), 
        .B2(n15636), .ZN(n15638) );
  OAI211_X1 U18868 ( .C1(n19893), .C2(n15640), .A(n15639), .B(n15638), .ZN(
        P1_U2818) );
  INV_X1 U18869 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15641) );
  NOR2_X1 U18870 ( .A1(n19855), .A2(n15641), .ZN(n15646) );
  INV_X1 U18871 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20738) );
  NAND2_X1 U18872 ( .A1(n15642), .A2(n20738), .ZN(n15643) );
  OAI22_X1 U18873 ( .A1(n15644), .A2(n15643), .B1(n15652), .B2(n20738), .ZN(
        n15645) );
  NOR2_X1 U18874 ( .A1(n15646), .A2(n15645), .ZN(n15647) );
  OAI21_X1 U18875 ( .B1(n15749), .B2(n15712), .A(n15647), .ZN(n15648) );
  AOI21_X1 U18876 ( .B1(n19879), .B2(P1_EBX_REG_21__SCAN_IN), .A(n15648), .ZN(
        n15651) );
  AOI22_X1 U18877 ( .A1(n15745), .A2(n19847), .B1(n15649), .B2(n19860), .ZN(
        n15650) );
  NAND2_X1 U18878 ( .A1(n15651), .A2(n15650), .ZN(P1_U2819) );
  AOI21_X1 U18879 ( .B1(n14728), .B2(n15653), .A(n15652), .ZN(n15657) );
  AOI22_X1 U18880 ( .A1(n19884), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19883), .B2(n15750), .ZN(n15654) );
  OAI21_X1 U18881 ( .B1(n19833), .B2(n15655), .A(n15654), .ZN(n15656) );
  AOI211_X1 U18882 ( .C1(n15751), .C2(n19847), .A(n15657), .B(n15656), .ZN(
        n15658) );
  OAI21_X1 U18883 ( .B1(n19893), .B2(n15659), .A(n15658), .ZN(P1_U2820) );
  NAND3_X1 U18884 ( .A1(n15660), .A2(n15701), .A3(n14744), .ZN(n15665) );
  INV_X1 U18885 ( .A(n15759), .ZN(n15663) );
  INV_X1 U18886 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15661) );
  NOR2_X1 U18887 ( .A1(n19855), .A2(n15661), .ZN(n15662) );
  AOI211_X1 U18888 ( .C1(n19883), .C2(n15663), .A(n19868), .B(n15662), .ZN(
        n15664) );
  OAI211_X1 U18889 ( .C1(n20829), .C2(n19833), .A(n15665), .B(n15664), .ZN(
        n15666) );
  AOI21_X1 U18890 ( .B1(n15755), .B2(n19847), .A(n15666), .ZN(n15670) );
  OAI21_X1 U18891 ( .B1(n15668), .B2(n15667), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15669) );
  OAI211_X1 U18892 ( .C1(n15671), .C2(n19893), .A(n15670), .B(n15669), .ZN(
        P1_U2821) );
  OAI22_X1 U18893 ( .A1(n15673), .A2(n19893), .B1(n15672), .B2(n19833), .ZN(
        n15674) );
  AOI211_X1 U18894 ( .C1(n19884), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19868), .B(n15674), .ZN(n15679) );
  INV_X1 U18895 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20729) );
  NOR3_X1 U18896 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n20729), .A3(n15675), 
        .ZN(n15677) );
  OR2_X1 U18897 ( .A1(n15675), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15689) );
  AOI21_X1 U18898 ( .B1(n15700), .B2(n15689), .A(n14773), .ZN(n15676) );
  AOI211_X1 U18899 ( .C1(n15767), .C2(n19847), .A(n15677), .B(n15676), .ZN(
        n15678) );
  OAI211_X1 U18900 ( .C1(n15765), .C2(n15712), .A(n15679), .B(n15678), .ZN(
        P1_U2824) );
  INV_X1 U18901 ( .A(n15680), .ZN(n15776) );
  NOR2_X1 U18902 ( .A1(n15682), .A2(n15681), .ZN(n15683) );
  OR2_X1 U18903 ( .A1(n15684), .A2(n15683), .ZN(n15720) );
  INV_X1 U18904 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15722) );
  AOI21_X1 U18905 ( .B1(n19884), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n19868), .ZN(n15685) );
  OAI21_X1 U18906 ( .B1(n19833), .B2(n15722), .A(n15685), .ZN(n15686) );
  AOI21_X1 U18907 ( .B1(n19883), .B2(n15775), .A(n15686), .ZN(n15687) );
  OAI21_X1 U18908 ( .B1(n15720), .B2(n19893), .A(n15687), .ZN(n15688) );
  AOI21_X1 U18909 ( .B1(n15776), .B2(n19847), .A(n15688), .ZN(n15690) );
  OAI211_X1 U18910 ( .C1(n15700), .C2(n20729), .A(n15690), .B(n15689), .ZN(
        P1_U2825) );
  NOR2_X1 U18911 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15691), .ZN(n15699) );
  INV_X1 U18912 ( .A(n15692), .ZN(n15693) );
  AOI22_X1 U18913 ( .A1(n19879), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n15693), 
        .B2(n19883), .ZN(n15698) );
  AOI21_X1 U18914 ( .B1(n19884), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n19868), .ZN(n15694) );
  OAI21_X1 U18915 ( .B1(n15847), .B2(n19893), .A(n15694), .ZN(n15695) );
  AOI21_X1 U18916 ( .B1(n15696), .B2(n19847), .A(n15695), .ZN(n15697) );
  OAI211_X1 U18917 ( .C1(n15700), .C2(n15699), .A(n15698), .B(n15697), .ZN(
        P1_U2826) );
  AOI21_X1 U18918 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15701), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15706) );
  AOI22_X1 U18919 ( .A1(n15780), .A2(n19883), .B1(n19860), .B2(n15723), .ZN(
        n15705) );
  INV_X1 U18920 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15725) );
  OAI22_X1 U18921 ( .A1(n19833), .A2(n15725), .B1(n15702), .B2(n19855), .ZN(
        n15703) );
  AOI211_X1 U18922 ( .C1(n15779), .C2(n19847), .A(n19868), .B(n15703), .ZN(
        n15704) );
  OAI211_X1 U18923 ( .C1(n15707), .C2(n15706), .A(n15705), .B(n15704), .ZN(
        P1_U2828) );
  OAI21_X1 U18924 ( .B1(n15709), .B2(n15708), .A(n14123), .ZN(n15710) );
  INV_X1 U18925 ( .A(n15710), .ZN(n15865) );
  INV_X1 U18926 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15711) );
  OAI21_X1 U18927 ( .B1(n19855), .B2(n15711), .A(n19839), .ZN(n15714) );
  INV_X1 U18928 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15727) );
  OAI22_X1 U18929 ( .A1(n19833), .A2(n15727), .B1(n15712), .B2(n15792), .ZN(
        n15713) );
  AOI211_X1 U18930 ( .C1(n19860), .C2(n15865), .A(n15714), .B(n15713), .ZN(
        n15717) );
  AOI22_X1 U18931 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15715), .B1(n19847), 
        .B2(n15789), .ZN(n15716) );
  OAI211_X1 U18932 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15718), .A(n15717), 
        .B(n15716), .ZN(P1_U2829) );
  AOI22_X1 U18933 ( .A1(n15732), .A2(n19900), .B1(n19899), .B2(n15814), .ZN(
        n15719) );
  OAI21_X1 U18934 ( .B1(n19904), .B2(n15618), .A(n15719), .ZN(P1_U2847) );
  INV_X1 U18935 ( .A(n15720), .ZN(n15840) );
  AOI22_X1 U18936 ( .A1(n15776), .A2(n19900), .B1(n19899), .B2(n15840), .ZN(
        n15721) );
  OAI21_X1 U18937 ( .B1(n19904), .B2(n15722), .A(n15721), .ZN(P1_U2857) );
  AOI22_X1 U18938 ( .A1(n15779), .A2(n19900), .B1(n19899), .B2(n15723), .ZN(
        n15724) );
  OAI21_X1 U18939 ( .B1(n19904), .B2(n15725), .A(n15724), .ZN(P1_U2860) );
  AOI22_X1 U18940 ( .A1(n15789), .A2(n19900), .B1(n19899), .B2(n15865), .ZN(
        n15726) );
  OAI21_X1 U18941 ( .B1(n19904), .B2(n15727), .A(n15726), .ZN(P1_U2861) );
  AOI22_X1 U18942 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n15734) );
  NOR2_X1 U18943 ( .A1(n15772), .A2(n15739), .ZN(n15728) );
  AOI21_X1 U18944 ( .B1(n12646), .B2(n15772), .A(n15728), .ZN(n15729) );
  OAI211_X1 U18945 ( .C1(n15730), .C2(n12646), .A(n15729), .B(n15740), .ZN(
        n15731) );
  XNOR2_X1 U18946 ( .A(n15731), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15813) );
  AOI22_X1 U18947 ( .A1(n19947), .A2(n15732), .B1(n15813), .B2(n19948), .ZN(
        n15733) );
  OAI211_X1 U18948 ( .C1(n19953), .C2(n15735), .A(n15734), .B(n15733), .ZN(
        P1_U2974) );
  AOI22_X1 U18949 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15743) );
  MUX2_X1 U18950 ( .A(n15739), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .S(
        n9588), .Z(n15737) );
  NAND2_X1 U18951 ( .A1(n15772), .A2(n15739), .ZN(n15736) );
  MUX2_X1 U18952 ( .A(n15737), .B(n15736), .S(n14591), .Z(n15738) );
  OAI21_X1 U18953 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(n15819) );
  AOI22_X1 U18954 ( .A1(n15819), .A2(n19948), .B1(n15741), .B2(n19947), .ZN(
        n15742) );
  OAI211_X1 U18955 ( .C1(n19953), .C2(n15744), .A(n15743), .B(n15742), .ZN(
        P1_U2976) );
  AOI22_X1 U18956 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U18957 ( .A1(n15746), .A2(n19948), .B1(n19947), .B2(n15745), .ZN(
        n15747) );
  OAI211_X1 U18958 ( .C1(n19953), .C2(n15749), .A(n15748), .B(n15747), .ZN(
        P1_U2978) );
  AOI22_X1 U18959 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15753) );
  AOI22_X1 U18960 ( .A1(n15751), .A2(n19947), .B1(n15781), .B2(n15750), .ZN(
        n15752) );
  OAI211_X1 U18961 ( .C1(n15754), .C2(n19803), .A(n15753), .B(n15752), .ZN(
        P1_U2979) );
  AOI22_X1 U18962 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15758) );
  AOI22_X1 U18963 ( .A1(n15756), .A2(n19948), .B1(n19947), .B2(n15755), .ZN(
        n15757) );
  OAI211_X1 U18964 ( .C1(n19953), .C2(n15759), .A(n15758), .B(n15757), .ZN(
        P1_U2980) );
  AOI22_X1 U18965 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15763) );
  AOI22_X1 U18966 ( .A1(n15761), .A2(n19947), .B1(n15781), .B2(n15760), .ZN(
        n15762) );
  OAI211_X1 U18967 ( .C1(n19803), .C2(n15764), .A(n15763), .B(n15762), .ZN(
        P1_U2982) );
  AOI22_X1 U18968 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15769) );
  INV_X1 U18969 ( .A(n15765), .ZN(n15766) );
  AOI22_X1 U18970 ( .A1(n15767), .A2(n19947), .B1(n15781), .B2(n15766), .ZN(
        n15768) );
  OAI211_X1 U18971 ( .C1(n19803), .C2(n15770), .A(n15769), .B(n15768), .ZN(
        P1_U2983) );
  AOI21_X1 U18972 ( .B1(n15842), .B2(n15772), .A(n15771), .ZN(n15773) );
  XNOR2_X1 U18973 ( .A(n15774), .B(n15773), .ZN(n15837) );
  AOI22_X1 U18974 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U18975 ( .A1(n15776), .A2(n19947), .B1(n15781), .B2(n15775), .ZN(
        n15777) );
  OAI211_X1 U18976 ( .C1(n15837), .C2(n19803), .A(n15778), .B(n15777), .ZN(
        P1_U2984) );
  AOI22_X1 U18977 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15783) );
  AOI22_X1 U18978 ( .A1(n15781), .A2(n15780), .B1(n19947), .B2(n15779), .ZN(
        n15782) );
  OAI211_X1 U18979 ( .C1(n15784), .C2(n19803), .A(n15783), .B(n15782), .ZN(
        P1_U2987) );
  AOI22_X1 U18980 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15791) );
  NOR3_X1 U18981 ( .A1(n14617), .A2(n15785), .A3(n11900), .ZN(n15787) );
  NOR2_X1 U18982 ( .A1(n15787), .A2(n15786), .ZN(n15788) );
  XNOR2_X1 U18983 ( .A(n15788), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15867) );
  AOI22_X1 U18984 ( .A1(n19948), .A2(n15867), .B1(n19947), .B2(n15789), .ZN(
        n15790) );
  OAI211_X1 U18985 ( .C1(n19953), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        P1_U2988) );
  AOI22_X1 U18986 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15798) );
  NAND2_X1 U18987 ( .A1(n15795), .A2(n15794), .ZN(n15796) );
  XNOR2_X1 U18988 ( .A(n15793), .B(n15796), .ZN(n15909) );
  AOI22_X1 U18989 ( .A1(n15909), .A2(n19948), .B1(n19947), .B2(n19895), .ZN(
        n15797) );
  OAI211_X1 U18990 ( .C1(n19953), .C2(n19830), .A(n15798), .B(n15797), .ZN(
        P1_U2992) );
  AOI22_X1 U18991 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15803) );
  XNOR2_X1 U18992 ( .A(n15800), .B(n15900), .ZN(n15801) );
  XNOR2_X1 U18993 ( .A(n15799), .B(n15801), .ZN(n15917) );
  AOI22_X1 U18994 ( .A1(n15917), .A2(n19948), .B1(n19947), .B2(n19901), .ZN(
        n15802) );
  OAI211_X1 U18995 ( .C1(n19953), .C2(n19843), .A(n15803), .B(n15802), .ZN(
        P1_U2993) );
  AOI22_X1 U18996 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15809) );
  OAI21_X1 U18997 ( .B1(n15806), .B2(n15805), .A(n15804), .ZN(n15928) );
  INV_X1 U18998 ( .A(n15928), .ZN(n15807) );
  AOI22_X1 U18999 ( .A1(n15807), .A2(n19948), .B1(n19947), .B2(n19862), .ZN(
        n15808) );
  OAI211_X1 U19000 ( .C1(n19953), .C2(n19852), .A(n15809), .B(n15808), .ZN(
        P1_U2994) );
  NOR4_X1 U19001 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n12646), .A3(
        n15739), .A4(n15810), .ZN(n15812) );
  NOR2_X1 U19002 ( .A1(n19957), .A2(n20745), .ZN(n15811) );
  AOI211_X1 U19003 ( .C1(n15813), .C2(n19970), .A(n15812), .B(n15811), .ZN(
        n15817) );
  AOI22_X1 U19004 ( .A1(n15815), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n19967), .B2(n15814), .ZN(n15816) );
  NAND2_X1 U19005 ( .A1(n15817), .A2(n15816), .ZN(P1_U3006) );
  AOI22_X1 U19006 ( .A1(n15819), .A2(n19970), .B1(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15818), .ZN(n15826) );
  INV_X1 U19007 ( .A(n15820), .ZN(n15824) );
  INV_X1 U19008 ( .A(n15821), .ZN(n15835) );
  OAI22_X1 U19009 ( .A1(n15822), .A2(n19983), .B1(n20741), .B2(n19957), .ZN(
        n15823) );
  AOI21_X1 U19010 ( .B1(n15824), .B2(n15835), .A(n15823), .ZN(n15825) );
  NAND2_X1 U19011 ( .A1(n15826), .A2(n15825), .ZN(P1_U3008) );
  OAI22_X1 U19012 ( .A1(n15828), .A2(n19977), .B1(n19983), .B2(n15827), .ZN(
        n15829) );
  AOI21_X1 U19013 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15830), .A(
        n15829), .ZN(n15834) );
  NAND3_X1 U19014 ( .A1(n15832), .A2(n15831), .A3(n15835), .ZN(n15833) );
  OAI211_X1 U19015 ( .C1(n20734), .C2(n19957), .A(n15834), .B(n15833), .ZN(
        P1_U3013) );
  NAND2_X1 U19016 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15835), .ZN(
        n15836) );
  OAI22_X1 U19017 ( .A1(n19957), .A2(n20729), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15836), .ZN(n15839) );
  NOR2_X1 U19018 ( .A1(n15837), .A2(n19977), .ZN(n15838) );
  AOI211_X1 U19019 ( .C1(n19967), .C2(n15840), .A(n15839), .B(n15838), .ZN(
        n15841) );
  OAI21_X1 U19020 ( .B1(n15843), .B2(n15842), .A(n15841), .ZN(P1_U3016) );
  INV_X1 U19021 ( .A(n15844), .ZN(n15850) );
  NAND2_X1 U19022 ( .A1(n15872), .A2(n15922), .ZN(n15920) );
  NOR4_X1 U19023 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15846), .A3(
        n15845), .A4(n15920), .ZN(n15849) );
  INV_X1 U19024 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20726) );
  OAI22_X1 U19025 ( .A1(n15847), .A2(n19983), .B1(n20726), .B2(n19957), .ZN(
        n15848) );
  AOI211_X1 U19026 ( .C1(n15850), .C2(n19970), .A(n15849), .B(n15848), .ZN(
        n15851) );
  OAI21_X1 U19027 ( .B1(n15853), .B2(n15852), .A(n15851), .ZN(P1_U3017) );
  AOI21_X1 U19028 ( .B1(n15856), .B2(n15855), .A(n15854), .ZN(n15864) );
  INV_X1 U19029 ( .A(n15857), .ZN(n15858) );
  AOI21_X1 U19030 ( .B1(n15859), .B2(n19967), .A(n15858), .ZN(n15863) );
  AOI22_X1 U19031 ( .A1(n15861), .A2(n19970), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15860), .ZN(n15862) );
  OAI211_X1 U19032 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15864), .A(
        n15863), .B(n15862), .ZN(P1_U3018) );
  AOI22_X1 U19033 ( .A1(n15865), .A2(n19967), .B1(n19940), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15869) );
  AOI22_X1 U19034 ( .A1(n15867), .A2(n19970), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15866), .ZN(n15868) );
  OAI211_X1 U19035 ( .C1(n15920), .C2(n15870), .A(n15869), .B(n15868), .ZN(
        P1_U3020) );
  AOI21_X1 U19036 ( .B1(n15893), .B2(n15872), .A(n15871), .ZN(n15873) );
  AOI221_X1 U19037 ( .B1(n15873), .B2(n15896), .C1(n15877), .C2(n15896), .A(
        n15887), .ZN(n15886) );
  OAI222_X1 U19038 ( .A1(n15875), .A2(n19983), .B1(n19957), .B2(n20720), .C1(
        n19977), .C2(n15874), .ZN(n15876) );
  INV_X1 U19039 ( .A(n15876), .ZN(n15879) );
  NOR2_X1 U19040 ( .A1(n15877), .A2(n15920), .ZN(n15882) );
  OAI221_X1 U19041 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n11900), .C2(n12632), .A(
        n15882), .ZN(n15878) );
  OAI211_X1 U19042 ( .C1(n15886), .C2(n11900), .A(n15879), .B(n15878), .ZN(
        P1_U3021) );
  INV_X1 U19043 ( .A(n15880), .ZN(n15881) );
  AOI21_X1 U19044 ( .B1(n19820), .B2(n19967), .A(n15881), .ZN(n15885) );
  AOI22_X1 U19045 ( .A1(n15883), .A2(n19970), .B1(n12632), .B2(n15882), .ZN(
        n15884) );
  OAI211_X1 U19046 ( .C1(n15886), .C2(n12632), .A(n15885), .B(n15884), .ZN(
        P1_U3022) );
  NAND2_X1 U19047 ( .A1(n19954), .A2(n15926), .ZN(n15932) );
  AOI21_X1 U19048 ( .B1(n15889), .B2(n15888), .A(n15887), .ZN(n19989) );
  NAND2_X1 U19049 ( .A1(n15890), .A2(n15921), .ZN(n19982) );
  OAI211_X1 U19050 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n15893), .A(
        n19989), .B(n19982), .ZN(n19972) );
  INV_X1 U19051 ( .A(n15891), .ZN(n15892) );
  OAI22_X1 U19052 ( .A1(n15893), .A2(n19954), .B1(n15892), .B2(n19981), .ZN(
        n15894) );
  NOR2_X1 U19053 ( .A1(n19972), .A2(n15894), .ZN(n15927) );
  OAI21_X1 U19054 ( .B1(n15895), .B2(n15932), .A(n15927), .ZN(n15916) );
  AOI21_X1 U19055 ( .B1(n15900), .B2(n15896), .A(n15916), .ZN(n15913) );
  OAI222_X1 U19056 ( .A1(n15898), .A2(n19983), .B1(n19957), .B2(n20717), .C1(
        n19977), .C2(n15897), .ZN(n15899) );
  INV_X1 U19057 ( .A(n15899), .ZN(n15902) );
  NOR2_X1 U19058 ( .A1(n15900), .A2(n15920), .ZN(n15908) );
  OAI221_X1 U19059 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12628), .C2(n15912), .A(
        n15908), .ZN(n15901) );
  OAI211_X1 U19060 ( .C1(n15913), .C2(n12628), .A(n15902), .B(n15901), .ZN(
        P1_U3023) );
  NAND2_X1 U19061 ( .A1(n15914), .A2(n15915), .ZN(n15905) );
  INV_X1 U19062 ( .A(n15903), .ZN(n15904) );
  NAND2_X1 U19063 ( .A1(n15905), .A2(n15904), .ZN(n15907) );
  AND2_X1 U19064 ( .A1(n15907), .A2(n15906), .ZN(n19894) );
  AOI22_X1 U19065 ( .A1(n19894), .A2(n19967), .B1(n19940), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n15911) );
  AOI22_X1 U19066 ( .A1(n15909), .A2(n19970), .B1(n15908), .B2(n15912), .ZN(
        n15910) );
  OAI211_X1 U19067 ( .C1(n15913), .C2(n15912), .A(n15911), .B(n15910), .ZN(
        P1_U3024) );
  XOR2_X1 U19068 ( .A(n15915), .B(n15914), .Z(n19898) );
  AOI22_X1 U19069 ( .A1(n19898), .A2(n19967), .B1(n19940), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15919) );
  AOI22_X1 U19070 ( .A1(n15917), .A2(n19970), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15916), .ZN(n15918) );
  OAI211_X1 U19071 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15920), .A(
        n15919), .B(n15918), .ZN(P1_U3025) );
  INV_X1 U19072 ( .A(n15921), .ZN(n15923) );
  NAND2_X1 U19073 ( .A1(n15923), .A2(n15922), .ZN(n19975) );
  INV_X1 U19074 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n15924) );
  OAI22_X1 U19075 ( .A1(n19854), .A2(n19983), .B1(n19957), .B2(n15924), .ZN(
        n15925) );
  INV_X1 U19076 ( .A(n15925), .ZN(n15931) );
  OAI22_X1 U19077 ( .A1(n15928), .A2(n19977), .B1(n15927), .B2(n15926), .ZN(
        n15929) );
  INV_X1 U19078 ( .A(n15929), .ZN(n15930) );
  OAI211_X1 U19079 ( .C1(n15932), .C2(n19975), .A(n15931), .B(n15930), .ZN(
        P1_U3026) );
  INV_X1 U19080 ( .A(n20781), .ZN(n20783) );
  NAND4_X1 U19081 ( .A1(n15936), .A2(n15935), .A3(n15934), .A4(n15933), .ZN(
        n15937) );
  OAI21_X1 U19082 ( .B1(n20783), .B2(n13828), .A(n15937), .ZN(P1_U3468) );
  NAND4_X1 U19083 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20689), .A4(n20797), .ZN(n15938) );
  AND2_X1 U19084 ( .A1(n15939), .A2(n15938), .ZN(n20688) );
  NAND2_X1 U19085 ( .A1(n20688), .A2(n15940), .ZN(n15941) );
  AOI22_X1 U19086 ( .A1(n15944), .A2(n15943), .B1(n15942), .B2(n15941), .ZN(
        P1_U3162) );
  OAI21_X1 U19087 ( .B1(n20690), .B2(n20323), .A(n15945), .ZN(P1_U3466) );
  AOI22_X1 U19088 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18912), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n9691), .ZN(n15957) );
  AOI22_X1 U19089 ( .A1(n15946), .A2(n13079), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n18927), .ZN(n15956) );
  INV_X1 U19090 ( .A(n15947), .ZN(n15949) );
  AOI22_X1 U19091 ( .A1(n15949), .A2(n18932), .B1(n15948), .B2(n18958), .ZN(
        n15955) );
  AOI21_X1 U19092 ( .B1(n15952), .B2(n15950), .A(n15951), .ZN(n15953) );
  NAND2_X1 U19093 ( .A1(n18933), .A2(n15953), .ZN(n15954) );
  NAND4_X1 U19094 ( .A1(n15957), .A2(n15956), .A3(n15955), .A4(n15954), .ZN(
        P2_U2826) );
  AOI22_X1 U19095 ( .A1(n15959), .A2(n18932), .B1(n15958), .B2(n18958), .ZN(
        n15968) );
  AOI211_X1 U19096 ( .C1(n15962), .C2(n15960), .A(n15961), .B(n19638), .ZN(
        n15966) );
  AOI22_X1 U19097 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n9691), .ZN(n15963) );
  OAI21_X1 U19098 ( .B1(n15964), .B2(n18924), .A(n15963), .ZN(n15965) );
  AOI211_X1 U19099 ( .C1(P2_EBX_REG_27__SCAN_IN), .C2(n18927), .A(n15966), .B(
        n15965), .ZN(n15967) );
  NAND2_X1 U19100 ( .A1(n15968), .A2(n15967), .ZN(P2_U2828) );
  AOI211_X1 U19101 ( .C1(n15971), .C2(n15969), .A(n15970), .B(n19638), .ZN(
        n15979) );
  NAND2_X1 U19102 ( .A1(n15972), .A2(n13079), .ZN(n15976) );
  AOI22_X1 U19103 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n9691), .ZN(n15973) );
  INV_X1 U19104 ( .A(n15973), .ZN(n15974) );
  AOI21_X1 U19105 ( .B1(n18927), .B2(P2_EBX_REG_26__SCAN_IN), .A(n15974), .ZN(
        n15975) );
  OAI211_X1 U19106 ( .C1(n18954), .C2(n15977), .A(n15976), .B(n15975), .ZN(
        n15978) );
  AOI211_X1 U19107 ( .C1(n18958), .C2(n15980), .A(n15979), .B(n15978), .ZN(
        n15981) );
  INV_X1 U19108 ( .A(n15981), .ZN(P2_U2829) );
  AOI22_X1 U19109 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n9691), .ZN(n15992) );
  AOI22_X1 U19110 ( .A1(n15982), .A2(n13079), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n18927), .ZN(n15991) );
  INV_X1 U19111 ( .A(n15983), .ZN(n16131) );
  AOI22_X1 U19112 ( .A1(n18932), .A2(n16131), .B1(n18958), .B2(n15984), .ZN(
        n15990) );
  AOI21_X1 U19113 ( .B1(n15987), .B2(n15986), .A(n15985), .ZN(n15988) );
  NAND2_X1 U19114 ( .A1(n18933), .A2(n15988), .ZN(n15989) );
  NAND4_X1 U19115 ( .A1(n15992), .A2(n15991), .A3(n15990), .A4(n15989), .ZN(
        P2_U2830) );
  AOI22_X1 U19116 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n9691), .ZN(n16002) );
  AOI22_X1 U19117 ( .A1(n15993), .A2(n13079), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n18927), .ZN(n16001) );
  AOI22_X1 U19118 ( .A1(n18932), .A2(n16144), .B1(n18958), .B2(n15994), .ZN(
        n16000) );
  AOI21_X1 U19119 ( .B1(n15997), .B2(n15996), .A(n15995), .ZN(n15998) );
  NAND2_X1 U19120 ( .A1(n18933), .A2(n15998), .ZN(n15999) );
  NAND4_X1 U19121 ( .A1(n16002), .A2(n16001), .A3(n16000), .A4(n15999), .ZN(
        P2_U2832) );
  INV_X1 U19122 ( .A(n16003), .ZN(n16005) );
  AOI22_X1 U19123 ( .A1(n16005), .A2(n16004), .B1(n18995), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16012) );
  AOI22_X1 U19124 ( .A1(n18962), .A2(BUF1_REG_19__SCAN_IN), .B1(n18963), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n16011) );
  INV_X1 U19125 ( .A(n16006), .ZN(n16007) );
  XNOR2_X1 U19126 ( .A(n16008), .B(n16007), .ZN(n18802) );
  AOI22_X1 U19127 ( .A1(n16009), .A2(n18998), .B1(n18996), .B2(n18802), .ZN(
        n16010) );
  NAND3_X1 U19128 ( .A1(n16012), .A2(n16011), .A3(n16010), .ZN(P2_U2900) );
  AOI22_X1 U19129 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19040), .ZN(n16020) );
  NAND2_X1 U19130 ( .A1(n16013), .A2(n19048), .ZN(n16016) );
  NAND2_X1 U19131 ( .A1(n19047), .A2(n16014), .ZN(n16015) );
  OAI211_X1 U19132 ( .C1(n16017), .C2(n16109), .A(n16016), .B(n16015), .ZN(
        n16018) );
  INV_X1 U19133 ( .A(n16018), .ZN(n16019) );
  OAI211_X1 U19134 ( .C1(n19052), .C2(n16021), .A(n16020), .B(n16019), .ZN(
        P2_U2990) );
  AOI22_X1 U19135 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19040), .ZN(n16029) );
  NAND2_X1 U19136 ( .A1(n16022), .A2(n19046), .ZN(n16025) );
  NAND2_X1 U19137 ( .A1(n16023), .A2(n19047), .ZN(n16024) );
  OAI211_X1 U19138 ( .C1(n16026), .C2(n16108), .A(n16025), .B(n16024), .ZN(
        n16027) );
  INV_X1 U19139 ( .A(n16027), .ZN(n16028) );
  OAI211_X1 U19140 ( .C1(n19052), .C2(n16030), .A(n16029), .B(n16028), .ZN(
        P2_U2992) );
  AOI22_X1 U19141 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19040), .ZN(n16039) );
  AOI211_X1 U19142 ( .C1(n16032), .C2(n15307), .A(n16031), .B(n16108), .ZN(
        n16037) );
  OAI22_X1 U19143 ( .A1(n16035), .A2(n16109), .B1(n16034), .B2(n16033), .ZN(
        n16036) );
  NOR2_X1 U19144 ( .A1(n16037), .A2(n16036), .ZN(n16038) );
  OAI211_X1 U19145 ( .C1(n19052), .C2(n16040), .A(n16039), .B(n16038), .ZN(
        P2_U2998) );
  AOI22_X1 U19146 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19040), .B1(n16115), 
        .B2(n18836), .ZN(n16045) );
  OAI22_X1 U19147 ( .A1(n16042), .A2(n16108), .B1(n16041), .B2(n16109), .ZN(
        n16043) );
  AOI21_X1 U19148 ( .B1(n19047), .B2(n18837), .A(n16043), .ZN(n16044) );
  OAI211_X1 U19149 ( .C1(n16124), .C2(n18830), .A(n16045), .B(n16044), .ZN(
        P2_U2999) );
  AOI22_X1 U19150 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19040), .ZN(n16054) );
  OAI21_X1 U19151 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16047), .A(
        n16046), .ZN(n16171) );
  OR2_X1 U19152 ( .A1(n16171), .A2(n16108), .ZN(n16053) );
  NAND2_X1 U19153 ( .A1(n16049), .A2(n16048), .ZN(n16050) );
  XNOR2_X1 U19154 ( .A(n16051), .B(n16050), .ZN(n16168) );
  AOI22_X1 U19155 ( .A1(n16168), .A2(n19046), .B1(n19047), .B2(n18850), .ZN(
        n16052) );
  OAI211_X1 U19156 ( .C1(n19052), .C2(n18843), .A(n16054), .B(n9912), .ZN(
        P2_U3000) );
  AOI22_X1 U19157 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19040), .ZN(n16059) );
  AOI222_X1 U19158 ( .A1(n16057), .A2(n19046), .B1(n19047), .B2(n16056), .C1(
        n16055), .C2(n19048), .ZN(n16058) );
  OAI211_X1 U19159 ( .C1(n19052), .C2(n18870), .A(n16059), .B(n16058), .ZN(
        P2_U3002) );
  AOI22_X1 U19160 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19040), .B1(n16115), 
        .B2(n18890), .ZN(n16072) );
  NOR2_X1 U19161 ( .A1(n16183), .A2(n16082), .ZN(n16081) );
  OAI21_X1 U19162 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16081), .A(
        n16060), .ZN(n16176) );
  NAND2_X1 U19163 ( .A1(n16061), .A2(n16062), .ZN(n16065) );
  INV_X1 U19164 ( .A(n16063), .ZN(n16064) );
  NAND2_X1 U19165 ( .A1(n16065), .A2(n16064), .ZN(n16069) );
  NOR2_X1 U19166 ( .A1(n16067), .A2(n16066), .ZN(n16068) );
  XNOR2_X1 U19167 ( .A(n16069), .B(n16068), .ZN(n16180) );
  OAI22_X1 U19168 ( .A1(n16176), .A2(n16108), .B1(n16180), .B2(n16109), .ZN(
        n16070) );
  AOI21_X1 U19169 ( .B1(n19047), .B2(n18889), .A(n16070), .ZN(n16071) );
  OAI211_X1 U19170 ( .C1(n16124), .C2(n16073), .A(n16072), .B(n16071), .ZN(
        P2_U3003) );
  AOI22_X1 U19171 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19040), .ZN(n16085) );
  AND2_X1 U19172 ( .A1(n16061), .A2(n16074), .ZN(n16076) );
  NOR2_X1 U19173 ( .A1(n16076), .A2(n16075), .ZN(n16080) );
  NAND2_X1 U19174 ( .A1(n16078), .A2(n16077), .ZN(n16079) );
  XNOR2_X1 U19175 ( .A(n16080), .B(n16079), .ZN(n16192) );
  INV_X1 U19176 ( .A(n16192), .ZN(n16083) );
  AOI21_X1 U19177 ( .B1(n16183), .B2(n16082), .A(n16081), .ZN(n16188) );
  AOI222_X1 U19178 ( .A1(n16083), .A2(n19046), .B1(n19047), .B2(n16187), .C1(
        n19048), .C2(n16188), .ZN(n16084) );
  OAI211_X1 U19179 ( .C1(n19052), .C2(n16086), .A(n16085), .B(n16084), .ZN(
        P2_U3004) );
  AOI22_X1 U19180 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19040), .B1(n16115), 
        .B2(n18900), .ZN(n16091) );
  OAI22_X1 U19181 ( .A1(n16088), .A2(n16108), .B1(n16109), .B2(n16087), .ZN(
        n16089) );
  AOI21_X1 U19182 ( .B1(n19047), .B2(n18901), .A(n16089), .ZN(n16090) );
  OAI211_X1 U19183 ( .C1(n16124), .C2(n18894), .A(n16091), .B(n16090), .ZN(
        P2_U3005) );
  AOI22_X1 U19184 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19040), .ZN(n16105) );
  OAI21_X1 U19185 ( .B1(n16094), .B2(n16093), .A(n16092), .ZN(n16205) );
  AOI21_X1 U19186 ( .B1(n15161), .B2(n16096), .A(n16095), .ZN(n16101) );
  INV_X1 U19187 ( .A(n16097), .ZN(n16099) );
  NOR2_X1 U19188 ( .A1(n16099), .A2(n16098), .ZN(n16100) );
  XNOR2_X1 U19189 ( .A(n16101), .B(n16100), .ZN(n16202) );
  AOI22_X1 U19190 ( .A1(n16202), .A2(n19046), .B1(n19047), .B2(n16201), .ZN(
        n16102) );
  OAI21_X1 U19191 ( .B1(n16205), .B2(n16108), .A(n16102), .ZN(n16103) );
  INV_X1 U19192 ( .A(n16103), .ZN(n16104) );
  OAI211_X1 U19193 ( .C1(n19052), .C2(n16106), .A(n16105), .B(n16104), .ZN(
        P2_U3006) );
  AOI22_X1 U19194 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19040), .B1(n16115), 
        .B2(n18930), .ZN(n16113) );
  OAI22_X1 U19195 ( .A1(n16110), .A2(n16109), .B1(n16108), .B2(n16107), .ZN(
        n16111) );
  AOI21_X1 U19196 ( .B1(n19047), .B2(n18931), .A(n16111), .ZN(n16112) );
  OAI211_X1 U19197 ( .C1(n16124), .C2(n20875), .A(n16113), .B(n16112), .ZN(
        P2_U3009) );
  AOI22_X1 U19198 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19040), .B1(n16115), 
        .B2(n16114), .ZN(n16123) );
  XNOR2_X1 U19199 ( .A(n16116), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16117) );
  XNOR2_X1 U19200 ( .A(n16118), .B(n16117), .ZN(n16211) );
  OAI21_X1 U19201 ( .B1(n16120), .B2(n16119), .A(n12490), .ZN(n16208) );
  INV_X1 U19202 ( .A(n16208), .ZN(n16121) );
  AOI222_X1 U19203 ( .A1(n19046), .A2(n16211), .B1(n16121), .B2(n19048), .C1(
        n16232), .C2(n19047), .ZN(n16122) );
  OAI211_X1 U19204 ( .C1(n16125), .C2(n16124), .A(n16123), .B(n16122), .ZN(
        P2_U3011) );
  OAI22_X1 U19205 ( .A1(n19058), .A2(n16126), .B1(n19691), .B2(n18920), .ZN(
        n16127) );
  AOI221_X1 U19206 ( .B1(n16130), .B2(n16129), .C1(n16128), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n16127), .ZN(n16134) );
  AOI22_X1 U19207 ( .A1(n16132), .A2(n19064), .B1(n19053), .B2(n16131), .ZN(
        n16133) );
  OAI211_X1 U19208 ( .C1(n16207), .C2(n16135), .A(n16134), .B(n16133), .ZN(
        P2_U3021) );
  NOR2_X1 U19209 ( .A1(n19688), .A2(n18920), .ZN(n16141) );
  OAI21_X1 U19210 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16136), .ZN(n16138) );
  OAI22_X1 U19211 ( .A1(n16139), .A2(n16138), .B1(n19058), .B2(n16137), .ZN(
        n16140) );
  AOI211_X1 U19212 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16142), .A(
        n16141), .B(n16140), .ZN(n16147) );
  INV_X1 U19213 ( .A(n16143), .ZN(n16145) );
  AOI22_X1 U19214 ( .A1(n16145), .A2(n19064), .B1(n19053), .B2(n16144), .ZN(
        n16146) );
  OAI211_X1 U19215 ( .C1(n16207), .C2(n16148), .A(n16147), .B(n16146), .ZN(
        P2_U3023) );
  NAND2_X1 U19216 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19040), .ZN(n16149) );
  OAI221_X1 U19217 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16152), 
        .C1(n16151), .C2(n16150), .A(n16149), .ZN(n16153) );
  AOI21_X1 U19218 ( .B1(n16199), .B2(n18802), .A(n16153), .ZN(n16156) );
  AOI22_X1 U19219 ( .A1(n16154), .A2(n19064), .B1(n19053), .B2(n18803), .ZN(
        n16155) );
  OAI211_X1 U19220 ( .C1(n16207), .C2(n16157), .A(n16156), .B(n16155), .ZN(
        P2_U3027) );
  NOR2_X1 U19221 ( .A1(n16158), .A2(n16159), .ZN(n16164) );
  INV_X1 U19222 ( .A(n16159), .ZN(n16161) );
  AOI221_X1 U19223 ( .B1(n12377), .B2(n16161), .C1(n12325), .C2(n16161), .A(
        n16160), .ZN(n16162) );
  INV_X1 U19224 ( .A(n16162), .ZN(n16163) );
  MUX2_X1 U19225 ( .A(n16164), .B(n16163), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16167) );
  AOI21_X1 U19226 ( .B1(n16165), .B2(n13847), .A(n13956), .ZN(n18849) );
  INV_X1 U19227 ( .A(n18849), .ZN(n18968) );
  OAI22_X1 U19228 ( .A1(n19058), .A2(n18968), .B1(n12951), .B2(n18920), .ZN(
        n16166) );
  NOR2_X1 U19229 ( .A1(n16167), .A2(n16166), .ZN(n16170) );
  AOI22_X1 U19230 ( .A1(n16168), .A2(n19064), .B1(n19053), .B2(n18850), .ZN(
        n16169) );
  OAI211_X1 U19231 ( .C1(n16207), .C2(n16171), .A(n16170), .B(n16169), .ZN(
        P2_U3032) );
  NAND2_X1 U19232 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16172), .ZN(
        n16184) );
  AOI211_X1 U19233 ( .C1(n16183), .C2(n12317), .A(n16173), .B(n16184), .ZN(
        n16175) );
  OAI22_X1 U19234 ( .A1(n16182), .A2(n12317), .B1(n19058), .B2(n18882), .ZN(
        n16174) );
  AOI211_X1 U19235 ( .C1(n19040), .C2(P2_REIP_REG_11__SCAN_IN), .A(n16175), 
        .B(n16174), .ZN(n16179) );
  INV_X1 U19236 ( .A(n16176), .ZN(n16177) );
  AOI22_X1 U19237 ( .A1(n19063), .A2(n16177), .B1(n19053), .B2(n18889), .ZN(
        n16178) );
  OAI211_X1 U19238 ( .C1(n16180), .C2(n16191), .A(n16179), .B(n16178), .ZN(
        P2_U3035) );
  NAND2_X1 U19239 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19040), .ZN(n16181) );
  OAI221_X1 U19240 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16184), 
        .C1(n16183), .C2(n16182), .A(n16181), .ZN(n16185) );
  AOI21_X1 U19241 ( .B1(n16186), .B2(n16199), .A(n16185), .ZN(n16190) );
  AOI22_X1 U19242 ( .A1(n16188), .A2(n19063), .B1(n19053), .B2(n16187), .ZN(
        n16189) );
  OAI211_X1 U19243 ( .C1(n16192), .C2(n16191), .A(n16190), .B(n16189), .ZN(
        P2_U3036) );
  NOR2_X1 U19244 ( .A1(n18920), .A2(n12929), .ZN(n16198) );
  OAI21_X1 U19245 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16193), .ZN(n16194) );
  OAI22_X1 U19246 ( .A1(n12302), .A2(n16196), .B1(n16195), .B2(n16194), .ZN(
        n16197) );
  AOI211_X1 U19247 ( .C1(n16200), .C2(n16199), .A(n16198), .B(n16197), .ZN(
        n16204) );
  AOI22_X1 U19248 ( .A1(n16202), .A2(n19064), .B1(n19053), .B2(n16201), .ZN(
        n16203) );
  OAI211_X1 U19249 ( .C1(n16207), .C2(n16205), .A(n16204), .B(n16203), .ZN(
        P2_U3038) );
  AOI22_X1 U19250 ( .A1(n16232), .A2(n19053), .B1(P2_REIP_REG_3__SCAN_IN), 
        .B2(n19040), .ZN(n16206) );
  OAI21_X1 U19251 ( .B1(n19728), .B2(n19058), .A(n16206), .ZN(n16210) );
  NOR2_X1 U19252 ( .A1(n16208), .A2(n16207), .ZN(n16209) );
  AOI211_X1 U19253 ( .C1(n16211), .C2(n19064), .A(n16210), .B(n16209), .ZN(
        n16212) );
  OAI221_X1 U19254 ( .B1(n16214), .B2(n9705), .C1(n16214), .C2(n16213), .A(
        n16212), .ZN(P2_U3043) );
  NOR2_X1 U19255 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19780), .ZN(n19636) );
  NAND3_X1 U19256 ( .A1(n16215), .A2(n13145), .A3(n19776), .ZN(n16216) );
  NAND2_X1 U19257 ( .A1(n16216), .A2(n19633), .ZN(n16277) );
  INV_X1 U19258 ( .A(n16277), .ZN(n16217) );
  AOI211_X1 U19259 ( .C1(n19785), .C2(n19636), .A(n16218), .B(n16217), .ZN(
        n16283) );
  NAND2_X1 U19260 ( .A1(n16262), .A2(n16219), .ZN(n16234) );
  NOR2_X1 U19261 ( .A1(n16220), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16241) );
  INV_X1 U19262 ( .A(n16241), .ZN(n16221) );
  NAND2_X1 U19263 ( .A1(n16234), .A2(n16221), .ZN(n16223) );
  AOI21_X1 U19264 ( .B1(n13210), .B2(n12445), .A(n16235), .ZN(n16222) );
  NAND2_X1 U19265 ( .A1(n16223), .A2(n16222), .ZN(n16230) );
  NAND2_X1 U19266 ( .A1(n16234), .A2(n16241), .ZN(n16228) );
  NAND2_X1 U19267 ( .A1(n13209), .A2(n16224), .ZN(n16225) );
  NAND2_X1 U19268 ( .A1(n16225), .A2(n12802), .ZN(n16240) );
  INV_X1 U19269 ( .A(n12445), .ZN(n16226) );
  NAND2_X1 U19270 ( .A1(n13210), .A2(n16226), .ZN(n16227) );
  NAND3_X1 U19271 ( .A1(n16228), .A2(n16240), .A3(n16227), .ZN(n16229) );
  MUX2_X1 U19272 ( .A(n16230), .B(n16229), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n16231) );
  AOI21_X1 U19273 ( .B1(n16232), .B2(n16243), .A(n16231), .ZN(n19712) );
  INV_X1 U19274 ( .A(n19712), .ZN(n16233) );
  INV_X1 U19275 ( .A(n16271), .ZN(n16249) );
  MUX2_X1 U19276 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16233), .S(
        n16249), .Z(n16273) );
  OAI21_X1 U19277 ( .B1(n16235), .B2(n16241), .A(n16234), .ZN(n16239) );
  NOR2_X1 U19278 ( .A1(n16236), .A2(n12445), .ZN(n16237) );
  NAND2_X1 U19279 ( .A1(n13210), .A2(n16237), .ZN(n16238) );
  OAI211_X1 U19280 ( .C1(n16241), .C2(n16240), .A(n16239), .B(n16238), .ZN(
        n16242) );
  AOI21_X1 U19281 ( .B1(n11973), .B2(n16243), .A(n16242), .ZN(n19718) );
  AND2_X1 U19282 ( .A1(n16271), .A2(n9883), .ZN(n16244) );
  AOI21_X1 U19283 ( .B1(n19718), .B2(n16249), .A(n16244), .ZN(n16272) );
  AND2_X1 U19284 ( .A1(n16272), .A2(n19734), .ZN(n16252) );
  INV_X1 U19285 ( .A(n16252), .ZN(n16245) );
  NOR2_X1 U19286 ( .A1(n16245), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16256) );
  NAND2_X1 U19287 ( .A1(n16246), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16251) );
  NAND2_X1 U19288 ( .A1(n16251), .A2(n19751), .ZN(n16247) );
  NAND2_X1 U19289 ( .A1(n16248), .A2(n16247), .ZN(n16250) );
  OAI211_X1 U19290 ( .C1(n19751), .C2(n16251), .A(n16250), .B(n16249), .ZN(
        n16254) );
  NOR2_X1 U19291 ( .A1(n16252), .A2(n19742), .ZN(n16253) );
  AOI211_X1 U19292 ( .C1(n19712), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16254), .B(n16253), .ZN(n16255) );
  AOI211_X1 U19293 ( .C1(n16273), .C2(n19734), .A(n16256), .B(n16255), .ZN(
        n16276) );
  NAND2_X1 U19294 ( .A1(n16263), .A2(n16257), .ZN(n16261) );
  NAND2_X1 U19295 ( .A1(n16259), .A2(n16258), .ZN(n16260) );
  OAI211_X1 U19296 ( .C1(n16263), .C2(n16262), .A(n16261), .B(n16260), .ZN(
        n19767) );
  OAI21_X1 U19297 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16264), .ZN(n16267) );
  NAND2_X1 U19298 ( .A1(n12449), .A2(n9609), .ZN(n16266) );
  OAI211_X1 U19299 ( .C1(n16269), .C2(n16268), .A(n16267), .B(n16266), .ZN(
        n16270) );
  AOI211_X1 U19300 ( .C1(n16271), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19767), .B(n16270), .ZN(n16275) );
  NAND2_X1 U19301 ( .A1(n16273), .A2(n16272), .ZN(n16274) );
  OAI211_X1 U19302 ( .C1(n16276), .C2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16275), .B(n16274), .ZN(n16281) );
  OR2_X1 U19303 ( .A1(n16281), .A2(n16277), .ZN(n16286) );
  NAND2_X1 U19304 ( .A1(n16286), .A2(n16278), .ZN(n19639) );
  AOI21_X1 U19305 ( .B1(n19780), .B2(n19719), .A(n19778), .ZN(n16279) );
  AOI21_X1 U19306 ( .B1(n19785), .B2(n19639), .A(n16279), .ZN(n16280) );
  AOI21_X1 U19307 ( .B1(n19633), .B2(n16281), .A(n16280), .ZN(n16282) );
  OAI211_X1 U19308 ( .C1(n19766), .C2(n16285), .A(n16283), .B(n16282), .ZN(
        P2_U3176) );
  INV_X1 U19309 ( .A(n19075), .ZN(n16284) );
  OAI211_X1 U19310 ( .C1(n20926), .C2(n16286), .A(n16285), .B(n16284), .ZN(
        P2_U3593) );
  NOR2_X1 U19311 ( .A1(n9624), .A2(n16287), .ZN(n16296) );
  INV_X1 U19312 ( .A(n16288), .ZN(n16290) );
  OAI21_X1 U19313 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n9624), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16289) );
  OAI221_X1 U19314 ( .B1(n20944), .B2(n16290), .C1(n9624), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16289), .ZN(n16295) );
  OAI21_X1 U19315 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n20944), .A(
        n16290), .ZN(n16293) );
  NAND2_X1 U19316 ( .A1(n9624), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16291) );
  OAI22_X1 U19317 ( .A1(n9624), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n16291), .B2(n20944), .ZN(n16292) );
  OAI21_X1 U19318 ( .B1(n16296), .B2(n16293), .A(n16292), .ZN(n16294) );
  OAI21_X1 U19319 ( .B1(n16296), .B2(n16295), .A(n16294), .ZN(n16334) );
  INV_X1 U19320 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18688) );
  NOR2_X1 U19321 ( .A1(n9600), .A2(n18688), .ZN(n16331) );
  INV_X1 U19322 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16465) );
  XOR2_X1 U19323 ( .A(n16465), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16299) );
  OAI22_X1 U19324 ( .A1(n16300), .A2(n16299), .B1(n16298), .B2(n16465), .ZN(
        n16301) );
  AOI211_X1 U19325 ( .C1(n17615), .C2(n16297), .A(n16331), .B(n16301), .ZN(
        n16306) );
  NAND2_X1 U19326 ( .A1(n16302), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16303) );
  XNOR2_X1 U19327 ( .A(n16303), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16324) );
  NAND2_X1 U19328 ( .A1(n16307), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16304) );
  XNOR2_X1 U19329 ( .A(n16304), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16325) );
  AOI22_X1 U19330 ( .A1(n17749), .A2(n16324), .B1(n17627), .B2(n16325), .ZN(
        n16305) );
  OAI211_X1 U19331 ( .C1(n17622), .C2(n16334), .A(n16306), .B(n16305), .ZN(
        P3_U2799) );
  AOI211_X1 U19332 ( .C1(n16309), .C2(n16308), .A(n16307), .B(n17674), .ZN(
        n16316) );
  OAI21_X1 U19333 ( .B1(n17615), .B2(n16311), .A(n16468), .ZN(n16312) );
  OAI211_X1 U19334 ( .C1(n16314), .C2(n9758), .A(n16313), .B(n16312), .ZN(
        n16315) );
  AOI211_X1 U19335 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16317), .A(
        n16316), .B(n16315), .ZN(n16321) );
  OAI211_X1 U19336 ( .C1(n16319), .C2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17749), .B(n16318), .ZN(n16320) );
  OAI211_X1 U19337 ( .C1(n16322), .C2(n17622), .A(n16321), .B(n16320), .ZN(
        P3_U2801) );
  OAI21_X1 U19338 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18076), .A(
        n16323), .ZN(n16332) );
  AOI22_X1 U19339 ( .A1(n18000), .A2(n16325), .B1(n17966), .B2(n16324), .ZN(
        n16329) );
  INV_X1 U19340 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18715) );
  NAND4_X1 U19341 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16327), .A3(
        n16326), .A4(n18715), .ZN(n16328) );
  AOI21_X1 U19342 ( .B1(n16329), .B2(n16328), .A(n18090), .ZN(n16330) );
  AOI211_X1 U19343 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16332), .A(
        n16331), .B(n16330), .ZN(n16333) );
  OAI21_X1 U19344 ( .B1(n17960), .B2(n16334), .A(n16333), .ZN(P3_U2831) );
  NOR3_X1 U19345 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16336) );
  NOR4_X1 U19346 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16335) );
  NAND4_X1 U19347 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16336), .A3(n16335), .A4(
        U215), .ZN(U213) );
  INV_X1 U19348 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16426) );
  INV_X1 U19349 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16427) );
  OAI222_X1 U19350 ( .A1(U212), .A2(n16426), .B1(n16391), .B2(n16338), .C1(
        U214), .C2(n16427), .ZN(U216) );
  INV_X1 U19351 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16424) );
  INV_X1 U19352 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16339) );
  INV_X1 U19353 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n20844) );
  OAI222_X1 U19354 ( .A1(U212), .A2(n16424), .B1(n16391), .B2(n16339), .C1(
        U214), .C2(n20844), .ZN(U217) );
  INV_X1 U19355 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16341) );
  AOI22_X1 U19356 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16388), .ZN(n16340) );
  OAI21_X1 U19357 ( .B1(n16341), .B2(n16391), .A(n16340), .ZN(U218) );
  INV_X1 U19358 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16343) );
  AOI22_X1 U19359 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16388), .ZN(n16342) );
  OAI21_X1 U19360 ( .B1(n16343), .B2(n16391), .A(n16342), .ZN(U219) );
  INV_X1 U19361 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16345) );
  AOI22_X1 U19362 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16388), .ZN(n16344) );
  OAI21_X1 U19363 ( .B1(n16345), .B2(n16391), .A(n16344), .ZN(U220) );
  INV_X1 U19364 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16347) );
  AOI22_X1 U19365 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16388), .ZN(n16346) );
  OAI21_X1 U19366 ( .B1(n16347), .B2(n16391), .A(n16346), .ZN(U221) );
  AOI22_X1 U19367 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16388), .ZN(n16348) );
  OAI21_X1 U19368 ( .B1(n16349), .B2(n16391), .A(n16348), .ZN(U222) );
  INV_X1 U19369 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16351) );
  AOI22_X1 U19370 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16388), .ZN(n16350) );
  OAI21_X1 U19371 ( .B1(n16351), .B2(n16391), .A(n16350), .ZN(U223) );
  AOI22_X1 U19372 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16388), .ZN(n16352) );
  OAI21_X1 U19373 ( .B1(n14998), .B2(n16391), .A(n16352), .ZN(U224) );
  AOI22_X1 U19374 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16388), .ZN(n16353) );
  OAI21_X1 U19375 ( .B1(n15007), .B2(n16391), .A(n16353), .ZN(U225) );
  AOI22_X1 U19376 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16388), .ZN(n16354) );
  OAI21_X1 U19377 ( .B1(n15015), .B2(n16391), .A(n16354), .ZN(U226) );
  AOI22_X1 U19378 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16388), .ZN(n16355) );
  OAI21_X1 U19379 ( .B1(n19101), .B2(n16391), .A(n16355), .ZN(U227) );
  AOI22_X1 U19380 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16388), .ZN(n16356) );
  OAI21_X1 U19381 ( .B1(n14517), .B2(n16391), .A(n16356), .ZN(U228) );
  INV_X1 U19382 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n19093) );
  AOI22_X1 U19383 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16388), .ZN(n16357) );
  OAI21_X1 U19384 ( .B1(n19093), .B2(n16391), .A(n16357), .ZN(U229) );
  AOI22_X1 U19385 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16388), .ZN(n16358) );
  OAI21_X1 U19386 ( .B1(n15039), .B2(n16391), .A(n16358), .ZN(U230) );
  INV_X1 U19387 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n19073) );
  AOI22_X1 U19388 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16388), .ZN(n16359) );
  OAI21_X1 U19389 ( .B1(n19073), .B2(n16391), .A(n16359), .ZN(U231) );
  AOI22_X1 U19390 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16388), .ZN(n16360) );
  OAI21_X1 U19391 ( .B1(n13744), .B2(n16391), .A(n16360), .ZN(U232) );
  AOI22_X1 U19392 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16388), .ZN(n16361) );
  OAI21_X1 U19393 ( .B1(n13006), .B2(n16391), .A(n16361), .ZN(U233) );
  INV_X1 U19394 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16363) );
  AOI22_X1 U19395 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16388), .ZN(n16362) );
  OAI21_X1 U19396 ( .B1(n16363), .B2(n16391), .A(n16362), .ZN(U234) );
  AOI22_X1 U19397 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16388), .ZN(n16364) );
  OAI21_X1 U19398 ( .B1(n16365), .B2(n16391), .A(n16364), .ZN(U235) );
  INV_X1 U19399 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19400 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16388), .ZN(n16366) );
  OAI21_X1 U19401 ( .B1(n16367), .B2(n16391), .A(n16366), .ZN(U236) );
  INV_X1 U19402 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16369) );
  AOI22_X1 U19403 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16388), .ZN(n16368) );
  OAI21_X1 U19404 ( .B1(n16369), .B2(n16391), .A(n16368), .ZN(U237) );
  INV_X1 U19405 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16371) );
  AOI22_X1 U19406 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16388), .ZN(n16370) );
  OAI21_X1 U19407 ( .B1(n16371), .B2(n16391), .A(n16370), .ZN(U238) );
  INV_X1 U19408 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16373) );
  AOI22_X1 U19409 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16388), .ZN(n16372) );
  OAI21_X1 U19410 ( .B1(n16373), .B2(n16391), .A(n16372), .ZN(U239) );
  INV_X1 U19411 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16375) );
  AOI22_X1 U19412 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16388), .ZN(n16374) );
  OAI21_X1 U19413 ( .B1(n16375), .B2(n16391), .A(n16374), .ZN(U240) );
  INV_X1 U19414 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16377) );
  AOI22_X1 U19415 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16388), .ZN(n16376) );
  OAI21_X1 U19416 ( .B1(n16377), .B2(n16391), .A(n16376), .ZN(U241) );
  INV_X1 U19417 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16379) );
  AOI22_X1 U19418 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16388), .ZN(n16378) );
  OAI21_X1 U19419 ( .B1(n16379), .B2(n16391), .A(n16378), .ZN(U242) );
  INV_X1 U19420 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16381) );
  AOI22_X1 U19421 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16388), .ZN(n16380) );
  OAI21_X1 U19422 ( .B1(n16381), .B2(n16391), .A(n16380), .ZN(U243) );
  INV_X1 U19423 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16383) );
  AOI22_X1 U19424 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16388), .ZN(n16382) );
  OAI21_X1 U19425 ( .B1(n16383), .B2(n16391), .A(n16382), .ZN(U244) );
  INV_X1 U19426 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16385) );
  AOI22_X1 U19427 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16388), .ZN(n16384) );
  OAI21_X1 U19428 ( .B1(n16385), .B2(n16391), .A(n16384), .ZN(U245) );
  INV_X1 U19429 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16387) );
  AOI22_X1 U19430 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16388), .ZN(n16386) );
  OAI21_X1 U19431 ( .B1(n16387), .B2(n16391), .A(n16386), .ZN(U246) );
  INV_X1 U19432 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16392) );
  AOI22_X1 U19433 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16389), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16388), .ZN(n16390) );
  OAI21_X1 U19434 ( .B1(n16392), .B2(n16391), .A(n16390), .ZN(U247) );
  OAI22_X1 U19435 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16425), .ZN(n16393) );
  INV_X1 U19436 ( .A(n16393), .ZN(U251) );
  OAI22_X1 U19437 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16425), .ZN(n16394) );
  INV_X1 U19438 ( .A(n16394), .ZN(U252) );
  INV_X1 U19439 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16395) );
  INV_X1 U19440 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18109) );
  AOI22_X1 U19441 ( .A1(n16425), .A2(n16395), .B1(n18109), .B2(U215), .ZN(U253) );
  INV_X1 U19442 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16396) );
  INV_X1 U19443 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18114) );
  AOI22_X1 U19444 ( .A1(n16420), .A2(n16396), .B1(n18114), .B2(U215), .ZN(U254) );
  INV_X1 U19445 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16397) );
  INV_X1 U19446 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U19447 ( .A1(n16425), .A2(n16397), .B1(n18118), .B2(U215), .ZN(U255) );
  OAI22_X1 U19448 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16425), .ZN(n16398) );
  INV_X1 U19449 ( .A(n16398), .ZN(U256) );
  INV_X1 U19450 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16399) );
  INV_X1 U19451 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18126) );
  AOI22_X1 U19452 ( .A1(n16425), .A2(n16399), .B1(n18126), .B2(U215), .ZN(U257) );
  INV_X1 U19453 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16400) );
  INV_X1 U19454 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18131) );
  AOI22_X1 U19455 ( .A1(n16425), .A2(n16400), .B1(n18131), .B2(U215), .ZN(U258) );
  OAI22_X1 U19456 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16425), .ZN(n16401) );
  INV_X1 U19457 ( .A(n16401), .ZN(U259) );
  INV_X1 U19458 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16402) );
  INV_X1 U19459 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U19460 ( .A1(n16420), .A2(n16402), .B1(n17253), .B2(U215), .ZN(U260) );
  INV_X1 U19461 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16403) );
  INV_X1 U19462 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U19463 ( .A1(n16425), .A2(n16403), .B1(n17249), .B2(U215), .ZN(U261) );
  OAI22_X1 U19464 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16425), .ZN(n16404) );
  INV_X1 U19465 ( .A(n16404), .ZN(U262) );
  INV_X1 U19466 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16405) );
  INV_X1 U19467 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U19468 ( .A1(n16425), .A2(n16405), .B1(n17242), .B2(U215), .ZN(U263) );
  OAI22_X1 U19469 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16425), .ZN(n16406) );
  INV_X1 U19470 ( .A(n16406), .ZN(U264) );
  OAI22_X1 U19471 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16425), .ZN(n16407) );
  INV_X1 U19472 ( .A(n16407), .ZN(U265) );
  INV_X1 U19473 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16408) );
  INV_X1 U19474 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n20889) );
  AOI22_X1 U19475 ( .A1(n16420), .A2(n16408), .B1(n20889), .B2(U215), .ZN(U266) );
  INV_X1 U19476 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n16409) );
  INV_X1 U19477 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19072) );
  AOI22_X1 U19478 ( .A1(n16425), .A2(n16409), .B1(n19072), .B2(U215), .ZN(U267) );
  INV_X1 U19479 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16410) );
  AOI22_X1 U19480 ( .A1(n16420), .A2(n16410), .B1(n15041), .B2(U215), .ZN(U268) );
  INV_X1 U19481 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16411) );
  INV_X1 U19482 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19092) );
  AOI22_X1 U19483 ( .A1(n16420), .A2(n16411), .B1(n19092), .B2(U215), .ZN(U269) );
  INV_X1 U19484 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16412) );
  INV_X1 U19485 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19097) );
  AOI22_X1 U19486 ( .A1(n16420), .A2(n16412), .B1(n19097), .B2(U215), .ZN(U270) );
  INV_X1 U19487 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16413) );
  AOI22_X1 U19488 ( .A1(n16420), .A2(n16413), .B1(n15022), .B2(U215), .ZN(U271) );
  INV_X1 U19489 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16414) );
  AOI22_X1 U19490 ( .A1(n16425), .A2(n16414), .B1(n15016), .B2(U215), .ZN(U272) );
  INV_X1 U19491 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16415) );
  AOI22_X1 U19492 ( .A1(n16425), .A2(n16415), .B1(n15008), .B2(U215), .ZN(U273) );
  INV_X1 U19493 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16416) );
  AOI22_X1 U19494 ( .A1(n16425), .A2(n16416), .B1(n14999), .B2(U215), .ZN(U274) );
  INV_X1 U19495 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16417) );
  INV_X1 U19496 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n20807) );
  AOI22_X1 U19497 ( .A1(n16425), .A2(n16417), .B1(n20807), .B2(U215), .ZN(U275) );
  OAI22_X1 U19498 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16420), .ZN(n16418) );
  INV_X1 U19499 ( .A(n16418), .ZN(U276) );
  OAI22_X1 U19500 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16420), .ZN(n16419) );
  INV_X1 U19501 ( .A(n16419), .ZN(U277) );
  OAI22_X1 U19502 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16420), .ZN(n16421) );
  INV_X1 U19503 ( .A(n16421), .ZN(U278) );
  OAI22_X1 U19504 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16425), .ZN(n16422) );
  INV_X1 U19505 ( .A(n16422), .ZN(U279) );
  OAI22_X1 U19506 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16425), .ZN(n16423) );
  INV_X1 U19507 ( .A(n16423), .ZN(U280) );
  INV_X1 U19508 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18125) );
  AOI22_X1 U19509 ( .A1(n16425), .A2(n16424), .B1(n18125), .B2(U215), .ZN(U281) );
  INV_X1 U19510 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18130) );
  AOI22_X1 U19511 ( .A1(n16425), .A2(n16426), .B1(n18130), .B2(U215), .ZN(U282) );
  INV_X1 U19512 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20892) );
  AOI222_X1 U19513 ( .A1(n16427), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16426), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n20892), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16428) );
  INV_X1 U19514 ( .A(n16430), .ZN(n16429) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18648) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19672) );
  AOI22_X1 U19517 ( .A1(n16429), .A2(n18648), .B1(n19672), .B2(n16430), .ZN(
        U347) );
  INV_X1 U19518 ( .A(n16430), .ZN(n16431) );
  INV_X1 U19519 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18646) );
  INV_X1 U19520 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19671) );
  AOI22_X1 U19521 ( .A1(n16431), .A2(n18646), .B1(n19671), .B2(n16430), .ZN(
        U348) );
  INV_X1 U19522 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18644) );
  INV_X1 U19523 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19670) );
  AOI22_X1 U19524 ( .A1(n16429), .A2(n18644), .B1(n19670), .B2(n16430), .ZN(
        U349) );
  INV_X1 U19525 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18642) );
  INV_X1 U19526 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19669) );
  AOI22_X1 U19527 ( .A1(n16429), .A2(n18642), .B1(n19669), .B2(n16430), .ZN(
        U350) );
  INV_X1 U19528 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18640) );
  INV_X1 U19529 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19667) );
  AOI22_X1 U19530 ( .A1(n16429), .A2(n18640), .B1(n19667), .B2(n16430), .ZN(
        U351) );
  INV_X1 U19531 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18637) );
  INV_X1 U19532 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19665) );
  AOI22_X1 U19533 ( .A1(n16429), .A2(n18637), .B1(n19665), .B2(n16430), .ZN(
        U352) );
  INV_X1 U19534 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18636) );
  INV_X1 U19535 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19664) );
  AOI22_X1 U19536 ( .A1(n16431), .A2(n18636), .B1(n19664), .B2(n16430), .ZN(
        U353) );
  INV_X1 U19537 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18634) );
  AOI22_X1 U19538 ( .A1(n16429), .A2(n18634), .B1(n19663), .B2(n16430), .ZN(
        U354) );
  INV_X1 U19539 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18687) );
  INV_X1 U19540 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19701) );
  AOI22_X1 U19541 ( .A1(n16429), .A2(n18687), .B1(n19701), .B2(n16430), .ZN(
        U355) );
  INV_X1 U19542 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18684) );
  INV_X1 U19543 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19698) );
  AOI22_X1 U19544 ( .A1(n16429), .A2(n18684), .B1(n19698), .B2(n16430), .ZN(
        U356) );
  INV_X1 U19545 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18681) );
  INV_X1 U19546 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19696) );
  AOI22_X1 U19547 ( .A1(n16429), .A2(n18681), .B1(n19696), .B2(n16430), .ZN(
        U357) );
  INV_X1 U19548 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18680) );
  INV_X1 U19549 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19693) );
  AOI22_X1 U19550 ( .A1(n16429), .A2(n18680), .B1(n19693), .B2(n16430), .ZN(
        U358) );
  INV_X1 U19551 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18678) );
  INV_X1 U19552 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20943) );
  AOI22_X1 U19553 ( .A1(n16429), .A2(n18678), .B1(n20943), .B2(n16430), .ZN(
        U359) );
  INV_X1 U19554 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18676) );
  INV_X1 U19555 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19692) );
  AOI22_X1 U19556 ( .A1(n16429), .A2(n18676), .B1(n19692), .B2(n16430), .ZN(
        U360) );
  INV_X1 U19557 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18674) );
  INV_X1 U19558 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19690) );
  AOI22_X1 U19559 ( .A1(n16429), .A2(n18674), .B1(n19690), .B2(n16430), .ZN(
        U361) );
  INV_X1 U19560 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18672) );
  INV_X1 U19561 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19689) );
  AOI22_X1 U19562 ( .A1(n16429), .A2(n18672), .B1(n19689), .B2(n16430), .ZN(
        U362) );
  INV_X1 U19563 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18670) );
  INV_X1 U19564 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19687) );
  AOI22_X1 U19565 ( .A1(n16429), .A2(n18670), .B1(n19687), .B2(n16430), .ZN(
        U363) );
  INV_X1 U19566 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18668) );
  INV_X1 U19567 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20888) );
  AOI22_X1 U19568 ( .A1(n16429), .A2(n18668), .B1(n20888), .B2(n16430), .ZN(
        U364) );
  INV_X1 U19569 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18632) );
  INV_X1 U19570 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U19571 ( .A1(n16429), .A2(n18632), .B1(n19662), .B2(n16430), .ZN(
        U365) );
  INV_X1 U19572 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18667) );
  INV_X1 U19573 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19685) );
  AOI22_X1 U19574 ( .A1(n16429), .A2(n18667), .B1(n19685), .B2(n16430), .ZN(
        U366) );
  INV_X1 U19575 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18665) );
  INV_X1 U19576 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19683) );
  AOI22_X1 U19577 ( .A1(n16429), .A2(n18665), .B1(n19683), .B2(n16430), .ZN(
        U367) );
  INV_X1 U19578 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18664) );
  INV_X1 U19579 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19682) );
  AOI22_X1 U19580 ( .A1(n16429), .A2(n18664), .B1(n19682), .B2(n16430), .ZN(
        U368) );
  INV_X1 U19581 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18661) );
  INV_X1 U19582 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19681) );
  AOI22_X1 U19583 ( .A1(n16429), .A2(n18661), .B1(n19681), .B2(n16430), .ZN(
        U369) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18660) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19679) );
  AOI22_X1 U19586 ( .A1(n16429), .A2(n18660), .B1(n19679), .B2(n16430), .ZN(
        U370) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18658) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19678) );
  AOI22_X1 U19589 ( .A1(n16431), .A2(n18658), .B1(n19678), .B2(n16430), .ZN(
        U371) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18655) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19677) );
  AOI22_X1 U19592 ( .A1(n16431), .A2(n18655), .B1(n19677), .B2(n16430), .ZN(
        U372) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18654) );
  INV_X1 U19594 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19676) );
  AOI22_X1 U19595 ( .A1(n16431), .A2(n18654), .B1(n19676), .B2(n16430), .ZN(
        U373) );
  INV_X1 U19596 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18652) );
  INV_X1 U19597 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19675) );
  AOI22_X1 U19598 ( .A1(n16431), .A2(n18652), .B1(n19675), .B2(n16430), .ZN(
        U374) );
  INV_X1 U19599 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18650) );
  INV_X1 U19600 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19674) );
  AOI22_X1 U19601 ( .A1(n16431), .A2(n18650), .B1(n19674), .B2(n16430), .ZN(
        U375) );
  INV_X1 U19602 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18630) );
  INV_X1 U19603 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19660) );
  AOI22_X1 U19604 ( .A1(n16431), .A2(n18630), .B1(n19660), .B2(n16430), .ZN(
        U376) );
  INV_X1 U19605 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16432) );
  NAND2_X1 U19606 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18629), .ZN(n18616) );
  AOI22_X1 U19607 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18616), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18626), .ZN(n18701) );
  INV_X1 U19608 ( .A(n18701), .ZN(n18698) );
  OAI21_X1 U19609 ( .B1(n18626), .B2(n16432), .A(n18698), .ZN(P3_U2633) );
  NAND2_X1 U19610 ( .A1(n18765), .A2(n18704), .ZN(n16434) );
  INV_X1 U19611 ( .A(n17760), .ZN(n18607) );
  OAI21_X1 U19612 ( .B1(n16439), .B2(n17330), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16433) );
  OAI21_X1 U19613 ( .B1(n16434), .B2(n18607), .A(n16433), .ZN(P3_U2634) );
  AOI21_X1 U19614 ( .B1(n18626), .B2(n18629), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16435) );
  AOI22_X1 U19615 ( .A1(n18745), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16435), 
        .B2(n18763), .ZN(P3_U2635) );
  OAI21_X1 U19616 ( .B1(n18613), .B2(BS16), .A(n18701), .ZN(n18699) );
  OAI21_X1 U19617 ( .B1(n18701), .B2(n16436), .A(n18699), .ZN(P3_U2636) );
  INV_X1 U19618 ( .A(n16437), .ZN(n16438) );
  NOR3_X1 U19619 ( .A1(n16439), .A2(n18535), .A3(n16438), .ZN(n18542) );
  NOR2_X1 U19620 ( .A1(n18542), .A2(n18603), .ZN(n18746) );
  OAI21_X1 U19621 ( .B1(n18746), .B2(n18096), .A(n16440), .ZN(P3_U2637) );
  NOR4_X1 U19622 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16444) );
  NOR4_X1 U19623 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16443) );
  NOR4_X1 U19624 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16442) );
  NOR4_X1 U19625 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16441) );
  NAND4_X1 U19626 ( .A1(n16444), .A2(n16443), .A3(n16442), .A4(n16441), .ZN(
        n16450) );
  NOR4_X1 U19627 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16448) );
  AOI211_X1 U19628 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16447) );
  NOR4_X1 U19629 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16446) );
  NOR4_X1 U19630 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16445) );
  NAND4_X1 U19631 ( .A1(n16448), .A2(n16447), .A3(n16446), .A4(n16445), .ZN(
        n16449) );
  NOR2_X1 U19632 ( .A1(n16450), .A2(n16449), .ZN(n18739) );
  INV_X1 U19633 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18694) );
  NOR3_X1 U19634 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16452) );
  OAI21_X1 U19635 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16452), .A(n18739), .ZN(
        n16451) );
  OAI21_X1 U19636 ( .B1(n18739), .B2(n18694), .A(n16451), .ZN(P3_U2638) );
  INV_X1 U19637 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18735) );
  INV_X1 U19638 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18700) );
  AOI21_X1 U19639 ( .B1(n18735), .B2(n18700), .A(n16452), .ZN(n16453) );
  INV_X1 U19640 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18691) );
  INV_X1 U19641 ( .A(n18739), .ZN(n18742) );
  AOI22_X1 U19642 ( .A1(n18739), .A2(n16453), .B1(n18691), .B2(n18742), .ZN(
        P3_U2639) );
  NOR3_X1 U19643 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18686), .A3(n16454), 
        .ZN(n16455) );
  AOI21_X1 U19644 ( .B1(n16794), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16455), .ZN(
        n16464) );
  INV_X1 U19645 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16804) );
  NAND2_X1 U19646 ( .A1(n16297), .A2(n16743), .ZN(n16707) );
  NOR3_X1 U19647 ( .A1(n16457), .A2(n16456), .A3(n16707), .ZN(n16461) );
  INV_X1 U19648 ( .A(n16458), .ZN(n16459) );
  AOI21_X1 U19649 ( .B1(n16477), .B2(n16459), .A(n18688), .ZN(n16460) );
  AOI211_X1 U19650 ( .C1(n16462), .C2(n16804), .A(n16461), .B(n16460), .ZN(
        n16463) );
  INV_X1 U19651 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18683) );
  AOI211_X1 U19652 ( .C1(n16468), .C2(n16467), .A(n16466), .B(n18610), .ZN(
        n16472) );
  NAND3_X1 U19653 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16491), .ZN(n16470) );
  OAI22_X1 U19654 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16470), .B1(n16469), 
        .B2(n16724), .ZN(n16471) );
  INV_X1 U19655 ( .A(n16473), .ZN(n16474) );
  OAI21_X1 U19656 ( .B1(n16478), .B2(n16835), .A(n16474), .ZN(n16475) );
  OAI211_X1 U19657 ( .C1(n16477), .C2(n18683), .A(n16476), .B(n16475), .ZN(
        P3_U2642) );
  AOI22_X1 U19658 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16779), .B1(
        n16794), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16485) );
  AOI211_X1 U19659 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16492), .A(n16478), .B(
        n16786), .ZN(n16481) );
  AOI211_X1 U19660 ( .C1(n17411), .C2(n16479), .A(n9764), .B(n18610), .ZN(
        n16480) );
  AOI211_X1 U19661 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16503), .A(n16481), 
        .B(n16480), .ZN(n16484) );
  NAND2_X1 U19662 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16482) );
  OAI211_X1 U19663 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16491), .B(n16482), .ZN(n16483) );
  NAND3_X1 U19664 ( .A1(n16485), .A2(n16484), .A3(n16483), .ZN(P3_U2643) );
  INV_X1 U19665 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18679) );
  AOI211_X1 U19666 ( .C1(n16488), .C2(n16487), .A(n16486), .B(n18610), .ZN(
        n16490) );
  OAI22_X1 U19667 ( .A1(n9757), .A2(n16724), .B1(n16783), .B2(n16846), .ZN(
        n16489) );
  AOI211_X1 U19668 ( .C1(n16491), .C2(n18679), .A(n16490), .B(n16489), .ZN(
        n16494) );
  OAI211_X1 U19669 ( .C1(n16498), .C2(n16846), .A(n16793), .B(n16492), .ZN(
        n16493) );
  OAI211_X1 U19670 ( .C1(n16495), .C2(n18679), .A(n16494), .B(n16493), .ZN(
        P3_U2644) );
  AOI22_X1 U19671 ( .A1(n16794), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16497), 
        .B2(n16496), .ZN(n16505) );
  AOI211_X1 U19672 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16514), .A(n16498), .B(
        n16786), .ZN(n16502) );
  AOI211_X1 U19673 ( .C1(n17434), .C2(n16500), .A(n16499), .B(n18610), .ZN(
        n16501) );
  AOI211_X1 U19674 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16503), .A(n16502), 
        .B(n16501), .ZN(n16504) );
  OAI211_X1 U19675 ( .C1(n17432), .C2(n16724), .A(n16505), .B(n16504), .ZN(
        P3_U2645) );
  INV_X1 U19676 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18673) );
  OAI21_X1 U19677 ( .B1(n16519), .B2(n16784), .A(n16795), .ZN(n16530) );
  AOI21_X1 U19678 ( .B1(n16766), .B2(n18673), .A(n16530), .ZN(n16517) );
  AOI211_X1 U19679 ( .C1(n16508), .C2(n16507), .A(n16506), .B(n18610), .ZN(
        n16513) );
  NOR3_X1 U19680 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16784), .A3(n16509), 
        .ZN(n16512) );
  INV_X1 U19681 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16510) );
  OAI22_X1 U19682 ( .A1(n16510), .A2(n16724), .B1(n16783), .B2(n16852), .ZN(
        n16511) );
  NOR3_X1 U19683 ( .A1(n16513), .A2(n16512), .A3(n16511), .ZN(n16516) );
  OAI211_X1 U19684 ( .C1(n16520), .C2(n16852), .A(n16793), .B(n16514), .ZN(
        n16515) );
  OAI211_X1 U19685 ( .C1(n16517), .C2(n18675), .A(n16516), .B(n16515), .ZN(
        P3_U2646) );
  NOR2_X1 U19686 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16784), .ZN(n16518) );
  AOI22_X1 U19687 ( .A1(n16794), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16519), 
        .B2(n16518), .ZN(n16526) );
  AOI211_X1 U19688 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16531), .A(n16520), .B(
        n16786), .ZN(n16524) );
  AOI211_X1 U19689 ( .C1(n17459), .C2(n16522), .A(n16521), .B(n18610), .ZN(
        n16523) );
  AOI211_X1 U19690 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16530), .A(n16524), 
        .B(n16523), .ZN(n16525) );
  OAI211_X1 U19691 ( .C1(n17463), .C2(n16724), .A(n16526), .B(n16525), .ZN(
        P3_U2647) );
  NAND2_X1 U19692 ( .A1(n16591), .A2(n18671), .ZN(n16537) );
  AOI211_X1 U19693 ( .C1(n17473), .C2(n9652), .A(n16527), .B(n18610), .ZN(
        n16529) );
  OAI22_X1 U19694 ( .A1(n17469), .A2(n16724), .B1(n16783), .B2(n16532), .ZN(
        n16528) );
  AOI211_X1 U19695 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16530), .A(n16529), 
        .B(n16528), .ZN(n16535) );
  OAI211_X1 U19696 ( .C1(n16533), .C2(n16532), .A(n16793), .B(n16531), .ZN(
        n16534) );
  OAI211_X1 U19697 ( .C1(n16537), .C2(n16536), .A(n16535), .B(n16534), .ZN(
        P3_U2648) );
  INV_X1 U19698 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20839) );
  AOI211_X1 U19699 ( .C1(n17499), .C2(n16539), .A(n16538), .B(n18610), .ZN(
        n16544) );
  OAI211_X1 U19700 ( .C1(n16541), .C2(n16900), .A(n16793), .B(n16540), .ZN(
        n16542) );
  OAI21_X1 U19701 ( .B1(n16900), .B2(n16783), .A(n16542), .ZN(n16543) );
  AOI211_X1 U19702 ( .C1(n16779), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16544), .B(n16543), .ZN(n16545) );
  OAI221_X1 U19703 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16547), .C1(n20839), 
        .C2(n16546), .A(n16545), .ZN(P3_U2650) );
  INV_X1 U19704 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17534) );
  NAND2_X1 U19705 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16548), .ZN(
        n17519) );
  NOR2_X1 U19706 ( .A1(n17534), .A2(n17519), .ZN(n16558) );
  OAI21_X1 U19707 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16558), .A(
        n17485), .ZN(n17521) );
  NOR2_X1 U19708 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17755), .ZN(
        n16775) );
  AOI21_X1 U19709 ( .B1(n16548), .B2(n16775), .A(n9763), .ZN(n16561) );
  AOI21_X1 U19710 ( .B1(n16297), .B2(n17534), .A(n16561), .ZN(n16549) );
  XNOR2_X1 U19711 ( .A(n17521), .B(n16549), .ZN(n16557) );
  OAI211_X1 U19712 ( .C1(n16562), .C2(n16918), .A(n16793), .B(n16550), .ZN(
        n16551) );
  OAI211_X1 U19713 ( .C1(n16783), .C2(n16918), .A(n9600), .B(n16551), .ZN(
        n16555) );
  INV_X1 U19714 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20812) );
  XOR2_X1 U19715 ( .A(n20812), .B(P3_REIP_REG_18__SCAN_IN), .Z(n16553) );
  OAI21_X1 U19716 ( .B1(n16552), .B2(n16603), .A(n16792), .ZN(n16573) );
  OAI22_X1 U19717 ( .A1(n16568), .A2(n16553), .B1(n16573), .B2(n20812), .ZN(
        n16554) );
  AOI211_X1 U19718 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n16779), .A(
        n16555), .B(n16554), .ZN(n16556) );
  OAI21_X1 U19719 ( .B1(n16557), .B2(n18610), .A(n16556), .ZN(P3_U2652) );
  INV_X1 U19720 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18663) );
  AOI21_X1 U19721 ( .B1(n17534), .B2(n17519), .A(n16558), .ZN(n17537) );
  INV_X1 U19722 ( .A(n17537), .ZN(n16560) );
  INV_X1 U19723 ( .A(n16561), .ZN(n16559) );
  AOI221_X1 U19724 ( .B1(n17537), .B2(n16561), .C1(n16560), .C2(n16559), .A(
        n18610), .ZN(n16566) );
  AOI211_X1 U19725 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16570), .A(n16562), .B(
        n16786), .ZN(n16565) );
  INV_X1 U19726 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16563) );
  OAI22_X1 U19727 ( .A1(n17534), .A2(n16724), .B1(n16783), .B2(n16563), .ZN(
        n16564) );
  NOR4_X1 U19728 ( .A1(n13104), .A2(n16566), .A3(n16565), .A4(n16564), .ZN(
        n16567) );
  OAI221_X1 U19729 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16568), .C1(n18663), 
        .C2(n16573), .A(n16567), .ZN(P3_U2653) );
  INV_X1 U19730 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17573) );
  INV_X1 U19731 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16585) );
  INV_X1 U19732 ( .A(n17555), .ZN(n16593) );
  NOR3_X1 U19733 ( .A1(n17573), .A2(n16585), .A3(n16593), .ZN(n16580) );
  OAI21_X1 U19734 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16580), .A(
        n17519), .ZN(n17545) );
  INV_X1 U19735 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16772) );
  AOI21_X1 U19736 ( .B1(n16772), .B2(n16580), .A(n9763), .ZN(n16569) );
  XOR2_X1 U19737 ( .A(n17545), .B(n16569), .Z(n16579) );
  OAI211_X1 U19738 ( .C1(n16583), .C2(n16572), .A(n16793), .B(n16570), .ZN(
        n16571) );
  OAI211_X1 U19739 ( .C1(n16783), .C2(n16572), .A(n9600), .B(n16571), .ZN(
        n16577) );
  INV_X1 U19740 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18659) );
  NAND2_X1 U19741 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16591), .ZN(n16590) );
  NOR2_X1 U19742 ( .A1(n18659), .A2(n16590), .ZN(n16575) );
  INV_X1 U19743 ( .A(n16573), .ZN(n16574) );
  MUX2_X1 U19744 ( .A(n16575), .B(n16574), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n16576) );
  AOI211_X1 U19745 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n16779), .A(
        n16577), .B(n16576), .ZN(n16578) );
  OAI21_X1 U19746 ( .B1(n18610), .B2(n16579), .A(n16578), .ZN(P3_U2654) );
  INV_X1 U19747 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18657) );
  OAI21_X1 U19748 ( .B1(n18657), .B2(n16603), .A(n16792), .ZN(n16602) );
  INV_X1 U19749 ( .A(n16581), .ZN(n16598) );
  AOI21_X1 U19750 ( .B1(n16585), .B2(n16592), .A(n16580), .ZN(n16582) );
  INV_X1 U19751 ( .A(n16582), .ZN(n17561) );
  AOI221_X1 U19752 ( .B1(n16598), .B2(n16582), .C1(n16581), .C2(n17561), .A(
        n18610), .ZN(n16588) );
  AOI211_X1 U19753 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16594), .A(n16583), .B(
        n16786), .ZN(n16587) );
  INV_X1 U19754 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16584) );
  OAI22_X1 U19755 ( .A1(n16585), .A2(n16724), .B1(n16783), .B2(n16584), .ZN(
        n16586) );
  NOR4_X1 U19756 ( .A1(n17892), .A2(n16588), .A3(n16587), .A4(n16586), .ZN(
        n16589) );
  OAI221_X1 U19757 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16590), .C1(n18659), 
        .C2(n16602), .A(n16589), .ZN(P3_U2655) );
  NOR2_X1 U19758 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16591), .ZN(n16601) );
  NOR2_X1 U19759 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18610), .ZN(
        n16701) );
  NAND2_X1 U19760 ( .A1(n16743), .A2(n9763), .ZN(n16778) );
  INV_X1 U19761 ( .A(n16778), .ZN(n16700) );
  NOR2_X1 U19762 ( .A1(n16701), .A2(n16700), .ZN(n16791) );
  OAI21_X1 U19763 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17555), .A(
        n16592), .ZN(n17570) );
  AOI211_X1 U19764 ( .C1(n16297), .C2(n16593), .A(n16791), .B(n17570), .ZN(
        n16597) );
  OAI211_X1 U19765 ( .C1(n16604), .C2(n16972), .A(n16793), .B(n16594), .ZN(
        n16595) );
  OAI211_X1 U19766 ( .C1(n16783), .C2(n16972), .A(n9600), .B(n16595), .ZN(
        n16596) );
  AOI211_X1 U19767 ( .C1(n16779), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16597), .B(n16596), .ZN(n16600) );
  NAND3_X1 U19768 ( .A1(n16598), .A2(n16743), .A3(n17570), .ZN(n16599) );
  OAI211_X1 U19769 ( .C1(n16602), .C2(n16601), .A(n16600), .B(n16599), .ZN(
        P3_U2656) );
  NAND2_X1 U19770 ( .A1(n16792), .A2(n16603), .ZN(n16615) );
  AOI211_X1 U19771 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16623), .A(n16604), .B(
        n16786), .ZN(n16612) );
  INV_X1 U19772 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16605) );
  OAI22_X1 U19773 ( .A1(n17586), .A2(n16724), .B1(n16783), .B2(n16605), .ZN(
        n16611) );
  NAND2_X1 U19774 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16606), .ZN(
        n16644) );
  INV_X1 U19775 ( .A(n16644), .ZN(n17596) );
  NAND2_X1 U19776 ( .A1(n17600), .A2(n17596), .ZN(n16619) );
  AOI21_X1 U19777 ( .B1(n17586), .B2(n16619), .A(n17555), .ZN(n17589) );
  NAND2_X1 U19778 ( .A1(n16606), .A2(n16775), .ZN(n16632) );
  OAI21_X1 U19779 ( .B1(n16607), .B2(n16632), .A(n16297), .ZN(n16618) );
  INV_X1 U19780 ( .A(n16618), .ZN(n16609) );
  INV_X1 U19781 ( .A(n17589), .ZN(n16608) );
  AOI221_X1 U19782 ( .B1(n17589), .B2(n16609), .C1(n16608), .C2(n16618), .A(
        n18610), .ZN(n16610) );
  NOR4_X1 U19783 ( .A1(n13104), .A2(n16612), .A3(n16611), .A4(n16610), .ZN(
        n16613) );
  OAI221_X1 U19784 ( .B1(n16615), .B2(n18656), .C1(n16615), .C2(n16614), .A(
        n16613), .ZN(P3_U2657) );
  OR2_X1 U19785 ( .A1(n16764), .A2(n16616), .ZN(n16687) );
  OAI21_X1 U19786 ( .B1(n16617), .B2(n16687), .A(n16792), .ZN(n16647) );
  INV_X1 U19787 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18651) );
  NAND2_X1 U19788 ( .A1(n16766), .A2(n18651), .ZN(n16636) );
  NOR2_X1 U19789 ( .A1(n18610), .A2(n16618), .ZN(n16628) );
  INV_X1 U19790 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16631) );
  NOR2_X1 U19791 ( .A1(n16631), .A2(n16644), .ZN(n16630) );
  OAI21_X1 U19792 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16630), .A(
        n16619), .ZN(n17597) );
  INV_X1 U19793 ( .A(n16630), .ZN(n16620) );
  AOI211_X1 U19794 ( .C1(n16297), .C2(n16620), .A(n16791), .B(n17597), .ZN(
        n16627) );
  NOR3_X1 U19795 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16784), .A3(n16621), 
        .ZN(n16622) );
  AOI211_X1 U19796 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16779), .A(
        n17892), .B(n16622), .ZN(n16625) );
  OAI211_X1 U19797 ( .C1(n16634), .C2(n20860), .A(n16793), .B(n16623), .ZN(
        n16624) );
  OAI211_X1 U19798 ( .C1(n20860), .C2(n16783), .A(n16625), .B(n16624), .ZN(
        n16626) );
  AOI211_X1 U19799 ( .C1(n16628), .C2(n17597), .A(n16627), .B(n16626), .ZN(
        n16629) );
  OAI221_X1 U19800 ( .B1(n18653), .B2(n16647), .C1(n18653), .C2(n16636), .A(
        n16629), .ZN(P3_U2658) );
  AOI22_X1 U19801 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16779), .B1(
        n16794), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16642) );
  AOI21_X1 U19802 ( .B1(n16631), .B2(n16644), .A(n16630), .ZN(n17614) );
  NAND2_X1 U19803 ( .A1(n16297), .A2(n16632), .ZN(n16633) );
  XNOR2_X1 U19804 ( .A(n17614), .B(n16633), .ZN(n16640) );
  AOI211_X1 U19805 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16650), .A(n16634), .B(
        n16786), .ZN(n16639) );
  INV_X1 U19806 ( .A(n16635), .ZN(n16637) );
  OAI21_X1 U19807 ( .B1(n16637), .B2(n16636), .A(n9600), .ZN(n16638) );
  AOI211_X1 U19808 ( .C1(n16640), .C2(n16743), .A(n16639), .B(n16638), .ZN(
        n16641) );
  OAI211_X1 U19809 ( .C1(n18651), .C2(n16647), .A(n16642), .B(n16641), .ZN(
        P3_U2659) );
  NAND3_X1 U19810 ( .A1(n16766), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n16715), 
        .ZN(n16681) );
  INV_X1 U19811 ( .A(n16681), .ZN(n16710) );
  AOI21_X1 U19812 ( .B1(n16643), .B2(n16710), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16648) );
  INV_X1 U19813 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16657) );
  INV_X1 U19814 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17664) );
  INV_X1 U19815 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17676) );
  NOR2_X1 U19816 ( .A1(n17658), .A2(n17676), .ZN(n17661) );
  NAND2_X1 U19817 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17661), .ZN(
        n16689) );
  NOR2_X1 U19818 ( .A1(n17664), .A2(n16689), .ZN(n16679) );
  NAND2_X1 U19819 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16679), .ZN(
        n16666) );
  NOR2_X1 U19820 ( .A1(n16657), .A2(n16666), .ZN(n16654) );
  OAI21_X1 U19821 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16654), .A(
        n16644), .ZN(n17624) );
  INV_X1 U19822 ( .A(n16775), .ZN(n16736) );
  NOR2_X1 U19823 ( .A1(n17658), .A2(n16736), .ZN(n16708) );
  INV_X1 U19824 ( .A(n16708), .ZN(n16690) );
  OAI21_X1 U19825 ( .B1(n17623), .B2(n16690), .A(n16297), .ZN(n16645) );
  XNOR2_X1 U19826 ( .A(n17624), .B(n16645), .ZN(n16646) );
  OAI22_X1 U19827 ( .A1(n16648), .A2(n16647), .B1(n18610), .B2(n16646), .ZN(
        n16649) );
  AOI211_X1 U19828 ( .C1(n16794), .C2(P3_EBX_REG_11__SCAN_IN), .A(n17892), .B(
        n16649), .ZN(n16653) );
  OAI211_X1 U19829 ( .C1(n16656), .C2(n16651), .A(n16793), .B(n16650), .ZN(
        n16652) );
  OAI211_X1 U19830 ( .C1(n16724), .C2(n17626), .A(n16653), .B(n16652), .ZN(
        P3_U2660) );
  AOI21_X1 U19831 ( .B1(n16657), .B2(n16666), .A(n16654), .ZN(n17642) );
  OAI21_X1 U19832 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16666), .A(
        n16297), .ZN(n16655) );
  XOR2_X1 U19833 ( .A(n17642), .B(n16655), .Z(n16665) );
  AOI211_X1 U19834 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16667), .A(n16656), .B(
        n16786), .ZN(n16659) );
  OAI21_X1 U19835 ( .B1(n16657), .B2(n16724), .A(n9600), .ZN(n16658) );
  AOI211_X1 U19836 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16794), .A(n16659), .B(
        n16658), .ZN(n16664) );
  OAI21_X1 U19837 ( .B1(n16661), .B2(n16687), .A(n16792), .ZN(n16660) );
  INV_X1 U19838 ( .A(n16660), .ZN(n16684) );
  NOR2_X1 U19839 ( .A1(n16661), .A2(n16681), .ZN(n16672) );
  XNOR2_X1 U19840 ( .A(P3_REIP_REG_10__SCAN_IN), .B(n18645), .ZN(n16662) );
  AOI22_X1 U19841 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16684), .B1(n16672), 
        .B2(n16662), .ZN(n16663) );
  OAI211_X1 U19842 ( .C1(n18610), .C2(n16665), .A(n16664), .B(n16663), .ZN(
        P3_U2661) );
  NOR2_X1 U19843 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16666), .ZN(
        n16676) );
  INV_X1 U19844 ( .A(n16707), .ZN(n16780) );
  OAI21_X1 U19845 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16679), .A(
        n16666), .ZN(n17653) );
  AOI22_X1 U19846 ( .A1(n16780), .A2(n17653), .B1(n16679), .B2(n16701), .ZN(
        n16675) );
  OAI211_X1 U19847 ( .C1(n16677), .C2(n16669), .A(n16793), .B(n16667), .ZN(
        n16668) );
  OAI211_X1 U19848 ( .C1(n16783), .C2(n16669), .A(n9600), .B(n16668), .ZN(
        n16670) );
  AOI21_X1 U19849 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16779), .A(
        n16670), .ZN(n16674) );
  NOR2_X1 U19850 ( .A1(n17653), .A2(n16778), .ZN(n16671) );
  AOI221_X1 U19851 ( .B1(n16684), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n16672), 
        .C2(n18645), .A(n16671), .ZN(n16673) );
  OAI211_X1 U19852 ( .C1(n16676), .C2(n16675), .A(n16674), .B(n16673), .ZN(
        P3_U2662) );
  AOI211_X1 U19853 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16694), .A(n16677), .B(
        n16786), .ZN(n16678) );
  AOI211_X1 U19854 ( .C1(n16794), .C2(P3_EBX_REG_8__SCAN_IN), .A(n17892), .B(
        n16678), .ZN(n16686) );
  AOI21_X1 U19855 ( .B1(n17664), .B2(n16689), .A(n16679), .ZN(n17666) );
  AOI21_X1 U19856 ( .B1(n17661), .B2(n16775), .A(n9763), .ZN(n16692) );
  OAI21_X1 U19857 ( .B1(n17666), .B2(n16692), .A(n16743), .ZN(n16680) );
  AOI21_X1 U19858 ( .B1(n17666), .B2(n16692), .A(n16680), .ZN(n16683) );
  NAND2_X1 U19859 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16688) );
  NOR3_X1 U19860 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16688), .A3(n16681), .ZN(
        n16682) );
  AOI211_X1 U19861 ( .C1(n16684), .C2(P3_REIP_REG_8__SCAN_IN), .A(n16683), .B(
        n16682), .ZN(n16685) );
  OAI211_X1 U19862 ( .C1(n17664), .C2(n16724), .A(n16686), .B(n16685), .ZN(
        P3_U2663) );
  AND2_X1 U19863 ( .A1(n16792), .A2(n16687), .ZN(n16727) );
  AOI22_X1 U19864 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16727), .B1(n16710), 
        .B2(n16688), .ZN(n16699) );
  INV_X1 U19865 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18641) );
  INV_X1 U19866 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18639) );
  INV_X1 U19867 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17700) );
  NAND2_X1 U19868 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17688), .ZN(
        n16716) );
  NOR2_X1 U19869 ( .A1(n17700), .A2(n16716), .ZN(n16702) );
  OAI21_X1 U19870 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16702), .A(
        n16689), .ZN(n17687) );
  INV_X1 U19871 ( .A(n17687), .ZN(n16693) );
  NAND2_X1 U19872 ( .A1(n16297), .A2(n16690), .ZN(n16691) );
  OAI221_X1 U19873 ( .B1(n16693), .B2(n16692), .C1(n17687), .C2(n16691), .A(
        n16743), .ZN(n16696) );
  OAI211_X1 U19874 ( .C1(n16703), .C2(n17105), .A(n16793), .B(n16694), .ZN(
        n16695) );
  OAI211_X1 U19875 ( .C1(n16724), .C2(n17676), .A(n16696), .B(n16695), .ZN(
        n16697) );
  AOI211_X1 U19876 ( .C1(n16794), .C2(P3_EBX_REG_7__SCAN_IN), .A(n17892), .B(
        n16697), .ZN(n16698) );
  OAI221_X1 U19877 ( .B1(n16699), .B2(n18641), .C1(n16699), .C2(n18639), .A(
        n16698), .ZN(P3_U2664) );
  AOI21_X1 U19878 ( .B1(n16701), .B2(n17700), .A(n16700), .ZN(n16714) );
  AOI21_X1 U19879 ( .B1(n17700), .B2(n16716), .A(n16702), .ZN(n17697) );
  INV_X1 U19880 ( .A(n17697), .ZN(n16713) );
  AOI211_X1 U19881 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16720), .A(n16703), .B(
        n16786), .ZN(n16706) );
  OAI22_X1 U19882 ( .A1(n17700), .A2(n16724), .B1(n16783), .B2(n16704), .ZN(
        n16705) );
  NOR3_X1 U19883 ( .A1(n17892), .A2(n16706), .A3(n16705), .ZN(n16712) );
  NOR3_X1 U19884 ( .A1(n17697), .A2(n16708), .A3(n16707), .ZN(n16709) );
  AOI221_X1 U19885 ( .B1(n16727), .B2(P3_REIP_REG_6__SCAN_IN), .C1(n16710), 
        .C2(n18639), .A(n16709), .ZN(n16711) );
  OAI211_X1 U19886 ( .C1(n16714), .C2(n16713), .A(n16712), .B(n16711), .ZN(
        P3_U2665) );
  AND2_X1 U19887 ( .A1(n16766), .A2(n16715), .ZN(n16726) );
  INV_X1 U19888 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16723) );
  AND2_X1 U19889 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17701), .ZN(
        n16734) );
  OAI21_X1 U19890 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16734), .A(
        n16716), .ZN(n16718) );
  INV_X1 U19891 ( .A(n16718), .ZN(n17709) );
  AOI21_X1 U19892 ( .B1(n16772), .B2(n16734), .A(n9763), .ZN(n16719) );
  INV_X1 U19893 ( .A(n16719), .ZN(n16737) );
  OAI221_X1 U19894 ( .B1(n17709), .B2(n16719), .C1(n16718), .C2(n16737), .A(
        n16743), .ZN(n16722) );
  OAI211_X1 U19895 ( .C1(n16738), .C2(n16729), .A(n16793), .B(n16720), .ZN(
        n16721) );
  OAI211_X1 U19896 ( .C1(n16724), .C2(n16723), .A(n16722), .B(n16721), .ZN(
        n16725) );
  AOI221_X1 U19897 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n16727), .C1(n16726), 
        .C2(n16727), .A(n16725), .ZN(n16728) );
  OAI211_X1 U19898 ( .C1(n16783), .C2(n16729), .A(n16728), .B(n9600), .ZN(
        P3_U2666) );
  AOI21_X1 U19899 ( .B1(n16766), .B2(n16746), .A(n16764), .ZN(n16752) );
  NOR3_X1 U19900 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16784), .A3(n16746), .ZN(
        n16732) );
  NAND2_X1 U19901 ( .A1(n16730), .A2(n18768), .ZN(n16782) );
  OAI221_X1 U19902 ( .B1(n16782), .B2(n17011), .C1(n16782), .C2(n18545), .A(
        n9600), .ZN(n16731) );
  AOI211_X1 U19903 ( .C1(n16779), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16732), .B(n16731), .ZN(n16745) );
  INV_X1 U19904 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16735) );
  NAND2_X1 U19905 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16733), .ZN(
        n16749) );
  AOI21_X1 U19906 ( .B1(n16735), .B2(n16749), .A(n16734), .ZN(n16739) );
  NAND2_X1 U19907 ( .A1(n16733), .A2(n16735), .ZN(n17716) );
  OAI22_X1 U19908 ( .A1(n16739), .A2(n16737), .B1(n16736), .B2(n17716), .ZN(
        n16742) );
  AOI211_X1 U19909 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16755), .A(n16738), .B(
        n16786), .ZN(n16741) );
  INV_X1 U19910 ( .A(n16739), .ZN(n17724) );
  OAI22_X1 U19911 ( .A1(n16783), .A2(n17116), .B1(n17724), .B2(n16778), .ZN(
        n16740) );
  AOI211_X1 U19912 ( .C1(n16743), .C2(n16742), .A(n16741), .B(n16740), .ZN(
        n16744) );
  OAI211_X1 U19913 ( .C1(n16752), .C2(n18635), .A(n16745), .B(n16744), .ZN(
        P3_U2667) );
  NOR2_X1 U19914 ( .A1(n18733), .A2(n18562), .ZN(n18552) );
  OAI21_X1 U19915 ( .B1(n18711), .B2(n18552), .A(n17087), .ZN(n18707) );
  INV_X1 U19916 ( .A(n18707), .ZN(n16748) );
  NAND2_X1 U19917 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16765) );
  NAND2_X1 U19918 ( .A1(n16766), .A2(n16746), .ZN(n16747) );
  OAI22_X1 U19919 ( .A1(n16748), .A2(n16782), .B1(n16765), .B2(n16747), .ZN(
        n16754) );
  INV_X1 U19920 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18633) );
  NOR2_X1 U19921 ( .A1(n17755), .A2(n17747), .ZN(n16773) );
  OAI21_X1 U19922 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16773), .A(
        n16749), .ZN(n17737) );
  INV_X1 U19923 ( .A(n16773), .ZN(n16759) );
  OAI21_X1 U19924 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16759), .A(
        n16297), .ZN(n16750) );
  XNOR2_X1 U19925 ( .A(n17737), .B(n16750), .ZN(n16751) );
  OAI22_X1 U19926 ( .A1(n16752), .A2(n18633), .B1(n18610), .B2(n16751), .ZN(
        n16753) );
  AOI211_X1 U19927 ( .C1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n16779), .A(
        n16754), .B(n16753), .ZN(n16757) );
  OAI211_X1 U19928 ( .C1(n16760), .C2(n16758), .A(n16793), .B(n16755), .ZN(
        n16756) );
  OAI211_X1 U19929 ( .C1(n16758), .C2(n16783), .A(n16757), .B(n16756), .ZN(
        P3_U2668) );
  OAI21_X1 U19930 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16759), .ZN(n17743) );
  INV_X1 U19931 ( .A(n16760), .ZN(n16771) );
  NOR2_X1 U19932 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16761) );
  INV_X1 U19933 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16762) );
  NOR2_X1 U19934 ( .A1(n16761), .A2(n16762), .ZN(n16763) );
  OAI22_X1 U19935 ( .A1(n16786), .A2(n16763), .B1(n16783), .B2(n16762), .ZN(
        n16770) );
  NAND2_X1 U19936 ( .A1(n10651), .A2(n9915), .ZN(n18551) );
  OAI21_X1 U19937 ( .B1(n18562), .B2(n18733), .A(n18551), .ZN(n18716) );
  AOI22_X1 U19938 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16779), .B1(
        n16764), .B2(P3_REIP_REG_2__SCAN_IN), .ZN(n16768) );
  OAI211_X1 U19939 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16766), .B(n16765), .ZN(n16767) );
  OAI211_X1 U19940 ( .C1(n16782), .C2(n18716), .A(n16768), .B(n16767), .ZN(
        n16769) );
  AOI21_X1 U19941 ( .B1(n16771), .B2(n16770), .A(n16769), .ZN(n16777) );
  NAND2_X1 U19942 ( .A1(n16773), .A2(n16772), .ZN(n16774) );
  OAI211_X1 U19943 ( .C1(n16775), .C2(n17743), .A(n16780), .B(n16774), .ZN(
        n16776) );
  OAI211_X1 U19944 ( .C1(n16778), .C2(n17743), .A(n16777), .B(n16776), .ZN(
        P3_U2669) );
  AOI21_X1 U19945 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16780), .A(
        n16779), .ZN(n16790) );
  NOR2_X1 U19946 ( .A1(n16781), .A2(n18556), .ZN(n18724) );
  INV_X1 U19947 ( .A(n16782), .ZN(n18770) );
  INV_X1 U19948 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17132) );
  OAI22_X1 U19949 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16784), .B1(n16783), 
        .B2(n17132), .ZN(n16788) );
  OAI21_X1 U19950 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n16785), .ZN(n17133) );
  OAI22_X1 U19951 ( .A1(n16786), .A2(n17133), .B1(n16795), .B2(n18735), .ZN(
        n16787) );
  AOI211_X1 U19952 ( .C1(n18724), .C2(n18770), .A(n16788), .B(n16787), .ZN(
        n16789) );
  OAI221_X1 U19953 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16791), .C1(
        n17755), .C2(n16790), .A(n16789), .ZN(P3_U2670) );
  AOI22_X1 U19954 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16792), .B1(n18770), 
        .B2(n18733), .ZN(n16798) );
  OAI21_X1 U19955 ( .B1(n16794), .B2(n16793), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16797) );
  NAND3_X1 U19956 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18708), .A3(
        n16795), .ZN(n16796) );
  NAND3_X1 U19957 ( .A1(n16798), .A2(n16797), .A3(n16796), .ZN(P3_U2671) );
  INV_X1 U19958 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16853) );
  NAND4_X1 U19959 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_20__SCAN_IN), .A4(n16899), .ZN(n16799) );
  NOR4_X1 U19960 ( .A1(n16835), .A2(n16853), .A3(n16852), .A4(n16799), .ZN(
        n16800) );
  NAND4_X1 U19961 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16836), .A4(n16800), .ZN(n16803) );
  NOR2_X1 U19962 ( .A1(n16804), .A2(n16803), .ZN(n16834) );
  NAND2_X1 U19963 ( .A1(n17129), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16802) );
  NAND2_X1 U19964 ( .A1(n16834), .A2(n18134), .ZN(n16801) );
  OAI22_X1 U19965 ( .A1(n16834), .A2(n16802), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16801), .ZN(P3_U2672) );
  NAND2_X1 U19966 ( .A1(n16804), .A2(n16803), .ZN(n16805) );
  NAND2_X1 U19967 ( .A1(n16805), .A2(n17121), .ZN(n16833) );
  AOI22_X1 U19968 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n15473), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16806) );
  OAI21_X1 U19969 ( .B1(n16807), .B2(n17061), .A(n16806), .ZN(n16817) );
  AOI22_X1 U19970 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n15471), .ZN(n16815) );
  OAI22_X1 U19971 ( .A1(n16957), .A2(n16995), .B1(n16808), .B2(n16821), .ZN(
        n16813) );
  AOI22_X1 U19972 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n17062), .ZN(n16811) );
  AOI22_X1 U19973 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n17082), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16810) );
  AOI22_X1 U19974 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n16828), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16809) );
  NAND3_X1 U19975 ( .A1(n16811), .A2(n16810), .A3(n16809), .ZN(n16812) );
  AOI211_X1 U19976 ( .C1(n10721), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n16813), .B(n16812), .ZN(n16814) );
  OAI211_X1 U19977 ( .C1(n10692), .C2(n16997), .A(n16815), .B(n16814), .ZN(
        n16816) );
  AOI211_X1 U19978 ( .C1(n9591), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n16817), .B(n16816), .ZN(n16839) );
  NOR2_X1 U19979 ( .A1(n16839), .A2(n16838), .ZN(n16837) );
  AOI22_X1 U19980 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16830) );
  AOI22_X1 U19981 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16819) );
  AOI22_X1 U19982 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16818) );
  OAI211_X1 U19983 ( .C1(n16821), .C2(n16820), .A(n16819), .B(n16818), .ZN(
        n16827) );
  AOI22_X1 U19984 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16825) );
  AOI22_X1 U19985 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16824) );
  AOI22_X1 U19986 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16823) );
  NAND2_X1 U19987 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n16822) );
  NAND4_X1 U19988 ( .A1(n16825), .A2(n16824), .A3(n16823), .A4(n16822), .ZN(
        n16826) );
  AOI211_X1 U19989 ( .C1(n16828), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n16827), .B(n16826), .ZN(n16829) );
  OAI211_X1 U19990 ( .C1(n10714), .C2(n16831), .A(n16830), .B(n16829), .ZN(
        n16832) );
  XNOR2_X1 U19991 ( .A(n16837), .B(n16832), .ZN(n17148) );
  OAI22_X1 U19992 ( .A1(n16834), .A2(n16833), .B1(n17148), .B2(n17121), .ZN(
        P3_U2673) );
  NAND2_X1 U19993 ( .A1(n16836), .A2(n16835), .ZN(n16842) );
  AOI21_X1 U19994 ( .B1(n16839), .B2(n16838), .A(n16837), .ZN(n17152) );
  AOI22_X1 U19995 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16840), .B1(n17152), 
        .B2(n17114), .ZN(n16841) );
  OAI21_X1 U19996 ( .B1(n16847), .B2(n16842), .A(n16841), .ZN(P3_U2674) );
  AOI21_X1 U19997 ( .B1(n16844), .B2(n16848), .A(n16843), .ZN(n17162) );
  NAND2_X1 U19998 ( .A1(n17162), .A2(n17114), .ZN(n16845) );
  OAI221_X1 U19999 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16847), .C1(n16846), 
        .C2(n16850), .A(n16845), .ZN(P3_U2676) );
  OAI21_X1 U20000 ( .B1(n16856), .B2(n16849), .A(n16848), .ZN(n17168) );
  INV_X1 U20001 ( .A(n16850), .ZN(n16854) );
  NOR2_X1 U20002 ( .A1(n16852), .A2(n16851), .ZN(n16860) );
  AOI22_X1 U20003 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16854), .B1(n16860), 
        .B2(n16853), .ZN(n16855) );
  OAI21_X1 U20004 ( .B1(n17168), .B2(n17121), .A(n16855), .ZN(P3_U2677) );
  AOI21_X1 U20005 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17129), .A(n16864), .ZN(
        n16859) );
  AOI21_X1 U20006 ( .B1(n16857), .B2(n16861), .A(n16856), .ZN(n17172) );
  INV_X1 U20007 ( .A(n17172), .ZN(n16858) );
  OAI22_X1 U20008 ( .A1(n16860), .A2(n16859), .B1(n16858), .B2(n17121), .ZN(
        P3_U2678) );
  AOI21_X1 U20009 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17129), .A(n16871), .ZN(
        n16863) );
  OAI21_X1 U20010 ( .B1(n16866), .B2(n16862), .A(n16861), .ZN(n17179) );
  OAI22_X1 U20011 ( .A1(n16864), .A2(n16863), .B1(n17129), .B2(n17179), .ZN(
        P3_U2679) );
  AOI21_X1 U20012 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17129), .A(n16865), .ZN(
        n16870) );
  AOI21_X1 U20013 ( .B1(n16868), .B2(n16867), .A(n16866), .ZN(n17180) );
  INV_X1 U20014 ( .A(n17180), .ZN(n16869) );
  OAI22_X1 U20015 ( .A1(n16871), .A2(n16870), .B1(n17129), .B2(n16869), .ZN(
        P3_U2680) );
  AOI22_X1 U20016 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n9595), .B1(
        P3_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n15471), .ZN(n16882) );
  AOI22_X1 U20017 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16872) );
  OAI21_X1 U20018 ( .B1(n16997), .B2(n17061), .A(n16872), .ZN(n16880) );
  AOI22_X1 U20019 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n17082), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16878) );
  INV_X1 U20020 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U20021 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U20022 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n9591), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16873) );
  OAI211_X1 U20023 ( .C1(n17065), .C2(n16875), .A(n16874), .B(n16873), .ZN(
        n16876) );
  AOI21_X1 U20024 ( .B1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n17091), .A(
        n16876), .ZN(n16877) );
  OAI211_X1 U20025 ( .C1(n16995), .C2(n10732), .A(n16878), .B(n16877), .ZN(
        n16879) );
  AOI211_X1 U20026 ( .C1(n9599), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n16880), .B(n16879), .ZN(n16881) );
  OAI211_X1 U20027 ( .C1(n17109), .C2(n16957), .A(n16882), .B(n16881), .ZN(
        n17185) );
  INV_X1 U20028 ( .A(n17185), .ZN(n16884) );
  NAND3_X1 U20029 ( .A1(n16885), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17121), 
        .ZN(n16883) );
  OAI221_X1 U20030 ( .B1(n16885), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17129), 
        .C2(n16884), .A(n16883), .ZN(P3_U2681) );
  INV_X1 U20031 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20032 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16886) );
  OAI21_X1 U20033 ( .B1(n9598), .B2(n16887), .A(n16886), .ZN(n16898) );
  AOI22_X1 U20034 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16896) );
  OAI22_X1 U20035 ( .A1(n17065), .A2(n16889), .B1(n10692), .B2(n16888), .ZN(
        n16894) );
  AOI22_X1 U20036 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16892) );
  AOI22_X1 U20037 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20038 ( .A1(n16828), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16890) );
  NAND3_X1 U20039 ( .A1(n16892), .A2(n16891), .A3(n16890), .ZN(n16893) );
  AOI211_X1 U20040 ( .C1(n10721), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n16894), .B(n16893), .ZN(n16895) );
  OAI211_X1 U20041 ( .C1(n16957), .C2(n17113), .A(n16896), .B(n16895), .ZN(
        n16897) );
  AOI211_X1 U20042 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n16898), .B(n16897), .ZN(n17192) );
  AOI21_X1 U20043 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16899), .A(n17114), .ZN(
        n16915) );
  AOI22_X1 U20044 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16915), .B1(n16901), 
        .B2(n16900), .ZN(n16902) );
  OAI21_X1 U20045 ( .B1(n17192), .B2(n17129), .A(n16902), .ZN(P3_U2682) );
  AOI22_X1 U20046 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16903), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16904) );
  OAI21_X1 U20047 ( .B1(n9644), .B2(n16905), .A(n16904), .ZN(n16914) );
  AOI22_X1 U20048 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20049 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16906) );
  OAI21_X1 U20050 ( .B1(n10692), .B2(n17013), .A(n16906), .ZN(n16910) );
  AOI22_X1 U20051 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16908) );
  AOI22_X1 U20052 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16907) );
  OAI211_X1 U20053 ( .C1(n10732), .C2(n17010), .A(n16908), .B(n16907), .ZN(
        n16909) );
  AOI211_X1 U20054 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n16910), .B(n16909), .ZN(n16911) );
  OAI211_X1 U20055 ( .C1(n16957), .C2(n17120), .A(n16912), .B(n16911), .ZN(
        n16913) );
  AOI211_X1 U20056 ( .C1(n17014), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n16914), .B(n16913), .ZN(n17199) );
  OAI21_X1 U20057 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16916), .A(n16915), .ZN(
        n16917) );
  OAI21_X1 U20058 ( .B1(n17199), .B2(n17129), .A(n16917), .ZN(P3_U2683) );
  AOI21_X1 U20059 ( .B1(n16918), .B2(n16944), .A(n17114), .ZN(n16930) );
  AOI22_X1 U20060 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20061 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16928) );
  AOI22_X1 U20062 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16828), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16927) );
  OAI22_X1 U20063 ( .A1(n16957), .A2(n17122), .B1(n17087), .B2(n16919), .ZN(
        n16925) );
  AOI22_X1 U20064 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20065 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20066 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16921) );
  NAND2_X1 U20067 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n16920) );
  NAND4_X1 U20068 ( .A1(n16923), .A2(n16922), .A3(n16921), .A4(n16920), .ZN(
        n16924) );
  AOI211_X1 U20069 ( .C1(n10721), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n16925), .B(n16924), .ZN(n16926) );
  NAND4_X1 U20070 ( .A1(n16929), .A2(n16928), .A3(n16927), .A4(n16926), .ZN(
        n17200) );
  AOI22_X1 U20071 ( .A1(n16931), .A2(n16930), .B1(n17200), .B2(n17114), .ZN(
        n16932) );
  INV_X1 U20072 ( .A(n16932), .ZN(P3_U2684) );
  AOI22_X1 U20073 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20074 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20075 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16933) );
  OAI211_X1 U20076 ( .C1(n10732), .C2(n16935), .A(n16934), .B(n16933), .ZN(
        n16941) );
  AOI22_X1 U20077 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20078 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16938) );
  AOI22_X1 U20079 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16937) );
  NAND2_X1 U20080 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n16936) );
  NAND4_X1 U20081 ( .A1(n16939), .A2(n16938), .A3(n16937), .A4(n16936), .ZN(
        n16940) );
  AOI211_X1 U20082 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n16941), .B(n16940), .ZN(n16942) );
  OAI211_X1 U20083 ( .C1(n16957), .C2(n17128), .A(n16943), .B(n16942), .ZN(
        n17205) );
  INV_X1 U20084 ( .A(n17205), .ZN(n16946) );
  OAI21_X1 U20085 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16961), .A(n16944), .ZN(
        n16945) );
  AOI22_X1 U20086 ( .A1(n17114), .A2(n16946), .B1(n16945), .B2(n17121), .ZN(
        P3_U2685) );
  INV_X1 U20087 ( .A(n16973), .ZN(n16947) );
  OAI21_X1 U20088 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16947), .A(n17121), .ZN(
        n16960) );
  AOI22_X1 U20089 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16948) );
  OAI21_X1 U20090 ( .B1(n17087), .B2(n16949), .A(n16948), .ZN(n16959) );
  AOI22_X1 U20091 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16956) );
  INV_X1 U20092 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n20870) );
  OAI22_X1 U20093 ( .A1(n10692), .A2(n20870), .B1(n10732), .B2(n10674), .ZN(
        n16954) );
  AOI22_X1 U20094 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10721), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U20095 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16951) );
  AOI22_X1 U20096 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16950) );
  NAND3_X1 U20097 ( .A1(n16952), .A2(n16951), .A3(n16950), .ZN(n16953) );
  AOI211_X1 U20098 ( .C1(n17089), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n16954), .B(n16953), .ZN(n16955) );
  OAI211_X1 U20099 ( .C1(n16957), .C2(n17130), .A(n16956), .B(n16955), .ZN(
        n16958) );
  AOI211_X1 U20100 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n16959), .B(n16958), .ZN(n17215) );
  OAI22_X1 U20101 ( .A1(n16961), .A2(n16960), .B1(n17215), .B2(n17121), .ZN(
        P3_U2686) );
  AOI22_X1 U20102 ( .A1(n16828), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20103 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20104 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16962) );
  OAI211_X1 U20105 ( .C1(n17065), .C2(n17100), .A(n16963), .B(n16962), .ZN(
        n16969) );
  AOI22_X1 U20106 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10721), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U20107 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20108 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16965) );
  NAND2_X1 U20109 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n16964) );
  NAND4_X1 U20110 ( .A1(n16967), .A2(n16966), .A3(n16965), .A4(n16964), .ZN(
        n16968) );
  AOI211_X1 U20111 ( .C1(n17091), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n16969), .B(n16968), .ZN(n16970) );
  OAI211_X1 U20112 ( .C1(n16957), .C2(n17085), .A(n16971), .B(n16970), .ZN(
        n17216) );
  INV_X1 U20113 ( .A(n17216), .ZN(n16975) );
  NOR3_X1 U20114 ( .A1(n16972), .A2(n16990), .A3(n17040), .ZN(n16993) );
  OAI21_X1 U20115 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n16993), .A(n16973), .ZN(
        n16974) );
  AOI22_X1 U20116 ( .A1(n17114), .A2(n16975), .B1(n16974), .B2(n17121), .ZN(
        P3_U2687) );
  AOI22_X1 U20117 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16976) );
  OAI21_X1 U20118 ( .B1(n9644), .B2(n16977), .A(n16976), .ZN(n16989) );
  AOI22_X1 U20119 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20120 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16978) );
  OAI21_X1 U20121 ( .B1(n10692), .B2(n16979), .A(n16978), .ZN(n16984) );
  AOI22_X1 U20122 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20123 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16980) );
  OAI211_X1 U20124 ( .C1(n10732), .C2(n16982), .A(n16981), .B(n16980), .ZN(
        n16983) );
  AOI211_X1 U20125 ( .C1(n17091), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n16984), .B(n16983), .ZN(n16985) );
  OAI211_X1 U20126 ( .C1(n16957), .C2(n16987), .A(n16986), .B(n16985), .ZN(
        n16988) );
  AOI211_X1 U20127 ( .C1(n17090), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n16989), .B(n16988), .ZN(n17225) );
  NOR2_X1 U20128 ( .A1(n16990), .A2(n17040), .ZN(n16991) );
  OAI21_X1 U20129 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16991), .A(n17129), .ZN(
        n16992) );
  OAI22_X1 U20130 ( .A1(n17225), .A2(n17121), .B1(n16993), .B2(n16992), .ZN(
        P3_U2688) );
  NAND3_X1 U20131 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17025), .ZN(n17008) );
  AOI22_X1 U20132 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n17047), .B1(
        P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n9595), .ZN(n16994) );
  OAI21_X1 U20133 ( .B1(n16995), .B2(n17011), .A(n16994), .ZN(n17006) );
  INV_X1 U20134 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20135 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20136 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n17030), .B1(
        P3_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n17091), .ZN(n16996) );
  OAI21_X1 U20137 ( .B1(n17087), .B2(n16997), .A(n16996), .ZN(n17001) );
  AOI22_X1 U20138 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n15471), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20139 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10721), .B1(
        n17062), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16998) );
  OAI211_X1 U20140 ( .C1(n17109), .C2(n10732), .A(n16999), .B(n16998), .ZN(
        n17000) );
  AOI211_X1 U20141 ( .C1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .C2(n9596), .A(
        n17001), .B(n17000), .ZN(n17002) );
  OAI211_X1 U20142 ( .C1(n10714), .C2(n17004), .A(n17003), .B(n17002), .ZN(
        n17005) );
  AOI211_X1 U20143 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17006), .B(n17005), .ZN(n17233) );
  NAND3_X1 U20144 ( .A1(n17008), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n17121), 
        .ZN(n17007) );
  OAI221_X1 U20145 ( .B1(n17008), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17129), 
        .C2(n17233), .A(n17007), .ZN(P3_U2689) );
  AOI22_X1 U20146 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17009) );
  OAI21_X1 U20147 ( .B1(n17011), .B2(n17010), .A(n17009), .ZN(n17023) );
  AOI22_X1 U20148 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10657), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20149 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17012) );
  OAI21_X1 U20150 ( .B1(n17061), .B2(n17013), .A(n17012), .ZN(n17018) );
  AOI22_X1 U20151 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20152 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17015) );
  OAI211_X1 U20153 ( .C1(n10732), .C2(n17120), .A(n17016), .B(n17015), .ZN(
        n17017) );
  AOI211_X1 U20154 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17018), .B(n17017), .ZN(n17019) );
  OAI211_X1 U20155 ( .C1(n10811), .C2(n17021), .A(n17020), .B(n17019), .ZN(
        n17022) );
  AOI211_X1 U20156 ( .C1(n9591), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n17023), .B(n17022), .ZN(n17239) );
  OAI211_X1 U20157 ( .C1(n17025), .C2(P3_EBX_REG_12__SCAN_IN), .A(n17121), .B(
        n17024), .ZN(n17026) );
  OAI21_X1 U20158 ( .B1(n17239), .B2(n17129), .A(n17026), .ZN(P3_U2691) );
  INV_X1 U20159 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20160 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10657), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20161 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20162 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17028) );
  OAI211_X1 U20163 ( .C1(n10732), .C2(n17122), .A(n17029), .B(n17028), .ZN(
        n17036) );
  AOI22_X1 U20164 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20165 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20166 ( .A1(n17030), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17032) );
  NAND2_X1 U20167 ( .A1(n17091), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n17031) );
  NAND4_X1 U20168 ( .A1(n17034), .A2(n17033), .A3(n17032), .A4(n17031), .ZN(
        n17035) );
  AOI211_X1 U20169 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17036), .B(n17035), .ZN(n17037) );
  OAI211_X1 U20170 ( .C1(n10714), .C2(n17039), .A(n17038), .B(n17037), .ZN(
        n17243) );
  INV_X1 U20171 ( .A(n17243), .ZN(n17042) );
  AND2_X1 U20172 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17057), .ZN(n17059) );
  OAI21_X1 U20173 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17059), .A(n17040), .ZN(
        n17041) );
  AOI22_X1 U20174 ( .A1(n17114), .A2(n17042), .B1(n17041), .B2(n17121), .ZN(
        P3_U2692) );
  AOI22_X1 U20175 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17043) );
  OAI21_X1 U20176 ( .B1(n17087), .B2(n17044), .A(n17043), .ZN(n17056) );
  INV_X1 U20177 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20178 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20179 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17045) );
  OAI21_X1 U20180 ( .B1(n9586), .B2(n17046), .A(n17045), .ZN(n17051) );
  AOI22_X1 U20181 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20182 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17048) );
  OAI211_X1 U20183 ( .C1(n10732), .C2(n17128), .A(n17049), .B(n17048), .ZN(
        n17050) );
  AOI211_X1 U20184 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17051), .B(n17050), .ZN(n17052) );
  OAI211_X1 U20185 ( .C1(n10714), .C2(n17054), .A(n17053), .B(n17052), .ZN(
        n17055) );
  AOI211_X1 U20186 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17056), .B(n17055), .ZN(n17246) );
  OAI21_X1 U20187 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17057), .A(n17121), .ZN(
        n17058) );
  OAI22_X1 U20188 ( .A1(n17246), .A2(n17121), .B1(n17059), .B2(n17058), .ZN(
        P3_U2693) );
  AOI22_X1 U20189 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17060) );
  OAI21_X1 U20190 ( .B1(n17061), .B2(n20870), .A(n17060), .ZN(n17076) );
  AOI22_X1 U20191 ( .A1(n10657), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17072) );
  INV_X1 U20192 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20193 ( .A1(n17062), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17063) );
  OAI21_X1 U20194 ( .B1(n17065), .B2(n17064), .A(n17063), .ZN(n17070) );
  AOI22_X1 U20195 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15471), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20196 ( .A1(n10721), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17067) );
  OAI211_X1 U20197 ( .C1(n10732), .C2(n17130), .A(n17068), .B(n17067), .ZN(
        n17069) );
  AOI211_X1 U20198 ( .C1(n17091), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n17070), .B(n17069), .ZN(n17071) );
  OAI211_X1 U20199 ( .C1(n17074), .C2(n17073), .A(n17072), .B(n17071), .ZN(
        n17075) );
  AOI211_X1 U20200 ( .C1(n17077), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17076), .B(n17075), .ZN(n17250) );
  OAI21_X1 U20201 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17079), .A(n17078), .ZN(
        n17080) );
  AOI22_X1 U20202 ( .A1(n17114), .A2(n17250), .B1(n17080), .B2(n17121), .ZN(
        P3_U2694) );
  NOR2_X1 U20203 ( .A1(n17114), .A2(n17081), .ZN(n17103) );
  AOI22_X1 U20204 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17030), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20205 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17083) );
  OAI21_X1 U20206 ( .B1(n10811), .B2(n17084), .A(n17083), .ZN(n17097) );
  OAI22_X1 U20207 ( .A1(n17087), .A2(n17086), .B1(n10732), .B2(n17085), .ZN(
        n17088) );
  AOI21_X1 U20208 ( .B1(n10657), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n17088), .ZN(n17095) );
  AOI22_X1 U20209 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20210 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20211 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17091), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17092) );
  NAND4_X1 U20212 ( .A1(n17095), .A2(n17094), .A3(n17093), .A4(n17092), .ZN(
        n17096) );
  AOI211_X1 U20213 ( .C1(n10721), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17097), .B(n17096), .ZN(n17098) );
  OAI211_X1 U20214 ( .C1(n9587), .C2(n17100), .A(n17099), .B(n17098), .ZN(
        n17254) );
  AOI22_X1 U20215 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17103), .B1(n17114), .B2(
        n17254), .ZN(n17101) );
  OAI21_X1 U20216 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17102), .A(n17101), .ZN(
        P3_U2695) );
  AOI21_X1 U20217 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17107), .A(n17114), .ZN(
        n17106) );
  AOI21_X1 U20218 ( .B1(n17114), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n17103), .ZN(n17104) );
  AOI21_X1 U20219 ( .B1(n17106), .B2(n17105), .A(n17104), .ZN(P3_U2696) );
  OAI21_X1 U20220 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17107), .A(n17106), .ZN(
        n17108) );
  OAI21_X1 U20221 ( .B1(n17129), .B2(n17109), .A(n17108), .ZN(P3_U2697) );
  OAI21_X1 U20222 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17111), .A(n17110), .ZN(
        n17112) );
  AOI22_X1 U20223 ( .A1(n17114), .A2(n17113), .B1(n17112), .B2(n17121), .ZN(
        P3_U2698) );
  NOR2_X1 U20224 ( .A1(n17115), .A2(n17136), .ZN(n17126) );
  AND2_X1 U20225 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17126), .ZN(n17124) );
  NOR2_X1 U20226 ( .A1(n17114), .A2(n17116), .ZN(n17118) );
  OAI22_X1 U20227 ( .A1(n17124), .A2(n17118), .B1(n17117), .B2(n17136), .ZN(
        n17119) );
  OAI21_X1 U20228 ( .B1(n17129), .B2(n17120), .A(n17119), .ZN(P3_U2699) );
  AOI21_X1 U20229 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17129), .A(n17126), .ZN(
        n17123) );
  OAI22_X1 U20230 ( .A1(n17124), .A2(n17123), .B1(n17122), .B2(n17121), .ZN(
        P3_U2700) );
  AOI221_X1 U20231 ( .B1(n17125), .B2(n17131), .C1(n17259), .C2(n17131), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17127) );
  AOI211_X1 U20232 ( .C1(n17114), .C2(n17128), .A(n17127), .B(n17126), .ZN(
        P3_U2701) );
  OAI222_X1 U20233 ( .A1(n17133), .A2(n17136), .B1(n17132), .B2(n17131), .C1(
        n17130), .C2(n17129), .ZN(P3_U2702) );
  AOI22_X1 U20234 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17114), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17134), .ZN(n17135) );
  OAI21_X1 U20235 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17136), .A(n17135), .ZN(
        P3_U2703) );
  INV_X1 U20236 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17360) );
  INV_X1 U20237 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17352) );
  INV_X1 U20238 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17378) );
  INV_X1 U20239 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17372) );
  INV_X1 U20240 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17370) );
  INV_X1 U20241 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17368) );
  NOR4_X1 U20242 ( .A1(n17378), .A2(n17372), .A3(n17370), .A4(n17368), .ZN(
        n17137) );
  NAND4_X1 U20243 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(n17137), .ZN(n17226) );
  NOR2_X2 U20244 ( .A1(n17286), .A2(n17226), .ZN(n17255) );
  NAND2_X1 U20245 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .ZN(n17227) );
  NAND3_X1 U20246 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n17228) );
  NOR2_X1 U20247 ( .A1(n17227), .A2(n17228), .ZN(n17138) );
  AND2_X1 U20248 ( .A1(n17138), .A2(n9920), .ZN(n17139) );
  INV_X1 U20249 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17399) );
  NAND2_X1 U20250 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n17191) );
  NAND4_X1 U20251 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17140)
         );
  NOR3_X2 U20252 ( .A1(n17218), .A2(n17191), .A3(n17140), .ZN(n17182) );
  NAND2_X1 U20253 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17182), .ZN(n17181) );
  NOR2_X2 U20254 ( .A1(n17259), .A2(n17181), .ZN(n17176) );
  NAND2_X1 U20255 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17176), .ZN(n17175) );
  INV_X1 U20256 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17356) );
  NAND2_X1 U20257 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17159), .ZN(n17155) );
  NAND2_X1 U20258 ( .A1(n17149), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17145) );
  NAND2_X2 U20259 ( .A1(n17141), .A2(n17259), .ZN(n17287) );
  OAI22_X1 U20260 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17186), .B1(n17270), 
        .B2(n17149), .ZN(n17142) );
  AOI22_X1 U20261 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17209), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17142), .ZN(n17143) );
  OAI21_X1 U20262 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17145), .A(n17143), .ZN(
        P3_U2704) );
  NOR2_X2 U20263 ( .A1(n17144), .A2(n17287), .ZN(n17217) );
  AOI22_X1 U20264 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17217), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17209), .ZN(n17147) );
  OAI211_X1 U20265 ( .C1(n17149), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17287), .B(
        n17145), .ZN(n17146) );
  OAI211_X1 U20266 ( .C1(n17148), .C2(n17290), .A(n17147), .B(n17146), .ZN(
        P3_U2705) );
  INV_X1 U20267 ( .A(n17149), .ZN(n17151) );
  OAI21_X1 U20268 ( .B1(n17270), .B2(n17360), .A(n17155), .ZN(n17150) );
  AOI22_X1 U20269 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n17209), .B1(n17151), .B2(
        n17150), .ZN(n17154) );
  AOI22_X1 U20270 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17217), .B1(n17268), .B2(
        n17152), .ZN(n17153) );
  NAND2_X1 U20271 ( .A1(n17154), .A2(n17153), .ZN(P3_U2706) );
  AOI22_X1 U20272 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17217), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17209), .ZN(n17157) );
  OAI211_X1 U20273 ( .C1(n17159), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17287), .B(
        n17155), .ZN(n17156) );
  OAI211_X1 U20274 ( .C1(n17158), .C2(n17290), .A(n17157), .B(n17156), .ZN(
        P3_U2707) );
  INV_X1 U20275 ( .A(n17159), .ZN(n17161) );
  OAI21_X1 U20276 ( .B1(n17270), .B2(n17356), .A(n17165), .ZN(n17160) );
  AOI22_X1 U20277 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17209), .B1(n17161), .B2(
        n17160), .ZN(n17164) );
  AOI22_X1 U20278 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17217), .B1(n17268), .B2(
        n17162), .ZN(n17163) );
  NAND2_X1 U20279 ( .A1(n17164), .A2(n17163), .ZN(P3_U2708) );
  AOI22_X1 U20280 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17217), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17209), .ZN(n17167) );
  OAI211_X1 U20281 ( .C1(n17169), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17287), .B(
        n17165), .ZN(n17166) );
  OAI211_X1 U20282 ( .C1(n17168), .C2(n17290), .A(n17167), .B(n17166), .ZN(
        P3_U2709) );
  INV_X1 U20283 ( .A(n17169), .ZN(n17171) );
  OAI21_X1 U20284 ( .B1(n17270), .B2(n17352), .A(n17175), .ZN(n17170) );
  AOI22_X1 U20285 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n17209), .B1(n17171), .B2(
        n17170), .ZN(n17174) );
  AOI22_X1 U20286 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17217), .B1(n17268), .B2(
        n17172), .ZN(n17173) );
  NAND2_X1 U20287 ( .A1(n17174), .A2(n17173), .ZN(P3_U2710) );
  AOI22_X1 U20288 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17217), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17209), .ZN(n17178) );
  OAI211_X1 U20289 ( .C1(n17176), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17287), .B(
        n17175), .ZN(n17177) );
  OAI211_X1 U20290 ( .C1(n17179), .C2(n17290), .A(n17178), .B(n17177), .ZN(
        P3_U2711) );
  INV_X1 U20291 ( .A(n17209), .ZN(n17221) );
  AOI22_X1 U20292 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17217), .B1(n17268), .B2(
        n17180), .ZN(n17184) );
  OAI211_X1 U20293 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17182), .A(n17287), .B(
        n17181), .ZN(n17183) );
  OAI211_X1 U20294 ( .C1(n17221), .C2(n14999), .A(n17184), .B(n17183), .ZN(
        P3_U2712) );
  INV_X1 U20295 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17340) );
  INV_X1 U20296 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17336) );
  NAND2_X1 U20297 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17210), .ZN(n17206) );
  INV_X1 U20298 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17346) );
  NAND2_X1 U20299 ( .A1(n17201), .A2(n17346), .ZN(n17190) );
  AOI22_X1 U20300 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17209), .B1(n17268), .B2(
        n17185), .ZN(n17189) );
  NAND2_X1 U20301 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17201), .ZN(n17196) );
  NAND2_X1 U20302 ( .A1(n17287), .A2(n17196), .ZN(n17195) );
  OAI21_X1 U20303 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17186), .A(n17195), .ZN(
        n17187) );
  AOI22_X1 U20304 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17217), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17187), .ZN(n17188) );
  OAI211_X1 U20305 ( .C1(n17191), .C2(n17190), .A(n17189), .B(n17188), .ZN(
        P3_U2713) );
  INV_X1 U20306 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17344) );
  OAI22_X1 U20307 ( .A1(n17192), .A2(n17290), .B1(n15016), .B2(n17221), .ZN(
        n17193) );
  AOI21_X1 U20308 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17217), .A(n17193), .ZN(
        n17194) );
  OAI221_X1 U20309 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17196), .C1(n17344), 
        .C2(n17195), .A(n17194), .ZN(P3_U2714) );
  AOI22_X1 U20310 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17217), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17209), .ZN(n17198) );
  OAI211_X1 U20311 ( .C1(n17201), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17287), .B(
        n17196), .ZN(n17197) );
  OAI211_X1 U20312 ( .C1(n17199), .C2(n17290), .A(n17198), .B(n17197), .ZN(
        P3_U2715) );
  AOI22_X1 U20313 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17217), .B1(n17268), .B2(
        n17200), .ZN(n17204) );
  AOI211_X1 U20314 ( .C1(n17340), .C2(n17206), .A(n17201), .B(n17270), .ZN(
        n17202) );
  INV_X1 U20315 ( .A(n17202), .ZN(n17203) );
  OAI211_X1 U20316 ( .C1(n17221), .C2(n19097), .A(n17204), .B(n17203), .ZN(
        P3_U2716) );
  AOI22_X1 U20317 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17217), .B1(n17268), .B2(
        n17205), .ZN(n17208) );
  OAI211_X1 U20318 ( .C1(n17210), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17287), .B(
        n17206), .ZN(n17207) );
  OAI211_X1 U20319 ( .C1(n17221), .C2(n19092), .A(n17208), .B(n17207), .ZN(
        P3_U2717) );
  AOI22_X1 U20320 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17217), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17209), .ZN(n17214) );
  INV_X1 U20321 ( .A(n17218), .ZN(n17212) );
  INV_X1 U20322 ( .A(n17210), .ZN(n17211) );
  OAI211_X1 U20323 ( .C1(n17212), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17287), .B(
        n17211), .ZN(n17213) );
  OAI211_X1 U20324 ( .C1(n17215), .C2(n17290), .A(n17214), .B(n17213), .ZN(
        P3_U2718) );
  AOI22_X1 U20325 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17217), .B1(n17268), .B2(
        n17216), .ZN(n17220) );
  OAI211_X1 U20326 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17222), .A(n17287), .B(
        n17218), .ZN(n17219) );
  OAI211_X1 U20327 ( .C1(n17221), .C2(n19072), .A(n17220), .B(n17219), .ZN(
        P3_U2719) );
  AOI211_X1 U20328 ( .C1(n17399), .C2(n17230), .A(n17270), .B(n17222), .ZN(
        n17223) );
  AOI21_X1 U20329 ( .B1(n17285), .B2(BUF2_REG_15__SCAN_IN), .A(n17223), .ZN(
        n17224) );
  OAI21_X1 U20330 ( .B1(n17225), .B2(n17290), .A(n17224), .ZN(P3_U2720) );
  NOR3_X1 U20331 ( .A1(n17259), .A2(n17286), .A3(n17226), .ZN(n17263) );
  INV_X1 U20332 ( .A(n17263), .ZN(n17258) );
  NOR2_X1 U20333 ( .A1(n17227), .A2(n17258), .ZN(n17252) );
  NAND2_X1 U20334 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17252), .ZN(n17245) );
  NOR3_X1 U20335 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17228), .A3(n17245), .ZN(
        n17229) );
  AOI21_X1 U20336 ( .B1(n17285), .B2(BUF2_REG_14__SCAN_IN), .A(n17229), .ZN(
        n17232) );
  NAND3_X1 U20337 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17287), .A3(n17230), 
        .ZN(n17231) );
  OAI211_X1 U20338 ( .C1(n17233), .C2(n17290), .A(n17232), .B(n17231), .ZN(
        P3_U2721) );
  INV_X1 U20339 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17386) );
  NOR2_X1 U20340 ( .A1(n17386), .A2(n17245), .ZN(n17238) );
  NAND2_X1 U20341 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17238), .ZN(n17237) );
  NAND2_X1 U20342 ( .A1(n17237), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20343 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17285), .B1(n17268), .B2(
        n17234), .ZN(n17235) );
  OAI221_X1 U20344 ( .B1(n17237), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17236), 
        .C2(n17270), .A(n17235), .ZN(P3_U2722) );
  INV_X1 U20345 ( .A(n17237), .ZN(n17241) );
  AOI21_X1 U20346 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17287), .A(n17238), .ZN(
        n17240) );
  OAI222_X1 U20347 ( .A1(n17283), .A2(n17242), .B1(n17241), .B2(n17240), .C1(
        n17290), .C2(n17239), .ZN(P3_U2723) );
  NAND2_X1 U20348 ( .A1(n17287), .A2(n17245), .ZN(n17248) );
  AOI22_X1 U20349 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17285), .B1(n17268), .B2(
        n17243), .ZN(n17244) );
  OAI221_X1 U20350 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17245), .C1(n17386), 
        .C2(n17248), .A(n17244), .ZN(P3_U2724) );
  NOR2_X1 U20351 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17252), .ZN(n17247) );
  OAI222_X1 U20352 ( .A1(n17283), .A2(n17249), .B1(n17248), .B2(n17247), .C1(
        n17290), .C2(n17246), .ZN(P3_U2725) );
  AOI22_X1 U20353 ( .A1(n17263), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17287), .ZN(n17251) );
  OAI222_X1 U20354 ( .A1(n17283), .A2(n17253), .B1(n17252), .B2(n17251), .C1(
        n17290), .C2(n17250), .ZN(P3_U2726) );
  AOI22_X1 U20355 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17285), .B1(n17268), .B2(
        n17254), .ZN(n17257) );
  INV_X1 U20356 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17380) );
  OR3_X1 U20357 ( .A1(n17380), .A2(n17270), .A3(n17255), .ZN(n17256) );
  OAI211_X1 U20358 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n17258), .A(n17257), .B(
        n17256), .ZN(P3_U2727) );
  NAND2_X1 U20359 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17260) );
  NOR2_X1 U20360 ( .A1(n17259), .A2(n17286), .ZN(n17284) );
  NAND3_X1 U20361 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(n17284), .ZN(n17276) );
  NOR2_X1 U20362 ( .A1(n17370), .A2(n17276), .ZN(n17279) );
  NAND2_X1 U20363 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17279), .ZN(n17272) );
  NOR2_X1 U20364 ( .A1(n17260), .A2(n17272), .ZN(n17266) );
  AOI21_X1 U20365 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17287), .A(n17266), .ZN(
        n17262) );
  OAI222_X1 U20366 ( .A1(n17283), .A2(n18131), .B1(n17263), .B2(n17262), .C1(
        n17290), .C2(n17261), .ZN(P3_U2728) );
  INV_X1 U20367 ( .A(n17272), .ZN(n17275) );
  AOI22_X1 U20368 ( .A1(n17275), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17287), .ZN(n17265) );
  OAI222_X1 U20369 ( .A1(n18126), .A2(n17283), .B1(n17266), .B2(n17265), .C1(
        n17290), .C2(n17264), .ZN(P3_U2729) );
  NAND2_X1 U20370 ( .A1(n17272), .A2(P3_EAX_REG_5__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20371 ( .A1(n17285), .A2(BUF2_REG_5__SCAN_IN), .B1(n17268), .B2(
        n17267), .ZN(n17269) );
  OAI221_X1 U20372 ( .B1(n17272), .B2(P3_EAX_REG_5__SCAN_IN), .C1(n17271), 
        .C2(n17270), .A(n17269), .ZN(P3_U2730) );
  AOI21_X1 U20373 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17287), .A(n17279), .ZN(
        n17274) );
  OAI222_X1 U20374 ( .A1(n18118), .A2(n17283), .B1(n17275), .B2(n17274), .C1(
        n17290), .C2(n17273), .ZN(P3_U2731) );
  INV_X1 U20375 ( .A(n17276), .ZN(n17282) );
  AOI21_X1 U20376 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17287), .A(n17282), .ZN(
        n17278) );
  OAI222_X1 U20377 ( .A1(n18114), .A2(n17283), .B1(n17279), .B2(n17278), .C1(
        n17290), .C2(n17277), .ZN(P3_U2732) );
  AOI22_X1 U20378 ( .A1(n17284), .A2(P3_EAX_REG_1__SCAN_IN), .B1(
        P3_EAX_REG_2__SCAN_IN), .B2(n17287), .ZN(n17281) );
  OAI222_X1 U20379 ( .A1(n18109), .A2(n17283), .B1(n17282), .B2(n17281), .C1(
        n17290), .C2(n17280), .ZN(P3_U2733) );
  INV_X1 U20380 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U20381 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17285), .B1(n17284), .B2(
        n17366), .ZN(n17289) );
  NAND3_X1 U20382 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17287), .A3(n17286), .ZN(
        n17288) );
  OAI211_X1 U20383 ( .C1(n17291), .C2(n17290), .A(n17289), .B(n17288), .ZN(
        P3_U2734) );
  NOR2_X1 U20384 ( .A1(n18714), .A2(n17593), .ZN(n18760) );
  INV_X1 U20385 ( .A(n17330), .ZN(n17331) );
  AND2_X1 U20386 ( .A1(n17318), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20387 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17362) );
  NAND2_X1 U20388 ( .A1(n17293), .A2(n10901), .ZN(n17309) );
  AOI22_X1 U20389 ( .A1(n18760), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17294) );
  OAI21_X1 U20390 ( .B1(n17362), .B2(n17309), .A(n17294), .ZN(P3_U2737) );
  AOI22_X1 U20391 ( .A1(n18760), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17295) );
  OAI21_X1 U20392 ( .B1(n17360), .B2(n17309), .A(n17295), .ZN(P3_U2738) );
  INV_X1 U20393 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U20394 ( .A1(n18760), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17296) );
  OAI21_X1 U20395 ( .B1(n17358), .B2(n17309), .A(n17296), .ZN(P3_U2739) );
  AOI22_X1 U20396 ( .A1(n18760), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17297) );
  OAI21_X1 U20397 ( .B1(n17356), .B2(n17309), .A(n17297), .ZN(P3_U2740) );
  INV_X1 U20398 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17354) );
  AOI22_X1 U20399 ( .A1(n18760), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17298) );
  OAI21_X1 U20400 ( .B1(n17354), .B2(n17309), .A(n17298), .ZN(P3_U2741) );
  AOI22_X1 U20401 ( .A1(n18760), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17299) );
  OAI21_X1 U20402 ( .B1(n17352), .B2(n17309), .A(n17299), .ZN(P3_U2742) );
  INV_X1 U20403 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U20404 ( .A1(n18760), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17300) );
  OAI21_X1 U20405 ( .B1(n17350), .B2(n17309), .A(n17300), .ZN(P3_U2743) );
  INV_X1 U20406 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17348) );
  AOI22_X1 U20407 ( .A1(n17327), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17301) );
  OAI21_X1 U20408 ( .B1(n17348), .B2(n17309), .A(n17301), .ZN(P3_U2744) );
  AOI22_X1 U20409 ( .A1(n17327), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17302) );
  OAI21_X1 U20410 ( .B1(n17346), .B2(n17309), .A(n17302), .ZN(P3_U2745) );
  AOI22_X1 U20411 ( .A1(n17327), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17303) );
  OAI21_X1 U20412 ( .B1(n17344), .B2(n17309), .A(n17303), .ZN(P3_U2746) );
  INV_X1 U20413 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20414 ( .A1(n17327), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17304) );
  OAI21_X1 U20415 ( .B1(n17342), .B2(n17309), .A(n17304), .ZN(P3_U2747) );
  AOI22_X1 U20416 ( .A1(n17327), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17305) );
  OAI21_X1 U20417 ( .B1(n17340), .B2(n17309), .A(n17305), .ZN(P3_U2748) );
  INV_X1 U20418 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20419 ( .A1(n17327), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17306) );
  OAI21_X1 U20420 ( .B1(n17338), .B2(n17309), .A(n17306), .ZN(P3_U2749) );
  AOI22_X1 U20421 ( .A1(n17327), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17307) );
  OAI21_X1 U20422 ( .B1(n17336), .B2(n17309), .A(n17307), .ZN(P3_U2750) );
  INV_X1 U20423 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U20424 ( .A1(n17327), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17308) );
  OAI21_X1 U20425 ( .B1(n17334), .B2(n17309), .A(n17308), .ZN(P3_U2751) );
  AOI22_X1 U20426 ( .A1(n17327), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17310) );
  OAI21_X1 U20427 ( .B1(n17399), .B2(n17329), .A(n17310), .ZN(P3_U2752) );
  INV_X1 U20428 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U20429 ( .A1(n17327), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17311) );
  OAI21_X1 U20430 ( .B1(n17394), .B2(n17329), .A(n17311), .ZN(P3_U2753) );
  INV_X1 U20431 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20432 ( .A1(n17327), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17312) );
  OAI21_X1 U20433 ( .B1(n17392), .B2(n17329), .A(n17312), .ZN(P3_U2754) );
  INV_X1 U20434 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20435 ( .A1(n17327), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17313) );
  OAI21_X1 U20436 ( .B1(n17390), .B2(n17329), .A(n17313), .ZN(P3_U2755) );
  AOI22_X1 U20437 ( .A1(n17327), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17314) );
  OAI21_X1 U20438 ( .B1(n17386), .B2(n17329), .A(n17314), .ZN(P3_U2756) );
  INV_X1 U20439 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U20440 ( .A1(n17327), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17315) );
  OAI21_X1 U20441 ( .B1(n17384), .B2(n17329), .A(n17315), .ZN(P3_U2757) );
  INV_X1 U20442 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U20443 ( .A1(n17327), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17316) );
  OAI21_X1 U20444 ( .B1(n17382), .B2(n17329), .A(n17316), .ZN(P3_U2758) );
  AOI22_X1 U20445 ( .A1(n17327), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17317) );
  OAI21_X1 U20446 ( .B1(n17380), .B2(n17329), .A(n17317), .ZN(P3_U2759) );
  AOI22_X1 U20447 ( .A1(n17327), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17318), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17319) );
  OAI21_X1 U20448 ( .B1(n17378), .B2(n17329), .A(n17319), .ZN(P3_U2760) );
  INV_X1 U20449 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17376) );
  AOI22_X1 U20450 ( .A1(n17327), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17320) );
  OAI21_X1 U20451 ( .B1(n17376), .B2(n17329), .A(n17320), .ZN(P3_U2761) );
  INV_X1 U20452 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U20453 ( .A1(n17327), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17321) );
  OAI21_X1 U20454 ( .B1(n17374), .B2(n17329), .A(n17321), .ZN(P3_U2762) );
  AOI22_X1 U20455 ( .A1(n17327), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17322) );
  OAI21_X1 U20456 ( .B1(n17372), .B2(n17329), .A(n17322), .ZN(P3_U2763) );
  AOI22_X1 U20457 ( .A1(n17327), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17323) );
  OAI21_X1 U20458 ( .B1(n17370), .B2(n17329), .A(n17323), .ZN(P3_U2764) );
  AOI22_X1 U20459 ( .A1(n17327), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17324) );
  OAI21_X1 U20460 ( .B1(n17368), .B2(n17329), .A(n17324), .ZN(P3_U2765) );
  AOI22_X1 U20461 ( .A1(n17327), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17325) );
  OAI21_X1 U20462 ( .B1(n17366), .B2(n17329), .A(n17325), .ZN(P3_U2766) );
  AOI22_X1 U20463 ( .A1(n17327), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17326), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17328) );
  OAI21_X1 U20464 ( .B1(n17364), .B2(n17329), .A(n17328), .ZN(P3_U2767) );
  OAI211_X1 U20465 ( .C1(n17332), .C2(n18759), .A(n10902), .B(n17331), .ZN(
        n17395) );
  AOI22_X1 U20466 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17396), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17387), .ZN(n17333) );
  OAI21_X1 U20467 ( .B1(n17334), .B2(n17398), .A(n17333), .ZN(P3_U2768) );
  AOI22_X1 U20468 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17396), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17387), .ZN(n17335) );
  OAI21_X1 U20469 ( .B1(n17336), .B2(n17398), .A(n17335), .ZN(P3_U2769) );
  AOI22_X1 U20470 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17396), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17387), .ZN(n17337) );
  OAI21_X1 U20471 ( .B1(n17338), .B2(n17398), .A(n17337), .ZN(P3_U2770) );
  AOI22_X1 U20472 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17387), .ZN(n17339) );
  OAI21_X1 U20473 ( .B1(n17340), .B2(n17398), .A(n17339), .ZN(P3_U2771) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17387), .ZN(n17341) );
  OAI21_X1 U20475 ( .B1(n17342), .B2(n17398), .A(n17341), .ZN(P3_U2772) );
  AOI22_X1 U20476 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17387), .ZN(n17343) );
  OAI21_X1 U20477 ( .B1(n17344), .B2(n17398), .A(n17343), .ZN(P3_U2773) );
  AOI22_X1 U20478 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17387), .ZN(n17345) );
  OAI21_X1 U20479 ( .B1(n17346), .B2(n17398), .A(n17345), .ZN(P3_U2774) );
  AOI22_X1 U20480 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17387), .ZN(n17347) );
  OAI21_X1 U20481 ( .B1(n17348), .B2(n17398), .A(n17347), .ZN(P3_U2775) );
  AOI22_X1 U20482 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17387), .ZN(n17349) );
  OAI21_X1 U20483 ( .B1(n17350), .B2(n17398), .A(n17349), .ZN(P3_U2776) );
  AOI22_X1 U20484 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17387), .ZN(n17351) );
  OAI21_X1 U20485 ( .B1(n17352), .B2(n17398), .A(n17351), .ZN(P3_U2777) );
  AOI22_X1 U20486 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17387), .ZN(n17353) );
  OAI21_X1 U20487 ( .B1(n17354), .B2(n17398), .A(n17353), .ZN(P3_U2778) );
  AOI22_X1 U20488 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17388), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17387), .ZN(n17355) );
  OAI21_X1 U20489 ( .B1(n17356), .B2(n17398), .A(n17355), .ZN(P3_U2779) );
  AOI22_X1 U20490 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17396), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17387), .ZN(n17357) );
  OAI21_X1 U20491 ( .B1(n17358), .B2(n17398), .A(n17357), .ZN(P3_U2780) );
  AOI22_X1 U20492 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17396), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17387), .ZN(n17359) );
  OAI21_X1 U20493 ( .B1(n17360), .B2(n17398), .A(n17359), .ZN(P3_U2781) );
  AOI22_X1 U20494 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17396), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17387), .ZN(n17361) );
  OAI21_X1 U20495 ( .B1(n17362), .B2(n17398), .A(n17361), .ZN(P3_U2782) );
  AOI22_X1 U20496 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17387), .ZN(n17363) );
  OAI21_X1 U20497 ( .B1(n17364), .B2(n17398), .A(n17363), .ZN(P3_U2783) );
  AOI22_X1 U20498 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17387), .ZN(n17365) );
  OAI21_X1 U20499 ( .B1(n17366), .B2(n17398), .A(n17365), .ZN(P3_U2784) );
  AOI22_X1 U20500 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17387), .ZN(n17367) );
  OAI21_X1 U20501 ( .B1(n17368), .B2(n17398), .A(n17367), .ZN(P3_U2785) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17387), .ZN(n17369) );
  OAI21_X1 U20503 ( .B1(n17370), .B2(n17398), .A(n17369), .ZN(P3_U2786) );
  AOI22_X1 U20504 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17395), .ZN(n17371) );
  OAI21_X1 U20505 ( .B1(n17372), .B2(n17398), .A(n17371), .ZN(P3_U2787) );
  AOI22_X1 U20506 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17395), .ZN(n17373) );
  OAI21_X1 U20507 ( .B1(n17374), .B2(n17398), .A(n17373), .ZN(P3_U2788) );
  AOI22_X1 U20508 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17395), .ZN(n17375) );
  OAI21_X1 U20509 ( .B1(n17376), .B2(n17398), .A(n17375), .ZN(P3_U2789) );
  AOI22_X1 U20510 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17395), .ZN(n17377) );
  OAI21_X1 U20511 ( .B1(n17378), .B2(n17398), .A(n17377), .ZN(P3_U2790) );
  AOI22_X1 U20512 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17395), .ZN(n17379) );
  OAI21_X1 U20513 ( .B1(n17380), .B2(n17398), .A(n17379), .ZN(P3_U2791) );
  AOI22_X1 U20514 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17395), .ZN(n17381) );
  OAI21_X1 U20515 ( .B1(n17382), .B2(n17398), .A(n17381), .ZN(P3_U2792) );
  AOI22_X1 U20516 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17388), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17387), .ZN(n17383) );
  OAI21_X1 U20517 ( .B1(n17384), .B2(n17398), .A(n17383), .ZN(P3_U2793) );
  AOI22_X1 U20518 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17395), .ZN(n17385) );
  OAI21_X1 U20519 ( .B1(n17386), .B2(n17398), .A(n17385), .ZN(P3_U2794) );
  AOI22_X1 U20520 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17388), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17387), .ZN(n17389) );
  OAI21_X1 U20521 ( .B1(n17390), .B2(n17398), .A(n17389), .ZN(P3_U2795) );
  AOI22_X1 U20522 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17395), .ZN(n17391) );
  OAI21_X1 U20523 ( .B1(n17392), .B2(n17398), .A(n17391), .ZN(P3_U2796) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17395), .ZN(n17393) );
  OAI21_X1 U20525 ( .B1(n17394), .B2(n17398), .A(n17393), .ZN(P3_U2797) );
  AOI22_X1 U20526 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17396), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17395), .ZN(n17397) );
  OAI21_X1 U20527 ( .B1(n17399), .B2(n17398), .A(n17397), .ZN(P3_U2798) );
  NAND2_X1 U20528 ( .A1(n17401), .A2(n17402), .ZN(n17415) );
  NAND2_X1 U20529 ( .A1(n17403), .A2(n17612), .ZN(n17409) );
  NAND2_X1 U20530 ( .A1(n18050), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17408) );
  AND3_X1 U20531 ( .A1(n9757), .A2(n17612), .A3(n17404), .ZN(n17423) );
  OAI21_X1 U20532 ( .B1(n17404), .B2(n17721), .A(n17759), .ZN(n17405) );
  AOI21_X1 U20533 ( .B1(n17520), .B2(n17406), .A(n17405), .ZN(n17431) );
  OAI21_X1 U20534 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17446), .A(
        n17431), .ZN(n17424) );
  OAI21_X1 U20535 ( .B1(n17423), .B2(n17424), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17407) );
  OAI211_X1 U20536 ( .C1(n17410), .C2(n17409), .A(n17408), .B(n17407), .ZN(
        n17413) );
  AND2_X1 U20537 ( .A1(n17615), .A2(n17411), .ZN(n17412) );
  AOI22_X1 U20538 ( .A1(n17749), .A2(n17772), .B1(n17627), .B2(n17416), .ZN(
        n17436) );
  NAND2_X1 U20539 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17436), .ZN(
        n17425) );
  OAI211_X1 U20540 ( .C1(n17749), .C2(n17627), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17425), .ZN(n17417) );
  AOI21_X1 U20541 ( .B1(n10791), .B2(n17420), .A(n17419), .ZN(n17778) );
  OAI22_X1 U20542 ( .A1(n9600), .A2(n18679), .B1(n17598), .B2(n17421), .ZN(
        n17422) );
  AOI211_X1 U20543 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17424), .A(
        n17423), .B(n17422), .ZN(n17428) );
  OAI21_X1 U20544 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17426), .A(
        n17425), .ZN(n17427) );
  OAI211_X1 U20545 ( .C1(n17778), .C2(n17622), .A(n17428), .B(n17427), .ZN(
        P3_U2803) );
  AOI21_X1 U20546 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17430), .A(
        n17429), .ZN(n17784) );
  INV_X1 U20547 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18677) );
  NOR2_X1 U20548 ( .A1(n9600), .A2(n18677), .ZN(n17781) );
  AOI221_X1 U20549 ( .B1(n17433), .B2(n17432), .C1(n18201), .C2(n17432), .A(
        n17431), .ZN(n17441) );
  INV_X1 U20550 ( .A(n17434), .ZN(n17435) );
  AOI21_X1 U20551 ( .B1(n17598), .B2(n17446), .A(n17435), .ZN(n17440) );
  NOR2_X1 U20552 ( .A1(n17789), .A2(n17483), .ZN(n17438) );
  INV_X1 U20553 ( .A(n17436), .ZN(n17437) );
  MUX2_X1 U20554 ( .A(n17438), .B(n17437), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17439) );
  NOR4_X1 U20555 ( .A1(n17781), .A2(n17441), .A3(n17440), .A4(n17439), .ZN(
        n17442) );
  OAI21_X1 U20556 ( .B1(n17784), .B2(n17622), .A(n17442), .ZN(P3_U2804) );
  OR2_X1 U20557 ( .A1(n10800), .A2(n17465), .ZN(n17785) );
  NOR2_X1 U20558 ( .A1(n17785), .A2(n17909), .ZN(n17443) );
  XNOR2_X1 U20559 ( .A(n17443), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17795) );
  INV_X1 U20560 ( .A(n17759), .ZN(n17732) );
  NOR2_X1 U20561 ( .A1(n17458), .A2(n18201), .ZN(n17444) );
  AOI211_X1 U20562 ( .C1(n17520), .C2(n17445), .A(n17732), .B(n17444), .ZN(
        n17468) );
  OAI21_X1 U20563 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17446), .A(
        n17468), .ZN(n17462) );
  NOR2_X1 U20564 ( .A1(n9600), .A2(n18675), .ZN(n17798) );
  OAI211_X1 U20565 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17458), .B(n17612), .ZN(n17448) );
  OAI22_X1 U20566 ( .A1(n9919), .A2(n17448), .B1(n17598), .B2(n17447), .ZN(
        n17449) );
  AOI211_X1 U20567 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17462), .A(
        n17798), .B(n17449), .ZN(n17454) );
  INV_X1 U20568 ( .A(n17827), .ZN(n17918) );
  NOR2_X1 U20569 ( .A1(n17918), .A2(n17785), .ZN(n17450) );
  XNOR2_X1 U20570 ( .A(n17450), .B(n17801), .ZN(n17794) );
  AOI21_X1 U20571 ( .B1(n17455), .B2(n10791), .A(n17451), .ZN(n17452) );
  XNOR2_X1 U20572 ( .A(n17452), .B(n17801), .ZN(n17799) );
  AOI22_X1 U20573 ( .A1(n17749), .A2(n17794), .B1(n17671), .B2(n17799), .ZN(
        n17453) );
  OAI211_X1 U20574 ( .C1(n17674), .C2(n17795), .A(n17454), .B(n17453), .ZN(
        P3_U2805) );
  INV_X1 U20575 ( .A(n17455), .ZN(n17456) );
  AOI21_X1 U20576 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17457), .A(
        n17456), .ZN(n17817) );
  AND2_X1 U20577 ( .A1(n17612), .A2(n17458), .ZN(n17464) );
  INV_X1 U20578 ( .A(n17459), .ZN(n17460) );
  OAI22_X1 U20579 ( .A1(n9600), .A2(n18673), .B1(n17598), .B2(n17460), .ZN(
        n17461) );
  AOI221_X1 U20580 ( .B1(n17464), .B2(n17463), .C1(n17462), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17461), .ZN(n17467) );
  NOR2_X1 U20581 ( .A1(n17909), .A2(n17465), .ZN(n17806) );
  NOR2_X1 U20582 ( .A1(n17918), .A2(n17465), .ZN(n17805) );
  OAI22_X1 U20583 ( .A1(n17806), .A2(n17674), .B1(n17805), .B2(n17764), .ZN(
        n17480) );
  NOR2_X1 U20584 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17465), .ZN(
        n17814) );
  AOI22_X1 U20585 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17480), .B1(
        n17549), .B2(n17814), .ZN(n17466) );
  OAI211_X1 U20586 ( .C1(n17817), .C2(n17622), .A(n17467), .B(n17466), .ZN(
        P3_U2806) );
  AOI221_X1 U20587 ( .B1(n17470), .B2(n17469), .C1(n18201), .C2(n17469), .A(
        n17468), .ZN(n17471) );
  NOR2_X1 U20588 ( .A1(n9600), .A2(n18671), .ZN(n17820) );
  AOI211_X1 U20589 ( .C1(n17473), .C2(n17472), .A(n17471), .B(n17820), .ZN(
        n17482) );
  OAI221_X1 U20590 ( .B1(n17476), .B2(n17475), .C1(n17476), .C2(n17500), .A(
        n17474), .ZN(n17484) );
  AOI221_X1 U20591 ( .B1(n10791), .B2(n17477), .C1(n17839), .C2(n17477), .A(
        n17484), .ZN(n17479) );
  INV_X1 U20592 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17478) );
  XNOR2_X1 U20593 ( .A(n17479), .B(n17478), .ZN(n17821) );
  AOI22_X1 U20594 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17480), .B1(
        n17671), .B2(n17821), .ZN(n17481) );
  OAI211_X1 U20595 ( .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17483), .A(
        n17482), .B(n17481), .ZN(P3_U2807) );
  XNOR2_X1 U20596 ( .A(n17839), .B(n17484), .ZN(n17843) );
  INV_X1 U20597 ( .A(n17832), .ZN(n17826) );
  NOR2_X1 U20598 ( .A1(n17749), .A2(n17627), .ZN(n17514) );
  AOI22_X1 U20599 ( .A1(n17749), .A2(n17918), .B1(n17627), .B2(n17909), .ZN(
        n17564) );
  OAI21_X1 U20600 ( .B1(n17826), .B2(n17514), .A(n17564), .ZN(n17503) );
  NAND2_X1 U20601 ( .A1(n17487), .A2(n17612), .ZN(n17497) );
  AOI221_X1 U20602 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17496), .C2(n17490), .A(
        n17497), .ZN(n17492) );
  AOI21_X1 U20603 ( .B1(n17520), .B2(n17485), .A(n17732), .ZN(n17486) );
  OAI21_X1 U20604 ( .B1(n17487), .B2(n17721), .A(n17486), .ZN(n17513) );
  AOI21_X1 U20605 ( .B1(n17508), .B2(n17506), .A(n17513), .ZN(n17495) );
  INV_X1 U20606 ( .A(n9600), .ZN(n18050) );
  AOI22_X1 U20607 ( .A1(n18050), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17615), 
        .B2(n17488), .ZN(n17489) );
  OAI21_X1 U20608 ( .B1(n17495), .B2(n17490), .A(n17489), .ZN(n17491) );
  AOI211_X1 U20609 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17503), .A(
        n17492), .B(n17491), .ZN(n17494) );
  NAND3_X1 U20610 ( .A1(n17826), .A2(n17549), .A3(n17839), .ZN(n17493) );
  OAI211_X1 U20611 ( .C1(n17622), .C2(n17843), .A(n17494), .B(n17493), .ZN(
        P3_U2808) );
  OR2_X1 U20612 ( .A1(n17849), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17856) );
  INV_X1 U20613 ( .A(n17549), .ZN(n17565) );
  NAND2_X1 U20614 ( .A1(n17879), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17846) );
  NAND2_X1 U20615 ( .A1(n18050), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17854) );
  OAI221_X1 U20616 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17497), .C1(
        n17496), .C2(n17495), .A(n17854), .ZN(n17498) );
  AOI21_X1 U20617 ( .B1(n17615), .B2(n17499), .A(n17498), .ZN(n17505) );
  NAND3_X1 U20618 ( .A1(n9624), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17500), .ZN(n17525) );
  OAI22_X1 U20619 ( .A1(n17849), .A2(n17525), .B1(n9645), .B2(n17501), .ZN(
        n17502) );
  XOR2_X1 U20620 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17502), .Z(
        n17853) );
  AOI22_X1 U20621 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17503), .B1(
        n17671), .B2(n17853), .ZN(n17504) );
  OAI211_X1 U20622 ( .C1(n17856), .C2(n17530), .A(n17505), .B(n17504), .ZN(
        P3_U2809) );
  NAND2_X1 U20623 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17861), .ZN(
        n17867) );
  OAI21_X1 U20624 ( .B1(n17507), .B2(n18201), .A(n17506), .ZN(n17512) );
  INV_X1 U20625 ( .A(n17509), .ZN(n17510) );
  AOI21_X1 U20626 ( .B1(n17598), .B2(n17446), .A(n17510), .ZN(n17511) );
  NOR2_X1 U20627 ( .A1(n9600), .A2(n18666), .ZN(n17864) );
  AOI211_X1 U20628 ( .C1(n17513), .C2(n17512), .A(n17511), .B(n17864), .ZN(
        n17518) );
  INV_X1 U20629 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17871) );
  NOR2_X1 U20630 ( .A1(n17871), .A2(n17846), .ZN(n17858) );
  OAI21_X1 U20631 ( .B1(n17514), .B2(n17858), .A(n17564), .ZN(n17527) );
  AOI221_X1 U20632 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17525), 
        .C1(n17871), .C2(n17531), .A(n17515), .ZN(n17516) );
  XNOR2_X1 U20633 ( .A(n17516), .B(n17861), .ZN(n17865) );
  AOI22_X1 U20634 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17527), .B1(
        n17671), .B2(n17865), .ZN(n17517) );
  OAI211_X1 U20635 ( .C1(n17530), .C2(n17867), .A(n17518), .B(n17517), .ZN(
        P3_U2810) );
  INV_X1 U20636 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17522) );
  NAND2_X1 U20637 ( .A1(n16548), .A2(n17612), .ZN(n17535) );
  AOI221_X1 U20638 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n17534), .C2(n17522), .A(
        n17535), .ZN(n17524) );
  OAI21_X1 U20639 ( .B1(n16548), .B2(n17721), .A(n17759), .ZN(n17548) );
  AOI21_X1 U20640 ( .B1(n17520), .B2(n17519), .A(n17548), .ZN(n17533) );
  OAI22_X1 U20641 ( .A1(n17533), .A2(n17522), .B1(n17598), .B2(n17521), .ZN(
        n17523) );
  AOI211_X1 U20642 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n18050), .A(n17524), 
        .B(n17523), .ZN(n17529) );
  OAI21_X1 U20643 ( .B1(n9645), .B2(n17531), .A(n17525), .ZN(n17526) );
  XNOR2_X1 U20644 ( .A(n17526), .B(n17871), .ZN(n17868) );
  AOI22_X1 U20645 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17527), .B1(
        n17671), .B2(n17868), .ZN(n17528) );
  OAI211_X1 U20646 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17530), .A(
        n17529), .B(n17528), .ZN(P3_U2811) );
  OAI21_X1 U20647 ( .B1(n17884), .B2(n10791), .A(n17531), .ZN(n17532) );
  XNOR2_X1 U20648 ( .A(n17532), .B(n9645), .ZN(n17889) );
  NAND2_X1 U20649 ( .A1(n18050), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17887) );
  OAI221_X1 U20650 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17535), .C1(
        n17534), .C2(n17533), .A(n17887), .ZN(n17536) );
  AOI21_X1 U20651 ( .B1(n17615), .B2(n17537), .A(n17536), .ZN(n17540) );
  OAI21_X1 U20652 ( .B1(n17879), .B2(n17565), .A(n17564), .ZN(n17550) );
  NOR2_X1 U20653 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17538), .ZN(
        n17886) );
  AOI22_X1 U20654 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17550), .B1(
        n17549), .B2(n17886), .ZN(n17539) );
  OAI211_X1 U20655 ( .C1(n17622), .C2(n17889), .A(n17540), .B(n17539), .ZN(
        P3_U2812) );
  AOI21_X1 U20656 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17542), .A(
        n17541), .ZN(n17897) );
  OAI21_X1 U20657 ( .B1(n17544), .B2(n18201), .A(n17543), .ZN(n17547) );
  NAND2_X1 U20658 ( .A1(n18050), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17895) );
  OAI21_X1 U20659 ( .B1(n17744), .B2(n17545), .A(n17895), .ZN(n17546) );
  AOI21_X1 U20660 ( .B1(n17548), .B2(n17547), .A(n17546), .ZN(n17552) );
  NOR2_X1 U20661 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10794), .ZN(
        n17894) );
  AOI22_X1 U20662 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17550), .B1(
        n17549), .B2(n17894), .ZN(n17551) );
  OAI211_X1 U20663 ( .C1(n17897), .C2(n17622), .A(n17552), .B(n17551), .ZN(
        P3_U2813) );
  AOI22_X1 U20664 ( .A1(n17629), .A2(n17553), .B1(n9631), .B2(n10791), .ZN(
        n17554) );
  XNOR2_X1 U20665 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17554), .ZN(
        n17905) );
  OAI21_X1 U20666 ( .B1(n17732), .B2(n17556), .A(n17689), .ZN(n17585) );
  OAI21_X1 U20667 ( .B1(n17555), .B2(n17593), .A(n17585), .ZN(n17572) );
  AOI22_X1 U20668 ( .A1(n18050), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17572), .ZN(n17560) );
  NOR2_X1 U20669 ( .A1(n17557), .A2(n17556), .ZN(n17574) );
  OAI211_X1 U20670 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17574), .B(n17558), .ZN(n17559) );
  OAI211_X1 U20671 ( .C1(n17598), .C2(n17561), .A(n17560), .B(n17559), .ZN(
        n17562) );
  AOI21_X1 U20672 ( .B1(n17671), .B2(n17905), .A(n17562), .ZN(n17563) );
  OAI221_X1 U20673 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17565), 
        .C1(n10794), .C2(n17564), .A(n17563), .ZN(P3_U2814) );
  NOR2_X1 U20674 ( .A1(n17575), .A2(n17605), .ZN(n17567) );
  AOI21_X1 U20675 ( .B1(n17953), .B2(n17567), .A(n17566), .ZN(n17568) );
  AOI221_X1 U20676 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17945), 
        .C1(n10791), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17568), .ZN(
        n17569) );
  XNOR2_X1 U20677 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17569), .ZN(
        n17921) );
  OAI22_X1 U20678 ( .A1(n9600), .A2(n18657), .B1(n17598), .B2(n17570), .ZN(
        n17571) );
  AOI221_X1 U20679 ( .B1(n17574), .B2(n17573), .C1(n17572), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17571), .ZN(n17579) );
  NOR2_X1 U20680 ( .A1(n17827), .A2(n17764), .ZN(n17577) );
  NOR2_X1 U20681 ( .A1(n17965), .A2(n17926), .ZN(n17603) );
  INV_X1 U20682 ( .A(n17603), .ZN(n17941) );
  OR2_X1 U20683 ( .A1(n17575), .A2(n17941), .ZN(n17584) );
  NAND2_X1 U20684 ( .A1(n17899), .A2(n17584), .ZN(n17917) );
  INV_X1 U20685 ( .A(n17909), .ZN(n17828) );
  NOR2_X1 U20686 ( .A1(n17828), .A2(n17674), .ZN(n17576) );
  NAND2_X1 U20687 ( .A1(n17969), .A2(n17902), .ZN(n17580) );
  NAND2_X1 U20688 ( .A1(n17899), .A2(n17580), .ZN(n17908) );
  AOI22_X1 U20689 ( .A1(n17577), .A2(n17917), .B1(n17576), .B2(n17908), .ZN(
        n17578) );
  OAI211_X1 U20690 ( .C1(n17622), .C2(n17921), .A(n17579), .B(n17578), .ZN(
        P3_U2815) );
  OAI221_X1 U20691 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17944), .A(n17580), .ZN(
        n17929) );
  INV_X1 U20692 ( .A(n17629), .ZN(n17647) );
  INV_X1 U20693 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17581) );
  NOR2_X1 U20694 ( .A1(n17926), .A2(n17581), .ZN(n17922) );
  INV_X1 U20695 ( .A(n17922), .ZN(n17925) );
  OAI21_X1 U20696 ( .B1(n17647), .B2(n17925), .A(n17582), .ZN(n17583) );
  XNOR2_X1 U20697 ( .A(n17583), .B(n17932), .ZN(n17934) );
  OAI221_X1 U20698 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17603), .A(n17584), .ZN(
        n17928) );
  AOI221_X1 U20699 ( .B1(n17587), .B2(n17586), .C1(n18201), .C2(n17586), .A(
        n17585), .ZN(n17588) );
  AOI21_X1 U20700 ( .B1(n17589), .B2(n17472), .A(n17588), .ZN(n17590) );
  NAND2_X1 U20701 ( .A1(n18050), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n17935) );
  OAI211_X1 U20702 ( .C1(n17764), .C2(n17928), .A(n17590), .B(n17935), .ZN(
        n17591) );
  AOI21_X1 U20703 ( .B1(n17671), .B2(n17934), .A(n17591), .ZN(n17592) );
  OAI21_X1 U20704 ( .B1(n17674), .B2(n17929), .A(n17592), .ZN(P3_U2816) );
  OR2_X1 U20705 ( .A1(n17926), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17950) );
  OAI21_X1 U20706 ( .B1(n17721), .B2(n16606), .A(n17593), .ZN(n17594) );
  INV_X1 U20707 ( .A(n17594), .ZN(n17595) );
  OAI21_X1 U20708 ( .B1(n17596), .B2(n17595), .A(n17759), .ZN(n17613) );
  NOR2_X1 U20709 ( .A1(n9600), .A2(n18653), .ZN(n17602) );
  OAI211_X1 U20710 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n16606), .B(n17612), .ZN(n17599) );
  OAI22_X1 U20711 ( .A1(n17600), .A2(n17599), .B1(n17598), .B2(n17597), .ZN(
        n17601) );
  AOI211_X1 U20712 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17613), .A(
        n17602), .B(n17601), .ZN(n17609) );
  OAI22_X1 U20713 ( .A1(n17603), .A2(n17764), .B1(n17944), .B2(n17674), .ZN(
        n17619) );
  INV_X1 U20714 ( .A(n17604), .ZN(n17610) );
  OAI22_X1 U20715 ( .A1(n9624), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n17605), .B2(n17926), .ZN(n17606) );
  OAI21_X1 U20716 ( .B1(n9624), .B2(n17610), .A(n17606), .ZN(n17607) );
  XNOR2_X1 U20717 ( .A(n17607), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17938) );
  AOI22_X1 U20718 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17619), .B1(
        n17671), .B2(n17938), .ZN(n17608) );
  OAI211_X1 U20719 ( .C1(n17657), .C2(n17950), .A(n17609), .B(n17608), .ZN(
        P3_U2817) );
  AOI21_X1 U20720 ( .B1(n17629), .B2(n17953), .A(n17610), .ZN(n17611) );
  XNOR2_X1 U20721 ( .A(n17611), .B(n17945), .ZN(n17961) );
  NAND2_X1 U20722 ( .A1(n16606), .A2(n17612), .ZN(n17617) );
  AOI22_X1 U20723 ( .A1(n17615), .A2(n17614), .B1(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17613), .ZN(n17616) );
  NAND2_X1 U20724 ( .A1(n18050), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17958) );
  OAI211_X1 U20725 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17617), .A(
        n17616), .B(n17958), .ZN(n17618) );
  AOI21_X1 U20726 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17619), .A(
        n17618), .ZN(n17621) );
  INV_X1 U20727 ( .A(n17657), .ZN(n17635) );
  NAND3_X1 U20728 ( .A1(n17953), .A2(n17945), .A3(n17635), .ZN(n17620) );
  OAI211_X1 U20729 ( .C1(n17961), .C2(n17622), .A(n17621), .B(n17620), .ZN(
        P3_U2818) );
  INV_X1 U20730 ( .A(n17972), .ZN(n17630) );
  NAND2_X1 U20731 ( .A1(n17630), .A2(n17946), .ZN(n17977) );
  INV_X1 U20732 ( .A(n17689), .ZN(n17756) );
  NAND3_X1 U20733 ( .A1(n17688), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18477), .ZN(n17677) );
  NOR2_X1 U20734 ( .A1(n17623), .A2(n17677), .ZN(n17637) );
  NOR2_X1 U20735 ( .A1(n17756), .A2(n17637), .ZN(n17639) );
  INV_X1 U20736 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18649) );
  OAI22_X1 U20737 ( .A1(n17744), .A2(n17624), .B1(n9600), .B2(n18649), .ZN(
        n17625) );
  AOI221_X1 U20738 ( .B1(n17639), .B2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C1(
        n17637), .C2(n17626), .A(n17625), .ZN(n17634) );
  OAI21_X1 U20739 ( .B1(n17630), .B2(n17657), .A(n17656), .ZN(n17632) );
  AOI21_X1 U20740 ( .B1(n17630), .B2(n17629), .A(n17628), .ZN(n17631) );
  XNOR2_X1 U20741 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17631), .ZN(
        n17962) );
  AOI22_X1 U20742 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17632), .B1(
        n17671), .B2(n17962), .ZN(n17633) );
  OAI211_X1 U20743 ( .C1(n17657), .C2(n17977), .A(n17634), .B(n17633), .ZN(
        P3_U2819) );
  INV_X1 U20744 ( .A(n17656), .ZN(n17636) );
  AOI22_X1 U20745 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17636), .B1(
        n17972), .B2(n17635), .ZN(n17645) );
  NAND2_X1 U20746 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17660) );
  NOR2_X1 U20747 ( .A1(n17660), .A2(n17677), .ZN(n17650) );
  NAND2_X1 U20748 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17650), .ZN(
        n17649) );
  OAI22_X1 U20749 ( .A1(n17637), .A2(n17649), .B1(n9600), .B2(n18647), .ZN(
        n17638) );
  AOI21_X1 U20750 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17639), .A(
        n17638), .ZN(n17644) );
  INV_X1 U20751 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17995) );
  AOI22_X1 U20752 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17647), .B1(
        n17640), .B2(n17995), .ZN(n17641) );
  XOR2_X1 U20753 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17641), .Z(
        n17982) );
  AOI22_X1 U20754 ( .A1(n17671), .A2(n17982), .B1(n17642), .B2(n17472), .ZN(
        n17643) );
  OAI211_X1 U20755 ( .C1(n17646), .C2(n17645), .A(n17644), .B(n17643), .ZN(
        P3_U2820) );
  NAND2_X1 U20756 ( .A1(n17647), .A2(n17640), .ZN(n17648) );
  XNOR2_X1 U20757 ( .A(n17648), .B(n17995), .ZN(n17992) );
  OAI211_X1 U20758 ( .C1(n17650), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17689), .B(n17649), .ZN(n17652) );
  NAND2_X1 U20759 ( .A1(n18050), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17651) );
  OAI211_X1 U20760 ( .C1(n17744), .C2(n17653), .A(n17652), .B(n17651), .ZN(
        n17654) );
  AOI21_X1 U20761 ( .B1(n17671), .B2(n17992), .A(n17654), .ZN(n17655) );
  OAI221_X1 U20762 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17657), .C1(
        n17995), .C2(n17656), .A(n17655), .ZN(P3_U2821) );
  AOI21_X1 U20763 ( .B1(n17659), .B2(n17658), .A(n17732), .ZN(n17678) );
  OAI211_X1 U20764 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17661), .A(
        n18477), .B(n17660), .ZN(n17663) );
  NAND2_X1 U20765 ( .A1(n17892), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17662) );
  OAI211_X1 U20766 ( .C1(n17664), .C2(n17678), .A(n17663), .B(n17662), .ZN(
        n17665) );
  AOI21_X1 U20767 ( .B1(n17666), .B2(n17472), .A(n17665), .ZN(n17673) );
  AOI21_X1 U20768 ( .B1(n17668), .B2(n17997), .A(n17667), .ZN(n18007) );
  OAI21_X1 U20769 ( .B1(n9624), .B2(n17999), .A(n17669), .ZN(n18008) );
  AOI22_X1 U20770 ( .A1(n17749), .A2(n18007), .B1(n17671), .B2(n18008), .ZN(
        n17672) );
  OAI211_X1 U20771 ( .C1(n17675), .C2(n17674), .A(n17673), .B(n17672), .ZN(
        P3_U2822) );
  AOI22_X1 U20772 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17678), .B1(
        n17677), .B2(n17676), .ZN(n17679) );
  AOI21_X1 U20773 ( .B1(n13104), .B2(P3_REIP_REG_7__SCAN_IN), .A(n17679), .ZN(
        n17686) );
  NAND2_X1 U20774 ( .A1(n17681), .A2(n17680), .ZN(n17682) );
  XNOR2_X1 U20775 ( .A(n17682), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18018) );
  AOI21_X1 U20776 ( .B1(n18015), .B2(n17684), .A(n17683), .ZN(n18019) );
  AOI22_X1 U20777 ( .A1(n17749), .A2(n18018), .B1(n17752), .B2(n18019), .ZN(
        n17685) );
  OAI211_X1 U20778 ( .C1(n17744), .C2(n17687), .A(n17686), .B(n17685), .ZN(
        P3_U2823) );
  NAND2_X1 U20779 ( .A1(n17688), .A2(n18477), .ZN(n17693) );
  NAND2_X1 U20780 ( .A1(n17689), .A2(n17693), .ZN(n17712) );
  AOI21_X1 U20781 ( .B1(n17692), .B2(n17691), .A(n17690), .ZN(n18025) );
  OAI22_X1 U20782 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17693), .B1(
        n9600), .B2(n18639), .ZN(n17694) );
  AOI21_X1 U20783 ( .B1(n17752), .B2(n18025), .A(n17694), .ZN(n17699) );
  AOI21_X1 U20784 ( .B1(n18026), .B2(n17696), .A(n17695), .ZN(n18024) );
  AOI22_X1 U20785 ( .A1(n17749), .A2(n18024), .B1(n17697), .B2(n17472), .ZN(
        n17698) );
  OAI211_X1 U20786 ( .C1(n17700), .C2(n17712), .A(n17699), .B(n17698), .ZN(
        P3_U2824) );
  AOI21_X1 U20787 ( .B1(n17701), .B2(n17759), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17713) );
  AOI21_X1 U20788 ( .B1(n17704), .B2(n17703), .A(n17702), .ZN(n18032) );
  AOI22_X1 U20789 ( .A1(n18050), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17749), 
        .B2(n18032), .ZN(n17711) );
  AOI21_X1 U20790 ( .B1(n17707), .B2(n17706), .A(n17705), .ZN(n17708) );
  XNOR2_X1 U20791 ( .A(n17708), .B(n9789), .ZN(n18033) );
  AOI22_X1 U20792 ( .A1(n17752), .A2(n18033), .B1(n17709), .B2(n17472), .ZN(
        n17710) );
  OAI211_X1 U20793 ( .C1(n17713), .C2(n17712), .A(n17711), .B(n17710), .ZN(
        P3_U2825) );
  AOI21_X1 U20794 ( .B1(n9785), .B2(n17715), .A(n17714), .ZN(n18043) );
  OAI22_X1 U20795 ( .A1(n9600), .A2(n18635), .B1(n18201), .B2(n17716), .ZN(
        n17717) );
  AOI21_X1 U20796 ( .B1(n17749), .B2(n18043), .A(n17717), .ZN(n17723) );
  OAI21_X1 U20797 ( .B1(n17720), .B2(n17719), .A(n17718), .ZN(n18037) );
  OAI21_X1 U20798 ( .B1(n16733), .B2(n17721), .A(n17759), .ZN(n17734) );
  AOI22_X1 U20799 ( .A1(n17752), .A2(n18037), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17734), .ZN(n17722) );
  OAI211_X1 U20800 ( .C1(n17744), .C2(n17724), .A(n17723), .B(n17722), .ZN(
        P3_U2826) );
  AOI21_X1 U20801 ( .B1(n17727), .B2(n17726), .A(n17725), .ZN(n18049) );
  AOI22_X1 U20802 ( .A1(n17892), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n17752), 
        .B2(n18049), .ZN(n17736) );
  AOI21_X1 U20803 ( .B1(n17730), .B2(n17729), .A(n17728), .ZN(n18051) );
  OAI21_X1 U20804 ( .B1(n17732), .B2(n17747), .A(n17731), .ZN(n17733) );
  AOI22_X1 U20805 ( .A1(n17749), .A2(n18051), .B1(n17734), .B2(n17733), .ZN(
        n17735) );
  OAI211_X1 U20806 ( .C1(n17744), .C2(n17737), .A(n17736), .B(n17735), .ZN(
        P3_U2827) );
  AOI21_X1 U20807 ( .B1(n17740), .B2(n17739), .A(n17738), .ZN(n18058) );
  INV_X1 U20808 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18631) );
  NOR2_X1 U20809 ( .A1(n9600), .A2(n18631), .ZN(n18057) );
  XNOR2_X1 U20810 ( .A(n17742), .B(n17741), .ZN(n18065) );
  OAI22_X1 U20811 ( .A1(n17744), .A2(n17743), .B1(n17764), .B2(n18065), .ZN(
        n17745) );
  AOI211_X1 U20812 ( .C1(n17752), .C2(n18058), .A(n18057), .B(n17745), .ZN(
        n17746) );
  OAI221_X1 U20813 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18201), .C1(
        n17747), .C2(n17759), .A(n17746), .ZN(P3_U2828) );
  NOR2_X1 U20814 ( .A1(n17758), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17748) );
  XNOR2_X1 U20815 ( .A(n17748), .B(n17751), .ZN(n18080) );
  AOI22_X1 U20816 ( .A1(n18050), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17749), 
        .B2(n18080), .ZN(n17754) );
  AOI21_X1 U20817 ( .B1(n17757), .B2(n17751), .A(n17750), .ZN(n18072) );
  AOI22_X1 U20818 ( .A1(n17752), .A2(n18072), .B1(n17755), .B2(n17472), .ZN(
        n17753) );
  OAI211_X1 U20819 ( .C1(n17756), .C2(n17755), .A(n17754), .B(n17753), .ZN(
        P3_U2829) );
  OAI21_X1 U20820 ( .B1(n17758), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17757), .ZN(n18088) );
  INV_X1 U20821 ( .A(n18088), .ZN(n18086) );
  INV_X1 U20822 ( .A(n18752), .ZN(n18594) );
  OAI21_X1 U20823 ( .B1(n17760), .B2(n18594), .A(n17759), .ZN(n17761) );
  AOI22_X1 U20824 ( .A1(n17892), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17761), .ZN(n17762) );
  OAI221_X1 U20825 ( .B1(n18086), .B2(n17764), .C1(n18088), .C2(n17763), .A(
        n17762), .ZN(P3_U2830) );
  NAND3_X1 U20826 ( .A1(n17826), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n17825), .ZN(n17818) );
  NOR2_X1 U20827 ( .A1(n17765), .A2(n17818), .ZN(n17774) );
  AOI21_X1 U20828 ( .B1(n17768), .B2(n17767), .A(n17766), .ZN(n17769) );
  NAND2_X1 U20829 ( .A1(n18730), .A2(n17987), .ZN(n18038) );
  NAND2_X1 U20830 ( .A1(n17829), .A2(n18038), .ZN(n17803) );
  OAI21_X1 U20831 ( .B1(n17803), .B2(n17785), .A(n17768), .ZN(n17791) );
  OAI211_X1 U20832 ( .C1(n17770), .C2(n17968), .A(n17769), .B(n17791), .ZN(
        n17771) );
  AOI21_X1 U20833 ( .B1(n17966), .B2(n17772), .A(n17771), .ZN(n17779) );
  INV_X1 U20834 ( .A(n17779), .ZN(n17773) );
  MUX2_X1 U20835 ( .A(n17774), .B(n17773), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17775) );
  AOI22_X1 U20836 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18052), .B1(
        n18074), .B2(n17775), .ZN(n17777) );
  NAND2_X1 U20837 ( .A1(n13104), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17776) );
  OAI211_X1 U20838 ( .C1(n17778), .C2(n17960), .A(n17777), .B(n17776), .ZN(
        P3_U2835) );
  INV_X1 U20839 ( .A(n18052), .ZN(n18075) );
  OAI21_X1 U20840 ( .B1(n17779), .B2(n18090), .A(n18075), .ZN(n17782) );
  NOR4_X1 U20841 ( .A1(n17779), .A2(n18090), .A3(n17789), .A4(n17818), .ZN(
        n17780) );
  AOI211_X1 U20842 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17782), .A(
        n17781), .B(n17780), .ZN(n17783) );
  OAI21_X1 U20843 ( .B1(n17784), .B2(n17960), .A(n17783), .ZN(P3_U2836) );
  OAI21_X1 U20844 ( .B1(n17786), .B2(n17785), .A(n17801), .ZN(n17793) );
  AOI21_X1 U20845 ( .B1(n17804), .B2(n17787), .A(n18540), .ZN(n17788) );
  INV_X1 U20846 ( .A(n17788), .ZN(n17809) );
  OAI21_X1 U20847 ( .B1(n18559), .B2(n17801), .A(n17789), .ZN(n17790) );
  NAND3_X1 U20848 ( .A1(n17809), .A2(n17791), .A3(n17790), .ZN(n17792) );
  AOI22_X1 U20849 ( .A1(n17966), .A2(n17794), .B1(n17793), .B2(n17792), .ZN(
        n17796) );
  AOI221_X1 U20850 ( .B1(n17968), .B2(n17796), .C1(n17795), .C2(n17796), .A(
        n18090), .ZN(n17797) );
  AOI211_X1 U20851 ( .C1(n17799), .C2(n18009), .A(n17798), .B(n17797), .ZN(
        n17800) );
  OAI21_X1 U20852 ( .B1(n17801), .B2(n18075), .A(n17800), .ZN(P3_U2837) );
  INV_X1 U20853 ( .A(n17802), .ZN(n17844) );
  INV_X1 U20854 ( .A(n17803), .ZN(n17880) );
  AOI21_X1 U20855 ( .B1(n17804), .B2(n17880), .A(n18039), .ZN(n17808) );
  OAI22_X1 U20856 ( .A1(n17806), .A2(n17968), .B1(n17805), .B2(n18539), .ZN(
        n17807) );
  NOR3_X1 U20857 ( .A1(n18052), .A2(n17808), .A3(n17807), .ZN(n17812) );
  NAND3_X1 U20858 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17809), .A3(
        n17812), .ZN(n17810) );
  NAND2_X1 U20859 ( .A1(n9600), .A2(n17810), .ZN(n17823) );
  AOI211_X1 U20860 ( .C1(n17812), .C2(n17811), .A(n10800), .B(n17823), .ZN(
        n17813) );
  AOI21_X1 U20861 ( .B1(n17814), .B2(n17844), .A(n17813), .ZN(n17816) );
  NAND2_X1 U20862 ( .A1(n17892), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17815) );
  OAI211_X1 U20863 ( .C1(n17817), .C2(n17960), .A(n17816), .B(n17815), .ZN(
        P3_U2838) );
  INV_X1 U20864 ( .A(n17818), .ZN(n17819) );
  AOI21_X1 U20865 ( .B1(n17819), .B2(n18075), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17824) );
  AOI21_X1 U20866 ( .B1(n17821), .B2(n18009), .A(n17820), .ZN(n17822) );
  OAI21_X1 U20867 ( .B1(n17824), .B2(n17823), .A(n17822), .ZN(P3_U2839) );
  NAND2_X1 U20868 ( .A1(n17826), .A2(n17825), .ZN(n17838) );
  OAI22_X1 U20869 ( .A1(n17828), .A2(n17968), .B1(n17827), .B2(n18539), .ZN(
        n17845) );
  AOI21_X1 U20870 ( .B1(n17829), .B2(n17858), .A(n18546), .ZN(n17830) );
  AOI221_X1 U20871 ( .B1(n17831), .B2(n18559), .C1(n17846), .C2(n18559), .A(
        n17830), .ZN(n17857) );
  NAND2_X1 U20872 ( .A1(n17968), .A2(n18539), .ZN(n17971) );
  AOI22_X1 U20873 ( .A1(n17861), .A2(n18574), .B1(n17832), .B2(n17971), .ZN(
        n17833) );
  NAND2_X1 U20874 ( .A1(n17857), .A2(n17833), .ZN(n17848) );
  AOI22_X1 U20875 ( .A1(n18559), .A2(n17849), .B1(n17850), .B2(n17898), .ZN(
        n17834) );
  OAI211_X1 U20876 ( .C1(n18571), .C2(n17835), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17834), .ZN(n17836) );
  NOR3_X1 U20877 ( .A1(n17845), .A2(n17848), .A3(n17836), .ZN(n17837) );
  AOI211_X1 U20878 ( .C1(n17839), .C2(n17838), .A(n17837), .B(n18090), .ZN(
        n17840) );
  AOI21_X1 U20879 ( .B1(n18052), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17840), .ZN(n17842) );
  NAND2_X1 U20880 ( .A1(n17892), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17841) );
  OAI211_X1 U20881 ( .C1(n17843), .C2(n17960), .A(n17842), .B(n17841), .ZN(
        P3_U2840) );
  NAND2_X1 U20882 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17844), .ZN(
        n17872) );
  NAND2_X1 U20883 ( .A1(n18571), .A2(n18540), .ZN(n18073) );
  NOR2_X1 U20884 ( .A1(n18090), .A2(n17845), .ZN(n17881) );
  OAI21_X1 U20885 ( .B1(n17900), .B2(n17846), .A(n17987), .ZN(n17847) );
  NAND2_X1 U20886 ( .A1(n17881), .A2(n17847), .ZN(n17860) );
  AOI211_X1 U20887 ( .C1(n17849), .C2(n18073), .A(n17848), .B(n17860), .ZN(
        n17851) );
  NOR3_X1 U20888 ( .A1(n17892), .A2(n17851), .A3(n17850), .ZN(n17852) );
  AOI21_X1 U20889 ( .B1(n18009), .B2(n17853), .A(n17852), .ZN(n17855) );
  OAI211_X1 U20890 ( .C1(n17856), .C2(n17872), .A(n17855), .B(n17854), .ZN(
        P3_U2841) );
  INV_X1 U20891 ( .A(n17971), .ZN(n17877) );
  OAI21_X1 U20892 ( .B1(n17858), .B2(n17877), .A(n17857), .ZN(n17859) );
  OAI21_X1 U20893 ( .B1(n17860), .B2(n17859), .A(n9600), .ZN(n17870) );
  NAND3_X1 U20894 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n17871), .A3(n18073), 
        .ZN(n17862) );
  AOI21_X1 U20895 ( .B1(n17870), .B2(n17862), .A(n17861), .ZN(n17863) );
  AOI211_X1 U20896 ( .C1(n17865), .C2(n18009), .A(n17864), .B(n17863), .ZN(
        n17866) );
  OAI21_X1 U20897 ( .B1(n17867), .B2(n17872), .A(n17866), .ZN(P3_U2842) );
  AOI22_X1 U20898 ( .A1(n17892), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n18009), 
        .B2(n17868), .ZN(n17869) );
  OAI221_X1 U20899 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17872), 
        .C1(n17871), .C2(n17870), .A(n17869), .ZN(P3_U2843) );
  INV_X1 U20900 ( .A(n18066), .ZN(n18042) );
  INV_X1 U20901 ( .A(n18040), .ZN(n17874) );
  INV_X1 U20902 ( .A(n17873), .ZN(n18059) );
  OAI22_X1 U20903 ( .A1(n18042), .A2(n18540), .B1(n17874), .B2(n18059), .ZN(
        n18048) );
  NAND3_X1 U20904 ( .A1(n18027), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18048), .ZN(n18014) );
  NOR2_X1 U20905 ( .A1(n18015), .A2(n18014), .ZN(n17998) );
  NAND2_X1 U20906 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17998), .ZN(
        n17910) );
  NAND2_X1 U20907 ( .A1(n17875), .A2(n17910), .ZN(n17952) );
  NAND2_X1 U20908 ( .A1(n18074), .A2(n17952), .ZN(n17996) );
  NOR2_X1 U20909 ( .A1(n17876), .A2(n17996), .ZN(n17904) );
  AOI22_X1 U20910 ( .A1(n17879), .A2(n17878), .B1(n17877), .B2(n18540), .ZN(
        n17883) );
  AOI21_X1 U20911 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17880), .A(
        n18039), .ZN(n17882) );
  INV_X1 U20912 ( .A(n17881), .ZN(n17903) );
  NOR3_X1 U20913 ( .A1(n17883), .A2(n17882), .A3(n17903), .ZN(n17891) );
  AOI221_X1 U20914 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17891), 
        .C1(n18039), .C2(n17891), .A(n17884), .ZN(n17885) );
  AOI22_X1 U20915 ( .A1(n17904), .A2(n17886), .B1(n17885), .B2(n9600), .ZN(
        n17888) );
  OAI211_X1 U20916 ( .C1(n17889), .C2(n17960), .A(n17888), .B(n17887), .ZN(
        P3_U2844) );
  NOR3_X1 U20917 ( .A1(n17892), .A2(n17891), .A3(n17890), .ZN(n17893) );
  AOI21_X1 U20918 ( .B1(n17904), .B2(n17894), .A(n17893), .ZN(n17896) );
  OAI211_X1 U20919 ( .C1(n17897), .C2(n17960), .A(n17896), .B(n17895), .ZN(
        P3_U2845) );
  INV_X1 U20920 ( .A(n17898), .ZN(n17980) );
  NOR2_X1 U20921 ( .A1(n17923), .A2(n18540), .ZN(n17964) );
  AOI211_X1 U20922 ( .C1(n17900), .C2(n17987), .A(n17964), .B(n17899), .ZN(
        n17901) );
  NAND2_X1 U20923 ( .A1(n18574), .A2(n17939), .ZN(n17979) );
  OAI211_X1 U20924 ( .C1(n17902), .C2(n17980), .A(n17901), .B(n17979), .ZN(
        n17912) );
  OAI221_X1 U20925 ( .B1(n17903), .B2(n18004), .C1(n17903), .C2(n17912), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17907) );
  AOI22_X1 U20926 ( .A1(n18009), .A2(n17905), .B1(n17904), .B2(n10794), .ZN(
        n17906) );
  OAI221_X1 U20927 ( .B1(n18050), .B2(n17907), .C1(n9600), .C2(n18659), .A(
        n17906), .ZN(P3_U2846) );
  NOR2_X1 U20928 ( .A1(n9600), .A2(n18657), .ZN(n17916) );
  NAND3_X1 U20929 ( .A1(n18000), .A2(n17909), .A3(n17908), .ZN(n17914) );
  NOR2_X1 U20930 ( .A1(n17910), .A2(n17925), .ZN(n17933) );
  OAI211_X1 U20931 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n17933), .A(
        n17912), .B(n17911), .ZN(n17913) );
  AOI21_X1 U20932 ( .B1(n17914), .B2(n17913), .A(n18090), .ZN(n17915) );
  AOI211_X1 U20933 ( .C1(n18052), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17916), .B(n17915), .ZN(n17920) );
  NAND3_X1 U20934 ( .A1(n18089), .A2(n17918), .A3(n17917), .ZN(n17919) );
  OAI211_X1 U20935 ( .C1(n17921), .C2(n17960), .A(n17920), .B(n17919), .ZN(
        P3_U2847) );
  AOI21_X1 U20936 ( .B1(n17923), .B2(n17922), .A(n18540), .ZN(n17924) );
  AOI221_X1 U20937 ( .B1(n17939), .B2(n18574), .C1(n17925), .C2(n18574), .A(
        n17924), .ZN(n17927) );
  INV_X1 U20938 ( .A(n17963), .ZN(n17986) );
  OAI21_X1 U20939 ( .B1(n17926), .B2(n17986), .A(n17987), .ZN(n17942) );
  OAI211_X1 U20940 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18571), .A(
        n17927), .B(n17942), .ZN(n17931) );
  OAI22_X1 U20941 ( .A1(n17968), .A2(n17929), .B1(n18539), .B2(n17928), .ZN(
        n17930) );
  AOI221_X1 U20942 ( .B1(n17933), .B2(n17932), .C1(n17931), .C2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n17930), .ZN(n17937) );
  AOI22_X1 U20943 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18052), .B1(
        n18009), .B2(n17934), .ZN(n17936) );
  OAI211_X1 U20944 ( .C1(n17937), .C2(n18090), .A(n17936), .B(n17935), .ZN(
        P3_U2848) );
  AOI22_X1 U20945 ( .A1(n18050), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18009), 
        .B2(n17938), .ZN(n17949) );
  OAI21_X1 U20946 ( .B1(n17972), .B2(n17939), .A(n18574), .ZN(n17940) );
  OAI21_X1 U20947 ( .B1(n17953), .B2(n18540), .A(n17940), .ZN(n17974) );
  AOI211_X1 U20948 ( .C1(n17966), .C2(n17941), .A(n17964), .B(n17974), .ZN(
        n17943) );
  OAI211_X1 U20949 ( .C1(n17944), .C2(n17968), .A(n17943), .B(n17942), .ZN(
        n17951) );
  AOI21_X1 U20950 ( .B1(n17946), .B2(n18574), .A(n17945), .ZN(n17955) );
  OAI21_X1 U20951 ( .B1(n17980), .B2(n17955), .A(n18074), .ZN(n17947) );
  OAI211_X1 U20952 ( .C1(n17951), .C2(n17947), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n9600), .ZN(n17948) );
  OAI211_X1 U20953 ( .C1(n17996), .C2(n17950), .A(n17949), .B(n17948), .ZN(
        P3_U2849) );
  INV_X1 U20954 ( .A(n17951), .ZN(n17956) );
  AOI21_X1 U20955 ( .B1(n17953), .B2(n17952), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17954) );
  AOI211_X1 U20956 ( .C1(n17956), .C2(n17955), .A(n17954), .B(n18090), .ZN(
        n17957) );
  AOI21_X1 U20957 ( .B1(n18052), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17957), .ZN(n17959) );
  OAI211_X1 U20958 ( .C1(n17961), .C2(n17960), .A(n17959), .B(n17958), .ZN(
        P3_U2850) );
  AOI22_X1 U20959 ( .A1(n18050), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18009), 
        .B2(n17962), .ZN(n17976) );
  AOI21_X1 U20960 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17963), .A(
        n18571), .ZN(n17970) );
  AOI211_X1 U20961 ( .C1(n17966), .C2(n17965), .A(n17964), .B(n18090), .ZN(
        n17967) );
  OAI21_X1 U20962 ( .B1(n17969), .B2(n17968), .A(n17967), .ZN(n17991) );
  AOI211_X1 U20963 ( .C1(n17972), .C2(n17971), .A(n17970), .B(n17991), .ZN(
        n17978) );
  OAI21_X1 U20964 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18571), .A(
        n17978), .ZN(n17973) );
  OAI211_X1 U20965 ( .C1(n17974), .C2(n17973), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n9600), .ZN(n17975) );
  OAI211_X1 U20966 ( .C1(n17977), .C2(n17996), .A(n17976), .B(n17975), .ZN(
        P3_U2851) );
  OAI211_X1 U20967 ( .C1(n17980), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17979), .B(n17978), .ZN(n17981) );
  NAND2_X1 U20968 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17981), .ZN(
        n17985) );
  NOR2_X1 U20969 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17996), .ZN(
        n17983) );
  AOI22_X1 U20970 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17983), .B1(
        n18009), .B2(n17982), .ZN(n17984) );
  OAI221_X1 U20971 ( .B1(n13104), .B2(n17985), .C1(n9600), .C2(n18647), .A(
        n17984), .ZN(P3_U2852) );
  NAND2_X1 U20972 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18005) );
  INV_X1 U20973 ( .A(n18005), .ZN(n17989) );
  OAI221_X1 U20974 ( .B1(n17987), .B2(n17997), .C1(n17987), .C2(n18574), .A(
        n17986), .ZN(n17988) );
  OAI221_X1 U20975 ( .B1(n18546), .B2(n17989), .C1(n18546), .C2(n18003), .A(
        n17988), .ZN(n17990) );
  OAI21_X1 U20976 ( .B1(n17991), .B2(n17990), .A(n9600), .ZN(n17994) );
  AOI22_X1 U20977 ( .A1(n18050), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18009), 
        .B2(n17992), .ZN(n17993) );
  OAI221_X1 U20978 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17996), .C1(
        n17995), .C2(n17994), .A(n17993), .ZN(P3_U2853) );
  AOI22_X1 U20979 ( .A1(n18000), .A2(n17999), .B1(n17998), .B2(n17997), .ZN(
        n18012) );
  NAND2_X1 U20980 ( .A1(n18559), .A2(n18001), .ZN(n18002) );
  OAI211_X1 U20981 ( .C1(n18003), .C2(n18039), .A(n18002), .B(n18038), .ZN(
        n18022) );
  AOI21_X1 U20982 ( .B1(n18005), .B2(n18004), .A(n18022), .ZN(n18013) );
  OAI21_X1 U20983 ( .B1(n18013), .B2(n18076), .A(n18075), .ZN(n18006) );
  AOI22_X1 U20984 ( .A1(n18050), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18006), .ZN(n18011) );
  AOI22_X1 U20985 ( .A1(n18009), .A2(n18008), .B1(n18089), .B2(n18007), .ZN(
        n18010) );
  OAI211_X1 U20986 ( .C1(n18012), .C2(n18090), .A(n18011), .B(n18010), .ZN(
        P3_U2854) );
  NOR2_X1 U20987 ( .A1(n9600), .A2(n18641), .ZN(n18017) );
  AOI211_X1 U20988 ( .C1(n18015), .C2(n18014), .A(n18013), .B(n18090), .ZN(
        n18016) );
  AOI211_X1 U20989 ( .C1(n18052), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18017), .B(n18016), .ZN(n18021) );
  INV_X1 U20990 ( .A(n18083), .ZN(n18087) );
  AOI22_X1 U20991 ( .A1(n18087), .A2(n18019), .B1(n18089), .B2(n18018), .ZN(
        n18020) );
  NAND2_X1 U20992 ( .A1(n18021), .A2(n18020), .ZN(P3_U2855) );
  AOI21_X1 U20993 ( .B1(n18022), .B2(n18074), .A(n18052), .ZN(n18023) );
  INV_X1 U20994 ( .A(n18023), .ZN(n18031) );
  AOI22_X1 U20995 ( .A1(n18050), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18031), .ZN(n18030) );
  AOI22_X1 U20996 ( .A1(n18087), .A2(n18025), .B1(n18089), .B2(n18024), .ZN(
        n18029) );
  NAND4_X1 U20997 ( .A1(n18074), .A2(n18027), .A3(n18026), .A4(n18048), .ZN(
        n18028) );
  NAND3_X1 U20998 ( .A1(n18030), .A2(n18029), .A3(n18028), .ZN(P3_U2856) );
  NAND4_X1 U20999 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18074), .A3(
        n9789), .A4(n18048), .ZN(n18036) );
  AOI22_X1 U21000 ( .A1(n18050), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18031), .ZN(n18035) );
  AOI22_X1 U21001 ( .A1(n18087), .A2(n18033), .B1(n18089), .B2(n18032), .ZN(
        n18034) );
  OAI211_X1 U21002 ( .C1(n9785), .C2(n18036), .A(n18035), .B(n18034), .ZN(
        P3_U2857) );
  NAND3_X1 U21003 ( .A1(n18074), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18048), .ZN(n18047) );
  AOI22_X1 U21004 ( .A1(n18050), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18087), 
        .B2(n18037), .ZN(n18046) );
  OAI21_X1 U21005 ( .B1(n18040), .B2(n18039), .A(n18038), .ZN(n18060) );
  AOI211_X1 U21006 ( .C1(n18042), .C2(n18559), .A(n18041), .B(n18060), .ZN(
        n18056) );
  OAI21_X1 U21007 ( .B1(n18056), .B2(n18076), .A(n18075), .ZN(n18044) );
  AOI22_X1 U21008 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18044), .B1(
        n18089), .B2(n18043), .ZN(n18045) );
  OAI211_X1 U21009 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18047), .A(
        n18046), .B(n18045), .ZN(P3_U2858) );
  OAI21_X1 U21010 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18048), .A(
        n18074), .ZN(n18055) );
  AOI22_X1 U21011 ( .A1(n18050), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18087), 
        .B2(n18049), .ZN(n18054) );
  AOI22_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18052), .B1(
        n18089), .B2(n18051), .ZN(n18053) );
  OAI211_X1 U21013 ( .C1(n18056), .C2(n18055), .A(n18054), .B(n18053), .ZN(
        P3_U2859) );
  AOI21_X1 U21014 ( .B1(n18087), .B2(n18058), .A(n18057), .ZN(n18070) );
  NOR2_X1 U21015 ( .A1(n10690), .A2(n18059), .ZN(n18064) );
  NOR2_X1 U21016 ( .A1(n10690), .A2(n18730), .ZN(n18061) );
  AOI21_X1 U21017 ( .B1(n18559), .B2(n18061), .A(n18060), .ZN(n18062) );
  INV_X1 U21018 ( .A(n18062), .ZN(n18063) );
  MUX2_X1 U21019 ( .A(n18064), .B(n18063), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18068) );
  OAI22_X1 U21020 ( .A1(n18540), .A2(n18066), .B1(n18539), .B2(n18065), .ZN(
        n18067) );
  OAI21_X1 U21021 ( .B1(n18068), .B2(n18067), .A(n18074), .ZN(n18069) );
  OAI211_X1 U21022 ( .C1(n18075), .C2(n18071), .A(n18070), .B(n18069), .ZN(
        P3_U2860) );
  INV_X1 U21023 ( .A(n18072), .ZN(n18084) );
  NAND3_X1 U21024 ( .A1(n18074), .A2(n18730), .A3(n18073), .ZN(n18092) );
  AOI21_X1 U21025 ( .B1(n18075), .B2(n18092), .A(n10690), .ZN(n18079) );
  NOR3_X1 U21026 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18077), .A3(
        n18076), .ZN(n18078) );
  AOI211_X1 U21027 ( .C1(n18089), .C2(n18080), .A(n18079), .B(n18078), .ZN(
        n18082) );
  NAND2_X1 U21028 ( .A1(n17892), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18081) );
  OAI211_X1 U21029 ( .C1(n18084), .C2(n18083), .A(n18082), .B(n18081), .ZN(
        P3_U2861) );
  INV_X1 U21030 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18741) );
  NOR2_X1 U21031 ( .A1(n9600), .A2(n18741), .ZN(n18085) );
  AOI221_X1 U21032 ( .B1(n18089), .B2(n18088), .C1(n18087), .C2(n18086), .A(
        n18085), .ZN(n18093) );
  OAI211_X1 U21033 ( .C1(n18574), .C2(n18090), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n9600), .ZN(n18091) );
  NAND3_X1 U21034 ( .A1(n18093), .A2(n18092), .A3(n18091), .ZN(P3_U2862) );
  INV_X1 U21035 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18575) );
  AOI21_X1 U21036 ( .B1(n18096), .B2(n18095), .A(n18094), .ZN(n18598) );
  OAI21_X1 U21037 ( .B1(n18598), .B2(n18138), .A(n18101), .ZN(n18097) );
  OAI221_X1 U21038 ( .B1(n18575), .B2(n18756), .C1(n18575), .C2(n18101), .A(
        n18097), .ZN(P3_U2863) );
  NOR2_X1 U21039 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18585), .ZN(
        n18315) );
  NOR2_X1 U21040 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18411), .ZN(
        n18270) );
  NOR2_X1 U21041 ( .A1(n18315), .A2(n18270), .ZN(n18099) );
  OAI22_X1 U21042 ( .A1(n18100), .A2(n18585), .B1(n18099), .B2(n18098), .ZN(
        P3_U2866) );
  INV_X1 U21043 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18583) );
  NOR2_X1 U21044 ( .A1(n18583), .A2(n18101), .ZN(P3_U2867) );
  NOR2_X1 U21045 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18579) );
  NOR2_X1 U21046 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18179) );
  NAND2_X1 U21047 ( .A1(n18579), .A2(n18179), .ZN(n18192) );
  NOR2_X1 U21048 ( .A1(n18103), .A2(n18102), .ZN(n18110) );
  NAND2_X1 U21049 ( .A1(n18110), .A2(n10901), .ZN(n18481) );
  NAND3_X1 U21050 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18576), .ZN(n18410) );
  NOR2_X2 U21051 ( .A1(n18575), .A2(n18410), .ZN(n18509) );
  NOR2_X2 U21052 ( .A1(n20807), .A2(n18201), .ZN(n18473) );
  AND2_X1 U21053 ( .A1(n18385), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18472) );
  NOR2_X1 U21054 ( .A1(n18585), .A2(n18246), .ZN(n18475) );
  INV_X1 U21055 ( .A(n18475), .ZN(n18471) );
  NOR2_X2 U21056 ( .A1(n18575), .A2(n18471), .ZN(n18526) );
  INV_X1 U21057 ( .A(n18192), .ZN(n18196) );
  NOR2_X1 U21058 ( .A1(n18526), .A2(n18196), .ZN(n18158) );
  NOR2_X1 U21059 ( .A1(n18605), .A2(n18158), .ZN(n18132) );
  AOI22_X1 U21060 ( .A1(n18509), .A2(n18473), .B1(n18472), .B2(n18132), .ZN(
        n18106) );
  INV_X1 U21061 ( .A(n18509), .ZN(n18531) );
  NAND2_X1 U21062 ( .A1(n18475), .A2(n18575), .ZN(n18449) );
  NAND2_X1 U21063 ( .A1(n18531), .A2(n18449), .ZN(n18442) );
  AOI21_X1 U21064 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18200), .ZN(n18439) );
  INV_X1 U21065 ( .A(n18158), .ZN(n18104) );
  AOI22_X1 U21066 ( .A1(n18477), .A2(n18442), .B1(n18439), .B2(n18104), .ZN(
        n18135) );
  INV_X1 U21067 ( .A(n18449), .ZN(n18467) );
  NOR2_X2 U21068 ( .A1(n18201), .A2(n19072), .ZN(n18478) );
  AOI22_X1 U21069 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18135), .B1(
        n18467), .B2(n18478), .ZN(n18105) );
  OAI211_X1 U21070 ( .C1(n18192), .C2(n18481), .A(n18106), .B(n18105), .ZN(
        P3_U2868) );
  NAND2_X1 U21071 ( .A1(n18110), .A2(n18749), .ZN(n18487) );
  AND2_X1 U21072 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18477), .ZN(n18483) );
  AND2_X1 U21073 ( .A1(n18385), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18482) );
  AOI22_X1 U21074 ( .A1(n18509), .A2(n18483), .B1(n18132), .B2(n18482), .ZN(
        n18108) );
  NOR2_X2 U21075 ( .A1(n18201), .A2(n15041), .ZN(n18484) );
  AOI22_X1 U21076 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18135), .B1(
        n18467), .B2(n18484), .ZN(n18107) );
  OAI211_X1 U21077 ( .C1(n18192), .C2(n18487), .A(n18108), .B(n18107), .ZN(
        P3_U2869) );
  NAND2_X1 U21078 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18477), .ZN(n18393) );
  NOR2_X2 U21079 ( .A1(n18201), .A2(n19092), .ZN(n18490) );
  NOR2_X2 U21080 ( .A1(n18200), .A2(n18109), .ZN(n18488) );
  AOI22_X1 U21081 ( .A1(n18467), .A2(n18490), .B1(n18132), .B2(n18488), .ZN(
        n18113) );
  INV_X1 U21082 ( .A(n18110), .ZN(n18133) );
  NOR2_X1 U21083 ( .A1(n18111), .A2(n18133), .ZN(n18390) );
  AOI22_X1 U21084 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18135), .B1(
        n18196), .B2(n18390), .ZN(n18112) );
  OAI211_X1 U21085 ( .C1(n18531), .C2(n18393), .A(n18113), .B(n18112), .ZN(
        P3_U2870) );
  NAND2_X1 U21086 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18477), .ZN(n18453) );
  NOR2_X2 U21087 ( .A1(n18201), .A2(n19097), .ZN(n18496) );
  NOR2_X2 U21088 ( .A1(n18200), .A2(n18114), .ZN(n18494) );
  AOI22_X1 U21089 ( .A1(n18467), .A2(n18496), .B1(n18132), .B2(n18494), .ZN(
        n18117) );
  NOR2_X1 U21090 ( .A1(n18115), .A2(n18133), .ZN(n18450) );
  AOI22_X1 U21091 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18135), .B1(
        n18196), .B2(n18450), .ZN(n18116) );
  OAI211_X1 U21092 ( .C1(n18531), .C2(n18453), .A(n18117), .B(n18116), .ZN(
        P3_U2871) );
  NAND2_X1 U21093 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18477), .ZN(n18457) );
  NOR2_X2 U21094 ( .A1(n18201), .A2(n15022), .ZN(n18502) );
  NOR2_X2 U21095 ( .A1(n18200), .A2(n18118), .ZN(n18500) );
  AOI22_X1 U21096 ( .A1(n18467), .A2(n18502), .B1(n18132), .B2(n18500), .ZN(
        n18121) );
  NOR2_X1 U21097 ( .A1(n18119), .A2(n18133), .ZN(n18454) );
  AOI22_X1 U21098 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18135), .B1(
        n18196), .B2(n18454), .ZN(n18120) );
  OAI211_X1 U21099 ( .C1(n18531), .C2(n18457), .A(n18121), .B(n18120), .ZN(
        P3_U2872) );
  NAND2_X1 U21100 ( .A1(n18477), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18428) );
  NAND2_X1 U21101 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18477), .ZN(n18514) );
  INV_X1 U21102 ( .A(n18514), .ZN(n18425) );
  AND2_X1 U21103 ( .A1(n18385), .A2(BUF2_REG_5__SCAN_IN), .ZN(n18507) );
  AOI22_X1 U21104 ( .A1(n18509), .A2(n18425), .B1(n18132), .B2(n18507), .ZN(
        n18124) );
  NOR2_X2 U21105 ( .A1(n18122), .A2(n18133), .ZN(n18510) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18135), .B1(
        n18196), .B2(n18510), .ZN(n18123) );
  OAI211_X1 U21107 ( .C1(n18449), .C2(n18428), .A(n18124), .B(n18123), .ZN(
        P3_U2873) );
  NAND2_X1 U21108 ( .A1(n18477), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18520) );
  NOR2_X1 U21109 ( .A1(n18125), .A2(n18201), .ZN(n18515) );
  NOR2_X2 U21110 ( .A1(n18200), .A2(n18126), .ZN(n18516) );
  AOI22_X1 U21111 ( .A1(n18509), .A2(n18515), .B1(n18132), .B2(n18516), .ZN(
        n18129) );
  NOR2_X2 U21112 ( .A1(n18127), .A2(n18133), .ZN(n18517) );
  AOI22_X1 U21113 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18135), .B1(
        n18196), .B2(n18517), .ZN(n18128) );
  OAI211_X1 U21114 ( .C1(n18449), .C2(n18520), .A(n18129), .B(n18128), .ZN(
        P3_U2874) );
  NAND2_X1 U21115 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18477), .ZN(n18530) );
  NOR2_X1 U21116 ( .A1(n18201), .A2(n18130), .ZN(n18524) );
  NOR2_X2 U21117 ( .A1(n18131), .A2(n18200), .ZN(n18522) );
  AOI22_X1 U21118 ( .A1(n18509), .A2(n18524), .B1(n18132), .B2(n18522), .ZN(
        n18137) );
  NOR2_X2 U21119 ( .A1(n18134), .A2(n18133), .ZN(n18525) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18135), .B1(
        n18196), .B2(n18525), .ZN(n18136) );
  OAI211_X1 U21121 ( .C1(n18449), .C2(n18530), .A(n18137), .B(n18136), .ZN(
        P3_U2875) );
  NOR2_X1 U21122 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18575), .ZN(
        n18314) );
  NAND2_X1 U21123 ( .A1(n18179), .A2(n18314), .ZN(n18212) );
  INV_X1 U21124 ( .A(n18179), .ZN(n18157) );
  INV_X1 U21125 ( .A(n18605), .ZN(n18437) );
  NAND2_X1 U21126 ( .A1(n18576), .A2(n18437), .ZN(n18316) );
  NOR2_X1 U21127 ( .A1(n18157), .A2(n18316), .ZN(n18153) );
  AOI22_X1 U21128 ( .A1(n18467), .A2(n18473), .B1(n18472), .B2(n18153), .ZN(
        n18140) );
  NOR2_X1 U21129 ( .A1(n18200), .A2(n18138), .ZN(n18474) );
  INV_X1 U21130 ( .A(n18474), .ZN(n18178) );
  NOR2_X1 U21131 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18178), .ZN(
        n18412) );
  AOI22_X1 U21132 ( .A1(n18477), .A2(n18475), .B1(n18179), .B2(n18412), .ZN(
        n18154) );
  AOI22_X1 U21133 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18154), .B1(
        n18526), .B2(n18478), .ZN(n18139) );
  OAI211_X1 U21134 ( .C1(n18481), .C2(n18212), .A(n18140), .B(n18139), .ZN(
        P3_U2876) );
  AOI22_X1 U21135 ( .A1(n18526), .A2(n18484), .B1(n18482), .B2(n18153), .ZN(
        n18142) );
  AOI22_X1 U21136 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18154), .B1(
        n18467), .B2(n18483), .ZN(n18141) );
  OAI211_X1 U21137 ( .C1(n18487), .C2(n18212), .A(n18142), .B(n18141), .ZN(
        P3_U2877) );
  INV_X1 U21138 ( .A(n18390), .ZN(n18493) );
  INV_X1 U21139 ( .A(n18393), .ZN(n18489) );
  AOI22_X1 U21140 ( .A1(n18467), .A2(n18489), .B1(n18488), .B2(n18153), .ZN(
        n18144) );
  AOI22_X1 U21141 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18154), .B1(
        n18526), .B2(n18490), .ZN(n18143) );
  OAI211_X1 U21142 ( .C1(n18493), .C2(n18212), .A(n18144), .B(n18143), .ZN(
        P3_U2878) );
  AOI22_X1 U21143 ( .A1(n18526), .A2(n18496), .B1(n18494), .B2(n18153), .ZN(
        n18146) );
  INV_X1 U21144 ( .A(n18212), .ZN(n18220) );
  AOI22_X1 U21145 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18154), .B1(
        n18450), .B2(n18220), .ZN(n18145) );
  OAI211_X1 U21146 ( .C1(n18449), .C2(n18453), .A(n18146), .B(n18145), .ZN(
        P3_U2879) );
  INV_X1 U21147 ( .A(n18454), .ZN(n18505) );
  INV_X1 U21148 ( .A(n18457), .ZN(n18501) );
  AOI22_X1 U21149 ( .A1(n18467), .A2(n18501), .B1(n18500), .B2(n18153), .ZN(
        n18148) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18154), .B1(
        n18526), .B2(n18502), .ZN(n18147) );
  OAI211_X1 U21151 ( .C1(n18505), .C2(n18212), .A(n18148), .B(n18147), .ZN(
        P3_U2880) );
  INV_X1 U21152 ( .A(n18428), .ZN(n18508) );
  AOI22_X1 U21153 ( .A1(n18526), .A2(n18508), .B1(n18507), .B2(n18153), .ZN(
        n18150) );
  AOI22_X1 U21154 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18154), .B1(
        n18510), .B2(n18220), .ZN(n18149) );
  OAI211_X1 U21155 ( .C1(n18449), .C2(n18514), .A(n18150), .B(n18149), .ZN(
        P3_U2881) );
  INV_X1 U21156 ( .A(n18515), .ZN(n18464) );
  INV_X1 U21157 ( .A(n18520), .ZN(n18460) );
  AOI22_X1 U21158 ( .A1(n18526), .A2(n18460), .B1(n18516), .B2(n18153), .ZN(
        n18152) );
  AOI22_X1 U21159 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18154), .B1(
        n18517), .B2(n18220), .ZN(n18151) );
  OAI211_X1 U21160 ( .C1(n18449), .C2(n18464), .A(n18152), .B(n18151), .ZN(
        P3_U2882) );
  INV_X1 U21161 ( .A(n18524), .ZN(n18409) );
  INV_X1 U21162 ( .A(n18530), .ZN(n18404) );
  AOI22_X1 U21163 ( .A1(n18526), .A2(n18404), .B1(n18522), .B2(n18153), .ZN(
        n18156) );
  AOI22_X1 U21164 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18154), .B1(
        n18525), .B2(n18220), .ZN(n18155) );
  OAI211_X1 U21165 ( .C1(n18449), .C2(n18409), .A(n18156), .B(n18155), .ZN(
        P3_U2883) );
  NOR2_X1 U21166 ( .A1(n18576), .A2(n18157), .ZN(n18226) );
  NAND2_X1 U21167 ( .A1(n18226), .A2(n18575), .ZN(n18224) );
  INV_X1 U21168 ( .A(n18224), .ZN(n18242) );
  NOR2_X1 U21169 ( .A1(n18220), .A2(n18242), .ZN(n18202) );
  NOR2_X1 U21170 ( .A1(n18605), .A2(n18202), .ZN(n18174) );
  AOI22_X1 U21171 ( .A1(n18526), .A2(n18473), .B1(n18472), .B2(n18174), .ZN(
        n18161) );
  INV_X1 U21172 ( .A(n18441), .ZN(n18382) );
  OAI21_X1 U21173 ( .B1(n18158), .B2(n18382), .A(n18202), .ZN(n18159) );
  OAI211_X1 U21174 ( .C1(n18242), .C2(n18704), .A(n18385), .B(n18159), .ZN(
        n18175) );
  AOI22_X1 U21175 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18175), .B1(
        n18196), .B2(n18478), .ZN(n18160) );
  OAI211_X1 U21176 ( .C1(n18481), .C2(n18224), .A(n18161), .B(n18160), .ZN(
        P3_U2884) );
  AOI22_X1 U21177 ( .A1(n18526), .A2(n18483), .B1(n18482), .B2(n18174), .ZN(
        n18163) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18175), .B1(
        n18196), .B2(n18484), .ZN(n18162) );
  OAI211_X1 U21179 ( .C1(n18487), .C2(n18224), .A(n18163), .B(n18162), .ZN(
        P3_U2885) );
  AOI22_X1 U21180 ( .A1(n18526), .A2(n18489), .B1(n18488), .B2(n18174), .ZN(
        n18165) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18175), .B1(
        n18196), .B2(n18490), .ZN(n18164) );
  OAI211_X1 U21182 ( .C1(n18493), .C2(n18224), .A(n18165), .B(n18164), .ZN(
        P3_U2886) );
  INV_X1 U21183 ( .A(n18526), .ZN(n18506) );
  AOI22_X1 U21184 ( .A1(n18196), .A2(n18496), .B1(n18494), .B2(n18174), .ZN(
        n18167) );
  AOI22_X1 U21185 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18175), .B1(
        n18450), .B2(n18242), .ZN(n18166) );
  OAI211_X1 U21186 ( .C1(n18506), .C2(n18453), .A(n18167), .B(n18166), .ZN(
        P3_U2887) );
  AOI22_X1 U21187 ( .A1(n18526), .A2(n18501), .B1(n18500), .B2(n18174), .ZN(
        n18169) );
  AOI22_X1 U21188 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18175), .B1(
        n18196), .B2(n18502), .ZN(n18168) );
  OAI211_X1 U21189 ( .C1(n18505), .C2(n18224), .A(n18169), .B(n18168), .ZN(
        P3_U2888) );
  AOI22_X1 U21190 ( .A1(n18196), .A2(n18508), .B1(n18507), .B2(n18174), .ZN(
        n18171) );
  AOI22_X1 U21191 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18175), .B1(
        n18510), .B2(n18242), .ZN(n18170) );
  OAI211_X1 U21192 ( .C1(n18506), .C2(n18514), .A(n18171), .B(n18170), .ZN(
        P3_U2889) );
  AOI22_X1 U21193 ( .A1(n18196), .A2(n18460), .B1(n18516), .B2(n18174), .ZN(
        n18173) );
  AOI22_X1 U21194 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18175), .B1(
        n18517), .B2(n18242), .ZN(n18172) );
  OAI211_X1 U21195 ( .C1(n18506), .C2(n18464), .A(n18173), .B(n18172), .ZN(
        P3_U2890) );
  AOI22_X1 U21196 ( .A1(n18196), .A2(n18404), .B1(n18522), .B2(n18174), .ZN(
        n18177) );
  AOI22_X1 U21197 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18175), .B1(
        n18525), .B2(n18242), .ZN(n18176) );
  OAI211_X1 U21198 ( .C1(n18506), .C2(n18409), .A(n18177), .B(n18176), .ZN(
        P3_U2891) );
  NAND2_X1 U21199 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18226), .ZN(
        n18268) );
  AND2_X1 U21200 ( .A1(n18437), .A2(n18226), .ZN(n18195) );
  AOI22_X1 U21201 ( .A1(n18478), .A2(n18220), .B1(n18472), .B2(n18195), .ZN(
        n18181) );
  AOI21_X1 U21202 ( .B1(n18576), .B2(n18382), .A(n18178), .ZN(n18269) );
  NAND2_X1 U21203 ( .A1(n18179), .A2(n18269), .ZN(n18197) );
  AOI22_X1 U21204 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18473), .ZN(n18180) );
  OAI211_X1 U21205 ( .C1(n18481), .C2(n18268), .A(n18181), .B(n18180), .ZN(
        P3_U2892) );
  AOI22_X1 U21206 ( .A1(n18484), .A2(n18220), .B1(n18482), .B2(n18195), .ZN(
        n18183) );
  AOI22_X1 U21207 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18483), .ZN(n18182) );
  OAI211_X1 U21208 ( .C1(n18487), .C2(n18268), .A(n18183), .B(n18182), .ZN(
        P3_U2893) );
  AOI22_X1 U21209 ( .A1(n18490), .A2(n18220), .B1(n18488), .B2(n18195), .ZN(
        n18185) );
  AOI22_X1 U21210 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18489), .ZN(n18184) );
  OAI211_X1 U21211 ( .C1(n18493), .C2(n18268), .A(n18185), .B(n18184), .ZN(
        P3_U2894) );
  INV_X1 U21212 ( .A(n18450), .ZN(n18499) );
  INV_X1 U21213 ( .A(n18453), .ZN(n18495) );
  AOI22_X1 U21214 ( .A1(n18196), .A2(n18495), .B1(n18494), .B2(n18195), .ZN(
        n18187) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18197), .B1(
        n18496), .B2(n18220), .ZN(n18186) );
  OAI211_X1 U21216 ( .C1(n18499), .C2(n18268), .A(n18187), .B(n18186), .ZN(
        P3_U2895) );
  AOI22_X1 U21217 ( .A1(n18502), .A2(n18220), .B1(n18500), .B2(n18195), .ZN(
        n18189) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18197), .B1(
        n18196), .B2(n18501), .ZN(n18188) );
  OAI211_X1 U21219 ( .C1(n18505), .C2(n18268), .A(n18189), .B(n18188), .ZN(
        P3_U2896) );
  AOI22_X1 U21220 ( .A1(n18508), .A2(n18220), .B1(n18507), .B2(n18195), .ZN(
        n18191) );
  INV_X1 U21221 ( .A(n18268), .ZN(n18261) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18197), .B1(
        n18510), .B2(n18261), .ZN(n18190) );
  OAI211_X1 U21223 ( .C1(n18192), .C2(n18514), .A(n18191), .B(n18190), .ZN(
        P3_U2897) );
  AOI22_X1 U21224 ( .A1(n18196), .A2(n18515), .B1(n18516), .B2(n18195), .ZN(
        n18194) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18197), .B1(
        n18517), .B2(n18261), .ZN(n18193) );
  OAI211_X1 U21226 ( .C1(n18520), .C2(n18212), .A(n18194), .B(n18193), .ZN(
        P3_U2898) );
  AOI22_X1 U21227 ( .A1(n18196), .A2(n18524), .B1(n18522), .B2(n18195), .ZN(
        n18199) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18197), .B1(
        n18525), .B2(n18261), .ZN(n18198) );
  OAI211_X1 U21229 ( .C1(n18530), .C2(n18212), .A(n18199), .B(n18198), .ZN(
        P3_U2899) );
  NAND2_X1 U21230 ( .A1(n18579), .A2(n18270), .ZN(n18290) );
  INV_X1 U21231 ( .A(n18290), .ZN(n18279) );
  NOR2_X1 U21232 ( .A1(n18261), .A2(n18279), .ZN(n18247) );
  NOR2_X1 U21233 ( .A1(n18605), .A2(n18247), .ZN(n18219) );
  AOI22_X1 U21234 ( .A1(n18478), .A2(n18242), .B1(n18472), .B2(n18219), .ZN(
        n18205) );
  OAI22_X1 U21235 ( .A1(n18202), .A2(n18201), .B1(n18247), .B2(n18200), .ZN(
        n18203) );
  OAI21_X1 U21236 ( .B1(n18279), .B2(n18704), .A(n18203), .ZN(n18221) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18221), .B1(
        n18473), .B2(n18220), .ZN(n18204) );
  OAI211_X1 U21238 ( .C1(n18481), .C2(n18290), .A(n18205), .B(n18204), .ZN(
        P3_U2900) );
  AOI22_X1 U21239 ( .A1(n18484), .A2(n18242), .B1(n18482), .B2(n18219), .ZN(
        n18207) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18221), .B1(
        n18483), .B2(n18220), .ZN(n18206) );
  OAI211_X1 U21241 ( .C1(n18487), .C2(n18290), .A(n18207), .B(n18206), .ZN(
        P3_U2901) );
  AOI22_X1 U21242 ( .A1(n18490), .A2(n18242), .B1(n18488), .B2(n18219), .ZN(
        n18209) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18221), .B1(
        n18390), .B2(n18279), .ZN(n18208) );
  OAI211_X1 U21244 ( .C1(n18393), .C2(n18212), .A(n18209), .B(n18208), .ZN(
        P3_U2902) );
  AOI22_X1 U21245 ( .A1(n18494), .A2(n18219), .B1(n18496), .B2(n18242), .ZN(
        n18211) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18221), .B1(
        n18450), .B2(n18279), .ZN(n18210) );
  OAI211_X1 U21247 ( .C1(n18453), .C2(n18212), .A(n18211), .B(n18210), .ZN(
        P3_U2903) );
  AOI22_X1 U21248 ( .A1(n18501), .A2(n18220), .B1(n18500), .B2(n18219), .ZN(
        n18214) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18221), .B1(
        n18502), .B2(n18242), .ZN(n18213) );
  OAI211_X1 U21250 ( .C1(n18505), .C2(n18290), .A(n18214), .B(n18213), .ZN(
        P3_U2904) );
  AOI22_X1 U21251 ( .A1(n18425), .A2(n18220), .B1(n18507), .B2(n18219), .ZN(
        n18216) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18221), .B1(
        n18510), .B2(n18279), .ZN(n18215) );
  OAI211_X1 U21253 ( .C1(n18428), .C2(n18224), .A(n18216), .B(n18215), .ZN(
        P3_U2905) );
  AOI22_X1 U21254 ( .A1(n18516), .A2(n18219), .B1(n18515), .B2(n18220), .ZN(
        n18218) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18221), .B1(
        n18517), .B2(n18279), .ZN(n18217) );
  OAI211_X1 U21256 ( .C1(n18520), .C2(n18224), .A(n18218), .B(n18217), .ZN(
        P3_U2906) );
  AOI22_X1 U21257 ( .A1(n18524), .A2(n18220), .B1(n18522), .B2(n18219), .ZN(
        n18223) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18221), .B1(
        n18525), .B2(n18279), .ZN(n18222) );
  OAI211_X1 U21259 ( .C1(n18530), .C2(n18224), .A(n18223), .B(n18222), .ZN(
        P3_U2907) );
  NAND2_X1 U21260 ( .A1(n18270), .A2(n18314), .ZN(n18313) );
  INV_X1 U21261 ( .A(n18270), .ZN(n18225) );
  NOR2_X1 U21262 ( .A1(n18225), .A2(n18316), .ZN(n18241) );
  AOI22_X1 U21263 ( .A1(n18473), .A2(n18242), .B1(n18472), .B2(n18241), .ZN(
        n18228) );
  AOI22_X1 U21264 ( .A1(n18477), .A2(n18226), .B1(n18270), .B2(n18412), .ZN(
        n18243) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18243), .B1(
        n18478), .B2(n18261), .ZN(n18227) );
  OAI211_X1 U21266 ( .C1(n18481), .C2(n18313), .A(n18228), .B(n18227), .ZN(
        P3_U2908) );
  AOI22_X1 U21267 ( .A1(n18483), .A2(n18242), .B1(n18482), .B2(n18241), .ZN(
        n18230) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18243), .B1(
        n18484), .B2(n18261), .ZN(n18229) );
  OAI211_X1 U21269 ( .C1(n18487), .C2(n18313), .A(n18230), .B(n18229), .ZN(
        P3_U2909) );
  AOI22_X1 U21270 ( .A1(n18490), .A2(n18261), .B1(n18488), .B2(n18241), .ZN(
        n18232) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18243), .B1(
        n18489), .B2(n18242), .ZN(n18231) );
  OAI211_X1 U21272 ( .C1(n18493), .C2(n18313), .A(n18232), .B(n18231), .ZN(
        P3_U2910) );
  AOI22_X1 U21273 ( .A1(n18495), .A2(n18242), .B1(n18494), .B2(n18241), .ZN(
        n18234) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18243), .B1(
        n18496), .B2(n18261), .ZN(n18233) );
  OAI211_X1 U21275 ( .C1(n18499), .C2(n18313), .A(n18234), .B(n18233), .ZN(
        P3_U2911) );
  AOI22_X1 U21276 ( .A1(n18502), .A2(n18261), .B1(n18500), .B2(n18241), .ZN(
        n18236) );
  AOI22_X1 U21277 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18243), .B1(
        n18501), .B2(n18242), .ZN(n18235) );
  OAI211_X1 U21278 ( .C1(n18505), .C2(n18313), .A(n18236), .B(n18235), .ZN(
        P3_U2912) );
  AOI22_X1 U21279 ( .A1(n18425), .A2(n18242), .B1(n18507), .B2(n18241), .ZN(
        n18238) );
  INV_X1 U21280 ( .A(n18313), .ZN(n18304) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18243), .B1(
        n18510), .B2(n18304), .ZN(n18237) );
  OAI211_X1 U21282 ( .C1(n18428), .C2(n18268), .A(n18238), .B(n18237), .ZN(
        P3_U2913) );
  AOI22_X1 U21283 ( .A1(n18516), .A2(n18241), .B1(n18515), .B2(n18242), .ZN(
        n18240) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18243), .B1(
        n18517), .B2(n18304), .ZN(n18239) );
  OAI211_X1 U21285 ( .C1(n18520), .C2(n18268), .A(n18240), .B(n18239), .ZN(
        P3_U2914) );
  AOI22_X1 U21286 ( .A1(n18524), .A2(n18242), .B1(n18522), .B2(n18241), .ZN(
        n18245) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18243), .B1(
        n18525), .B2(n18304), .ZN(n18244) );
  OAI211_X1 U21288 ( .C1(n18530), .C2(n18268), .A(n18245), .B(n18244), .ZN(
        P3_U2915) );
  NOR2_X1 U21289 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18246), .ZN(
        n18317) );
  NAND2_X1 U21290 ( .A1(n18317), .A2(n18575), .ZN(n18330) );
  INV_X1 U21291 ( .A(n18330), .ZN(n18334) );
  NOR2_X1 U21292 ( .A1(n18304), .A2(n18334), .ZN(n18292) );
  NOR2_X1 U21293 ( .A1(n18605), .A2(n18292), .ZN(n18264) );
  AOI22_X1 U21294 ( .A1(n18473), .A2(n18261), .B1(n18472), .B2(n18264), .ZN(
        n18250) );
  OAI21_X1 U21295 ( .B1(n18247), .B2(n18382), .A(n18292), .ZN(n18248) );
  OAI211_X1 U21296 ( .C1(n18334), .C2(n18704), .A(n18385), .B(n18248), .ZN(
        n18265) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18265), .B1(
        n18478), .B2(n18279), .ZN(n18249) );
  OAI211_X1 U21298 ( .C1(n18481), .C2(n18330), .A(n18250), .B(n18249), .ZN(
        P3_U2916) );
  AOI22_X1 U21299 ( .A1(n18484), .A2(n18279), .B1(n18482), .B2(n18264), .ZN(
        n18252) );
  AOI22_X1 U21300 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18265), .B1(
        n18483), .B2(n18261), .ZN(n18251) );
  OAI211_X1 U21301 ( .C1(n18487), .C2(n18330), .A(n18252), .B(n18251), .ZN(
        P3_U2917) );
  AOI22_X1 U21302 ( .A1(n18490), .A2(n18279), .B1(n18488), .B2(n18264), .ZN(
        n18254) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18265), .B1(
        n18390), .B2(n18334), .ZN(n18253) );
  OAI211_X1 U21304 ( .C1(n18393), .C2(n18268), .A(n18254), .B(n18253), .ZN(
        P3_U2918) );
  AOI22_X1 U21305 ( .A1(n18495), .A2(n18261), .B1(n18494), .B2(n18264), .ZN(
        n18256) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18265), .B1(
        n18496), .B2(n18279), .ZN(n18255) );
  OAI211_X1 U21307 ( .C1(n18499), .C2(n18330), .A(n18256), .B(n18255), .ZN(
        P3_U2919) );
  AOI22_X1 U21308 ( .A1(n18501), .A2(n18261), .B1(n18500), .B2(n18264), .ZN(
        n18258) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18265), .B1(
        n18502), .B2(n18279), .ZN(n18257) );
  OAI211_X1 U21310 ( .C1(n18505), .C2(n18330), .A(n18258), .B(n18257), .ZN(
        P3_U2920) );
  AOI22_X1 U21311 ( .A1(n18425), .A2(n18261), .B1(n18507), .B2(n18264), .ZN(
        n18260) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18265), .B1(
        n18510), .B2(n18334), .ZN(n18259) );
  OAI211_X1 U21313 ( .C1(n18428), .C2(n18290), .A(n18260), .B(n18259), .ZN(
        P3_U2921) );
  AOI22_X1 U21314 ( .A1(n18516), .A2(n18264), .B1(n18515), .B2(n18261), .ZN(
        n18263) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18265), .B1(
        n18517), .B2(n18334), .ZN(n18262) );
  OAI211_X1 U21316 ( .C1(n18520), .C2(n18290), .A(n18263), .B(n18262), .ZN(
        P3_U2922) );
  AOI22_X1 U21317 ( .A1(n18404), .A2(n18279), .B1(n18522), .B2(n18264), .ZN(
        n18267) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18265), .B1(
        n18525), .B2(n18334), .ZN(n18266) );
  OAI211_X1 U21319 ( .C1(n18409), .C2(n18268), .A(n18267), .B(n18266), .ZN(
        P3_U2923) );
  NAND2_X1 U21320 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18317), .ZN(
        n18355) );
  AND2_X1 U21321 ( .A1(n18437), .A2(n18317), .ZN(n18286) );
  AOI22_X1 U21322 ( .A1(n18473), .A2(n18279), .B1(n18472), .B2(n18286), .ZN(
        n18272) );
  NAND2_X1 U21323 ( .A1(n18270), .A2(n18269), .ZN(n18287) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18287), .B1(
        n18478), .B2(n18304), .ZN(n18271) );
  OAI211_X1 U21325 ( .C1(n18481), .C2(n18355), .A(n18272), .B(n18271), .ZN(
        P3_U2924) );
  AOI22_X1 U21326 ( .A1(n18483), .A2(n18279), .B1(n18482), .B2(n18286), .ZN(
        n18274) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18287), .B1(
        n18484), .B2(n18304), .ZN(n18273) );
  OAI211_X1 U21328 ( .C1(n18487), .C2(n18355), .A(n18274), .B(n18273), .ZN(
        P3_U2925) );
  AOI22_X1 U21329 ( .A1(n18489), .A2(n18279), .B1(n18488), .B2(n18286), .ZN(
        n18276) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18287), .B1(
        n18490), .B2(n18304), .ZN(n18275) );
  OAI211_X1 U21331 ( .C1(n18493), .C2(n18355), .A(n18276), .B(n18275), .ZN(
        P3_U2926) );
  AOI22_X1 U21332 ( .A1(n18494), .A2(n18286), .B1(n18496), .B2(n18304), .ZN(
        n18278) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18287), .B1(
        n18495), .B2(n18279), .ZN(n18277) );
  OAI211_X1 U21334 ( .C1(n18499), .C2(n18355), .A(n18278), .B(n18277), .ZN(
        P3_U2927) );
  AOI22_X1 U21335 ( .A1(n18502), .A2(n18304), .B1(n18500), .B2(n18286), .ZN(
        n18281) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18287), .B1(
        n18501), .B2(n18279), .ZN(n18280) );
  OAI211_X1 U21337 ( .C1(n18505), .C2(n18355), .A(n18281), .B(n18280), .ZN(
        P3_U2928) );
  AOI22_X1 U21338 ( .A1(n18508), .A2(n18304), .B1(n18507), .B2(n18286), .ZN(
        n18283) );
  INV_X1 U21339 ( .A(n18355), .ZN(n18357) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18287), .B1(
        n18510), .B2(n18357), .ZN(n18282) );
  OAI211_X1 U21341 ( .C1(n18514), .C2(n18290), .A(n18283), .B(n18282), .ZN(
        P3_U2929) );
  AOI22_X1 U21342 ( .A1(n18460), .A2(n18304), .B1(n18516), .B2(n18286), .ZN(
        n18285) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18287), .B1(
        n18517), .B2(n18357), .ZN(n18284) );
  OAI211_X1 U21344 ( .C1(n18464), .C2(n18290), .A(n18285), .B(n18284), .ZN(
        P3_U2930) );
  AOI22_X1 U21345 ( .A1(n18404), .A2(n18304), .B1(n18522), .B2(n18286), .ZN(
        n18289) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18287), .B1(
        n18525), .B2(n18357), .ZN(n18288) );
  OAI211_X1 U21347 ( .C1(n18409), .C2(n18290), .A(n18289), .B(n18288), .ZN(
        P3_U2931) );
  NAND2_X1 U21348 ( .A1(n18579), .A2(n18315), .ZN(n18381) );
  INV_X1 U21349 ( .A(n18381), .ZN(n18370) );
  NOR2_X1 U21350 ( .A1(n18357), .A2(n18370), .ZN(n18339) );
  NOR2_X1 U21351 ( .A1(n18605), .A2(n18339), .ZN(n18309) );
  AOI22_X1 U21352 ( .A1(n18478), .A2(n18334), .B1(n18472), .B2(n18309), .ZN(
        n18295) );
  INV_X1 U21353 ( .A(n18439), .ZN(n18291) );
  AOI221_X1 U21354 ( .B1(n18339), .B2(n18382), .C1(n18339), .C2(n18292), .A(
        n18291), .ZN(n18293) );
  INV_X1 U21355 ( .A(n18293), .ZN(n18310) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18310), .B1(
        n18473), .B2(n18304), .ZN(n18294) );
  OAI211_X1 U21357 ( .C1(n18481), .C2(n18381), .A(n18295), .B(n18294), .ZN(
        P3_U2932) );
  AOI22_X1 U21358 ( .A1(n18483), .A2(n18304), .B1(n18482), .B2(n18309), .ZN(
        n18297) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18310), .B1(
        n18484), .B2(n18334), .ZN(n18296) );
  OAI211_X1 U21360 ( .C1(n18487), .C2(n18381), .A(n18297), .B(n18296), .ZN(
        P3_U2933) );
  AOI22_X1 U21361 ( .A1(n18490), .A2(n18334), .B1(n18488), .B2(n18309), .ZN(
        n18299) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18310), .B1(
        n18390), .B2(n18370), .ZN(n18298) );
  OAI211_X1 U21363 ( .C1(n18393), .C2(n18313), .A(n18299), .B(n18298), .ZN(
        P3_U2934) );
  AOI22_X1 U21364 ( .A1(n18495), .A2(n18304), .B1(n18494), .B2(n18309), .ZN(
        n18301) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18310), .B1(
        n18496), .B2(n18334), .ZN(n18300) );
  OAI211_X1 U21366 ( .C1(n18499), .C2(n18381), .A(n18301), .B(n18300), .ZN(
        P3_U2935) );
  AOI22_X1 U21367 ( .A1(n18501), .A2(n18304), .B1(n18500), .B2(n18309), .ZN(
        n18303) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18310), .B1(
        n18502), .B2(n18334), .ZN(n18302) );
  OAI211_X1 U21369 ( .C1(n18505), .C2(n18381), .A(n18303), .B(n18302), .ZN(
        P3_U2936) );
  AOI22_X1 U21370 ( .A1(n18425), .A2(n18304), .B1(n18507), .B2(n18309), .ZN(
        n18306) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18310), .B1(
        n18510), .B2(n18370), .ZN(n18305) );
  OAI211_X1 U21372 ( .C1(n18428), .C2(n18330), .A(n18306), .B(n18305), .ZN(
        P3_U2937) );
  AOI22_X1 U21373 ( .A1(n18460), .A2(n18334), .B1(n18516), .B2(n18309), .ZN(
        n18308) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18310), .B1(
        n18517), .B2(n18370), .ZN(n18307) );
  OAI211_X1 U21375 ( .C1(n18464), .C2(n18313), .A(n18308), .B(n18307), .ZN(
        P3_U2938) );
  AOI22_X1 U21376 ( .A1(n18404), .A2(n18334), .B1(n18522), .B2(n18309), .ZN(
        n18312) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18310), .B1(
        n18525), .B2(n18370), .ZN(n18311) );
  OAI211_X1 U21378 ( .C1(n18409), .C2(n18313), .A(n18312), .B(n18311), .ZN(
        P3_U2939) );
  NAND2_X1 U21379 ( .A1(n18315), .A2(n18314), .ZN(n18408) );
  INV_X1 U21380 ( .A(n18315), .ZN(n18338) );
  NOR2_X1 U21381 ( .A1(n18338), .A2(n18316), .ZN(n18333) );
  AOI22_X1 U21382 ( .A1(n18478), .A2(n18357), .B1(n18472), .B2(n18333), .ZN(
        n18319) );
  NOR2_X1 U21383 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18338), .ZN(
        n18361) );
  AOI22_X1 U21384 ( .A1(n18477), .A2(n18317), .B1(n18474), .B2(n18361), .ZN(
        n18335) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18335), .B1(
        n18473), .B2(n18334), .ZN(n18318) );
  OAI211_X1 U21386 ( .C1(n18481), .C2(n18408), .A(n18319), .B(n18318), .ZN(
        P3_U2940) );
  AOI22_X1 U21387 ( .A1(n18483), .A2(n18334), .B1(n18482), .B2(n18333), .ZN(
        n18321) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18335), .B1(
        n18484), .B2(n18357), .ZN(n18320) );
  OAI211_X1 U21389 ( .C1(n18487), .C2(n18408), .A(n18321), .B(n18320), .ZN(
        P3_U2941) );
  AOI22_X1 U21390 ( .A1(n18489), .A2(n18334), .B1(n18488), .B2(n18333), .ZN(
        n18323) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18335), .B1(
        n18490), .B2(n18357), .ZN(n18322) );
  OAI211_X1 U21392 ( .C1(n18493), .C2(n18408), .A(n18323), .B(n18322), .ZN(
        P3_U2942) );
  AOI22_X1 U21393 ( .A1(n18494), .A2(n18333), .B1(n18496), .B2(n18357), .ZN(
        n18325) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18335), .B1(
        n18495), .B2(n18334), .ZN(n18324) );
  OAI211_X1 U21395 ( .C1(n18499), .C2(n18408), .A(n18325), .B(n18324), .ZN(
        P3_U2943) );
  AOI22_X1 U21396 ( .A1(n18502), .A2(n18357), .B1(n18500), .B2(n18333), .ZN(
        n18327) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18335), .B1(
        n18501), .B2(n18334), .ZN(n18326) );
  OAI211_X1 U21398 ( .C1(n18505), .C2(n18408), .A(n18327), .B(n18326), .ZN(
        P3_U2944) );
  AOI22_X1 U21399 ( .A1(n18508), .A2(n18357), .B1(n18507), .B2(n18333), .ZN(
        n18329) );
  INV_X1 U21400 ( .A(n18408), .ZN(n18400) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18335), .B1(
        n18510), .B2(n18400), .ZN(n18328) );
  OAI211_X1 U21402 ( .C1(n18514), .C2(n18330), .A(n18329), .B(n18328), .ZN(
        P3_U2945) );
  AOI22_X1 U21403 ( .A1(n18516), .A2(n18333), .B1(n18515), .B2(n18334), .ZN(
        n18332) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18335), .B1(
        n18517), .B2(n18400), .ZN(n18331) );
  OAI211_X1 U21405 ( .C1(n18520), .C2(n18355), .A(n18332), .B(n18331), .ZN(
        P3_U2946) );
  AOI22_X1 U21406 ( .A1(n18524), .A2(n18334), .B1(n18522), .B2(n18333), .ZN(
        n18337) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18335), .B1(
        n18525), .B2(n18400), .ZN(n18336) );
  OAI211_X1 U21408 ( .C1(n18530), .C2(n18355), .A(n18337), .B(n18336), .ZN(
        P3_U2947) );
  NOR2_X1 U21409 ( .A1(n18576), .A2(n18338), .ZN(n18414) );
  NAND2_X1 U21410 ( .A1(n18414), .A2(n18575), .ZN(n18431) );
  INV_X1 U21411 ( .A(n18431), .ZN(n18433) );
  NOR2_X1 U21412 ( .A1(n18400), .A2(n18433), .ZN(n18383) );
  NOR2_X1 U21413 ( .A1(n18605), .A2(n18383), .ZN(n18356) );
  AOI22_X1 U21414 ( .A1(n18478), .A2(n18370), .B1(n18472), .B2(n18356), .ZN(
        n18342) );
  OAI21_X1 U21415 ( .B1(n18339), .B2(n18382), .A(n18383), .ZN(n18340) );
  OAI211_X1 U21416 ( .C1(n18433), .C2(n18704), .A(n18385), .B(n18340), .ZN(
        n18358) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18358), .B1(
        n18473), .B2(n18357), .ZN(n18341) );
  OAI211_X1 U21418 ( .C1(n18481), .C2(n18431), .A(n18342), .B(n18341), .ZN(
        P3_U2948) );
  AOI22_X1 U21419 ( .A1(n18483), .A2(n18357), .B1(n18482), .B2(n18356), .ZN(
        n18344) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18358), .B1(
        n18484), .B2(n18370), .ZN(n18343) );
  OAI211_X1 U21421 ( .C1(n18487), .C2(n18431), .A(n18344), .B(n18343), .ZN(
        P3_U2949) );
  AOI22_X1 U21422 ( .A1(n18490), .A2(n18370), .B1(n18488), .B2(n18356), .ZN(
        n18346) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18358), .B1(
        n18390), .B2(n18433), .ZN(n18345) );
  OAI211_X1 U21424 ( .C1(n18393), .C2(n18355), .A(n18346), .B(n18345), .ZN(
        P3_U2950) );
  AOI22_X1 U21425 ( .A1(n18495), .A2(n18357), .B1(n18494), .B2(n18356), .ZN(
        n18348) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18358), .B1(
        n18496), .B2(n18370), .ZN(n18347) );
  OAI211_X1 U21427 ( .C1(n18499), .C2(n18431), .A(n18348), .B(n18347), .ZN(
        P3_U2951) );
  AOI22_X1 U21428 ( .A1(n18502), .A2(n18370), .B1(n18500), .B2(n18356), .ZN(
        n18350) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18358), .B1(
        n18454), .B2(n18433), .ZN(n18349) );
  OAI211_X1 U21430 ( .C1(n18457), .C2(n18355), .A(n18350), .B(n18349), .ZN(
        P3_U2952) );
  AOI22_X1 U21431 ( .A1(n18508), .A2(n18370), .B1(n18507), .B2(n18356), .ZN(
        n18352) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18358), .B1(
        n18510), .B2(n18433), .ZN(n18351) );
  OAI211_X1 U21433 ( .C1(n18514), .C2(n18355), .A(n18352), .B(n18351), .ZN(
        P3_U2953) );
  AOI22_X1 U21434 ( .A1(n18460), .A2(n18370), .B1(n18516), .B2(n18356), .ZN(
        n18354) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18358), .B1(
        n18517), .B2(n18433), .ZN(n18353) );
  OAI211_X1 U21436 ( .C1(n18464), .C2(n18355), .A(n18354), .B(n18353), .ZN(
        P3_U2954) );
  AOI22_X1 U21437 ( .A1(n18524), .A2(n18357), .B1(n18522), .B2(n18356), .ZN(
        n18360) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18358), .B1(
        n18525), .B2(n18433), .ZN(n18359) );
  OAI211_X1 U21439 ( .C1(n18530), .C2(n18381), .A(n18360), .B(n18359), .ZN(
        P3_U2955) );
  NAND2_X1 U21440 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18414), .ZN(
        n18463) );
  AND2_X1 U21441 ( .A1(n18437), .A2(n18414), .ZN(n18377) );
  AOI22_X1 U21442 ( .A1(n18478), .A2(n18400), .B1(n18472), .B2(n18377), .ZN(
        n18363) );
  AOI22_X1 U21443 ( .A1(n18477), .A2(n18361), .B1(n18474), .B2(n18414), .ZN(
        n18378) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18378), .B1(
        n18473), .B2(n18370), .ZN(n18362) );
  OAI211_X1 U21445 ( .C1(n18481), .C2(n18463), .A(n18363), .B(n18362), .ZN(
        P3_U2956) );
  AOI22_X1 U21446 ( .A1(n18483), .A2(n18370), .B1(n18482), .B2(n18377), .ZN(
        n18365) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18378), .B1(
        n18484), .B2(n18400), .ZN(n18364) );
  OAI211_X1 U21448 ( .C1(n18487), .C2(n18463), .A(n18365), .B(n18364), .ZN(
        P3_U2957) );
  AOI22_X1 U21449 ( .A1(n18490), .A2(n18400), .B1(n18488), .B2(n18377), .ZN(
        n18367) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18378), .B1(
        n18489), .B2(n18370), .ZN(n18366) );
  OAI211_X1 U21451 ( .C1(n18493), .C2(n18463), .A(n18367), .B(n18366), .ZN(
        P3_U2958) );
  AOI22_X1 U21452 ( .A1(n18495), .A2(n18370), .B1(n18494), .B2(n18377), .ZN(
        n18369) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18378), .B1(
        n18496), .B2(n18400), .ZN(n18368) );
  OAI211_X1 U21454 ( .C1(n18499), .C2(n18463), .A(n18369), .B(n18368), .ZN(
        P3_U2959) );
  AOI22_X1 U21455 ( .A1(n18502), .A2(n18400), .B1(n18500), .B2(n18377), .ZN(
        n18372) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18378), .B1(
        n18501), .B2(n18370), .ZN(n18371) );
  OAI211_X1 U21457 ( .C1(n18505), .C2(n18463), .A(n18372), .B(n18371), .ZN(
        P3_U2960) );
  AOI22_X1 U21458 ( .A1(n18508), .A2(n18400), .B1(n18507), .B2(n18377), .ZN(
        n18374) );
  INV_X1 U21459 ( .A(n18463), .ZN(n18466) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18378), .B1(
        n18510), .B2(n18466), .ZN(n18373) );
  OAI211_X1 U21461 ( .C1(n18514), .C2(n18381), .A(n18374), .B(n18373), .ZN(
        P3_U2961) );
  AOI22_X1 U21462 ( .A1(n18460), .A2(n18400), .B1(n18516), .B2(n18377), .ZN(
        n18376) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18378), .B1(
        n18517), .B2(n18466), .ZN(n18375) );
  OAI211_X1 U21464 ( .C1(n18464), .C2(n18381), .A(n18376), .B(n18375), .ZN(
        P3_U2962) );
  AOI22_X1 U21465 ( .A1(n18404), .A2(n18400), .B1(n18522), .B2(n18377), .ZN(
        n18380) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18378), .B1(
        n18525), .B2(n18466), .ZN(n18379) );
  OAI211_X1 U21467 ( .C1(n18409), .C2(n18381), .A(n18380), .B(n18379), .ZN(
        P3_U2963) );
  INV_X1 U21468 ( .A(n18410), .ZN(n18476) );
  NAND2_X1 U21469 ( .A1(n18476), .A2(n18575), .ZN(n18513) );
  INV_X1 U21470 ( .A(n18513), .ZN(n18523) );
  NOR2_X1 U21471 ( .A1(n18466), .A2(n18523), .ZN(n18438) );
  NOR2_X1 U21472 ( .A1(n18605), .A2(n18438), .ZN(n18403) );
  AOI22_X1 U21473 ( .A1(n18473), .A2(n18400), .B1(n18472), .B2(n18403), .ZN(
        n18387) );
  OAI21_X1 U21474 ( .B1(n18383), .B2(n18382), .A(n18438), .ZN(n18384) );
  OAI211_X1 U21475 ( .C1(n18523), .C2(n18704), .A(n18385), .B(n18384), .ZN(
        n18405) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18405), .B1(
        n18478), .B2(n18433), .ZN(n18386) );
  OAI211_X1 U21477 ( .C1(n18481), .C2(n18513), .A(n18387), .B(n18386), .ZN(
        P3_U2964) );
  AOI22_X1 U21478 ( .A1(n18483), .A2(n18400), .B1(n18482), .B2(n18403), .ZN(
        n18389) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18405), .B1(
        n18484), .B2(n18433), .ZN(n18388) );
  OAI211_X1 U21480 ( .C1(n18487), .C2(n18513), .A(n18389), .B(n18388), .ZN(
        P3_U2965) );
  AOI22_X1 U21481 ( .A1(n18490), .A2(n18433), .B1(n18488), .B2(n18403), .ZN(
        n18392) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18405), .B1(
        n18390), .B2(n18523), .ZN(n18391) );
  OAI211_X1 U21483 ( .C1(n18393), .C2(n18408), .A(n18392), .B(n18391), .ZN(
        P3_U2966) );
  AOI22_X1 U21484 ( .A1(n18495), .A2(n18400), .B1(n18494), .B2(n18403), .ZN(
        n18395) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18405), .B1(
        n18496), .B2(n18433), .ZN(n18394) );
  OAI211_X1 U21486 ( .C1(n18499), .C2(n18513), .A(n18395), .B(n18394), .ZN(
        P3_U2967) );
  AOI22_X1 U21487 ( .A1(n18502), .A2(n18433), .B1(n18500), .B2(n18403), .ZN(
        n18397) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18405), .B1(
        n18454), .B2(n18523), .ZN(n18396) );
  OAI211_X1 U21489 ( .C1(n18457), .C2(n18408), .A(n18397), .B(n18396), .ZN(
        P3_U2968) );
  AOI22_X1 U21490 ( .A1(n18508), .A2(n18433), .B1(n18507), .B2(n18403), .ZN(
        n18399) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18405), .B1(
        n18510), .B2(n18523), .ZN(n18398) );
  OAI211_X1 U21492 ( .C1(n18514), .C2(n18408), .A(n18399), .B(n18398), .ZN(
        P3_U2969) );
  AOI22_X1 U21493 ( .A1(n18516), .A2(n18403), .B1(n18515), .B2(n18400), .ZN(
        n18402) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18405), .B1(
        n18517), .B2(n18523), .ZN(n18401) );
  OAI211_X1 U21495 ( .C1(n18520), .C2(n18431), .A(n18402), .B(n18401), .ZN(
        P3_U2970) );
  AOI22_X1 U21496 ( .A1(n18404), .A2(n18433), .B1(n18522), .B2(n18403), .ZN(
        n18407) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18405), .B1(
        n18525), .B2(n18523), .ZN(n18406) );
  OAI211_X1 U21498 ( .C1(n18409), .C2(n18408), .A(n18407), .B(n18406), .ZN(
        P3_U2971) );
  NOR2_X1 U21499 ( .A1(n18605), .A2(n18410), .ZN(n18432) );
  AOI22_X1 U21500 ( .A1(n18478), .A2(n18466), .B1(n18472), .B2(n18432), .ZN(
        n18416) );
  NOR2_X1 U21501 ( .A1(n18411), .A2(n18585), .ZN(n18413) );
  AOI22_X1 U21502 ( .A1(n18477), .A2(n18414), .B1(n18413), .B2(n18412), .ZN(
        n18434) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18434), .B1(
        n18473), .B2(n18433), .ZN(n18415) );
  OAI211_X1 U21504 ( .C1(n18531), .C2(n18481), .A(n18416), .B(n18415), .ZN(
        P3_U2972) );
  AOI22_X1 U21505 ( .A1(n18483), .A2(n18433), .B1(n18482), .B2(n18432), .ZN(
        n18418) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18434), .B1(
        n18484), .B2(n18466), .ZN(n18417) );
  OAI211_X1 U21507 ( .C1(n18531), .C2(n18487), .A(n18418), .B(n18417), .ZN(
        P3_U2973) );
  AOI22_X1 U21508 ( .A1(n18489), .A2(n18433), .B1(n18488), .B2(n18432), .ZN(
        n18420) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18434), .B1(
        n18490), .B2(n18466), .ZN(n18419) );
  OAI211_X1 U21510 ( .C1(n18531), .C2(n18493), .A(n18420), .B(n18419), .ZN(
        P3_U2974) );
  AOI22_X1 U21511 ( .A1(n18495), .A2(n18433), .B1(n18494), .B2(n18432), .ZN(
        n18422) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18434), .B1(
        n18496), .B2(n18466), .ZN(n18421) );
  OAI211_X1 U21513 ( .C1(n18531), .C2(n18499), .A(n18422), .B(n18421), .ZN(
        P3_U2975) );
  AOI22_X1 U21514 ( .A1(n18502), .A2(n18466), .B1(n18500), .B2(n18432), .ZN(
        n18424) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18434), .B1(
        n18509), .B2(n18454), .ZN(n18423) );
  OAI211_X1 U21516 ( .C1(n18457), .C2(n18431), .A(n18424), .B(n18423), .ZN(
        P3_U2976) );
  AOI22_X1 U21517 ( .A1(n18425), .A2(n18433), .B1(n18507), .B2(n18432), .ZN(
        n18427) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18434), .B1(
        n18509), .B2(n18510), .ZN(n18426) );
  OAI211_X1 U21519 ( .C1(n18428), .C2(n18463), .A(n18427), .B(n18426), .ZN(
        P3_U2977) );
  AOI22_X1 U21520 ( .A1(n18460), .A2(n18466), .B1(n18516), .B2(n18432), .ZN(
        n18430) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18434), .B1(
        n18509), .B2(n18517), .ZN(n18429) );
  OAI211_X1 U21522 ( .C1(n18464), .C2(n18431), .A(n18430), .B(n18429), .ZN(
        P3_U2978) );
  AOI22_X1 U21523 ( .A1(n18524), .A2(n18433), .B1(n18522), .B2(n18432), .ZN(
        n18436) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18434), .B1(
        n18509), .B2(n18525), .ZN(n18435) );
  OAI211_X1 U21525 ( .C1(n18530), .C2(n18463), .A(n18436), .B(n18435), .ZN(
        P3_U2979) );
  AND2_X1 U21526 ( .A1(n18437), .A2(n18442), .ZN(n18465) );
  AOI22_X1 U21527 ( .A1(n18478), .A2(n18523), .B1(n18472), .B2(n18465), .ZN(
        n18444) );
  INV_X1 U21528 ( .A(n18438), .ZN(n18440) );
  OAI221_X1 U21529 ( .B1(n18442), .B2(n18441), .C1(n18442), .C2(n18440), .A(
        n18439), .ZN(n18468) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18468), .B1(
        n18473), .B2(n18466), .ZN(n18443) );
  OAI211_X1 U21531 ( .C1(n18449), .C2(n18481), .A(n18444), .B(n18443), .ZN(
        P3_U2980) );
  AOI22_X1 U21532 ( .A1(n18483), .A2(n18466), .B1(n18482), .B2(n18465), .ZN(
        n18446) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18468), .B1(
        n18484), .B2(n18523), .ZN(n18445) );
  OAI211_X1 U21534 ( .C1(n18449), .C2(n18487), .A(n18446), .B(n18445), .ZN(
        P3_U2981) );
  AOI22_X1 U21535 ( .A1(n18489), .A2(n18466), .B1(n18488), .B2(n18465), .ZN(
        n18448) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18468), .B1(
        n18490), .B2(n18523), .ZN(n18447) );
  OAI211_X1 U21537 ( .C1(n18449), .C2(n18493), .A(n18448), .B(n18447), .ZN(
        P3_U2982) );
  AOI22_X1 U21538 ( .A1(n18494), .A2(n18465), .B1(n18496), .B2(n18523), .ZN(
        n18452) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18468), .B1(
        n18467), .B2(n18450), .ZN(n18451) );
  OAI211_X1 U21540 ( .C1(n18453), .C2(n18463), .A(n18452), .B(n18451), .ZN(
        P3_U2983) );
  AOI22_X1 U21541 ( .A1(n18502), .A2(n18523), .B1(n18500), .B2(n18465), .ZN(
        n18456) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18468), .B1(
        n18467), .B2(n18454), .ZN(n18455) );
  OAI211_X1 U21543 ( .C1(n18457), .C2(n18463), .A(n18456), .B(n18455), .ZN(
        P3_U2984) );
  AOI22_X1 U21544 ( .A1(n18508), .A2(n18523), .B1(n18507), .B2(n18465), .ZN(
        n18459) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18468), .B1(
        n18467), .B2(n18510), .ZN(n18458) );
  OAI211_X1 U21546 ( .C1(n18514), .C2(n18463), .A(n18459), .B(n18458), .ZN(
        P3_U2985) );
  AOI22_X1 U21547 ( .A1(n18460), .A2(n18523), .B1(n18516), .B2(n18465), .ZN(
        n18462) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18468), .B1(
        n18467), .B2(n18517), .ZN(n18461) );
  OAI211_X1 U21549 ( .C1(n18464), .C2(n18463), .A(n18462), .B(n18461), .ZN(
        P3_U2986) );
  AOI22_X1 U21550 ( .A1(n18524), .A2(n18466), .B1(n18522), .B2(n18465), .ZN(
        n18470) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18468), .B1(
        n18467), .B2(n18525), .ZN(n18469) );
  OAI211_X1 U21552 ( .C1(n18530), .C2(n18513), .A(n18470), .B(n18469), .ZN(
        P3_U2987) );
  NOR2_X1 U21553 ( .A1(n18605), .A2(n18471), .ZN(n18521) );
  AOI22_X1 U21554 ( .A1(n18473), .A2(n18523), .B1(n18472), .B2(n18521), .ZN(
        n18480) );
  AOI22_X1 U21555 ( .A1(n18477), .A2(n18476), .B1(n18475), .B2(n18474), .ZN(
        n18527) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18527), .B1(
        n18509), .B2(n18478), .ZN(n18479) );
  OAI211_X1 U21557 ( .C1(n18506), .C2(n18481), .A(n18480), .B(n18479), .ZN(
        P3_U2988) );
  AOI22_X1 U21558 ( .A1(n18483), .A2(n18523), .B1(n18482), .B2(n18521), .ZN(
        n18486) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18527), .B1(
        n18509), .B2(n18484), .ZN(n18485) );
  OAI211_X1 U21560 ( .C1(n18506), .C2(n18487), .A(n18486), .B(n18485), .ZN(
        P3_U2989) );
  AOI22_X1 U21561 ( .A1(n18489), .A2(n18523), .B1(n18488), .B2(n18521), .ZN(
        n18492) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18527), .B1(
        n18509), .B2(n18490), .ZN(n18491) );
  OAI211_X1 U21563 ( .C1(n18506), .C2(n18493), .A(n18492), .B(n18491), .ZN(
        P3_U2990) );
  AOI22_X1 U21564 ( .A1(n18495), .A2(n18523), .B1(n18494), .B2(n18521), .ZN(
        n18498) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18527), .B1(
        n18509), .B2(n18496), .ZN(n18497) );
  OAI211_X1 U21566 ( .C1(n18506), .C2(n18499), .A(n18498), .B(n18497), .ZN(
        P3_U2991) );
  AOI22_X1 U21567 ( .A1(n18501), .A2(n18523), .B1(n18500), .B2(n18521), .ZN(
        n18504) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18527), .B1(
        n18509), .B2(n18502), .ZN(n18503) );
  OAI211_X1 U21569 ( .C1(n18506), .C2(n18505), .A(n18504), .B(n18503), .ZN(
        P3_U2992) );
  AOI22_X1 U21570 ( .A1(n18509), .A2(n18508), .B1(n18507), .B2(n18521), .ZN(
        n18512) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18527), .B1(
        n18526), .B2(n18510), .ZN(n18511) );
  OAI211_X1 U21572 ( .C1(n18514), .C2(n18513), .A(n18512), .B(n18511), .ZN(
        P3_U2993) );
  AOI22_X1 U21573 ( .A1(n18516), .A2(n18521), .B1(n18515), .B2(n18523), .ZN(
        n18519) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18527), .B1(
        n18526), .B2(n18517), .ZN(n18518) );
  OAI211_X1 U21575 ( .C1(n18531), .C2(n18520), .A(n18519), .B(n18518), .ZN(
        P3_U2994) );
  AOI22_X1 U21576 ( .A1(n18524), .A2(n18523), .B1(n18522), .B2(n18521), .ZN(
        n18529) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18527), .B1(
        n18526), .B2(n18525), .ZN(n18528) );
  OAI211_X1 U21578 ( .C1(n18531), .C2(n18530), .A(n18529), .B(n18528), .ZN(
        P3_U2995) );
  NAND2_X1 U21579 ( .A1(n18533), .A2(n18532), .ZN(n18534) );
  AOI22_X1 U21580 ( .A1(n18537), .A2(n18536), .B1(n18535), .B2(n18534), .ZN(
        n18538) );
  OAI221_X1 U21581 ( .B1(n18541), .B2(n18540), .C1(n18541), .C2(n18539), .A(
        n18538), .ZN(n18747) );
  OAI21_X1 U21582 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18542), .ZN(n18543) );
  OAI211_X1 U21583 ( .C1(n18580), .C2(n18545), .A(n18544), .B(n18543), .ZN(
        n18592) );
  INV_X1 U21584 ( .A(n18562), .ZN(n18547) );
  NAND2_X1 U21585 ( .A1(n18546), .A2(n18733), .ZN(n18572) );
  AOI22_X1 U21586 ( .A1(n18547), .A2(n18572), .B1(n18559), .B2(n18551), .ZN(
        n18705) );
  NOR2_X1 U21587 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18705), .ZN(
        n18555) );
  AOI21_X1 U21588 ( .B1(n18550), .B2(n18549), .A(n18548), .ZN(n18557) );
  OAI21_X1 U21589 ( .B1(n18552), .B2(n18557), .A(n18551), .ZN(n18553) );
  AOI21_X1 U21590 ( .B1(n18562), .B2(n18574), .A(n18553), .ZN(n18709) );
  NAND2_X1 U21591 ( .A1(n18580), .A2(n18709), .ZN(n18554) );
  AOI22_X1 U21592 ( .A1(n18580), .A2(n18555), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18554), .ZN(n18590) );
  NOR2_X1 U21593 ( .A1(n18556), .A2(n10651), .ZN(n18561) );
  OAI21_X1 U21594 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18558), .A(
        n18557), .ZN(n18560) );
  AOI22_X1 U21595 ( .A1(n18561), .A2(n18560), .B1(n18559), .B2(n18716), .ZN(
        n18568) );
  OAI211_X1 U21596 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18563), .B(n18562), .ZN(
        n18567) );
  NOR2_X1 U21597 ( .A1(n18571), .A2(n18733), .ZN(n18565) );
  OAI211_X1 U21598 ( .C1(n18565), .C2(n18564), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n10651), .ZN(n18566) );
  NAND3_X1 U21599 ( .A1(n18568), .A2(n18567), .A3(n18566), .ZN(n18718) );
  AOI22_X1 U21600 ( .A1(n18569), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18718), .B2(n18580), .ZN(n18589) );
  NAND2_X1 U21601 ( .A1(n18583), .A2(n18585), .ZN(n18588) );
  INV_X1 U21602 ( .A(n18590), .ZN(n18586) );
  NAND2_X1 U21603 ( .A1(n18571), .A2(n18570), .ZN(n18573) );
  AOI22_X1 U21604 ( .A1(n18724), .A2(n18573), .B1(n18727), .B2(n18572), .ZN(
        n18720) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18574), .B1(
        n18573), .B2(n18733), .ZN(n18577) );
  INV_X1 U21606 ( .A(n18577), .ZN(n18729) );
  NOR3_X1 U21607 ( .A1(n18576), .A2(n18575), .A3(n18729), .ZN(n18578) );
  OAI22_X1 U21608 ( .A1(n18720), .A2(n18578), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18577), .ZN(n18581) );
  AOI21_X1 U21609 ( .B1(n18581), .B2(n18580), .A(n18579), .ZN(n18582) );
  AOI222_X1 U21610 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18589), 
        .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18582), .C1(n18589), 
        .C2(n18582), .ZN(n18584) );
  OAI211_X1 U21611 ( .C1(n18586), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        n18587) );
  OAI221_X1 U21612 ( .B1(n18590), .B2(n18589), .C1(n18590), .C2(n18588), .A(
        n18587), .ZN(n18591) );
  NOR4_X1 U21613 ( .A1(n18593), .A2(n18747), .A3(n18592), .A4(n18591), .ZN(
        n18604) );
  AOI22_X1 U21614 ( .A1(n18750), .A2(n18760), .B1(n18728), .B2(n18594), .ZN(
        n18595) );
  INV_X1 U21615 ( .A(n18595), .ZN(n18600) );
  OAI211_X1 U21616 ( .C1(n18597), .C2(n18596), .A(n18757), .B(n18604), .ZN(
        n18703) );
  OAI21_X1 U21617 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18759), .A(n18703), 
        .ZN(n18606) );
  NOR2_X1 U21618 ( .A1(n18598), .A2(n18606), .ZN(n18599) );
  MUX2_X1 U21619 ( .A(n18600), .B(n18599), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18602) );
  OAI211_X1 U21620 ( .C1(n18604), .C2(n18603), .A(n18602), .B(n18601), .ZN(
        P3_U2996) );
  NAND2_X1 U21621 ( .A1(n18750), .A2(n18760), .ZN(n18609) );
  NAND4_X1 U21622 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18750), .A4(n18765), .ZN(n18611) );
  OR3_X1 U21623 ( .A1(n18607), .A2(n18606), .A3(n18605), .ZN(n18608) );
  NAND4_X1 U21624 ( .A1(n18610), .A2(n18609), .A3(n18611), .A4(n18608), .ZN(
        P3_U2997) );
  AND4_X1 U21625 ( .A1(n18752), .A2(n18612), .A3(n18611), .A4(n18702), .ZN(
        P3_U2998) );
  AND2_X1 U21626 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18698), .ZN(
        P3_U2999) );
  AND2_X1 U21627 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18698), .ZN(
        P3_U3000) );
  AND2_X1 U21628 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18698), .ZN(
        P3_U3001) );
  AND2_X1 U21629 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18698), .ZN(
        P3_U3002) );
  AND2_X1 U21630 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18698), .ZN(
        P3_U3003) );
  AND2_X1 U21631 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18698), .ZN(
        P3_U3004) );
  AND2_X1 U21632 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18698), .ZN(
        P3_U3005) );
  AND2_X1 U21633 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18698), .ZN(
        P3_U3006) );
  AND2_X1 U21634 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18698), .ZN(
        P3_U3007) );
  AND2_X1 U21635 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18698), .ZN(
        P3_U3008) );
  AND2_X1 U21636 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18698), .ZN(
        P3_U3009) );
  AND2_X1 U21637 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18698), .ZN(
        P3_U3010) );
  AND2_X1 U21638 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18698), .ZN(
        P3_U3011) );
  AND2_X1 U21639 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18698), .ZN(
        P3_U3012) );
  AND2_X1 U21640 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18698), .ZN(
        P3_U3013) );
  AND2_X1 U21641 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18698), .ZN(
        P3_U3014) );
  AND2_X1 U21642 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18698), .ZN(
        P3_U3015) );
  AND2_X1 U21643 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18698), .ZN(
        P3_U3016) );
  AND2_X1 U21644 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18698), .ZN(
        P3_U3017) );
  AND2_X1 U21645 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18698), .ZN(
        P3_U3018) );
  AND2_X1 U21646 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18698), .ZN(
        P3_U3019) );
  AND2_X1 U21647 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18698), .ZN(
        P3_U3020) );
  AND2_X1 U21648 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18698), .ZN(P3_U3021) );
  AND2_X1 U21649 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18698), .ZN(P3_U3022) );
  AND2_X1 U21650 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18698), .ZN(P3_U3023) );
  AND2_X1 U21651 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18698), .ZN(P3_U3024) );
  AND2_X1 U21652 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18698), .ZN(P3_U3025) );
  AND2_X1 U21653 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18698), .ZN(P3_U3026) );
  AND2_X1 U21654 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18698), .ZN(P3_U3027) );
  AND2_X1 U21655 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18698), .ZN(P3_U3028) );
  OAI21_X1 U21656 ( .B1(n18613), .B2(n20692), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18614) );
  AOI22_X1 U21657 ( .A1(n18626), .A2(n18629), .B1(n18763), .B2(n18614), .ZN(
        n18615) );
  INV_X1 U21658 ( .A(NA), .ZN(n20696) );
  OR3_X1 U21659 ( .A1(n20696), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18621) );
  OAI211_X1 U21660 ( .C1(n18616), .C2(n18759), .A(n18615), .B(n18621), .ZN(
        P3_U3029) );
  AOI21_X1 U21661 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18617) );
  AOI21_X1 U21662 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18617), .ZN(
        n18618) );
  AOI22_X1 U21663 ( .A1(n18750), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18618), .ZN(n18620) );
  NAND2_X1 U21664 ( .A1(n18620), .A2(n18619), .ZN(P3_U3030) );
  AOI22_X1 U21665 ( .A1(n18750), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18626), 
        .B2(n18621), .ZN(n18627) );
  NOR2_X1 U21666 ( .A1(n18629), .A2(n20692), .ZN(n18624) );
  NAND2_X1 U21667 ( .A1(n18750), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18622) );
  OAI22_X1 U21668 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18622), .ZN(n18623) );
  OAI22_X1 U21669 ( .A1(n18624), .A2(n18623), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18625) );
  OAI22_X1 U21670 ( .A1(n18627), .A2(n18629), .B1(n18626), .B2(n18625), .ZN(
        P3_U3031) );
  OAI222_X1 U21671 ( .A1(n18735), .A2(n18685), .B1(n18630), .B2(n18745), .C1(
        n18631), .C2(n18689), .ZN(P3_U3032) );
  OAI222_X1 U21672 ( .A1(n18689), .A2(n18633), .B1(n18632), .B2(n18745), .C1(
        n18631), .C2(n18685), .ZN(P3_U3033) );
  OAI222_X1 U21673 ( .A1(n18689), .A2(n18635), .B1(n18634), .B2(n18745), .C1(
        n18633), .C2(n18685), .ZN(P3_U3034) );
  INV_X1 U21674 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18638) );
  OAI222_X1 U21675 ( .A1(n18689), .A2(n18638), .B1(n18636), .B2(n18745), .C1(
        n18635), .C2(n18685), .ZN(P3_U3035) );
  OAI222_X1 U21676 ( .A1(n18638), .A2(n18685), .B1(n18637), .B2(n18745), .C1(
        n18639), .C2(n18689), .ZN(P3_U3036) );
  OAI222_X1 U21677 ( .A1(n18689), .A2(n18641), .B1(n18640), .B2(n18745), .C1(
        n18639), .C2(n18685), .ZN(P3_U3037) );
  INV_X1 U21678 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18643) );
  OAI222_X1 U21679 ( .A1(n18689), .A2(n18643), .B1(n18642), .B2(n18745), .C1(
        n18641), .C2(n18685), .ZN(P3_U3038) );
  OAI222_X1 U21680 ( .A1(n18689), .A2(n18645), .B1(n18644), .B2(n18745), .C1(
        n18643), .C2(n18685), .ZN(P3_U3039) );
  OAI222_X1 U21681 ( .A1(n18689), .A2(n18647), .B1(n18646), .B2(n18745), .C1(
        n18645), .C2(n18685), .ZN(P3_U3040) );
  OAI222_X1 U21682 ( .A1(n18689), .A2(n18649), .B1(n18648), .B2(n18745), .C1(
        n18647), .C2(n18685), .ZN(P3_U3041) );
  OAI222_X1 U21683 ( .A1(n18689), .A2(n18651), .B1(n18650), .B2(n18745), .C1(
        n18649), .C2(n18685), .ZN(P3_U3042) );
  OAI222_X1 U21684 ( .A1(n18689), .A2(n18653), .B1(n18652), .B2(n18745), .C1(
        n18651), .C2(n18685), .ZN(P3_U3043) );
  OAI222_X1 U21685 ( .A1(n18689), .A2(n18656), .B1(n18654), .B2(n18745), .C1(
        n18653), .C2(n18685), .ZN(P3_U3044) );
  OAI222_X1 U21686 ( .A1(n18656), .A2(n18685), .B1(n18655), .B2(n18745), .C1(
        n18657), .C2(n18689), .ZN(P3_U3045) );
  OAI222_X1 U21687 ( .A1(n18689), .A2(n18659), .B1(n18658), .B2(n18745), .C1(
        n18657), .C2(n18685), .ZN(P3_U3046) );
  INV_X1 U21688 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18662) );
  OAI222_X1 U21689 ( .A1(n18689), .A2(n18662), .B1(n18660), .B2(n18745), .C1(
        n18659), .C2(n18685), .ZN(P3_U3047) );
  OAI222_X1 U21690 ( .A1(n18662), .A2(n18685), .B1(n18661), .B2(n18745), .C1(
        n18663), .C2(n18689), .ZN(P3_U3048) );
  OAI222_X1 U21691 ( .A1(n18689), .A2(n20812), .B1(n18664), .B2(n18745), .C1(
        n18663), .C2(n18685), .ZN(P3_U3049) );
  OAI222_X1 U21692 ( .A1(n18689), .A2(n18666), .B1(n18665), .B2(n18745), .C1(
        n20812), .C2(n18685), .ZN(P3_U3050) );
  OAI222_X1 U21693 ( .A1(n18689), .A2(n20839), .B1(n18667), .B2(n18745), .C1(
        n18666), .C2(n18685), .ZN(P3_U3051) );
  OAI222_X1 U21694 ( .A1(n20839), .A2(n18685), .B1(n18668), .B2(n18745), .C1(
        n18669), .C2(n18689), .ZN(P3_U3052) );
  OAI222_X1 U21695 ( .A1(n18689), .A2(n18671), .B1(n18670), .B2(n18745), .C1(
        n18669), .C2(n18685), .ZN(P3_U3053) );
  OAI222_X1 U21696 ( .A1(n18689), .A2(n18673), .B1(n18672), .B2(n18745), .C1(
        n18671), .C2(n18685), .ZN(P3_U3054) );
  OAI222_X1 U21697 ( .A1(n18689), .A2(n18675), .B1(n18674), .B2(n18745), .C1(
        n18673), .C2(n18685), .ZN(P3_U3055) );
  OAI222_X1 U21698 ( .A1(n18689), .A2(n18677), .B1(n18676), .B2(n18745), .C1(
        n18675), .C2(n18685), .ZN(P3_U3056) );
  OAI222_X1 U21699 ( .A1(n18689), .A2(n18679), .B1(n18678), .B2(n18745), .C1(
        n18677), .C2(n18685), .ZN(P3_U3057) );
  INV_X1 U21700 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18682) );
  OAI222_X1 U21701 ( .A1(n18689), .A2(n18682), .B1(n18680), .B2(n18745), .C1(
        n18679), .C2(n18685), .ZN(P3_U3058) );
  OAI222_X1 U21702 ( .A1(n18682), .A2(n18685), .B1(n18681), .B2(n18745), .C1(
        n18683), .C2(n18689), .ZN(P3_U3059) );
  OAI222_X1 U21703 ( .A1(n18689), .A2(n18686), .B1(n18684), .B2(n18745), .C1(
        n18683), .C2(n18685), .ZN(P3_U3060) );
  OAI222_X1 U21704 ( .A1(n18689), .A2(n18688), .B1(n18687), .B2(n18745), .C1(
        n18686), .C2(n18685), .ZN(P3_U3061) );
  INV_X1 U21705 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18690) );
  AOI22_X1 U21706 ( .A1(n18745), .A2(n18691), .B1(n18690), .B2(n18763), .ZN(
        P3_U3274) );
  INV_X1 U21707 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18737) );
  INV_X1 U21708 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18692) );
  AOI22_X1 U21709 ( .A1(n18745), .A2(n18737), .B1(n18692), .B2(n18763), .ZN(
        P3_U3275) );
  INV_X1 U21710 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18693) );
  AOI22_X1 U21711 ( .A1(n18745), .A2(n18694), .B1(n18693), .B2(n18763), .ZN(
        P3_U3276) );
  INV_X1 U21712 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18743) );
  INV_X1 U21713 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18695) );
  AOI22_X1 U21714 ( .A1(n18745), .A2(n18743), .B1(n18695), .B2(n18763), .ZN(
        P3_U3277) );
  INV_X1 U21715 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18697) );
  INV_X1 U21716 ( .A(n18699), .ZN(n18696) );
  AOI21_X1 U21717 ( .B1(n18698), .B2(n18697), .A(n18696), .ZN(P3_U3280) );
  OAI21_X1 U21718 ( .B1(n18701), .B2(n18700), .A(n18699), .ZN(P3_U3281) );
  OAI221_X1 U21719 ( .B1(n18704), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18704), 
        .C2(n18703), .A(n18702), .ZN(P3_U3282) );
  NOR3_X1 U21720 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18705), .A3(
        n18708), .ZN(n18706) );
  AOI21_X1 U21721 ( .B1(n18728), .B2(n18707), .A(n18706), .ZN(n18713) );
  INV_X1 U21722 ( .A(n18708), .ZN(n18766) );
  INV_X1 U21723 ( .A(n18709), .ZN(n18710) );
  AOI21_X1 U21724 ( .B1(n18766), .B2(n18710), .A(n18734), .ZN(n18712) );
  OAI22_X1 U21725 ( .A1(n18734), .A2(n18713), .B1(n18712), .B2(n18711), .ZN(
        P3_U3285) );
  NOR2_X1 U21726 ( .A1(n18714), .A2(n18730), .ZN(n18722) );
  AOI22_X1 U21727 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n18715), .B2(n10690), .ZN(
        n18721) );
  INV_X1 U21728 ( .A(n18716), .ZN(n18717) );
  AOI222_X1 U21729 ( .A1(n18718), .A2(n18766), .B1(n18722), .B2(n18721), .C1(
        n18728), .C2(n18717), .ZN(n18719) );
  AOI22_X1 U21730 ( .A1(n18734), .A2(n10651), .B1(n18719), .B2(n18731), .ZN(
        P3_U3288) );
  INV_X1 U21731 ( .A(n18720), .ZN(n18725) );
  INV_X1 U21732 ( .A(n18721), .ZN(n18723) );
  AOI222_X1 U21733 ( .A1(n18725), .A2(n18766), .B1(n18728), .B2(n18724), .C1(
        n18723), .C2(n18722), .ZN(n18726) );
  AOI22_X1 U21734 ( .A1(n18734), .A2(n18727), .B1(n18726), .B2(n18731), .ZN(
        P3_U3289) );
  AOI222_X1 U21735 ( .A1(n18730), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18766), 
        .B2(n18729), .C1(n18733), .C2(n18728), .ZN(n18732) );
  AOI22_X1 U21736 ( .A1(n18734), .A2(n18733), .B1(n18732), .B2(n18731), .ZN(
        P3_U3290) );
  AOI21_X1 U21737 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18736) );
  AOI22_X1 U21738 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18736), .B2(n18735), .ZN(n18738) );
  AOI22_X1 U21739 ( .A1(n18739), .A2(n18738), .B1(n18737), .B2(n18742), .ZN(
        P3_U3292) );
  NOR2_X1 U21740 ( .A1(n18742), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18740) );
  AOI22_X1 U21741 ( .A1(n18743), .A2(n18742), .B1(n18741), .B2(n18740), .ZN(
        P3_U3293) );
  INV_X1 U21742 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18744) );
  AOI22_X1 U21743 ( .A1(n18745), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18744), 
        .B2(n18763), .ZN(P3_U3294) );
  MUX2_X1 U21744 ( .A(P3_MORE_REG_SCAN_IN), .B(n18747), .S(n18746), .Z(
        P3_U3295) );
  OAI21_X1 U21745 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18749), .A(n18748), 
        .ZN(n18751) );
  AOI211_X1 U21746 ( .C1(n18767), .C2(n18751), .A(n18750), .B(n18765), .ZN(
        n18754) );
  OAI21_X1 U21747 ( .B1(n18754), .B2(n18753), .A(n18752), .ZN(n18762) );
  OAI21_X1 U21748 ( .B1(n18757), .B2(n18756), .A(n18755), .ZN(n18758) );
  AOI21_X1 U21749 ( .B1(n18760), .B2(n18759), .A(n18758), .ZN(n18761) );
  MUX2_X1 U21750 ( .A(n18762), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18761), 
        .Z(P3_U3296) );
  INV_X1 U21751 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18771) );
  INV_X1 U21752 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18764) );
  AOI22_X1 U21753 ( .A1(n18745), .A2(n18771), .B1(n18764), .B2(n18763), .ZN(
        P3_U3297) );
  AOI21_X1 U21754 ( .B1(n18766), .B2(n18765), .A(n18768), .ZN(n18772) );
  INV_X1 U21755 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18769) );
  AOI22_X1 U21756 ( .A1(n18772), .A2(n18769), .B1(n18768), .B2(n18767), .ZN(
        P3_U3298) );
  AOI21_X1 U21757 ( .B1(n18772), .B2(n18771), .A(n18770), .ZN(P3_U3299) );
  INV_X1 U21758 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18773) );
  INV_X1 U21759 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19658) );
  NAND2_X1 U21760 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19658), .ZN(n19649) );
  AOI22_X1 U21761 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19649), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19642), .ZN(n20961) );
  INV_X1 U21762 ( .A(n20961), .ZN(n19641) );
  OAI21_X1 U21763 ( .B1(n19642), .B2(n18773), .A(n19641), .ZN(P2_U2815) );
  INV_X1 U21764 ( .A(n19786), .ZN(n18775) );
  AOI22_X1 U21765 ( .A1(n18775), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_0__SCAN_IN), .B2(n18774), .ZN(n18776) );
  INV_X1 U21766 ( .A(n18776), .ZN(P2_U2816) );
  AOI21_X1 U21767 ( .B1(n19642), .B2(n19658), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18777) );
  AOI22_X1 U21768 ( .A1(n19792), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18777), 
        .B2(n19793), .ZN(P2_U2817) );
  NOR4_X1 U21769 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18781) );
  NOR4_X1 U21770 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18780) );
  NOR4_X1 U21771 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18779) );
  NOR4_X1 U21772 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18778) );
  NAND4_X1 U21773 ( .A1(n18781), .A2(n18780), .A3(n18779), .A4(n18778), .ZN(
        n18787) );
  NOR4_X1 U21774 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18785) );
  AOI211_X1 U21775 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_27__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18784) );
  NOR4_X1 U21776 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18783) );
  NOR4_X1 U21777 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18782) );
  NAND4_X1 U21778 ( .A1(n18785), .A2(n18784), .A3(n18783), .A4(n18782), .ZN(
        n18786) );
  NOR2_X1 U21779 ( .A1(n18787), .A2(n18786), .ZN(n18795) );
  INV_X1 U21780 ( .A(n18795), .ZN(n18794) );
  NOR2_X1 U21781 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18794), .ZN(n18788) );
  INV_X1 U21782 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19708) );
  AOI22_X1 U21783 ( .A1(n18788), .A2(n18789), .B1(n18794), .B2(n19708), .ZN(
        P2_U2820) );
  OR3_X1 U21784 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18793) );
  INV_X1 U21785 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19706) );
  AOI22_X1 U21786 ( .A1(n18788), .A2(n18793), .B1(n18794), .B2(n19706), .ZN(
        P2_U2821) );
  INV_X1 U21787 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19711) );
  NAND2_X1 U21788 ( .A1(n18788), .A2(n19711), .ZN(n18792) );
  OAI21_X1 U21789 ( .B1(n19659), .B2(n18789), .A(n18795), .ZN(n18790) );
  OAI21_X1 U21790 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18795), .A(n18790), 
        .ZN(n18791) );
  OAI221_X1 U21791 ( .B1(n18792), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18792), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18791), .ZN(P2_U2822) );
  INV_X1 U21792 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19704) );
  OAI221_X1 U21793 ( .B1(n18795), .B2(n19704), .C1(n18794), .C2(n18793), .A(
        n18792), .ZN(P2_U2823) );
  NAND2_X1 U21794 ( .A1(n14070), .A2(n18796), .ZN(n18797) );
  XOR2_X1 U21795 ( .A(n18798), .B(n18797), .Z(n18806) );
  AOI22_X1 U21796 ( .A1(n18799), .A2(n13079), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n18927), .ZN(n18800) );
  OAI211_X1 U21797 ( .C1(n20940), .C2(n18921), .A(n18800), .B(n18920), .ZN(
        n18801) );
  AOI21_X1 U21798 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18912), .A(
        n18801), .ZN(n18805) );
  AOI22_X1 U21799 ( .A1(n18932), .A2(n18803), .B1(n18958), .B2(n18802), .ZN(
        n18804) );
  OAI211_X1 U21800 ( .C1(n19638), .C2(n18806), .A(n18805), .B(n18804), .ZN(
        P2_U2836) );
  NOR2_X1 U21801 ( .A1(n18939), .A2(n18807), .ZN(n18808) );
  XOR2_X1 U21802 ( .A(n18809), .B(n18808), .Z(n18817) );
  AOI22_X1 U21803 ( .A1(n18810), .A2(n13079), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n18927), .ZN(n18811) );
  OAI211_X1 U21804 ( .C1(n12964), .C2(n18921), .A(n18811), .B(n18920), .ZN(
        n18815) );
  OAI22_X1 U21805 ( .A1(n18954), .A2(n18813), .B1(n18812), .B2(n18937), .ZN(
        n18814) );
  AOI211_X1 U21806 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18912), .A(
        n18815), .B(n18814), .ZN(n18816) );
  OAI21_X1 U21807 ( .B1(n19638), .B2(n18817), .A(n18816), .ZN(P2_U2837) );
  OAI21_X1 U21808 ( .B1(n19680), .B2(n18921), .A(n18920), .ZN(n18821) );
  OAI22_X1 U21809 ( .A1(n18819), .A2(n18924), .B1(n18818), .B2(n18952), .ZN(
        n18820) );
  AOI211_X1 U21810 ( .C1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n18947), .A(
        n18821), .B(n18820), .ZN(n18828) );
  NAND2_X1 U21811 ( .A1(n14070), .A2(n18822), .ZN(n18823) );
  XOR2_X1 U21812 ( .A(n18824), .B(n18823), .Z(n18826) );
  AOI22_X1 U21813 ( .A1(n18826), .A2(n18933), .B1(n18932), .B2(n18825), .ZN(
        n18827) );
  OAI211_X1 U21814 ( .C1(n18829), .C2(n18937), .A(n18828), .B(n18827), .ZN(
        P2_U2838) );
  OAI21_X1 U21815 ( .B1(n12959), .B2(n18921), .A(n18920), .ZN(n18833) );
  OAI22_X1 U21816 ( .A1(n18831), .A2(n18924), .B1(n18830), .B2(n18922), .ZN(
        n18832) );
  AOI211_X1 U21817 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n18927), .A(n18833), .B(
        n18832), .ZN(n18840) );
  NAND2_X1 U21818 ( .A1(n14070), .A2(n18834), .ZN(n18835) );
  XNOR2_X1 U21819 ( .A(n18836), .B(n18835), .ZN(n18838) );
  AOI22_X1 U21820 ( .A1(n18838), .A2(n18933), .B1(n18932), .B2(n18837), .ZN(
        n18839) );
  OAI211_X1 U21821 ( .C1(n18841), .C2(n18937), .A(n18840), .B(n18839), .ZN(
        P2_U2840) );
  NOR2_X1 U21822 ( .A1(n18939), .A2(n18842), .ZN(n18863) );
  XOR2_X1 U21823 ( .A(n18863), .B(n18843), .Z(n18853) );
  OAI21_X1 U21824 ( .B1(n12951), .B2(n18921), .A(n18920), .ZN(n18848) );
  INV_X1 U21825 ( .A(n18844), .ZN(n18846) );
  OAI22_X1 U21826 ( .A1(n18846), .A2(n18924), .B1(n18845), .B2(n18952), .ZN(
        n18847) );
  AOI211_X1 U21827 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n18947), .A(
        n18848), .B(n18847), .ZN(n18852) );
  AOI22_X1 U21828 ( .A1(n18850), .A2(n18932), .B1(n18958), .B2(n18849), .ZN(
        n18851) );
  OAI211_X1 U21829 ( .C1(n19638), .C2(n18853), .A(n18852), .B(n18851), .ZN(
        P2_U2841) );
  NOR2_X1 U21830 ( .A1(n18854), .A2(n18864), .ZN(n18861) );
  NOR2_X1 U21831 ( .A1(n18855), .A2(n18924), .ZN(n18860) );
  NOR2_X1 U21832 ( .A1(n18952), .A2(n12326), .ZN(n18859) );
  AOI22_X1 U21833 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n9691), .ZN(n18856) );
  OAI211_X1 U21834 ( .C1(n18954), .C2(n18857), .A(n18856), .B(n18920), .ZN(
        n18858) );
  NOR4_X1 U21835 ( .A1(n18861), .A2(n18860), .A3(n18859), .A4(n18858), .ZN(
        n18867) );
  INV_X1 U21836 ( .A(n18862), .ZN(n18865) );
  OAI211_X1 U21837 ( .C1(n18865), .C2(n18864), .A(n18933), .B(n18863), .ZN(
        n18866) );
  OAI211_X1 U21838 ( .C1(n18937), .C2(n18868), .A(n18867), .B(n18866), .ZN(
        P2_U2842) );
  NOR2_X1 U21839 ( .A1(n18939), .A2(n18879), .ZN(n18869) );
  XOR2_X1 U21840 ( .A(n18870), .B(n18869), .Z(n18878) );
  INV_X1 U21841 ( .A(n18871), .ZN(n18872) );
  AOI22_X1 U21842 ( .A1(n18872), .A2(n13079), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18947), .ZN(n18873) );
  OAI211_X1 U21843 ( .C1(n12945), .C2(n18921), .A(n18873), .B(n18920), .ZN(
        n18876) );
  OAI22_X1 U21844 ( .A1(n18954), .A2(n18874), .B1(n18937), .B2(n18972), .ZN(
        n18875) );
  AOI211_X1 U21845 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n18927), .A(n18876), .B(
        n18875), .ZN(n18877) );
  OAI21_X1 U21846 ( .B1(n19638), .B2(n18878), .A(n18877), .ZN(P2_U2843) );
  AOI21_X1 U21847 ( .B1(n18890), .B2(n18880), .A(n18879), .ZN(n18887) );
  AOI22_X1 U21848 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18947), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n9691), .ZN(n18881) );
  OAI211_X1 U21849 ( .C1(n18882), .C2(n18937), .A(n18881), .B(n18920), .ZN(
        n18886) );
  OAI22_X1 U21850 ( .A1(n18884), .A2(n18924), .B1(n18952), .B2(n18883), .ZN(
        n18885) );
  AOI211_X1 U21851 ( .C1(n18888), .C2(n18887), .A(n18886), .B(n18885), .ZN(
        n18893) );
  AOI22_X1 U21852 ( .A1(n18891), .A2(n18890), .B1(n18932), .B2(n18889), .ZN(
        n18892) );
  NAND2_X1 U21853 ( .A1(n18893), .A2(n18892), .ZN(P2_U2844) );
  OAI21_X1 U21854 ( .B1(n12936), .B2(n18921), .A(n18920), .ZN(n18897) );
  OAI22_X1 U21855 ( .A1(n18895), .A2(n18924), .B1(n18894), .B2(n18922), .ZN(
        n18896) );
  AOI211_X1 U21856 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n18927), .A(n18897), .B(
        n18896), .ZN(n18904) );
  NAND2_X1 U21857 ( .A1(n14070), .A2(n18898), .ZN(n18899) );
  XNOR2_X1 U21858 ( .A(n18900), .B(n18899), .ZN(n18902) );
  AOI22_X1 U21859 ( .A1(n18902), .A2(n18933), .B1(n18932), .B2(n18901), .ZN(
        n18903) );
  OAI211_X1 U21860 ( .C1(n18905), .C2(n18937), .A(n18904), .B(n18903), .ZN(
        P2_U2846) );
  NAND2_X1 U21861 ( .A1(n14070), .A2(n18906), .ZN(n18907) );
  XOR2_X1 U21862 ( .A(n18908), .B(n18907), .Z(n18919) );
  AOI22_X1 U21863 ( .A1(n18909), .A2(n13079), .B1(n18927), .B2(
        P2_EBX_REG_7__SCAN_IN), .ZN(n18910) );
  OAI211_X1 U21864 ( .C1(n19668), .C2(n18921), .A(n18910), .B(n18920), .ZN(
        n18911) );
  AOI21_X1 U21865 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18912), .A(
        n18911), .ZN(n18918) );
  INV_X1 U21866 ( .A(n18913), .ZN(n18916) );
  INV_X1 U21867 ( .A(n18914), .ZN(n18915) );
  AOI22_X1 U21868 ( .A1(n18932), .A2(n18916), .B1(n18958), .B2(n18915), .ZN(
        n18917) );
  OAI211_X1 U21869 ( .C1(n19638), .C2(n18919), .A(n18918), .B(n18917), .ZN(
        P2_U2848) );
  OAI21_X1 U21870 ( .B1(n12919), .B2(n18921), .A(n18920), .ZN(n18926) );
  OAI22_X1 U21871 ( .A1(n18924), .A2(n18923), .B1(n20875), .B2(n18922), .ZN(
        n18925) );
  AOI211_X1 U21872 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n18927), .A(n18926), .B(
        n18925), .ZN(n18936) );
  NAND2_X1 U21873 ( .A1(n14070), .A2(n18928), .ZN(n18929) );
  XNOR2_X1 U21874 ( .A(n18930), .B(n18929), .ZN(n18934) );
  AOI22_X1 U21875 ( .A1(n18934), .A2(n18933), .B1(n18932), .B2(n18931), .ZN(
        n18935) );
  OAI211_X1 U21876 ( .C1(n18937), .C2(n18981), .A(n18936), .B(n18935), .ZN(
        P2_U2850) );
  NOR2_X1 U21877 ( .A1(n18939), .A2(n18938), .ZN(n18940) );
  XOR2_X1 U21878 ( .A(n19051), .B(n18940), .Z(n18960) );
  NAND2_X1 U21879 ( .A1(n18942), .A2(n18941), .ZN(n18945) );
  INV_X1 U21880 ( .A(n18943), .ZN(n18944) );
  AND2_X1 U21881 ( .A1(n18945), .A2(n18944), .ZN(n19056) );
  INV_X1 U21882 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18951) );
  AOI21_X1 U21883 ( .B1(P2_REIP_REG_4__SCAN_IN), .B2(n9691), .A(n19040), .ZN(
        n18950) );
  AOI22_X1 U21884 ( .A1(n13079), .A2(n18948), .B1(n18947), .B2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18949) );
  OAI211_X1 U21885 ( .C1(n18952), .C2(n18951), .A(n18950), .B(n18949), .ZN(
        n18957) );
  OAI22_X1 U21886 ( .A1(n18984), .A2(n18955), .B1(n18954), .B2(n18953), .ZN(
        n18956) );
  AOI211_X1 U21887 ( .C1(n18958), .C2(n19056), .A(n18957), .B(n18956), .ZN(
        n18959) );
  OAI21_X1 U21888 ( .B1(n19638), .B2(n18960), .A(n18959), .ZN(P2_U2851) );
  AOI22_X1 U21889 ( .A1(n18962), .A2(BUF1_REG_31__SCAN_IN), .B1(n18996), .B2(
        n18961), .ZN(n18965) );
  AOI22_X1 U21890 ( .A1(n18963), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18995), .ZN(n18964) );
  NAND2_X1 U21891 ( .A1(n18965), .A2(n18964), .ZN(P2_U2888) );
  INV_X1 U21892 ( .A(n19002), .ZN(n18970) );
  AOI22_X1 U21893 ( .A1(n18970), .A2(n18966), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n18995), .ZN(n18967) );
  OAI21_X1 U21894 ( .B1(n18982), .B2(n18968), .A(n18967), .ZN(P2_U2905) );
  AOI22_X1 U21895 ( .A1(n18970), .A2(n18969), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n18995), .ZN(n18971) );
  OAI21_X1 U21896 ( .B1(n18982), .B2(n18972), .A(n18971), .ZN(P2_U2907) );
  INV_X1 U21897 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19026) );
  OAI22_X1 U21898 ( .A1(n19002), .A2(n19106), .B1(n18973), .B2(n19026), .ZN(
        n18974) );
  INV_X1 U21899 ( .A(n18974), .ZN(n18980) );
  NAND2_X1 U21900 ( .A1(n19730), .A2(n19728), .ZN(n18977) );
  XOR2_X1 U21901 ( .A(n19728), .B(n19730), .Z(n18990) );
  NAND2_X1 U21902 ( .A1(n19738), .A2(n19736), .ZN(n18976) );
  NAND2_X1 U21903 ( .A1(n18976), .A2(n18975), .ZN(n18989) );
  NAND2_X1 U21904 ( .A1(n18990), .A2(n18989), .ZN(n18988) );
  AOI21_X1 U21905 ( .B1(n18977), .B2(n18988), .A(n19056), .ZN(n18983) );
  OR3_X1 U21906 ( .A1(n18983), .A2(n18984), .A3(n18978), .ZN(n18979) );
  OAI211_X1 U21907 ( .C1(n18982), .C2(n18981), .A(n18980), .B(n18979), .ZN(
        P2_U2914) );
  AOI22_X1 U21908 ( .A1(n18996), .A2(n19056), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n18995), .ZN(n18987) );
  XOR2_X1 U21909 ( .A(n18984), .B(n18983), .Z(n18985) );
  NAND2_X1 U21910 ( .A1(n18985), .A2(n18998), .ZN(n18986) );
  OAI211_X1 U21911 ( .C1(n19103), .C2(n19002), .A(n18987), .B(n18986), .ZN(
        P2_U2915) );
  OAI21_X1 U21912 ( .B1(n18990), .B2(n18989), .A(n18988), .ZN(n18991) );
  NAND2_X1 U21913 ( .A1(n18991), .A2(n18998), .ZN(n18994) );
  INV_X1 U21914 ( .A(n19728), .ZN(n18992) );
  AOI22_X1 U21915 ( .A1(n18992), .A2(n18996), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n18995), .ZN(n18993) );
  OAI211_X1 U21916 ( .C1(n19098), .C2(n19002), .A(n18994), .B(n18993), .ZN(
        P2_U2916) );
  AOI22_X1 U21917 ( .A1(n18996), .A2(n18999), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n18995), .ZN(n19001) );
  OAI211_X1 U21918 ( .C1(n19507), .C2(n18999), .A(n18998), .B(n18997), .ZN(
        n19000) );
  OAI211_X1 U21919 ( .C1(n19081), .C2(n19002), .A(n19001), .B(n19000), .ZN(
        P2_U2919) );
  AND2_X1 U21920 ( .A1(n19027), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  INV_X1 U21921 ( .A(n19003), .ZN(n19039) );
  AOI22_X1 U21922 ( .A1(n19037), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19004) );
  OAI21_X1 U21923 ( .B1(n19005), .B2(n19039), .A(n19004), .ZN(P2_U2936) );
  AOI22_X1 U21924 ( .A1(n19037), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19006) );
  OAI21_X1 U21925 ( .B1(n19007), .B2(n19039), .A(n19006), .ZN(P2_U2937) );
  AOI22_X1 U21926 ( .A1(n19037), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19008) );
  OAI21_X1 U21927 ( .B1(n19009), .B2(n19039), .A(n19008), .ZN(P2_U2938) );
  AOI22_X1 U21928 ( .A1(n19037), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19010) );
  OAI21_X1 U21929 ( .B1(n19011), .B2(n19039), .A(n19010), .ZN(P2_U2939) );
  AOI22_X1 U21930 ( .A1(n19018), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19012) );
  OAI21_X1 U21931 ( .B1(n19013), .B2(n19039), .A(n19012), .ZN(P2_U2940) );
  AOI22_X1 U21932 ( .A1(n19018), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19014) );
  OAI21_X1 U21933 ( .B1(n19015), .B2(n19039), .A(n19014), .ZN(P2_U2941) );
  AOI22_X1 U21934 ( .A1(n19018), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19016) );
  OAI21_X1 U21935 ( .B1(n19017), .B2(n19039), .A(n19016), .ZN(P2_U2942) );
  AOI22_X1 U21936 ( .A1(n19018), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19019) );
  OAI21_X1 U21937 ( .B1(n19020), .B2(n19039), .A(n19019), .ZN(P2_U2943) );
  AOI22_X1 U21938 ( .A1(n19037), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19021) );
  OAI21_X1 U21939 ( .B1(n19022), .B2(n19039), .A(n19021), .ZN(P2_U2944) );
  AOI22_X1 U21940 ( .A1(n19037), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19023) );
  OAI21_X1 U21941 ( .B1(n19024), .B2(n19039), .A(n19023), .ZN(P2_U2945) );
  AOI22_X1 U21942 ( .A1(n19037), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19025) );
  OAI21_X1 U21943 ( .B1(n19026), .B2(n19039), .A(n19025), .ZN(P2_U2946) );
  INV_X1 U21944 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19029) );
  AOI22_X1 U21945 ( .A1(n19037), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19027), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19028) );
  OAI21_X1 U21946 ( .B1(n19029), .B2(n19039), .A(n19028), .ZN(P2_U2947) );
  INV_X1 U21947 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19031) );
  AOI22_X1 U21948 ( .A1(n19037), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19030) );
  OAI21_X1 U21949 ( .B1(n19031), .B2(n19039), .A(n19030), .ZN(P2_U2948) );
  AOI22_X1 U21950 ( .A1(n19037), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19032) );
  OAI21_X1 U21951 ( .B1(n19033), .B2(n19039), .A(n19032), .ZN(P2_U2949) );
  INV_X1 U21952 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19035) );
  AOI22_X1 U21953 ( .A1(n19037), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19034) );
  OAI21_X1 U21954 ( .B1(n19035), .B2(n19039), .A(n19034), .ZN(P2_U2950) );
  AOI22_X1 U21955 ( .A1(n19037), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19036), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19038) );
  OAI21_X1 U21956 ( .B1(n12885), .B2(n19039), .A(n19038), .ZN(P2_U2951) );
  AOI22_X1 U21957 ( .A1(n19041), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19040), .ZN(n19050) );
  OAI21_X1 U21958 ( .B1(n19043), .B2(n19059), .A(n19042), .ZN(n19062) );
  XOR2_X1 U21959 ( .A(n9608), .B(n19045), .Z(n19065) );
  AOI222_X1 U21960 ( .A1(n19062), .A2(n19048), .B1(n19047), .B2(n19054), .C1(
        n19046), .C2(n19065), .ZN(n19049) );
  OAI211_X1 U21961 ( .C1(n19052), .C2(n19051), .A(n19050), .B(n19049), .ZN(
        P2_U3010) );
  AOI22_X1 U21962 ( .A1(n19055), .A2(n19059), .B1(n19054), .B2(n19053), .ZN(
        n19069) );
  INV_X1 U21963 ( .A(n19056), .ZN(n19057) );
  OAI22_X1 U21964 ( .A1(n19060), .A2(n19059), .B1(n19058), .B2(n19057), .ZN(
        n19061) );
  INV_X1 U21965 ( .A(n19061), .ZN(n19068) );
  AOI22_X1 U21966 ( .A1(n19065), .A2(n19064), .B1(n19063), .B2(n19062), .ZN(
        n19067) );
  NAND2_X1 U21967 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19040), .ZN(n19066) );
  NAND4_X1 U21968 ( .A1(n19069), .A2(n19068), .A3(n19067), .A4(n19066), .ZN(
        P2_U3042) );
  OR2_X1 U21969 ( .A1(n19539), .A2(n19725), .ZN(n19747) );
  NOR3_X2 U21970 ( .A1(n19071), .A2(n19158), .A3(n19747), .ZN(n19113) );
  AOI22_X1 U21971 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19112), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19113), .ZN(n19473) );
  OAI22_X1 U21972 ( .A1(n19073), .A2(n19115), .B1(n19072), .B2(n19114), .ZN(
        n19470) );
  NAND2_X1 U21973 ( .A1(n19730), .A2(n19738), .ZN(n19153) );
  NAND2_X1 U21974 ( .A1(n19075), .A2(n19074), .ZN(n19117) );
  NOR2_X2 U21975 ( .A1(n19117), .A2(n19076), .ZN(n19573) );
  NAND2_X1 U21976 ( .A1(n19734), .A2(n19742), .ZN(n19187) );
  OR2_X1 U21977 ( .A1(n19187), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19128) );
  NOR2_X1 U21978 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19128), .ZN(
        n19118) );
  AOI22_X1 U21979 ( .A1(n19470), .A2(n19119), .B1(n19573), .B2(n19118), .ZN(
        n19088) );
  INV_X1 U21980 ( .A(n19569), .ZN(n19623) );
  NOR2_X1 U21981 ( .A1(n19086), .A2(n19623), .ZN(n19079) );
  AOI211_X1 U21982 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19082), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19079), .ZN(n19080) );
  NOR2_X2 U21983 ( .A1(n19081), .A2(n19158), .ZN(n19574) );
  NOR2_X1 U21984 ( .A1(n19623), .A2(n19118), .ZN(n19085) );
  INV_X1 U21985 ( .A(n19082), .ZN(n19083) );
  OAI21_X1 U21986 ( .B1(n19083), .B2(n19118), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19084) );
  AOI22_X1 U21987 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19122), .B1(
        n19574), .B2(n19121), .ZN(n19087) );
  OAI211_X1 U21988 ( .C1(n19473), .C2(n19631), .A(n19088), .B(n19087), .ZN(
        P2_U3048) );
  AOI22_X1 U21989 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19113), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19112), .ZN(n19477) );
  OAI22_X1 U21990 ( .A1(n15039), .A2(n19115), .B1(n15041), .B2(n19114), .ZN(
        n19474) );
  NOR2_X2 U21991 ( .A1(n19117), .A2(n13146), .ZN(n19586) );
  AOI22_X1 U21992 ( .A1(n19474), .A2(n19119), .B1(n19118), .B2(n19586), .ZN(
        n19091) );
  NOR2_X2 U21993 ( .A1(n19089), .A2(n19158), .ZN(n19587) );
  AOI22_X1 U21994 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19122), .B1(
        n19587), .B2(n19121), .ZN(n19090) );
  OAI211_X1 U21995 ( .C1(n19477), .C2(n19631), .A(n19091), .B(n19090), .ZN(
        P2_U3049) );
  AOI22_X1 U21996 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19112), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19113), .ZN(n19481) );
  OAI22_X1 U21997 ( .A1(n19093), .A2(n19115), .B1(n19092), .B2(n19114), .ZN(
        n19478) );
  NOR2_X2 U21998 ( .A1(n19117), .A2(n10061), .ZN(n19592) );
  AOI22_X1 U21999 ( .A1(n19478), .A2(n19119), .B1(n19118), .B2(n19592), .ZN(
        n19096) );
  NOR2_X2 U22000 ( .A1(n19094), .A2(n19158), .ZN(n19593) );
  AOI22_X1 U22001 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19122), .B1(
        n19593), .B2(n19121), .ZN(n19095) );
  OAI211_X1 U22002 ( .C1(n19481), .C2(n19631), .A(n19096), .B(n19095), .ZN(
        P2_U3050) );
  AOI22_X1 U22003 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19112), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19113), .ZN(n19485) );
  NOR2_X2 U22004 ( .A1(n19117), .A2(n10067), .ZN(n19598) );
  AOI22_X1 U22005 ( .A1(n19482), .A2(n19119), .B1(n19598), .B2(n19118), .ZN(
        n19100) );
  NOR2_X2 U22006 ( .A1(n19098), .A2(n19158), .ZN(n19599) );
  AOI22_X1 U22007 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19122), .B1(
        n19599), .B2(n19121), .ZN(n19099) );
  OAI211_X1 U22008 ( .C1(n19485), .C2(n19631), .A(n19100), .B(n19099), .ZN(
        P2_U3051) );
  AOI22_X1 U22009 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19112), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19113), .ZN(n19489) );
  NOR2_X2 U22010 ( .A1(n19117), .A2(n19102), .ZN(n19604) );
  AOI22_X1 U22011 ( .A1(n19486), .A2(n19119), .B1(n19118), .B2(n19604), .ZN(
        n19105) );
  NOR2_X2 U22012 ( .A1(n19103), .A2(n19158), .ZN(n19605) );
  AOI22_X1 U22013 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19122), .B1(
        n19605), .B2(n19121), .ZN(n19104) );
  OAI211_X1 U22014 ( .C1(n19489), .C2(n19631), .A(n19105), .B(n19104), .ZN(
        P2_U3052) );
  AOI22_X1 U22015 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19112), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19113), .ZN(n19493) );
  NOR2_X2 U22016 ( .A1(n19117), .A2(n9593), .ZN(n19610) );
  AOI22_X1 U22017 ( .A1(n19490), .A2(n19119), .B1(n19118), .B2(n19610), .ZN(
        n19108) );
  NOR2_X2 U22018 ( .A1(n19106), .A2(n19158), .ZN(n19611) );
  AOI22_X1 U22019 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19122), .B1(
        n19611), .B2(n19121), .ZN(n19107) );
  OAI211_X1 U22020 ( .C1(n19493), .C2(n19631), .A(n19108), .B(n19107), .ZN(
        P2_U3053) );
  AOI22_X1 U22021 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19113), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19112), .ZN(n19497) );
  OAI22_X1 U22022 ( .A1(n15007), .A2(n19115), .B1(n15008), .B2(n19114), .ZN(
        n19494) );
  NOR2_X2 U22023 ( .A1(n19117), .A2(n9996), .ZN(n19616) );
  AOI22_X1 U22024 ( .A1(n19494), .A2(n19119), .B1(n19118), .B2(n19616), .ZN(
        n19111) );
  NOR2_X2 U22025 ( .A1(n19109), .A2(n19158), .ZN(n19617) );
  AOI22_X1 U22026 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19122), .B1(
        n19617), .B2(n19121), .ZN(n19110) );
  OAI211_X1 U22027 ( .C1(n19497), .C2(n19631), .A(n19111), .B(n19110), .ZN(
        P2_U3054) );
  AOI22_X1 U22028 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19113), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19112), .ZN(n19505) );
  NOR2_X2 U22029 ( .A1(n19117), .A2(n19116), .ZN(n19622) );
  AOI22_X1 U22030 ( .A1(n19500), .A2(n19119), .B1(n19118), .B2(n19622), .ZN(
        n19124) );
  NOR2_X2 U22031 ( .A1(n19120), .A2(n19158), .ZN(n19624) );
  AOI22_X1 U22032 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19122), .B1(
        n19624), .B2(n19121), .ZN(n19123) );
  OAI211_X1 U22033 ( .C1(n19505), .C2(n19631), .A(n19124), .B(n19123), .ZN(
        P2_U3055) );
  NAND2_X1 U22034 ( .A1(n19751), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19367) );
  NOR2_X1 U22035 ( .A1(n19367), .A2(n19187), .ZN(n19147) );
  NOR2_X1 U22036 ( .A1(n19147), .A2(n19784), .ZN(n19125) );
  NAND2_X1 U22037 ( .A1(n19126), .A2(n19125), .ZN(n19129) );
  OAI21_X1 U22038 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19128), .A(n19784), 
        .ZN(n19127) );
  AOI22_X1 U22039 ( .A1(n19148), .A2(n19574), .B1(n19573), .B2(n19147), .ZN(
        n19134) );
  OAI21_X1 U22040 ( .B1(n19132), .B2(n19725), .A(n19128), .ZN(n19130) );
  AND2_X1 U22041 ( .A1(n19130), .A2(n19129), .ZN(n19131) );
  OAI211_X1 U22042 ( .C1(n19147), .C2(n20926), .A(n19576), .B(n19131), .ZN(
        n19149) );
  AOI22_X1 U22043 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19149), .B1(
        n19181), .B2(n19470), .ZN(n19133) );
  OAI211_X1 U22044 ( .C1(n19473), .C2(n19152), .A(n19134), .B(n19133), .ZN(
        P2_U3056) );
  AOI22_X1 U22045 ( .A1(n19148), .A2(n19587), .B1(n19586), .B2(n19147), .ZN(
        n19136) );
  AOI22_X1 U22046 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19149), .B1(
        n19181), .B2(n19474), .ZN(n19135) );
  OAI211_X1 U22047 ( .C1(n19477), .C2(n19152), .A(n19136), .B(n19135), .ZN(
        P2_U3057) );
  AOI22_X1 U22048 ( .A1(n19148), .A2(n19593), .B1(n19592), .B2(n19147), .ZN(
        n19138) );
  AOI22_X1 U22049 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19149), .B1(
        n19181), .B2(n19478), .ZN(n19137) );
  OAI211_X1 U22050 ( .C1(n19481), .C2(n19152), .A(n19138), .B(n19137), .ZN(
        P2_U3058) );
  AOI22_X1 U22051 ( .A1(n19148), .A2(n19599), .B1(n19598), .B2(n19147), .ZN(
        n19140) );
  AOI22_X1 U22052 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19149), .B1(
        n19181), .B2(n19482), .ZN(n19139) );
  OAI211_X1 U22053 ( .C1(n19485), .C2(n19152), .A(n19140), .B(n19139), .ZN(
        P2_U3059) );
  AOI22_X1 U22054 ( .A1(n19148), .A2(n19605), .B1(n19604), .B2(n19147), .ZN(
        n19142) );
  AOI22_X1 U22055 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19149), .B1(
        n19181), .B2(n19486), .ZN(n19141) );
  OAI211_X1 U22056 ( .C1(n19489), .C2(n19152), .A(n19142), .B(n19141), .ZN(
        P2_U3060) );
  AOI22_X1 U22057 ( .A1(n19148), .A2(n19611), .B1(n19610), .B2(n19147), .ZN(
        n19144) );
  AOI22_X1 U22058 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19149), .B1(
        n19181), .B2(n19490), .ZN(n19143) );
  OAI211_X1 U22059 ( .C1(n19493), .C2(n19152), .A(n19144), .B(n19143), .ZN(
        P2_U3061) );
  AOI22_X1 U22060 ( .A1(n19148), .A2(n19617), .B1(n19616), .B2(n19147), .ZN(
        n19146) );
  AOI22_X1 U22061 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19149), .B1(
        n19181), .B2(n19494), .ZN(n19145) );
  OAI211_X1 U22062 ( .C1(n19497), .C2(n19152), .A(n19146), .B(n19145), .ZN(
        P2_U3062) );
  AOI22_X1 U22063 ( .A1(n19148), .A2(n19624), .B1(n19622), .B2(n19147), .ZN(
        n19151) );
  AOI22_X1 U22064 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19149), .B1(
        n19181), .B2(n19500), .ZN(n19150) );
  OAI211_X1 U22065 ( .C1(n19505), .C2(n19152), .A(n19151), .B(n19150), .ZN(
        P2_U3063) );
  NAND2_X1 U22066 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19757), .ZN(
        n19398) );
  NOR2_X1 U22067 ( .A1(n19398), .A2(n19187), .ZN(n19179) );
  INV_X1 U22068 ( .A(n19179), .ZN(n19160) );
  INV_X1 U22069 ( .A(n12191), .ZN(n19161) );
  OAI21_X1 U22070 ( .B1(n19161), .B2(n19784), .A(n20926), .ZN(n19159) );
  NAND2_X1 U22071 ( .A1(n19216), .A2(n19154), .ZN(n19156) );
  NOR2_X1 U22072 ( .A1(n19401), .A2(n19187), .ZN(n19155) );
  AOI211_X1 U22073 ( .C1(n19156), .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19155), 
        .B(n19539), .ZN(n19157) );
  OAI21_X1 U22074 ( .B1(n19161), .B2(n19179), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19162) );
  OAI21_X1 U22075 ( .B1(n19187), .B2(n19401), .A(n19162), .ZN(n19180) );
  AOI22_X1 U22076 ( .A1(n19180), .A2(n19574), .B1(n19573), .B2(n19179), .ZN(
        n19164) );
  INV_X1 U22077 ( .A(n19473), .ZN(n19582) );
  AOI22_X1 U22078 ( .A1(n19202), .A2(n19470), .B1(n19181), .B2(n19582), .ZN(
        n19163) );
  OAI211_X1 U22079 ( .C1(n19185), .C2(n19165), .A(n19164), .B(n19163), .ZN(
        P2_U3064) );
  AOI22_X1 U22080 ( .A1(n19180), .A2(n19587), .B1(n19586), .B2(n19179), .ZN(
        n19167) );
  INV_X1 U22081 ( .A(n19477), .ZN(n19588) );
  AOI22_X1 U22082 ( .A1(n19202), .A2(n19474), .B1(n19181), .B2(n19588), .ZN(
        n19166) );
  OAI211_X1 U22083 ( .C1(n19185), .C2(n12036), .A(n19167), .B(n19166), .ZN(
        P2_U3065) );
  AOI22_X1 U22084 ( .A1(n19180), .A2(n19593), .B1(n19592), .B2(n19179), .ZN(
        n19169) );
  INV_X1 U22085 ( .A(n19481), .ZN(n19594) );
  AOI22_X1 U22086 ( .A1(n19202), .A2(n19478), .B1(n19181), .B2(n19594), .ZN(
        n19168) );
  OAI211_X1 U22087 ( .C1(n19185), .C2(n10353), .A(n19169), .B(n19168), .ZN(
        P2_U3066) );
  AOI22_X1 U22088 ( .A1(n19180), .A2(n19599), .B1(n19598), .B2(n19179), .ZN(
        n19171) );
  INV_X1 U22089 ( .A(n19485), .ZN(n19600) );
  AOI22_X1 U22090 ( .A1(n19202), .A2(n19482), .B1(n19181), .B2(n19600), .ZN(
        n19170) );
  OAI211_X1 U22091 ( .C1(n19185), .C2(n12000), .A(n19171), .B(n19170), .ZN(
        P2_U3067) );
  AOI22_X1 U22092 ( .A1(n19180), .A2(n19605), .B1(n19604), .B2(n19179), .ZN(
        n19173) );
  INV_X1 U22093 ( .A(n19489), .ZN(n19606) );
  AOI22_X1 U22094 ( .A1(n19202), .A2(n19486), .B1(n19181), .B2(n19606), .ZN(
        n19172) );
  OAI211_X1 U22095 ( .C1(n19185), .C2(n10324), .A(n19173), .B(n19172), .ZN(
        P2_U3068) );
  AOI22_X1 U22096 ( .A1(n19180), .A2(n19611), .B1(n19610), .B2(n19179), .ZN(
        n19175) );
  INV_X1 U22097 ( .A(n19493), .ZN(n19612) );
  AOI22_X1 U22098 ( .A1(n19202), .A2(n19490), .B1(n19181), .B2(n19612), .ZN(
        n19174) );
  OAI211_X1 U22099 ( .C1(n19185), .C2(n12192), .A(n19175), .B(n19174), .ZN(
        P2_U3069) );
  AOI22_X1 U22100 ( .A1(n19180), .A2(n19617), .B1(n19616), .B2(n19179), .ZN(
        n19177) );
  INV_X1 U22101 ( .A(n19497), .ZN(n19618) );
  AOI22_X1 U22102 ( .A1(n19202), .A2(n19494), .B1(n19181), .B2(n19618), .ZN(
        n19176) );
  OAI211_X1 U22103 ( .C1(n19185), .C2(n19178), .A(n19177), .B(n19176), .ZN(
        P2_U3070) );
  AOI22_X1 U22104 ( .A1(n19180), .A2(n19624), .B1(n19622), .B2(n19179), .ZN(
        n19183) );
  INV_X1 U22105 ( .A(n19505), .ZN(n19626) );
  AOI22_X1 U22106 ( .A1(n19202), .A2(n19500), .B1(n19181), .B2(n19626), .ZN(
        n19182) );
  OAI211_X1 U22107 ( .C1(n19185), .C2(n19184), .A(n19183), .B(n19182), .ZN(
        P2_U3071) );
  NOR2_X1 U22108 ( .A1(n19429), .A2(n19187), .ZN(n19211) );
  AOI22_X1 U22109 ( .A1(n19470), .A2(n19218), .B1(n19211), .B2(n19573), .ZN(
        n19197) );
  OAI21_X1 U22110 ( .B1(n19186), .B2(n19725), .A(n19724), .ZN(n19195) );
  NOR2_X1 U22111 ( .A1(n19751), .A2(n19187), .ZN(n19190) );
  INV_X1 U22112 ( .A(n19211), .ZN(n19188) );
  OAI211_X1 U22113 ( .C1(n19191), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19188), 
        .B(n19539), .ZN(n19189) );
  OAI211_X1 U22114 ( .C1(n19195), .C2(n19190), .A(n19576), .B(n19189), .ZN(
        n19213) );
  INV_X1 U22115 ( .A(n19190), .ZN(n19194) );
  INV_X1 U22116 ( .A(n19191), .ZN(n19192) );
  OAI21_X1 U22117 ( .B1(n19192), .B2(n19211), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19193) );
  OAI21_X1 U22118 ( .B1(n19195), .B2(n19194), .A(n19193), .ZN(n19212) );
  AOI22_X1 U22119 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19213), .B1(
        n19574), .B2(n19212), .ZN(n19196) );
  OAI211_X1 U22120 ( .C1(n19473), .C2(n19216), .A(n19197), .B(n19196), .ZN(
        P2_U3072) );
  INV_X1 U22121 ( .A(n19474), .ZN(n19591) );
  AOI22_X1 U22122 ( .A1(n19202), .A2(n19588), .B1(n19211), .B2(n19586), .ZN(
        n19199) );
  AOI22_X1 U22123 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19213), .B1(
        n19587), .B2(n19212), .ZN(n19198) );
  OAI211_X1 U22124 ( .C1(n19591), .C2(n19248), .A(n19199), .B(n19198), .ZN(
        P2_U3073) );
  INV_X1 U22125 ( .A(n19478), .ZN(n19597) );
  AOI22_X1 U22126 ( .A1(n19202), .A2(n19594), .B1(n19211), .B2(n19592), .ZN(
        n19201) );
  AOI22_X1 U22127 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19213), .B1(
        n19593), .B2(n19212), .ZN(n19200) );
  OAI211_X1 U22128 ( .C1(n19597), .C2(n19248), .A(n19201), .B(n19200), .ZN(
        P2_U3074) );
  INV_X1 U22129 ( .A(n19482), .ZN(n19603) );
  AOI22_X1 U22130 ( .A1(n19202), .A2(n19600), .B1(n19211), .B2(n19598), .ZN(
        n19204) );
  AOI22_X1 U22131 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19213), .B1(
        n19599), .B2(n19212), .ZN(n19203) );
  OAI211_X1 U22132 ( .C1(n19603), .C2(n19248), .A(n19204), .B(n19203), .ZN(
        P2_U3075) );
  AOI22_X1 U22133 ( .A1(n19486), .A2(n19218), .B1(n19211), .B2(n19604), .ZN(
        n19206) );
  AOI22_X1 U22134 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19213), .B1(
        n19605), .B2(n19212), .ZN(n19205) );
  OAI211_X1 U22135 ( .C1(n19489), .C2(n19216), .A(n19206), .B(n19205), .ZN(
        P2_U3076) );
  AOI22_X1 U22136 ( .A1(n19490), .A2(n19218), .B1(n19211), .B2(n19610), .ZN(
        n19208) );
  AOI22_X1 U22137 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19213), .B1(
        n19611), .B2(n19212), .ZN(n19207) );
  OAI211_X1 U22138 ( .C1(n19493), .C2(n19216), .A(n19208), .B(n19207), .ZN(
        P2_U3077) );
  AOI22_X1 U22139 ( .A1(n19494), .A2(n19218), .B1(n19211), .B2(n19616), .ZN(
        n19210) );
  AOI22_X1 U22140 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19213), .B1(
        n19617), .B2(n19212), .ZN(n19209) );
  OAI211_X1 U22141 ( .C1(n19497), .C2(n19216), .A(n19210), .B(n19209), .ZN(
        P2_U3078) );
  AOI22_X1 U22142 ( .A1(n19500), .A2(n19218), .B1(n19211), .B2(n19622), .ZN(
        n19215) );
  AOI22_X1 U22143 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19213), .B1(
        n19624), .B2(n19212), .ZN(n19214) );
  OAI211_X1 U22144 ( .C1(n19505), .C2(n19216), .A(n19215), .B(n19214), .ZN(
        P2_U3079) );
  NOR2_X1 U22145 ( .A1(n19464), .A2(n19507), .ZN(n19217) );
  NAND2_X1 U22146 ( .A1(n19217), .A2(n19730), .ZN(n19278) );
  NAND3_X1 U22147 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19734), .A3(
        n19751), .ZN(n19257) );
  NOR2_X1 U22148 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19257), .ZN(
        n19243) );
  AOI22_X1 U22149 ( .A1(n19470), .A2(n19271), .B1(n19573), .B2(n19243), .ZN(
        n19230) );
  NOR2_X1 U22150 ( .A1(n19218), .A2(n19271), .ZN(n19219) );
  OAI21_X1 U22151 ( .B1(n19219), .B2(n19725), .A(n19724), .ZN(n19228) );
  OR2_X1 U22152 ( .A1(n19221), .A2(n19220), .ZN(n19467) );
  NOR2_X1 U22153 ( .A1(n19467), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19224) );
  INV_X1 U22154 ( .A(n19243), .ZN(n19222) );
  OAI211_X1 U22155 ( .C1(n12181), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19222), 
        .B(n19539), .ZN(n19223) );
  INV_X1 U22156 ( .A(n19224), .ZN(n19227) );
  INV_X1 U22157 ( .A(n12181), .ZN(n19225) );
  OAI21_X1 U22158 ( .B1(n19225), .B2(n19243), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19226) );
  AOI22_X1 U22159 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19245), .B1(
        n19574), .B2(n19244), .ZN(n19229) );
  OAI211_X1 U22160 ( .C1(n19473), .C2(n19248), .A(n19230), .B(n19229), .ZN(
        P2_U3080) );
  AOI22_X1 U22161 ( .A1(n19474), .A2(n19271), .B1(n19586), .B2(n19243), .ZN(
        n19232) );
  AOI22_X1 U22162 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19245), .B1(
        n19587), .B2(n19244), .ZN(n19231) );
  OAI211_X1 U22163 ( .C1(n19477), .C2(n19248), .A(n19232), .B(n19231), .ZN(
        P2_U3081) );
  AOI22_X1 U22164 ( .A1(n19478), .A2(n19271), .B1(n19592), .B2(n19243), .ZN(
        n19234) );
  AOI22_X1 U22165 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19245), .B1(
        n19593), .B2(n19244), .ZN(n19233) );
  OAI211_X1 U22166 ( .C1(n19481), .C2(n19248), .A(n19234), .B(n19233), .ZN(
        P2_U3082) );
  AOI22_X1 U22167 ( .A1(n19482), .A2(n19271), .B1(n19598), .B2(n19243), .ZN(
        n19236) );
  AOI22_X1 U22168 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19245), .B1(
        n19599), .B2(n19244), .ZN(n19235) );
  OAI211_X1 U22169 ( .C1(n19485), .C2(n19248), .A(n19236), .B(n19235), .ZN(
        P2_U3083) );
  AOI22_X1 U22170 ( .A1(n19486), .A2(n19271), .B1(n19604), .B2(n19243), .ZN(
        n19238) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19245), .B1(
        n19605), .B2(n19244), .ZN(n19237) );
  OAI211_X1 U22172 ( .C1(n19489), .C2(n19248), .A(n19238), .B(n19237), .ZN(
        P2_U3084) );
  AOI22_X1 U22173 ( .A1(n19490), .A2(n19271), .B1(n19610), .B2(n19243), .ZN(
        n19240) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19245), .B1(
        n19611), .B2(n19244), .ZN(n19239) );
  OAI211_X1 U22175 ( .C1(n19493), .C2(n19248), .A(n19240), .B(n19239), .ZN(
        P2_U3085) );
  AOI22_X1 U22176 ( .A1(n19494), .A2(n19271), .B1(n19616), .B2(n19243), .ZN(
        n19242) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19245), .B1(
        n19617), .B2(n19244), .ZN(n19241) );
  OAI211_X1 U22178 ( .C1(n19497), .C2(n19248), .A(n19242), .B(n19241), .ZN(
        P2_U3086) );
  AOI22_X1 U22179 ( .A1(n19500), .A2(n19271), .B1(n19622), .B2(n19243), .ZN(
        n19247) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19245), .B1(
        n19624), .B2(n19244), .ZN(n19246) );
  OAI211_X1 U22181 ( .C1(n19505), .C2(n19248), .A(n19247), .B(n19246), .ZN(
        P2_U3087) );
  INV_X1 U22182 ( .A(n19470), .ZN(n19585) );
  NOR2_X1 U22183 ( .A1(n19464), .A2(n19752), .ZN(n19249) );
  NOR2_X1 U22184 ( .A1(n19757), .A2(n19257), .ZN(n19282) );
  AOI22_X1 U22185 ( .A1(n19582), .A2(n19271), .B1(n19573), .B2(n19282), .ZN(
        n19260) );
  INV_X1 U22186 ( .A(n19464), .ZN(n19250) );
  NAND3_X1 U22187 ( .A1(n19730), .A2(n19250), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19251) );
  NAND2_X1 U22188 ( .A1(n19251), .A2(n19724), .ZN(n19258) );
  INV_X1 U22189 ( .A(n19257), .ZN(n19254) );
  INV_X1 U22190 ( .A(n19282), .ZN(n19252) );
  OAI211_X1 U22191 ( .C1(n12182), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19252), 
        .B(n19539), .ZN(n19253) );
  OAI211_X1 U22192 ( .C1(n19258), .C2(n19254), .A(n19576), .B(n19253), .ZN(
        n19275) );
  INV_X1 U22193 ( .A(n12182), .ZN(n19255) );
  OAI21_X1 U22194 ( .B1(n19255), .B2(n19282), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19256) );
  OAI21_X1 U22195 ( .B1(n19258), .B2(n19257), .A(n19256), .ZN(n19274) );
  AOI22_X1 U22196 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19275), .B1(
        n19574), .B2(n19274), .ZN(n19259) );
  OAI211_X1 U22197 ( .C1(n19585), .C2(n19285), .A(n19260), .B(n19259), .ZN(
        P2_U3088) );
  AOI22_X1 U22198 ( .A1(n19474), .A2(n19307), .B1(n19586), .B2(n19282), .ZN(
        n19262) );
  AOI22_X1 U22199 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19275), .B1(
        n19587), .B2(n19274), .ZN(n19261) );
  OAI211_X1 U22200 ( .C1(n19477), .C2(n19278), .A(n19262), .B(n19261), .ZN(
        P2_U3089) );
  AOI22_X1 U22201 ( .A1(n19594), .A2(n19271), .B1(n19592), .B2(n19282), .ZN(
        n19264) );
  AOI22_X1 U22202 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19275), .B1(
        n19593), .B2(n19274), .ZN(n19263) );
  OAI211_X1 U22203 ( .C1(n19597), .C2(n19285), .A(n19264), .B(n19263), .ZN(
        P2_U3090) );
  AOI22_X1 U22204 ( .A1(n19482), .A2(n19307), .B1(n19598), .B2(n19282), .ZN(
        n19266) );
  AOI22_X1 U22205 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19275), .B1(
        n19599), .B2(n19274), .ZN(n19265) );
  OAI211_X1 U22206 ( .C1(n19485), .C2(n19278), .A(n19266), .B(n19265), .ZN(
        P2_U3091) );
  AOI22_X1 U22207 ( .A1(n19486), .A2(n19307), .B1(n19604), .B2(n19282), .ZN(
        n19268) );
  AOI22_X1 U22208 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19275), .B1(
        n19605), .B2(n19274), .ZN(n19267) );
  OAI211_X1 U22209 ( .C1(n19489), .C2(n19278), .A(n19268), .B(n19267), .ZN(
        P2_U3092) );
  AOI22_X1 U22210 ( .A1(n19490), .A2(n19307), .B1(n19610), .B2(n19282), .ZN(
        n19270) );
  AOI22_X1 U22211 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19275), .B1(
        n19611), .B2(n19274), .ZN(n19269) );
  OAI211_X1 U22212 ( .C1(n19493), .C2(n19278), .A(n19270), .B(n19269), .ZN(
        P2_U3093) );
  INV_X1 U22213 ( .A(n19494), .ZN(n19621) );
  AOI22_X1 U22214 ( .A1(n19618), .A2(n19271), .B1(n19616), .B2(n19282), .ZN(
        n19273) );
  AOI22_X1 U22215 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19275), .B1(
        n19617), .B2(n19274), .ZN(n19272) );
  OAI211_X1 U22216 ( .C1(n19621), .C2(n19285), .A(n19273), .B(n19272), .ZN(
        P2_U3094) );
  AOI22_X1 U22217 ( .A1(n19500), .A2(n19307), .B1(n19622), .B2(n19282), .ZN(
        n19277) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19275), .B1(
        n19624), .B2(n19274), .ZN(n19276) );
  OAI211_X1 U22219 ( .C1(n19505), .C2(n19278), .A(n19277), .B(n19276), .ZN(
        P2_U3095) );
  INV_X1 U22220 ( .A(n19279), .ZN(n19280) );
  NAND2_X1 U22221 ( .A1(n19730), .A2(n19280), .ZN(n19731) );
  INV_X1 U22222 ( .A(n19731), .ZN(n19281) );
  NAND2_X1 U22223 ( .A1(n19734), .A2(n19571), .ZN(n19313) );
  NOR2_X1 U22224 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19313), .ZN(
        n19305) );
  NOR2_X1 U22225 ( .A1(n19305), .A2(n19282), .ZN(n19286) );
  INV_X1 U22226 ( .A(n12187), .ZN(n19283) );
  OAI21_X1 U22227 ( .B1(n19283), .B2(n19305), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19284) );
  OAI21_X1 U22228 ( .B1(n19286), .B2(n19539), .A(n19284), .ZN(n19306) );
  AOI22_X1 U22229 ( .A1(n19306), .A2(n19574), .B1(n19573), .B2(n19305), .ZN(
        n19292) );
  AOI21_X1 U22230 ( .B1(n19335), .B2(n19285), .A(n19725), .ZN(n19290) );
  INV_X1 U22231 ( .A(n19286), .ZN(n19289) );
  INV_X1 U22232 ( .A(n19305), .ZN(n19287) );
  OAI211_X1 U22233 ( .C1(n12187), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19287), 
        .B(n19539), .ZN(n19288) );
  OAI211_X1 U22234 ( .C1(n19290), .C2(n19289), .A(n19576), .B(n19288), .ZN(
        n19308) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19582), .ZN(n19291) );
  OAI211_X1 U22236 ( .C1(n19585), .C2(n19335), .A(n19292), .B(n19291), .ZN(
        P2_U3096) );
  AOI22_X1 U22237 ( .A1(n19306), .A2(n19587), .B1(n19586), .B2(n19305), .ZN(
        n19294) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19588), .ZN(n19293) );
  OAI211_X1 U22239 ( .C1(n19591), .C2(n19335), .A(n19294), .B(n19293), .ZN(
        P2_U3097) );
  AOI22_X1 U22240 ( .A1(n19306), .A2(n19593), .B1(n19592), .B2(n19305), .ZN(
        n19296) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19594), .ZN(n19295) );
  OAI211_X1 U22242 ( .C1(n19597), .C2(n19335), .A(n19296), .B(n19295), .ZN(
        P2_U3098) );
  AOI22_X1 U22243 ( .A1(n19306), .A2(n19599), .B1(n19598), .B2(n19305), .ZN(
        n19298) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19600), .ZN(n19297) );
  OAI211_X1 U22245 ( .C1(n19603), .C2(n19335), .A(n19298), .B(n19297), .ZN(
        P2_U3099) );
  INV_X1 U22246 ( .A(n19486), .ZN(n19609) );
  AOI22_X1 U22247 ( .A1(n19306), .A2(n19605), .B1(n19604), .B2(n19305), .ZN(
        n19300) );
  AOI22_X1 U22248 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19606), .ZN(n19299) );
  OAI211_X1 U22249 ( .C1(n19609), .C2(n19335), .A(n19300), .B(n19299), .ZN(
        P2_U3100) );
  INV_X1 U22250 ( .A(n19490), .ZN(n19615) );
  AOI22_X1 U22251 ( .A1(n19306), .A2(n19611), .B1(n19610), .B2(n19305), .ZN(
        n19302) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19612), .ZN(n19301) );
  OAI211_X1 U22253 ( .C1(n19615), .C2(n19335), .A(n19302), .B(n19301), .ZN(
        P2_U3101) );
  AOI22_X1 U22254 ( .A1(n19306), .A2(n19617), .B1(n19616), .B2(n19305), .ZN(
        n19304) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19618), .ZN(n19303) );
  OAI211_X1 U22256 ( .C1(n19621), .C2(n19335), .A(n19304), .B(n19303), .ZN(
        P2_U3102) );
  INV_X1 U22257 ( .A(n19500), .ZN(n19632) );
  AOI22_X1 U22258 ( .A1(n19306), .A2(n19624), .B1(n19622), .B2(n19305), .ZN(
        n19310) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19626), .ZN(n19309) );
  OAI211_X1 U22260 ( .C1(n19632), .C2(n19335), .A(n19310), .B(n19309), .ZN(
        P2_U3103) );
  INV_X1 U22261 ( .A(n12185), .ZN(n19311) );
  NOR2_X1 U22262 ( .A1(n19757), .A2(n19313), .ZN(n19343) );
  OAI21_X1 U22263 ( .B1(n19311), .B2(n19343), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19312) );
  OAI21_X1 U22264 ( .B1(n19313), .B2(n19539), .A(n19312), .ZN(n19330) );
  AOI22_X1 U22265 ( .A1(n19330), .A2(n19574), .B1(n19573), .B2(n19343), .ZN(
        n19317) );
  OAI21_X1 U22266 ( .B1(n19731), .B2(n19725), .A(n19313), .ZN(n19315) );
  INV_X1 U22267 ( .A(n19343), .ZN(n19340) );
  OAI211_X1 U22268 ( .C1(n12185), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19340), 
        .B(n19539), .ZN(n19314) );
  NAND3_X1 U22269 ( .A1(n19315), .A2(n19576), .A3(n19314), .ZN(n19332) );
  AOI22_X1 U22270 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19470), .ZN(n19316) );
  OAI211_X1 U22271 ( .C1(n19473), .C2(n19335), .A(n19317), .B(n19316), .ZN(
        P2_U3104) );
  AOI22_X1 U22272 ( .A1(n19330), .A2(n19587), .B1(n19586), .B2(n19343), .ZN(
        n19319) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19474), .ZN(n19318) );
  OAI211_X1 U22274 ( .C1(n19477), .C2(n19335), .A(n19319), .B(n19318), .ZN(
        P2_U3105) );
  AOI22_X1 U22275 ( .A1(n19330), .A2(n19593), .B1(n19592), .B2(n19343), .ZN(
        n19321) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19478), .ZN(n19320) );
  OAI211_X1 U22277 ( .C1(n19481), .C2(n19335), .A(n19321), .B(n19320), .ZN(
        P2_U3106) );
  AOI22_X1 U22278 ( .A1(n19330), .A2(n19599), .B1(n19598), .B2(n19343), .ZN(
        n19323) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19482), .ZN(n19322) );
  OAI211_X1 U22280 ( .C1(n19485), .C2(n19335), .A(n19323), .B(n19322), .ZN(
        P2_U3107) );
  AOI22_X1 U22281 ( .A1(n19330), .A2(n19605), .B1(n19604), .B2(n19343), .ZN(
        n19325) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19486), .ZN(n19324) );
  OAI211_X1 U22283 ( .C1(n19489), .C2(n19335), .A(n19325), .B(n19324), .ZN(
        P2_U3108) );
  AOI22_X1 U22284 ( .A1(n19330), .A2(n19611), .B1(n19610), .B2(n19343), .ZN(
        n19327) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19490), .ZN(n19326) );
  OAI211_X1 U22286 ( .C1(n19493), .C2(n19335), .A(n19327), .B(n19326), .ZN(
        P2_U3109) );
  AOI22_X1 U22287 ( .A1(n19330), .A2(n19617), .B1(n19616), .B2(n19343), .ZN(
        n19329) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19494), .ZN(n19328) );
  OAI211_X1 U22289 ( .C1(n19497), .C2(n19335), .A(n19329), .B(n19328), .ZN(
        P2_U3110) );
  AOI22_X1 U22290 ( .A1(n19330), .A2(n19624), .B1(n19622), .B2(n19343), .ZN(
        n19334) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19332), .B1(
        n19331), .B2(n19500), .ZN(n19333) );
  OAI211_X1 U22292 ( .C1(n19505), .C2(n19335), .A(n19334), .B(n19333), .ZN(
        P2_U3111) );
  INV_X1 U22293 ( .A(n19738), .ZN(n19336) );
  NAND2_X1 U22294 ( .A1(n19744), .A2(n19752), .ZN(n19337) );
  NAND2_X1 U22295 ( .A1(n19742), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19432) );
  NOR2_X1 U22296 ( .A1(n19432), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19372) );
  INV_X1 U22297 ( .A(n19372), .ZN(n19375) );
  NOR2_X1 U22298 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19375), .ZN(
        n19361) );
  AOI22_X1 U22299 ( .A1(n19470), .A2(n19393), .B1(n19573), .B2(n19361), .ZN(
        n19348) );
  NAND2_X1 U22300 ( .A1(n19386), .A2(n19366), .ZN(n19338) );
  AOI21_X1 U22301 ( .B1(n19338), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19539), 
        .ZN(n19342) );
  INV_X1 U22302 ( .A(n12186), .ZN(n19344) );
  OAI21_X1 U22303 ( .B1(n19344), .B2(n19784), .A(n20926), .ZN(n19339) );
  AOI21_X1 U22304 ( .B1(n19342), .B2(n19340), .A(n19339), .ZN(n19341) );
  OAI21_X1 U22305 ( .B1(n19361), .B2(n19343), .A(n19342), .ZN(n19346) );
  OAI21_X1 U22306 ( .B1(n19344), .B2(n19361), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19345) );
  NAND2_X1 U22307 ( .A1(n19346), .A2(n19345), .ZN(n19362) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19363), .B1(
        n19574), .B2(n19362), .ZN(n19347) );
  OAI211_X1 U22309 ( .C1(n19473), .C2(n19366), .A(n19348), .B(n19347), .ZN(
        P2_U3112) );
  AOI22_X1 U22310 ( .A1(n19474), .A2(n19393), .B1(n19586), .B2(n19361), .ZN(
        n19350) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19363), .B1(
        n19362), .B2(n19587), .ZN(n19349) );
  OAI211_X1 U22312 ( .C1(n19477), .C2(n19366), .A(n19350), .B(n19349), .ZN(
        P2_U3113) );
  AOI22_X1 U22313 ( .A1(n19478), .A2(n19393), .B1(n19592), .B2(n19361), .ZN(
        n19352) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19363), .B1(
        n19362), .B2(n19593), .ZN(n19351) );
  OAI211_X1 U22315 ( .C1(n19481), .C2(n19366), .A(n19352), .B(n19351), .ZN(
        P2_U3114) );
  AOI22_X1 U22316 ( .A1(n19482), .A2(n19393), .B1(n19598), .B2(n19361), .ZN(
        n19354) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19363), .B1(
        n19362), .B2(n19599), .ZN(n19353) );
  OAI211_X1 U22318 ( .C1(n19485), .C2(n19366), .A(n19354), .B(n19353), .ZN(
        P2_U3115) );
  AOI22_X1 U22319 ( .A1(n19486), .A2(n19393), .B1(n19604), .B2(n19361), .ZN(
        n19356) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19363), .B1(
        n19362), .B2(n19605), .ZN(n19355) );
  OAI211_X1 U22321 ( .C1(n19489), .C2(n19366), .A(n19356), .B(n19355), .ZN(
        P2_U3116) );
  AOI22_X1 U22322 ( .A1(n19490), .A2(n19393), .B1(n19610), .B2(n19361), .ZN(
        n19358) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19363), .B1(
        n19362), .B2(n19611), .ZN(n19357) );
  OAI211_X1 U22324 ( .C1(n19493), .C2(n19366), .A(n19358), .B(n19357), .ZN(
        P2_U3117) );
  AOI22_X1 U22325 ( .A1(n19494), .A2(n19393), .B1(n19616), .B2(n19361), .ZN(
        n19360) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19363), .B1(
        n19362), .B2(n19617), .ZN(n19359) );
  OAI211_X1 U22327 ( .C1(n19497), .C2(n19366), .A(n19360), .B(n19359), .ZN(
        P2_U3118) );
  AOI22_X1 U22328 ( .A1(n19500), .A2(n19393), .B1(n19622), .B2(n19361), .ZN(
        n19365) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19363), .B1(
        n19362), .B2(n19624), .ZN(n19364) );
  OAI211_X1 U22330 ( .C1(n19505), .C2(n19366), .A(n19365), .B(n19364), .ZN(
        P2_U3119) );
  NOR2_X1 U22331 ( .A1(n19367), .A2(n19432), .ZN(n19404) );
  AOI22_X1 U22332 ( .A1(n19582), .A2(n19393), .B1(n19404), .B2(n19573), .ZN(
        n19378) );
  INV_X1 U22333 ( .A(n19368), .ZN(n19402) );
  NAND3_X1 U22334 ( .A1(n19402), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19744), 
        .ZN(n19369) );
  NAND2_X1 U22335 ( .A1(n19369), .A2(n19724), .ZN(n19376) );
  INV_X1 U22336 ( .A(n19404), .ZN(n19370) );
  OAI211_X1 U22337 ( .C1(n12196), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19370), 
        .B(n19539), .ZN(n19371) );
  OAI211_X1 U22338 ( .C1(n19376), .C2(n19372), .A(n19576), .B(n19371), .ZN(
        n19395) );
  INV_X1 U22339 ( .A(n12196), .ZN(n19373) );
  OAI21_X1 U22340 ( .B1(n19373), .B2(n19404), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19374) );
  OAI21_X1 U22341 ( .B1(n19376), .B2(n19375), .A(n19374), .ZN(n19394) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19395), .B1(
        n19574), .B2(n19394), .ZN(n19377) );
  OAI211_X1 U22343 ( .C1(n19585), .C2(n19427), .A(n19378), .B(n19377), .ZN(
        P2_U3120) );
  AOI22_X1 U22344 ( .A1(n19588), .A2(n19393), .B1(n19404), .B2(n19586), .ZN(
        n19380) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19395), .B1(
        n19587), .B2(n19394), .ZN(n19379) );
  OAI211_X1 U22346 ( .C1(n19591), .C2(n19427), .A(n19380), .B(n19379), .ZN(
        P2_U3121) );
  AOI22_X1 U22347 ( .A1(n19594), .A2(n19393), .B1(n19404), .B2(n19592), .ZN(
        n19382) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19395), .B1(
        n19593), .B2(n19394), .ZN(n19381) );
  OAI211_X1 U22349 ( .C1(n19597), .C2(n19427), .A(n19382), .B(n19381), .ZN(
        P2_U3122) );
  INV_X1 U22350 ( .A(n19427), .ZN(n19383) );
  AOI22_X1 U22351 ( .A1(n19383), .A2(n19482), .B1(n19598), .B2(n19404), .ZN(
        n19385) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19395), .B1(
        n19599), .B2(n19394), .ZN(n19384) );
  OAI211_X1 U22353 ( .C1(n19485), .C2(n19386), .A(n19385), .B(n19384), .ZN(
        P2_U3123) );
  AOI22_X1 U22354 ( .A1(n19606), .A2(n19393), .B1(n19404), .B2(n19604), .ZN(
        n19388) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19395), .B1(
        n19605), .B2(n19394), .ZN(n19387) );
  OAI211_X1 U22356 ( .C1(n19609), .C2(n19427), .A(n19388), .B(n19387), .ZN(
        P2_U3124) );
  AOI22_X1 U22357 ( .A1(n19612), .A2(n19393), .B1(n19404), .B2(n19610), .ZN(
        n19390) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19395), .B1(
        n19611), .B2(n19394), .ZN(n19389) );
  OAI211_X1 U22359 ( .C1(n19615), .C2(n19427), .A(n19390), .B(n19389), .ZN(
        P2_U3125) );
  AOI22_X1 U22360 ( .A1(n19618), .A2(n19393), .B1(n19404), .B2(n19616), .ZN(
        n19392) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19395), .B1(
        n19617), .B2(n19394), .ZN(n19391) );
  OAI211_X1 U22362 ( .C1(n19621), .C2(n19427), .A(n19392), .B(n19391), .ZN(
        P2_U3126) );
  AOI22_X1 U22363 ( .A1(n19626), .A2(n19393), .B1(n19404), .B2(n19622), .ZN(
        n19397) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19395), .B1(
        n19624), .B2(n19394), .ZN(n19396) );
  OAI211_X1 U22365 ( .C1(n19632), .C2(n19427), .A(n19397), .B(n19396), .ZN(
        P2_U3127) );
  INV_X1 U22366 ( .A(n12190), .ZN(n19399) );
  NOR2_X1 U22367 ( .A1(n19398), .A2(n19432), .ZN(n19422) );
  OAI21_X1 U22368 ( .B1(n19399), .B2(n19422), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19400) );
  OAI21_X1 U22369 ( .B1(n19432), .B2(n19401), .A(n19400), .ZN(n19423) );
  AOI22_X1 U22370 ( .A1(n19423), .A2(n19574), .B1(n19573), .B2(n19422), .ZN(
        n19409) );
  NAND2_X1 U22371 ( .A1(n19402), .A2(n19746), .ZN(n19435) );
  INV_X1 U22372 ( .A(n19455), .ZN(n19403) );
  NAND2_X1 U22373 ( .A1(n19403), .A2(n19427), .ZN(n19405) );
  AOI21_X1 U22374 ( .B1(n19405), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19404), 
        .ZN(n19406) );
  AOI211_X1 U22375 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n12190), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19406), .ZN(n19407) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19424), .B1(
        n19455), .B2(n19470), .ZN(n19408) );
  OAI211_X1 U22377 ( .C1(n19473), .C2(n19427), .A(n19409), .B(n19408), .ZN(
        P2_U3128) );
  AOI22_X1 U22378 ( .A1(n19423), .A2(n19587), .B1(n19586), .B2(n19422), .ZN(
        n19411) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19424), .B1(
        n19455), .B2(n19474), .ZN(n19410) );
  OAI211_X1 U22380 ( .C1(n19477), .C2(n19427), .A(n19411), .B(n19410), .ZN(
        P2_U3129) );
  AOI22_X1 U22381 ( .A1(n19423), .A2(n19593), .B1(n19592), .B2(n19422), .ZN(
        n19413) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19424), .B1(
        n19455), .B2(n19478), .ZN(n19412) );
  OAI211_X1 U22383 ( .C1(n19481), .C2(n19427), .A(n19413), .B(n19412), .ZN(
        P2_U3130) );
  AOI22_X1 U22384 ( .A1(n19423), .A2(n19599), .B1(n19598), .B2(n19422), .ZN(
        n19415) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19424), .B1(
        n19455), .B2(n19482), .ZN(n19414) );
  OAI211_X1 U22386 ( .C1(n19485), .C2(n19427), .A(n19415), .B(n19414), .ZN(
        P2_U3131) );
  AOI22_X1 U22387 ( .A1(n19423), .A2(n19605), .B1(n19604), .B2(n19422), .ZN(
        n19417) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19424), .B1(
        n19455), .B2(n19486), .ZN(n19416) );
  OAI211_X1 U22389 ( .C1(n19489), .C2(n19427), .A(n19417), .B(n19416), .ZN(
        P2_U3132) );
  AOI22_X1 U22390 ( .A1(n19423), .A2(n19611), .B1(n19610), .B2(n19422), .ZN(
        n19419) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19424), .B1(
        n19455), .B2(n19490), .ZN(n19418) );
  OAI211_X1 U22392 ( .C1(n19493), .C2(n19427), .A(n19419), .B(n19418), .ZN(
        P2_U3133) );
  AOI22_X1 U22393 ( .A1(n19423), .A2(n19617), .B1(n19616), .B2(n19422), .ZN(
        n19421) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19424), .B1(
        n19455), .B2(n19494), .ZN(n19420) );
  OAI211_X1 U22395 ( .C1(n19497), .C2(n19427), .A(n19421), .B(n19420), .ZN(
        P2_U3134) );
  AOI22_X1 U22396 ( .A1(n19423), .A2(n19624), .B1(n19622), .B2(n19422), .ZN(
        n19426) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19424), .B1(
        n19455), .B2(n19500), .ZN(n19425) );
  OAI211_X1 U22398 ( .C1(n19505), .C2(n19427), .A(n19426), .B(n19425), .ZN(
        P2_U3135) );
  NOR2_X1 U22399 ( .A1(n19429), .A2(n19432), .ZN(n19453) );
  INV_X1 U22400 ( .A(n19453), .ZN(n19430) );
  NAND3_X1 U22401 ( .A1(n19431), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19430), 
        .ZN(n19436) );
  OR2_X1 U22402 ( .A1(n19751), .A2(n19432), .ZN(n19434) );
  OAI21_X1 U22403 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19434), .A(n19784), 
        .ZN(n19433) );
  AND2_X1 U22404 ( .A1(n19436), .A2(n19433), .ZN(n19454) );
  AOI22_X1 U22405 ( .A1(n19454), .A2(n19574), .B1(n19573), .B2(n19453), .ZN(
        n19440) );
  OAI21_X1 U22406 ( .B1(n19435), .B2(n19725), .A(n19434), .ZN(n19437) );
  AND2_X1 U22407 ( .A1(n19437), .A2(n19436), .ZN(n19438) );
  OAI211_X1 U22408 ( .C1(n19453), .C2(n20926), .A(n19576), .B(n19438), .ZN(
        n19456) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19456), .B1(
        n19455), .B2(n19582), .ZN(n19439) );
  OAI211_X1 U22410 ( .C1(n19585), .C2(n19504), .A(n19440), .B(n19439), .ZN(
        P2_U3136) );
  AOI22_X1 U22411 ( .A1(n19454), .A2(n19587), .B1(n19586), .B2(n19453), .ZN(
        n19442) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19456), .B1(
        n19455), .B2(n19588), .ZN(n19441) );
  OAI211_X1 U22413 ( .C1(n19591), .C2(n19504), .A(n19442), .B(n19441), .ZN(
        P2_U3137) );
  AOI22_X1 U22414 ( .A1(n19454), .A2(n19593), .B1(n19592), .B2(n19453), .ZN(
        n19444) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19456), .B1(
        n19455), .B2(n19594), .ZN(n19443) );
  OAI211_X1 U22416 ( .C1(n19597), .C2(n19504), .A(n19444), .B(n19443), .ZN(
        P2_U3138) );
  AOI22_X1 U22417 ( .A1(n19454), .A2(n19599), .B1(n19598), .B2(n19453), .ZN(
        n19446) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19456), .B1(
        n19455), .B2(n19600), .ZN(n19445) );
  OAI211_X1 U22419 ( .C1(n19603), .C2(n19504), .A(n19446), .B(n19445), .ZN(
        P2_U3139) );
  AOI22_X1 U22420 ( .A1(n19454), .A2(n19605), .B1(n19604), .B2(n19453), .ZN(
        n19448) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19456), .B1(
        n19455), .B2(n19606), .ZN(n19447) );
  OAI211_X1 U22422 ( .C1(n19609), .C2(n19504), .A(n19448), .B(n19447), .ZN(
        P2_U3140) );
  AOI22_X1 U22423 ( .A1(n19454), .A2(n19611), .B1(n19610), .B2(n19453), .ZN(
        n19450) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19456), .B1(
        n19455), .B2(n19612), .ZN(n19449) );
  OAI211_X1 U22425 ( .C1(n19615), .C2(n19504), .A(n19450), .B(n19449), .ZN(
        P2_U3141) );
  AOI22_X1 U22426 ( .A1(n19454), .A2(n19617), .B1(n19616), .B2(n19453), .ZN(
        n19452) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19456), .B1(
        n19455), .B2(n19618), .ZN(n19451) );
  OAI211_X1 U22428 ( .C1(n19621), .C2(n19504), .A(n19452), .B(n19451), .ZN(
        P2_U3142) );
  AOI22_X1 U22429 ( .A1(n19454), .A2(n19624), .B1(n19622), .B2(n19453), .ZN(
        n19458) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19456), .B1(
        n19455), .B2(n19626), .ZN(n19457) );
  OAI211_X1 U22431 ( .C1(n19632), .C2(n19504), .A(n19458), .B(n19457), .ZN(
        P2_U3143) );
  INV_X1 U22432 ( .A(n19459), .ZN(n19462) );
  INV_X1 U22433 ( .A(n19463), .ZN(n19460) );
  NAND3_X1 U22434 ( .A1(n19751), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19513) );
  NOR2_X1 U22435 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19513), .ZN(
        n19498) );
  OAI21_X1 U22436 ( .B1(n19460), .B2(n19498), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19461) );
  OAI21_X1 U22437 ( .B1(n19467), .B2(n19462), .A(n19461), .ZN(n19499) );
  AOI22_X1 U22438 ( .A1(n19499), .A2(n19574), .B1(n19573), .B2(n19498), .ZN(
        n19472) );
  AOI21_X1 U22439 ( .B1(n19463), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19469) );
  NOR2_X2 U22440 ( .A1(n19506), .A2(n19507), .ZN(n19531) );
  OAI21_X1 U22441 ( .B1(n19465), .B2(n19531), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19466) );
  OAI21_X1 U22442 ( .B1(n19467), .B2(n19734), .A(n19466), .ZN(n19468) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19501), .B1(
        n19531), .B2(n19470), .ZN(n19471) );
  OAI211_X1 U22444 ( .C1(n19473), .C2(n19504), .A(n19472), .B(n19471), .ZN(
        P2_U3144) );
  AOI22_X1 U22445 ( .A1(n19499), .A2(n19587), .B1(n19586), .B2(n19498), .ZN(
        n19476) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19501), .B1(
        n19531), .B2(n19474), .ZN(n19475) );
  OAI211_X1 U22447 ( .C1(n19477), .C2(n19504), .A(n19476), .B(n19475), .ZN(
        P2_U3145) );
  AOI22_X1 U22448 ( .A1(n19499), .A2(n19593), .B1(n19592), .B2(n19498), .ZN(
        n19480) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19501), .B1(
        n19531), .B2(n19478), .ZN(n19479) );
  OAI211_X1 U22450 ( .C1(n19481), .C2(n19504), .A(n19480), .B(n19479), .ZN(
        P2_U3146) );
  AOI22_X1 U22451 ( .A1(n19499), .A2(n19599), .B1(n19598), .B2(n19498), .ZN(
        n19484) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19501), .B1(
        n19531), .B2(n19482), .ZN(n19483) );
  OAI211_X1 U22453 ( .C1(n19485), .C2(n19504), .A(n19484), .B(n19483), .ZN(
        P2_U3147) );
  AOI22_X1 U22454 ( .A1(n19499), .A2(n19605), .B1(n19604), .B2(n19498), .ZN(
        n19488) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19501), .B1(
        n19531), .B2(n19486), .ZN(n19487) );
  OAI211_X1 U22456 ( .C1(n19489), .C2(n19504), .A(n19488), .B(n19487), .ZN(
        P2_U3148) );
  AOI22_X1 U22457 ( .A1(n19499), .A2(n19611), .B1(n19610), .B2(n19498), .ZN(
        n19492) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19501), .B1(
        n19531), .B2(n19490), .ZN(n19491) );
  OAI211_X1 U22459 ( .C1(n19493), .C2(n19504), .A(n19492), .B(n19491), .ZN(
        P2_U3149) );
  AOI22_X1 U22460 ( .A1(n19499), .A2(n19617), .B1(n19616), .B2(n19498), .ZN(
        n19496) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19501), .B1(
        n19531), .B2(n19494), .ZN(n19495) );
  OAI211_X1 U22462 ( .C1(n19497), .C2(n19504), .A(n19496), .B(n19495), .ZN(
        P2_U3150) );
  AOI22_X1 U22463 ( .A1(n19499), .A2(n19624), .B1(n19622), .B2(n19498), .ZN(
        n19503) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19501), .B1(
        n19531), .B2(n19500), .ZN(n19502) );
  OAI211_X1 U22465 ( .C1(n19505), .C2(n19504), .A(n19503), .B(n19502), .ZN(
        P2_U3151) );
  NOR2_X1 U22466 ( .A1(n19757), .A2(n19513), .ZN(n19538) );
  NOR3_X1 U22467 ( .A1(n12027), .A2(n19538), .A3(n19784), .ZN(n19512) );
  INV_X1 U22468 ( .A(n19513), .ZN(n19509) );
  AOI21_X1 U22469 ( .B1(n20926), .B2(n19509), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19510) );
  NOR2_X1 U22470 ( .A1(n19512), .A2(n19510), .ZN(n19530) );
  AOI22_X1 U22471 ( .A1(n19530), .A2(n19574), .B1(n19573), .B2(n19538), .ZN(
        n19517) );
  NAND2_X1 U22472 ( .A1(n19511), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19514) );
  AOI21_X1 U22473 ( .B1(n19514), .B2(n19513), .A(n19512), .ZN(n19515) );
  OAI211_X1 U22474 ( .C1(n19538), .C2(n20926), .A(n19576), .B(n19515), .ZN(
        n19532) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19532), .B1(
        n19531), .B2(n19582), .ZN(n19516) );
  OAI211_X1 U22476 ( .C1(n19585), .C2(n19535), .A(n19517), .B(n19516), .ZN(
        P2_U3152) );
  AOI22_X1 U22477 ( .A1(n19530), .A2(n19587), .B1(n19586), .B2(n19538), .ZN(
        n19519) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19532), .B1(
        n19531), .B2(n19588), .ZN(n19518) );
  OAI211_X1 U22479 ( .C1(n19591), .C2(n19535), .A(n19519), .B(n19518), .ZN(
        P2_U3153) );
  AOI22_X1 U22480 ( .A1(n19530), .A2(n19593), .B1(n19592), .B2(n19538), .ZN(
        n19521) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19532), .B1(
        n19531), .B2(n19594), .ZN(n19520) );
  OAI211_X1 U22482 ( .C1(n19597), .C2(n19535), .A(n19521), .B(n19520), .ZN(
        P2_U3154) );
  AOI22_X1 U22483 ( .A1(n19530), .A2(n19599), .B1(n19598), .B2(n19538), .ZN(
        n19523) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19532), .B1(
        n19531), .B2(n19600), .ZN(n19522) );
  OAI211_X1 U22485 ( .C1(n19603), .C2(n19535), .A(n19523), .B(n19522), .ZN(
        P2_U3155) );
  AOI22_X1 U22486 ( .A1(n19530), .A2(n19605), .B1(n19604), .B2(n19538), .ZN(
        n19525) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19532), .B1(
        n19531), .B2(n19606), .ZN(n19524) );
  OAI211_X1 U22488 ( .C1(n19609), .C2(n19535), .A(n19525), .B(n19524), .ZN(
        P2_U3156) );
  AOI22_X1 U22489 ( .A1(n19530), .A2(n19611), .B1(n19610), .B2(n19538), .ZN(
        n19527) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19532), .B1(
        n19531), .B2(n19612), .ZN(n19526) );
  OAI211_X1 U22491 ( .C1(n19615), .C2(n19535), .A(n19527), .B(n19526), .ZN(
        P2_U3157) );
  AOI22_X1 U22492 ( .A1(n19530), .A2(n19617), .B1(n19616), .B2(n19538), .ZN(
        n19529) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19532), .B1(
        n19531), .B2(n19618), .ZN(n19528) );
  OAI211_X1 U22494 ( .C1(n19621), .C2(n19535), .A(n19529), .B(n19528), .ZN(
        P2_U3158) );
  AOI22_X1 U22495 ( .A1(n19530), .A2(n19624), .B1(n19622), .B2(n19538), .ZN(
        n19534) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19532), .B1(
        n19531), .B2(n19626), .ZN(n19533) );
  OAI211_X1 U22497 ( .C1(n19632), .C2(n19535), .A(n19534), .B(n19533), .ZN(
        P2_U3159) );
  NOR3_X2 U22498 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19734), .A3(
        n19536), .ZN(n19562) );
  AOI22_X1 U22499 ( .A1(n19563), .A2(n19582), .B1(n19573), .B2(n19562), .ZN(
        n19549) );
  NOR2_X1 U22500 ( .A1(n19627), .A2(n19563), .ZN(n19537) );
  OAI21_X1 U22501 ( .B1(n19537), .B2(n19725), .A(n19724), .ZN(n19547) );
  NOR2_X1 U22502 ( .A1(n19562), .A2(n19538), .ZN(n19546) );
  INV_X1 U22503 ( .A(n19546), .ZN(n19542) );
  INV_X1 U22504 ( .A(n19562), .ZN(n19540) );
  OAI211_X1 U22505 ( .C1(n19543), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19540), 
        .B(n19539), .ZN(n19541) );
  OAI211_X1 U22506 ( .C1(n19547), .C2(n19542), .A(n19576), .B(n19541), .ZN(
        n19565) );
  INV_X1 U22507 ( .A(n19543), .ZN(n19544) );
  OAI21_X1 U22508 ( .B1(n19544), .B2(n19562), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19545) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19565), .B1(
        n19574), .B2(n19564), .ZN(n19548) );
  OAI211_X1 U22510 ( .C1(n19585), .C2(n19568), .A(n19549), .B(n19548), .ZN(
        P2_U3160) );
  AOI22_X1 U22511 ( .A1(n19563), .A2(n19588), .B1(n19586), .B2(n19562), .ZN(
        n19551) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19565), .B1(
        n19587), .B2(n19564), .ZN(n19550) );
  OAI211_X1 U22513 ( .C1(n19591), .C2(n19568), .A(n19551), .B(n19550), .ZN(
        P2_U3161) );
  AOI22_X1 U22514 ( .A1(n19563), .A2(n19594), .B1(n19592), .B2(n19562), .ZN(
        n19553) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19565), .B1(
        n19593), .B2(n19564), .ZN(n19552) );
  OAI211_X1 U22516 ( .C1(n19597), .C2(n19568), .A(n19553), .B(n19552), .ZN(
        P2_U3162) );
  AOI22_X1 U22517 ( .A1(n19563), .A2(n19600), .B1(n19598), .B2(n19562), .ZN(
        n19555) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19565), .B1(
        n19599), .B2(n19564), .ZN(n19554) );
  OAI211_X1 U22519 ( .C1(n19603), .C2(n19568), .A(n19555), .B(n19554), .ZN(
        P2_U3163) );
  AOI22_X1 U22520 ( .A1(n19563), .A2(n19606), .B1(n19604), .B2(n19562), .ZN(
        n19557) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19565), .B1(
        n19605), .B2(n19564), .ZN(n19556) );
  OAI211_X1 U22522 ( .C1(n19609), .C2(n19568), .A(n19557), .B(n19556), .ZN(
        P2_U3164) );
  AOI22_X1 U22523 ( .A1(n19563), .A2(n19612), .B1(n19610), .B2(n19562), .ZN(
        n19559) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19565), .B1(
        n19611), .B2(n19564), .ZN(n19558) );
  OAI211_X1 U22525 ( .C1(n19615), .C2(n19568), .A(n19559), .B(n19558), .ZN(
        P2_U3165) );
  AOI22_X1 U22526 ( .A1(n19563), .A2(n19618), .B1(n19616), .B2(n19562), .ZN(
        n19561) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19565), .B1(
        n19617), .B2(n19564), .ZN(n19560) );
  OAI211_X1 U22528 ( .C1(n19621), .C2(n19568), .A(n19561), .B(n19560), .ZN(
        P2_U3166) );
  AOI22_X1 U22529 ( .A1(n19563), .A2(n19626), .B1(n19622), .B2(n19562), .ZN(
        n19567) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19565), .B1(
        n19624), .B2(n19564), .ZN(n19566) );
  OAI211_X1 U22531 ( .C1(n19632), .C2(n19568), .A(n19567), .B(n19566), .ZN(
        P2_U3167) );
  AND2_X1 U22532 ( .A1(n19569), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19570) );
  NAND2_X1 U22533 ( .A1(n12198), .A2(n19570), .ZN(n19577) );
  NAND2_X1 U22534 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19571), .ZN(
        n19575) );
  OAI21_X1 U22535 ( .B1(n19575), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19784), 
        .ZN(n19572) );
  AND2_X1 U22536 ( .A1(n19577), .A2(n19572), .ZN(n19625) );
  AOI22_X1 U22537 ( .A1(n19625), .A2(n19574), .B1(n19623), .B2(n19573), .ZN(
        n19584) );
  INV_X1 U22538 ( .A(n19575), .ZN(n19581) );
  OAI211_X1 U22539 ( .C1(n19623), .C2(n20926), .A(n19577), .B(n19576), .ZN(
        n19578) );
  INV_X1 U22540 ( .A(n19578), .ZN(n19579) );
  OAI221_X1 U22541 ( .B1(n19581), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19581), 
        .C2(n19580), .A(n19579), .ZN(n19628) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19628), .B1(
        n19627), .B2(n19582), .ZN(n19583) );
  OAI211_X1 U22543 ( .C1(n19585), .C2(n19631), .A(n19584), .B(n19583), .ZN(
        P2_U3168) );
  AOI22_X1 U22544 ( .A1(n19625), .A2(n19587), .B1(n19623), .B2(n19586), .ZN(
        n19590) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19628), .B1(
        n19627), .B2(n19588), .ZN(n19589) );
  OAI211_X1 U22546 ( .C1(n19591), .C2(n19631), .A(n19590), .B(n19589), .ZN(
        P2_U3169) );
  AOI22_X1 U22547 ( .A1(n19625), .A2(n19593), .B1(n19623), .B2(n19592), .ZN(
        n19596) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19628), .B1(
        n19627), .B2(n19594), .ZN(n19595) );
  OAI211_X1 U22549 ( .C1(n19597), .C2(n19631), .A(n19596), .B(n19595), .ZN(
        P2_U3170) );
  AOI22_X1 U22550 ( .A1(n19625), .A2(n19599), .B1(n19623), .B2(n19598), .ZN(
        n19602) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19628), .B1(
        n19627), .B2(n19600), .ZN(n19601) );
  OAI211_X1 U22552 ( .C1(n19603), .C2(n19631), .A(n19602), .B(n19601), .ZN(
        P2_U3171) );
  AOI22_X1 U22553 ( .A1(n19625), .A2(n19605), .B1(n19623), .B2(n19604), .ZN(
        n19608) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19628), .B1(
        n19627), .B2(n19606), .ZN(n19607) );
  OAI211_X1 U22555 ( .C1(n19609), .C2(n19631), .A(n19608), .B(n19607), .ZN(
        P2_U3172) );
  AOI22_X1 U22556 ( .A1(n19625), .A2(n19611), .B1(n19623), .B2(n19610), .ZN(
        n19614) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19628), .B1(
        n19627), .B2(n19612), .ZN(n19613) );
  OAI211_X1 U22558 ( .C1(n19615), .C2(n19631), .A(n19614), .B(n19613), .ZN(
        P2_U3173) );
  AOI22_X1 U22559 ( .A1(n19625), .A2(n19617), .B1(n19623), .B2(n19616), .ZN(
        n19620) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19628), .B1(
        n19627), .B2(n19618), .ZN(n19619) );
  OAI211_X1 U22561 ( .C1(n19621), .C2(n19631), .A(n19620), .B(n19619), .ZN(
        P2_U3174) );
  AOI22_X1 U22562 ( .A1(n19625), .A2(n19624), .B1(n19623), .B2(n19622), .ZN(
        n19630) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19628), .B1(
        n19627), .B2(n19626), .ZN(n19629) );
  OAI211_X1 U22564 ( .C1(n19632), .C2(n19631), .A(n19630), .B(n19629), .ZN(
        P2_U3175) );
  AOI21_X1 U22565 ( .B1(n19635), .B2(n19634), .A(n19633), .ZN(n19640) );
  OAI211_X1 U22566 ( .C1(n19636), .C2(n19639), .A(n19785), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19637) );
  OAI211_X1 U22567 ( .C1(n19640), .C2(n19639), .A(n19638), .B(n19637), .ZN(
        P2_U3177) );
  AND2_X1 U22568 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(
        P2_U3179) );
  AND2_X1 U22569 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(
        P2_U3180) );
  AND2_X1 U22570 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_29__SCAN_IN), .ZN(
        P2_U3181) );
  AND2_X1 U22571 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(
        P2_U3182) );
  AND2_X1 U22572 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19641), .ZN(
        P2_U3183) );
  AND2_X1 U22573 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(
        P2_U3184) );
  AND2_X1 U22574 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_25__SCAN_IN), .ZN(
        P2_U3185) );
  AND2_X1 U22575 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_24__SCAN_IN), .ZN(
        P2_U3186) );
  AND2_X1 U22576 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(
        P2_U3187) );
  AND2_X1 U22577 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(
        P2_U3188) );
  AND2_X1 U22578 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(
        P2_U3189) );
  AND2_X1 U22579 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_20__SCAN_IN), .ZN(
        P2_U3190) );
  AND2_X1 U22580 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(
        P2_U3191) );
  AND2_X1 U22581 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(
        P2_U3192) );
  AND2_X1 U22582 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(
        P2_U3193) );
  AND2_X1 U22583 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(
        P2_U3194) );
  AND2_X1 U22584 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(
        P2_U3195) );
  AND2_X1 U22585 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(
        P2_U3196) );
  AND2_X1 U22586 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(
        P2_U3197) );
  AND2_X1 U22587 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(
        P2_U3198) );
  AND2_X1 U22588 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        P2_U3199) );
  AND2_X1 U22589 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(
        P2_U3200) );
  AND2_X1 U22590 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(P2_U3201) );
  AND2_X1 U22591 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(P2_U3202) );
  AND2_X1 U22592 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(P2_U3203) );
  AND2_X1 U22593 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(P2_U3204) );
  AND2_X1 U22594 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(P2_U3205) );
  AND2_X1 U22595 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(P2_U3206) );
  AND2_X1 U22596 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(P2_U3207) );
  AND2_X1 U22597 ( .A1(n19641), .A2(P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(P2_U3208) );
  NAND2_X1 U22598 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19785), .ZN(n19650) );
  INV_X1 U22599 ( .A(n19650), .ZN(n19655) );
  INV_X1 U22600 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19645) );
  NOR3_X1 U22601 ( .A1(n19655), .A2(n19645), .A3(n19642), .ZN(n19644) );
  OAI211_X1 U22602 ( .C1(HOLD), .C2(n19645), .A(n19651), .B(n19793), .ZN(
        n19643) );
  NOR2_X1 U22603 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19646) );
  NAND2_X1 U22604 ( .A1(n19646), .A2(NA), .ZN(n19653) );
  OAI211_X1 U22605 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n19644), .A(n19643), 
        .B(n19653), .ZN(P2_U3209) );
  NAND2_X1 U22606 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20692), .ZN(n19654) );
  AOI211_X1 U22607 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n19654), .A(n19646), 
        .B(n19645), .ZN(n19647) );
  NOR3_X1 U22608 ( .A1(n19772), .A2(n19655), .A3(n19647), .ZN(n19648) );
  OAI21_X1 U22609 ( .B1(n19649), .B2(n20692), .A(n19648), .ZN(P2_U3210) );
  OAI22_X1 U22610 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19651), .B1(NA), 
        .B2(n19650), .ZN(n19652) );
  OAI211_X1 U22611 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19652), .ZN(n19657) );
  OAI211_X1 U22612 ( .C1(n19655), .C2(n19654), .A(P2_STATE_REG_2__SCAN_IN), 
        .B(n19653), .ZN(n19656) );
  NAND2_X1 U22613 ( .A1(n19657), .A2(n19656), .ZN(P2_U3211) );
  NAND2_X1 U22614 ( .A1(n19792), .A2(n19658), .ZN(n19702) );
  CLKBUF_X1 U22615 ( .A(n19702), .Z(n19699) );
  OAI222_X1 U22616 ( .A1(n19699), .A2(n19661), .B1(n19660), .B2(n19792), .C1(
        n19659), .C2(n19700), .ZN(P2_U3212) );
  OAI222_X1 U22617 ( .A1(n19702), .A2(n12910), .B1(n19662), .B2(n19792), .C1(
        n19661), .C2(n19700), .ZN(P2_U3213) );
  OAI222_X1 U22618 ( .A1(n19702), .A2(n12911), .B1(n19663), .B2(n19792), .C1(
        n12910), .C2(n19700), .ZN(P2_U3214) );
  OAI222_X1 U22619 ( .A1(n19702), .A2(n12919), .B1(n19664), .B2(n19792), .C1(
        n12911), .C2(n19700), .ZN(P2_U3215) );
  OAI222_X1 U22620 ( .A1(n19702), .A2(n19666), .B1(n19665), .B2(n19792), .C1(
        n12919), .C2(n19700), .ZN(P2_U3216) );
  OAI222_X1 U22621 ( .A1(n19702), .A2(n19668), .B1(n19667), .B2(n19792), .C1(
        n19666), .C2(n19700), .ZN(P2_U3217) );
  OAI222_X1 U22622 ( .A1(n19699), .A2(n12929), .B1(n19669), .B2(n19792), .C1(
        n19668), .C2(n19700), .ZN(P2_U3218) );
  OAI222_X1 U22623 ( .A1(n19699), .A2(n12936), .B1(n19670), .B2(n19792), .C1(
        n12929), .C2(n19700), .ZN(P2_U3219) );
  OAI222_X1 U22624 ( .A1(n19699), .A2(n12937), .B1(n19671), .B2(n19792), .C1(
        n12936), .C2(n19700), .ZN(P2_U3220) );
  INV_X1 U22625 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19673) );
  OAI222_X1 U22626 ( .A1(n19699), .A2(n19673), .B1(n19672), .B2(n19792), .C1(
        n12937), .C2(n19700), .ZN(P2_U3221) );
  OAI222_X1 U22627 ( .A1(n19699), .A2(n12945), .B1(n19674), .B2(n19792), .C1(
        n19673), .C2(n19700), .ZN(P2_U3222) );
  OAI222_X1 U22628 ( .A1(n19699), .A2(n15152), .B1(n19675), .B2(n19792), .C1(
        n12945), .C2(n19700), .ZN(P2_U3223) );
  OAI222_X1 U22629 ( .A1(n19702), .A2(n12951), .B1(n19676), .B2(n19792), .C1(
        n15152), .C2(n19700), .ZN(P2_U3224) );
  OAI222_X1 U22630 ( .A1(n19702), .A2(n12959), .B1(n19677), .B2(n19792), .C1(
        n12951), .C2(n19700), .ZN(P2_U3225) );
  OAI222_X1 U22631 ( .A1(n19702), .A2(n14159), .B1(n19678), .B2(n19792), .C1(
        n12959), .C2(n19700), .ZN(P2_U3226) );
  OAI222_X1 U22632 ( .A1(n19702), .A2(n19680), .B1(n19679), .B2(n19792), .C1(
        n14159), .C2(n19700), .ZN(P2_U3227) );
  OAI222_X1 U22633 ( .A1(n19702), .A2(n12964), .B1(n19681), .B2(n19792), .C1(
        n19680), .C2(n19700), .ZN(P2_U3228) );
  OAI222_X1 U22634 ( .A1(n19702), .A2(n20940), .B1(n19682), .B2(n19792), .C1(
        n12964), .C2(n19700), .ZN(P2_U3229) );
  OAI222_X1 U22635 ( .A1(n19699), .A2(n19684), .B1(n19683), .B2(n19792), .C1(
        n20940), .C2(n19700), .ZN(P2_U3230) );
  OAI222_X1 U22636 ( .A1(n19699), .A2(n19686), .B1(n19685), .B2(n19792), .C1(
        n19684), .C2(n19700), .ZN(P2_U3231) );
  OAI222_X1 U22637 ( .A1(n19699), .A2(n12973), .B1(n20888), .B2(n19792), .C1(
        n19686), .C2(n19700), .ZN(P2_U3232) );
  OAI222_X1 U22638 ( .A1(n19699), .A2(n19688), .B1(n19687), .B2(n19792), .C1(
        n12973), .C2(n19700), .ZN(P2_U3233) );
  OAI222_X1 U22639 ( .A1(n19699), .A2(n12978), .B1(n19689), .B2(n19792), .C1(
        n19688), .C2(n19700), .ZN(P2_U3234) );
  OAI222_X1 U22640 ( .A1(n19699), .A2(n19691), .B1(n19690), .B2(n19792), .C1(
        n12978), .C2(n19700), .ZN(P2_U3235) );
  OAI222_X1 U22641 ( .A1(n19699), .A2(n12983), .B1(n19692), .B2(n19792), .C1(
        n19691), .C2(n19700), .ZN(P2_U3236) );
  OAI222_X1 U22642 ( .A1(n19699), .A2(n19694), .B1(n20943), .B2(n19792), .C1(
        n12983), .C2(n19700), .ZN(P2_U3237) );
  OAI222_X1 U22643 ( .A1(n19700), .A2(n19694), .B1(n19693), .B2(n19792), .C1(
        n19695), .C2(n19699), .ZN(P2_U3238) );
  OAI222_X1 U22644 ( .A1(n19699), .A2(n19697), .B1(n19696), .B2(n19792), .C1(
        n19695), .C2(n19700), .ZN(P2_U3239) );
  OAI222_X1 U22645 ( .A1(n19699), .A2(n12992), .B1(n19698), .B2(n19792), .C1(
        n19697), .C2(n19700), .ZN(P2_U3240) );
  OAI222_X1 U22646 ( .A1(n19702), .A2(n13166), .B1(n19701), .B2(n19792), .C1(
        n12992), .C2(n19700), .ZN(P2_U3241) );
  INV_X1 U22647 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19703) );
  AOI22_X1 U22648 ( .A1(n19792), .A2(n19704), .B1(n19703), .B2(n19793), .ZN(
        P2_U3585) );
  MUX2_X1 U22649 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19792), .Z(P2_U3586) );
  INV_X1 U22650 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19705) );
  AOI22_X1 U22651 ( .A1(n19792), .A2(n19706), .B1(n19705), .B2(n19793), .ZN(
        P2_U3587) );
  INV_X1 U22652 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19707) );
  AOI22_X1 U22653 ( .A1(n19792), .A2(n19708), .B1(n19707), .B2(n19793), .ZN(
        P2_U3588) );
  OAI21_X1 U22654 ( .B1(n19709), .B2(BS16), .A(n20961), .ZN(n20960) );
  OAI21_X1 U22655 ( .B1(n20961), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20960), 
        .ZN(n19710) );
  INV_X1 U22656 ( .A(n19710), .ZN(P2_U3591) );
  OAI21_X1 U22657 ( .B1(n20961), .B2(n19711), .A(n20960), .ZN(P2_U3592) );
  OAI22_X1 U22658 ( .A1(n19730), .A2(n19719), .B1(n19726), .B2(n19712), .ZN(
        n19713) );
  OAI22_X1 U22659 ( .A1(n19714), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19713), .B2(n19720), .ZN(n19715) );
  INV_X1 U22660 ( .A(n19715), .ZN(P2_U3596) );
  OAI222_X1 U22661 ( .A1(n19719), .A2(n19738), .B1(n19726), .B2(n19718), .C1(
        n19717), .C2(n19716), .ZN(n19722) );
  MUX2_X1 U22662 ( .A(n19722), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19720), .Z(P2_U3599) );
  INV_X1 U22663 ( .A(n19747), .ZN(n19723) );
  NAND2_X1 U22664 ( .A1(n19738), .A2(n19723), .ZN(n19735) );
  OAI21_X1 U22665 ( .B1(n19744), .B2(n19725), .A(n19724), .ZN(n19727) );
  AND2_X1 U22666 ( .A1(n19727), .A2(n19726), .ZN(n19737) );
  AND2_X1 U22667 ( .A1(n19735), .A2(n19737), .ZN(n19729) );
  OAI222_X1 U22668 ( .A1(n19747), .A2(n19731), .B1(n19730), .B2(n19729), .C1(
        n20926), .C2(n19728), .ZN(n19732) );
  INV_X1 U22669 ( .A(n19732), .ZN(n19733) );
  AOI22_X1 U22670 ( .A1(n19758), .A2(n19734), .B1(n19733), .B2(n19755), .ZN(
        P2_U3602) );
  NOR2_X1 U22671 ( .A1(n19735), .A2(n19744), .ZN(n19740) );
  OAI22_X1 U22672 ( .A1(n19738), .A2(n19737), .B1(n19736), .B2(n20926), .ZN(
        n19739) );
  NOR2_X1 U22673 ( .A1(n19740), .A2(n19739), .ZN(n19741) );
  AOI22_X1 U22674 ( .A1(n19758), .A2(n19742), .B1(n19741), .B2(n19755), .ZN(
        P2_U3603) );
  OR3_X1 U22675 ( .A1(n19744), .A2(n19782), .A3(n19743), .ZN(n19745) );
  OAI21_X1 U22676 ( .B1(n19747), .B2(n19746), .A(n19745), .ZN(n19748) );
  AOI21_X1 U22677 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19749), .A(n19748), 
        .ZN(n19750) );
  AOI22_X1 U22678 ( .A1(n19758), .A2(n19751), .B1(n19750), .B2(n19755), .ZN(
        P2_U3604) );
  OAI22_X1 U22679 ( .A1(n19752), .A2(n19782), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20926), .ZN(n19753) );
  AOI21_X1 U22680 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19754), .A(n19753), 
        .ZN(n19756) );
  AOI22_X1 U22681 ( .A1(n19758), .A2(n19757), .B1(n19756), .B2(n19755), .ZN(
        P2_U3605) );
  INV_X1 U22682 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19759) );
  AOI22_X1 U22683 ( .A1(n19792), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19759), 
        .B2(n19793), .ZN(P2_U3608) );
  INV_X1 U22684 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19771) );
  INV_X1 U22685 ( .A(n19760), .ZN(n19770) );
  INV_X1 U22686 ( .A(n19761), .ZN(n19765) );
  INV_X1 U22687 ( .A(n19762), .ZN(n19764) );
  AOI22_X1 U22688 ( .A1(n19766), .A2(n19765), .B1(n19764), .B2(n19763), .ZN(
        n19769) );
  NOR2_X1 U22689 ( .A1(n19770), .A2(n19767), .ZN(n19768) );
  AOI22_X1 U22690 ( .A1(n19771), .A2(n19770), .B1(n19769), .B2(n19768), .ZN(
        P2_U3609) );
  NAND2_X1 U22691 ( .A1(n19772), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19777) );
  INV_X1 U22692 ( .A(n19773), .ZN(n19775) );
  AOI22_X1 U22693 ( .A1(n19777), .A2(n19776), .B1(n19775), .B2(n19774), .ZN(
        n19781) );
  NOR2_X1 U22694 ( .A1(n19785), .A2(n19784), .ZN(n19779) );
  OAI22_X1 U22695 ( .A1(n19781), .A2(n19780), .B1(n19779), .B2(n19778), .ZN(
        n19791) );
  INV_X1 U22696 ( .A(n19782), .ZN(n19788) );
  NOR3_X1 U22697 ( .A1(n19785), .A2(n19784), .A3(n19783), .ZN(n19787) );
  AOI211_X1 U22698 ( .C1(n19789), .C2(n19788), .A(n19787), .B(n19786), .ZN(
        n19790) );
  MUX2_X1 U22699 ( .A(n19791), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19790), 
        .Z(P2_U3610) );
  OAI22_X1 U22700 ( .A1(n19793), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19792), .ZN(n19794) );
  INV_X1 U22701 ( .A(n19794), .ZN(P2_U3611) );
  AOI21_X1 U22702 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20704), .A(n20701), 
        .ZN(n19801) );
  INV_X1 U22703 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19795) );
  NAND2_X1 U22704 ( .A1(n20701), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20792) );
  AOI21_X1 U22705 ( .B1(n19801), .B2(n19795), .A(n20794), .ZN(P1_U2802) );
  OAI21_X1 U22706 ( .B1(n19797), .B2(n19796), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19798) );
  OAI21_X1 U22707 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19799), .A(n19798), 
        .ZN(P1_U2803) );
  NOR2_X1 U22708 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19802) );
  OAI21_X1 U22709 ( .B1(n19802), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20792), .ZN(
        n19800) );
  OAI21_X1 U22710 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20792), .A(n19800), 
        .ZN(P1_U2804) );
  NOR2_X1 U22711 ( .A1(n20794), .A2(n19801), .ZN(n20770) );
  OAI21_X1 U22712 ( .B1(BS16), .B2(n19802), .A(n20770), .ZN(n20768) );
  OAI21_X1 U22713 ( .B1(n20770), .B2(n20359), .A(n20768), .ZN(P1_U2805) );
  OAI21_X1 U22714 ( .B1(n19805), .B2(n19804), .A(n19803), .ZN(P1_U2806) );
  NOR4_X1 U22715 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19809) );
  NOR4_X1 U22716 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19808) );
  NOR4_X1 U22717 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19807) );
  NOR4_X1 U22718 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19806) );
  NAND4_X1 U22719 ( .A1(n19809), .A2(n19808), .A3(n19807), .A4(n19806), .ZN(
        n19815) );
  NOR4_X1 U22720 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19813) );
  AOI211_X1 U22721 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_10__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19812) );
  NOR4_X1 U22722 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19811) );
  NOR4_X1 U22723 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19810) );
  NAND4_X1 U22724 ( .A1(n19813), .A2(n19812), .A3(n19811), .A4(n19810), .ZN(
        n19814) );
  NOR2_X1 U22725 ( .A1(n19815), .A2(n19814), .ZN(n20791) );
  INV_X1 U22726 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20763) );
  NOR3_X1 U22727 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19817) );
  OAI21_X1 U22728 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19817), .A(n20791), .ZN(
        n19816) );
  OAI21_X1 U22729 ( .B1(n20791), .B2(n20763), .A(n19816), .ZN(P1_U2807) );
  INV_X1 U22730 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20769) );
  AOI21_X1 U22731 ( .B1(n13525), .B2(n20769), .A(n19817), .ZN(n19818) );
  INV_X1 U22732 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20760) );
  INV_X1 U22733 ( .A(n20791), .ZN(n20786) );
  AOI22_X1 U22734 ( .A1(n20791), .A2(n19818), .B1(n20760), .B2(n20786), .ZN(
        P1_U2808) );
  AOI22_X1 U22735 ( .A1(n19879), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n19883), .B2(
        n19819), .ZN(n19829) );
  AOI22_X1 U22736 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19884), .B1(
        n19860), .B2(n19820), .ZN(n19828) );
  NOR2_X1 U22737 ( .A1(n19857), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n19822) );
  AOI21_X1 U22738 ( .B1(n19822), .B2(n19821), .A(n19868), .ZN(n19827) );
  INV_X1 U22739 ( .A(n19823), .ZN(n19825) );
  AOI22_X1 U22740 ( .A1(n19825), .A2(n19847), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n19824), .ZN(n19826) );
  NAND4_X1 U22741 ( .A1(n19829), .A2(n19828), .A3(n19827), .A4(n19826), .ZN(
        P1_U2831) );
  INV_X1 U22742 ( .A(n19830), .ZN(n19831) );
  AOI22_X1 U22743 ( .A1(n19831), .A2(n19883), .B1(n19860), .B2(n19894), .ZN(
        n19842) );
  NAND2_X1 U22744 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19836) );
  NOR3_X1 U22745 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19857), .A3(n19836), .ZN(
        n19835) );
  INV_X1 U22746 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19897) );
  INV_X1 U22747 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19832) );
  OAI22_X1 U22748 ( .A1(n19833), .A2(n19897), .B1(n19855), .B2(n19832), .ZN(
        n19834) );
  NOR2_X1 U22749 ( .A1(n19835), .A2(n19834), .ZN(n19841) );
  INV_X1 U22750 ( .A(n19836), .ZN(n19837) );
  OAI21_X1 U22751 ( .B1(n19838), .B2(n19837), .A(n19871), .ZN(n19846) );
  AOI22_X1 U22752 ( .A1(n19895), .A2(n19847), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19846), .ZN(n19840) );
  NAND4_X1 U22753 ( .A1(n19842), .A2(n19841), .A3(n19840), .A4(n19839), .ZN(
        P1_U2833) );
  INV_X1 U22754 ( .A(n19843), .ZN(n19844) );
  AOI22_X1 U22755 ( .A1(n19844), .A2(n19883), .B1(n19860), .B2(n19898), .ZN(
        n19851) );
  AOI22_X1 U22756 ( .A1(n19879), .A2(P1_EBX_REG_6__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19884), .ZN(n19850) );
  NOR2_X1 U22757 ( .A1(n19857), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n19845) );
  AOI21_X1 U22758 ( .B1(n19845), .B2(P1_REIP_REG_5__SCAN_IN), .A(n19868), .ZN(
        n19849) );
  AOI22_X1 U22759 ( .A1(n19901), .A2(n19847), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n19846), .ZN(n19848) );
  NAND4_X1 U22760 ( .A1(n19851), .A2(n19850), .A3(n19849), .A4(n19848), .ZN(
        P1_U2834) );
  INV_X1 U22761 ( .A(n19852), .ZN(n19853) );
  AOI22_X1 U22762 ( .A1(n19879), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n19853), .B2(
        n19883), .ZN(n19865) );
  INV_X1 U22763 ( .A(n19854), .ZN(n19859) );
  OAI22_X1 U22764 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19857), .B1(n19856), 
        .B2(n19855), .ZN(n19858) );
  AOI211_X1 U22765 ( .C1(n19860), .C2(n19859), .A(n19868), .B(n19858), .ZN(
        n19864) );
  NOR2_X1 U22766 ( .A1(n19871), .A2(n15924), .ZN(n19861) );
  AOI21_X1 U22767 ( .B1(n19862), .B2(n19889), .A(n19861), .ZN(n19863) );
  NAND3_X1 U22768 ( .A1(n19865), .A2(n19864), .A3(n19863), .ZN(P1_U2835) );
  NOR3_X1 U22769 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19877), .A3(n19866), .ZN(
        n19867) );
  AOI211_X1 U22770 ( .C1(n19884), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19868), .B(n19867), .ZN(n19875) );
  INV_X1 U22771 ( .A(n19952), .ZN(n19869) );
  AOI22_X1 U22772 ( .A1(n19879), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n19869), .B2(
        n19883), .ZN(n19870) );
  OAI21_X1 U22773 ( .B1(n19893), .B2(n19958), .A(n19870), .ZN(n19873) );
  NOR2_X1 U22774 ( .A1(n19871), .A2(n20711), .ZN(n19872) );
  AOI211_X1 U22775 ( .C1(n19946), .C2(n19889), .A(n19873), .B(n19872), .ZN(
        n19874) );
  OAI211_X1 U22776 ( .C1(n19876), .C2(n19887), .A(n19875), .B(n19874), .ZN(
        P1_U2836) );
  NOR3_X1 U22777 ( .A1(n19877), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n13525), .ZN(
        n19878) );
  AOI21_X1 U22778 ( .B1(n19879), .B2(P1_EBX_REG_2__SCAN_IN), .A(n19878), .ZN(
        n19892) );
  OAI21_X1 U22779 ( .B1(n19881), .B2(n19880), .A(P1_REIP_REG_2__SCAN_IN), .ZN(
        n19886) );
  AOI22_X1 U22780 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19884), .B1(
        n19883), .B2(n19882), .ZN(n19885) );
  OAI211_X1 U22781 ( .C1(n13583), .C2(n19887), .A(n19886), .B(n19885), .ZN(
        n19888) );
  AOI21_X1 U22782 ( .B1(n19890), .B2(n19889), .A(n19888), .ZN(n19891) );
  OAI211_X1 U22783 ( .C1(n19893), .C2(n19984), .A(n19892), .B(n19891), .ZN(
        P1_U2838) );
  AOI22_X1 U22784 ( .A1(n19895), .A2(n19900), .B1(n19899), .B2(n19894), .ZN(
        n19896) );
  OAI21_X1 U22785 ( .B1(n19904), .B2(n19897), .A(n19896), .ZN(P1_U2865) );
  INV_X1 U22786 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U22787 ( .A1(n19901), .A2(n19900), .B1(n19899), .B2(n19898), .ZN(
        n19902) );
  OAI21_X1 U22788 ( .B1(n19904), .B2(n19903), .A(n19902), .ZN(P1_U2866) );
  AOI22_X1 U22789 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19908), .B1(n19935), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19905) );
  OAI21_X1 U22790 ( .B1(n19907), .B2(n19906), .A(n19905), .ZN(P1_U2921) );
  AOI22_X1 U22791 ( .A1(n20798), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19909) );
  OAI21_X1 U22792 ( .B1(n19910), .B2(n19938), .A(n19909), .ZN(P1_U2922) );
  AOI22_X1 U22793 ( .A1(n20798), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19911) );
  OAI21_X1 U22794 ( .B1(n19912), .B2(n19938), .A(n19911), .ZN(P1_U2923) );
  AOI22_X1 U22795 ( .A1(n20798), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19913) );
  OAI21_X1 U22796 ( .B1(n14183), .B2(n19938), .A(n19913), .ZN(P1_U2924) );
  AOI22_X1 U22797 ( .A1(n19936), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19914) );
  OAI21_X1 U22798 ( .B1(n19915), .B2(n19938), .A(n19914), .ZN(P1_U2925) );
  AOI22_X1 U22799 ( .A1(n19936), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19916) );
  OAI21_X1 U22800 ( .B1(n19917), .B2(n19938), .A(n19916), .ZN(P1_U2926) );
  AOI22_X1 U22801 ( .A1(n19936), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19918) );
  OAI21_X1 U22802 ( .B1(n19919), .B2(n19938), .A(n19918), .ZN(P1_U2927) );
  AOI22_X1 U22803 ( .A1(n19936), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19920), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19921) );
  OAI21_X1 U22804 ( .B1(n19922), .B2(n19938), .A(n19921), .ZN(P1_U2928) );
  AOI22_X1 U22805 ( .A1(n20798), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19923) );
  OAI21_X1 U22806 ( .B1(n14540), .B2(n19938), .A(n19923), .ZN(P1_U2929) );
  AOI22_X1 U22807 ( .A1(n19936), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19924) );
  OAI21_X1 U22808 ( .B1(n13868), .B2(n19938), .A(n19924), .ZN(P1_U2930) );
  AOI22_X1 U22809 ( .A1(n19936), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19925) );
  OAI21_X1 U22810 ( .B1(n19926), .B2(n19938), .A(n19925), .ZN(P1_U2931) );
  AOI22_X1 U22811 ( .A1(n19936), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19927) );
  OAI21_X1 U22812 ( .B1(n19928), .B2(n19938), .A(n19927), .ZN(P1_U2932) );
  AOI22_X1 U22813 ( .A1(n19936), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19929) );
  OAI21_X1 U22814 ( .B1(n19930), .B2(n19938), .A(n19929), .ZN(P1_U2933) );
  AOI22_X1 U22815 ( .A1(n19936), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19931) );
  OAI21_X1 U22816 ( .B1(n19932), .B2(n19938), .A(n19931), .ZN(P1_U2934) );
  AOI22_X1 U22817 ( .A1(n19936), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19933) );
  OAI21_X1 U22818 ( .B1(n19934), .B2(n19938), .A(n19933), .ZN(P1_U2935) );
  AOI22_X1 U22819 ( .A1(n19936), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19935), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19937) );
  OAI21_X1 U22820 ( .B1(n19939), .B2(n19938), .A(n19937), .ZN(P1_U2936) );
  AOI22_X1 U22821 ( .A1(n19941), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19940), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19951) );
  OR2_X1 U22822 ( .A1(n19943), .A2(n19942), .ZN(n19944) );
  NAND2_X1 U22823 ( .A1(n19945), .A2(n19944), .ZN(n19956) );
  INV_X1 U22824 ( .A(n19956), .ZN(n19949) );
  AOI22_X1 U22825 ( .A1(n19949), .A2(n19948), .B1(n19947), .B2(n19946), .ZN(
        n19950) );
  OAI211_X1 U22826 ( .C1(n19953), .C2(n19952), .A(n19951), .B(n19950), .ZN(
        P1_U2995) );
  INV_X1 U22827 ( .A(n19972), .ZN(n19964) );
  AOI211_X1 U22828 ( .C1(n19963), .C2(n19955), .A(n19954), .B(n19975), .ZN(
        n19961) );
  NOR2_X1 U22829 ( .A1(n19956), .A2(n19977), .ZN(n19960) );
  OAI22_X1 U22830 ( .A1(n19958), .A2(n19983), .B1(n20711), .B2(n19957), .ZN(
        n19959) );
  NOR3_X1 U22831 ( .A1(n19961), .A2(n19960), .A3(n19959), .ZN(n19962) );
  OAI21_X1 U22832 ( .B1(n19964), .B2(n19963), .A(n19962), .ZN(P1_U3027) );
  INV_X1 U22833 ( .A(n19965), .ZN(n19966) );
  AOI21_X1 U22834 ( .B1(n19968), .B2(n19967), .A(n19966), .ZN(n19974) );
  INV_X1 U22835 ( .A(n19969), .ZN(n19971) );
  AOI22_X1 U22836 ( .A1(n19972), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n19971), .B2(n19970), .ZN(n19973) );
  OAI211_X1 U22837 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n19975), .A(
        n19974), .B(n19973), .ZN(P1_U3028) );
  INV_X1 U22838 ( .A(n19976), .ZN(n19991) );
  NOR2_X1 U22839 ( .A1(n19978), .A2(n19977), .ZN(n19987) );
  NAND3_X1 U22840 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U22841 ( .B1(n19981), .B2(n19980), .A(n19979), .ZN(n19986) );
  OAI21_X1 U22842 ( .B1(n19984), .B2(n19983), .A(n19982), .ZN(n19985) );
  AOI211_X1 U22843 ( .C1(n19987), .C2(n13664), .A(n19986), .B(n19985), .ZN(
        n19988) );
  OAI221_X1 U22844 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19991), .C1(
        n19990), .C2(n19989), .A(n19988), .ZN(P1_U3029) );
  NOR2_X1 U22845 ( .A1(n19993), .A2(n19992), .ZN(P1_U3032) );
  NOR2_X2 U22846 ( .A1(n19995), .A2(n19994), .ZN(n20036) );
  NOR2_X2 U22847 ( .A1(n19996), .A2(n19995), .ZN(n20037) );
  AOI22_X1 U22848 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20036), .B1(DATAI_16_), 
        .B2(n20037), .ZN(n20232) );
  INV_X1 U22849 ( .A(n12563), .ZN(n20528) );
  INV_X1 U22850 ( .A(n20622), .ZN(n20573) );
  NAND2_X1 U22851 ( .A1(n20039), .A2(n19999), .ZN(n20395) );
  NAND3_X1 U22852 ( .A1(n20435), .A2(n20394), .A3(n20482), .ZN(n20048) );
  NOR2_X1 U22853 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20048), .ZN(
        n20004) );
  INV_X1 U22854 ( .A(n20004), .ZN(n20040) );
  OAI22_X1 U22855 ( .A1(n20685), .A2(n20630), .B1(n20395), .B2(n20040), .ZN(
        n20000) );
  INV_X1 U22856 ( .A(n20000), .ZN(n20011) );
  AND2_X1 U22857 ( .A1(n20007), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20568) );
  NOR2_X1 U22858 ( .A1(n20568), .A2(n20165), .ZN(n20402) );
  NAND3_X1 U22859 ( .A1(n20077), .A2(n20625), .A3(n20685), .ZN(n20001) );
  NAND2_X1 U22860 ( .A1(n20625), .A2(n20359), .ZN(n20479) );
  NAND2_X1 U22861 ( .A1(n20001), .A2(n20479), .ZN(n20006) );
  OR2_X1 U22862 ( .A1(n20314), .A2(n20002), .ZN(n20047) );
  INV_X1 U22863 ( .A(n20047), .ZN(n20125) );
  NAND2_X1 U22864 ( .A1(n20125), .A2(n20315), .ZN(n20008) );
  INV_X1 U22865 ( .A(n20392), .ZN(n20091) );
  OR2_X1 U22866 ( .A1(n20316), .A2(n20091), .ZN(n20158) );
  AOI22_X1 U22867 ( .A1(n20006), .A2(n20008), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20158), .ZN(n20003) );
  OAI211_X1 U22868 ( .C1(n20004), .C2(n20323), .A(n20402), .B(n20003), .ZN(
        n20044) );
  NOR2_X2 U22869 ( .A1(n20005), .A2(n20165), .ZN(n20618) );
  INV_X1 U22870 ( .A(n20006), .ZN(n20009) );
  OR2_X1 U22871 ( .A1(n20007), .A2(n20689), .ZN(n20164) );
  OAI22_X1 U22872 ( .A1(n20009), .A2(n20008), .B1(n20164), .B2(n20158), .ZN(
        n20043) );
  AOI22_X1 U22873 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20044), .B1(
        n20618), .B2(n20043), .ZN(n20010) );
  OAI211_X1 U22874 ( .C1(n20232), .C2(n20077), .A(n20011), .B(n20010), .ZN(
        P1_U3033) );
  AOI22_X1 U22875 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20036), .B1(DATAI_17_), 
        .B2(n20037), .ZN(n20538) );
  AOI22_X1 U22876 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20036), .B1(DATAI_25_), 
        .B2(n20037), .ZN(n20637) );
  NAND2_X1 U22877 ( .A1(n20039), .A2(n11136), .ZN(n20632) );
  OAI22_X1 U22878 ( .A1(n20685), .A2(n20637), .B1(n20632), .B2(n20040), .ZN(
        n20012) );
  INV_X1 U22879 ( .A(n20012), .ZN(n20015) );
  NAND2_X1 U22880 ( .A1(n20013), .A2(n20051), .ZN(n20631) );
  INV_X1 U22881 ( .A(n20631), .ZN(n20245) );
  AOI22_X1 U22882 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20044), .B1(
        n20245), .B2(n20043), .ZN(n20014) );
  OAI211_X1 U22883 ( .C1(n20538), .C2(n20077), .A(n20015), .B(n20014), .ZN(
        P1_U3034) );
  AOI22_X1 U22884 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20036), .B1(DATAI_18_), 
        .B2(n20037), .ZN(n20543) );
  AOI22_X1 U22885 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20036), .B1(DATAI_26_), 
        .B2(n20037), .ZN(n20644) );
  NAND2_X1 U22886 ( .A1(n20039), .A2(n11123), .ZN(n20639) );
  OAI22_X1 U22887 ( .A1(n20685), .A2(n20644), .B1(n20639), .B2(n20040), .ZN(
        n20016) );
  INV_X1 U22888 ( .A(n20016), .ZN(n20019) );
  NAND2_X1 U22889 ( .A1(n20017), .A2(n20051), .ZN(n20638) );
  INV_X1 U22890 ( .A(n20638), .ZN(n20249) );
  AOI22_X1 U22891 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20044), .B1(
        n20249), .B2(n20043), .ZN(n20018) );
  OAI211_X1 U22892 ( .C1(n20543), .C2(n20077), .A(n20019), .B(n20018), .ZN(
        P1_U3035) );
  AOI22_X1 U22893 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20036), .B1(DATAI_19_), 
        .B2(n20037), .ZN(n20548) );
  NAND2_X1 U22894 ( .A1(n20039), .A2(n11120), .ZN(n20646) );
  OAI22_X1 U22895 ( .A1(n20685), .A2(n20651), .B1(n20646), .B2(n20040), .ZN(
        n20020) );
  INV_X1 U22896 ( .A(n20020), .ZN(n20023) );
  NAND2_X1 U22897 ( .A1(n20021), .A2(n20051), .ZN(n20645) );
  INV_X1 U22898 ( .A(n20645), .ZN(n20253) );
  AOI22_X1 U22899 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20044), .B1(
        n20253), .B2(n20043), .ZN(n20022) );
  OAI211_X1 U22900 ( .C1(n20548), .C2(n20077), .A(n20023), .B(n20022), .ZN(
        P1_U3036) );
  AOI22_X1 U22901 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20036), .B1(DATAI_28_), 
        .B2(n20037), .ZN(n20256) );
  NAND2_X1 U22902 ( .A1(n20039), .A2(n11046), .ZN(n20414) );
  OAI22_X1 U22903 ( .A1(n20685), .A2(n20256), .B1(n20414), .B2(n20040), .ZN(
        n20024) );
  INV_X1 U22904 ( .A(n20024), .ZN(n20027) );
  NOR2_X2 U22905 ( .A1(n20025), .A2(n20165), .ZN(n20653) );
  AOI22_X1 U22906 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20044), .B1(
        n20653), .B2(n20043), .ZN(n20026) );
  OAI211_X1 U22907 ( .C1(n20657), .C2(n20077), .A(n20027), .B(n20026), .ZN(
        P1_U3037) );
  AOI22_X1 U22908 ( .A1(DATAI_21_), .A2(n20037), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20036), .ZN(n20597) );
  AOI22_X1 U22909 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20036), .B1(DATAI_29_), 
        .B2(n20037), .ZN(n20667) );
  NAND2_X1 U22910 ( .A1(n20039), .A2(n11135), .ZN(n20418) );
  OAI22_X1 U22911 ( .A1(n20685), .A2(n20667), .B1(n20418), .B2(n20040), .ZN(
        n20028) );
  INV_X1 U22912 ( .A(n20028), .ZN(n20031) );
  NOR2_X2 U22913 ( .A1(n20029), .A2(n20165), .ZN(n20661) );
  AOI22_X1 U22914 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20044), .B1(
        n20661), .B2(n20043), .ZN(n20030) );
  OAI211_X1 U22915 ( .C1(n20597), .C2(n20077), .A(n20031), .B(n20030), .ZN(
        P1_U3038) );
  AOI22_X1 U22916 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20036), .B1(DATAI_22_), 
        .B2(n20037), .ZN(n20674) );
  AOI22_X1 U22917 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20036), .B1(DATAI_30_), 
        .B2(n20037), .ZN(n20468) );
  NAND2_X1 U22918 ( .A1(n20039), .A2(n11116), .ZN(n20669) );
  OAI22_X1 U22919 ( .A1(n20685), .A2(n20468), .B1(n20669), .B2(n20040), .ZN(
        n20032) );
  INV_X1 U22920 ( .A(n20032), .ZN(n20035) );
  NAND2_X1 U22921 ( .A1(n20033), .A2(n20051), .ZN(n20668) );
  INV_X1 U22922 ( .A(n20668), .ZN(n20264) );
  AOI22_X1 U22923 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20044), .B1(
        n20264), .B2(n20043), .ZN(n20034) );
  OAI211_X1 U22924 ( .C1(n20674), .C2(n20077), .A(n20035), .B(n20034), .ZN(
        P1_U3039) );
  AOI22_X1 U22925 ( .A1(DATAI_31_), .A2(n20037), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20036), .ZN(n20610) );
  NAND2_X1 U22926 ( .A1(n20039), .A2(n11129), .ZN(n20678) );
  OAI22_X1 U22927 ( .A1(n20685), .A2(n20610), .B1(n20678), .B2(n20040), .ZN(
        n20041) );
  INV_X1 U22928 ( .A(n20041), .ZN(n20046) );
  NAND2_X1 U22929 ( .A1(n20042), .A2(n20051), .ZN(n20675) );
  INV_X1 U22930 ( .A(n20675), .ZN(n20270) );
  AOI22_X1 U22931 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20044), .B1(
        n20270), .B2(n20043), .ZN(n20045) );
  OAI211_X1 U22932 ( .C1(n20686), .C2(n20077), .A(n20046), .B(n20045), .ZN(
        P1_U3040) );
  NOR2_X1 U22933 ( .A1(n13840), .A2(n12563), .ZN(n20362) );
  NOR2_X1 U22934 ( .A1(n20521), .A2(n20048), .ZN(n20069) );
  INV_X1 U22935 ( .A(n20069), .ZN(n20079) );
  OAI21_X1 U22936 ( .B1(n20047), .B2(n20522), .A(n20079), .ZN(n20052) );
  NAND2_X1 U22937 ( .A1(n20052), .A2(n20625), .ZN(n20050) );
  INV_X1 U22938 ( .A(n20048), .ZN(n20055) );
  NAND2_X1 U22939 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20055), .ZN(n20049) );
  NAND2_X1 U22940 ( .A1(n20050), .A2(n20049), .ZN(n20070) );
  AOI22_X1 U22941 ( .A1(n20618), .A2(n20070), .B1(n20617), .B2(n20069), .ZN(
        n20057) );
  OAI21_X1 U22942 ( .B1(n20323), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n20051), .ZN(n20519) );
  INV_X1 U22943 ( .A(n20121), .ZN(n20126) );
  INV_X1 U22944 ( .A(n20052), .ZN(n20053) );
  OAI211_X1 U22945 ( .C1(n20126), .C2(n20359), .A(n20625), .B(n20053), .ZN(
        n20054) );
  OAI211_X1 U22946 ( .C1(n20625), .C2(n20055), .A(n20624), .B(n20054), .ZN(
        n20082) );
  INV_X1 U22947 ( .A(n20077), .ZN(n20081) );
  INV_X1 U22948 ( .A(n20630), .ZN(n20530) );
  AOI22_X1 U22949 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20530), .ZN(n20056) );
  OAI211_X1 U22950 ( .C1(n20232), .C2(n20115), .A(n20057), .B(n20056), .ZN(
        P1_U3041) );
  INV_X1 U22951 ( .A(n20070), .ZN(n20078) );
  OAI22_X1 U22952 ( .A1(n20632), .A2(n20079), .B1(n20078), .B2(n20631), .ZN(
        n20058) );
  INV_X1 U22953 ( .A(n20058), .ZN(n20060) );
  INV_X1 U22954 ( .A(n20637), .ZN(n20535) );
  AOI22_X1 U22955 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20535), .ZN(n20059) );
  OAI211_X1 U22956 ( .C1(n20538), .C2(n20115), .A(n20060), .B(n20059), .ZN(
        P1_U3042) );
  OAI22_X1 U22957 ( .A1(n20639), .A2(n20079), .B1(n20078), .B2(n20638), .ZN(
        n20061) );
  INV_X1 U22958 ( .A(n20061), .ZN(n20063) );
  INV_X1 U22959 ( .A(n20644), .ZN(n20540) );
  AOI22_X1 U22960 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20540), .ZN(n20062) );
  OAI211_X1 U22961 ( .C1(n20543), .C2(n20115), .A(n20063), .B(n20062), .ZN(
        P1_U3043) );
  OAI22_X1 U22962 ( .A1(n20646), .A2(n20079), .B1(n20078), .B2(n20645), .ZN(
        n20064) );
  INV_X1 U22963 ( .A(n20064), .ZN(n20066) );
  INV_X1 U22964 ( .A(n20651), .ZN(n20545) );
  AOI22_X1 U22965 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20545), .ZN(n20065) );
  OAI211_X1 U22966 ( .C1(n20548), .C2(n20115), .A(n20066), .B(n20065), .ZN(
        P1_U3044) );
  AOI22_X1 U22967 ( .A1(n20653), .A2(n20070), .B1(n20652), .B2(n20069), .ZN(
        n20068) );
  INV_X1 U22968 ( .A(n20256), .ZN(n20654) );
  AOI22_X1 U22969 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20654), .ZN(n20067) );
  OAI211_X1 U22970 ( .C1(n20657), .C2(n20115), .A(n20068), .B(n20067), .ZN(
        P1_U3045) );
  AOI22_X1 U22971 ( .A1(n20661), .A2(n20070), .B1(n20659), .B2(n20069), .ZN(
        n20072) );
  INV_X1 U22972 ( .A(n20115), .ZN(n20074) );
  INV_X1 U22973 ( .A(n20597), .ZN(n20662) );
  AOI22_X1 U22974 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20082), .B1(
        n20074), .B2(n20662), .ZN(n20071) );
  OAI211_X1 U22975 ( .C1(n20667), .C2(n20077), .A(n20072), .B(n20071), .ZN(
        P1_U3046) );
  OAI22_X1 U22976 ( .A1(n20669), .A2(n20079), .B1(n20078), .B2(n20668), .ZN(
        n20073) );
  INV_X1 U22977 ( .A(n20073), .ZN(n20076) );
  INV_X1 U22978 ( .A(n20674), .ZN(n20508) );
  AOI22_X1 U22979 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20082), .B1(
        n20074), .B2(n20508), .ZN(n20075) );
  OAI211_X1 U22980 ( .C1(n20468), .C2(n20077), .A(n20076), .B(n20075), .ZN(
        P1_U3047) );
  OAI22_X1 U22981 ( .A1(n20678), .A2(n20079), .B1(n20078), .B2(n20675), .ZN(
        n20080) );
  INV_X1 U22982 ( .A(n20080), .ZN(n20084) );
  INV_X1 U22983 ( .A(n20610), .ZN(n20680) );
  AOI22_X1 U22984 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20082), .B1(
        n20081), .B2(n20680), .ZN(n20083) );
  OAI211_X1 U22985 ( .C1(n20686), .C2(n20115), .A(n20084), .B(n20083), .ZN(
        P1_U3048) );
  NAND3_X1 U22986 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20435), .A3(
        n20394), .ZN(n20129) );
  NOR2_X1 U22987 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20129), .ZN(
        n20087) );
  INV_X1 U22988 ( .A(n20087), .ZN(n20114) );
  OAI22_X1 U22989 ( .A1(n20151), .A2(n20232), .B1(n20395), .B2(n20114), .ZN(
        n20085) );
  INV_X1 U22990 ( .A(n20085), .ZN(n20095) );
  NAND2_X1 U22991 ( .A1(n20151), .A2(n20115), .ZN(n20086) );
  AOI21_X1 U22992 ( .B1(n20086), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20567), 
        .ZN(n20090) );
  NAND2_X1 U22993 ( .A1(n20125), .A2(n20565), .ZN(n20092) );
  NOR2_X1 U22994 ( .A1(n20087), .A2(n20323), .ZN(n20088) );
  AOI21_X1 U22995 ( .B1(n20090), .B2(n20092), .A(n20088), .ZN(n20089) );
  OAI21_X1 U22996 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20392), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20235) );
  NAND3_X1 U22997 ( .A1(n20402), .A2(n20089), .A3(n20235), .ZN(n20118) );
  INV_X1 U22998 ( .A(n20090), .ZN(n20093) );
  NAND2_X1 U22999 ( .A1(n20091), .A2(n20435), .ZN(n20239) );
  OAI22_X1 U23000 ( .A1(n20093), .A2(n20092), .B1(n20164), .B2(n20239), .ZN(
        n20117) );
  AOI22_X1 U23001 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20118), .B1(
        n20618), .B2(n20117), .ZN(n20094) );
  OAI211_X1 U23002 ( .C1(n20630), .C2(n20115), .A(n20095), .B(n20094), .ZN(
        P1_U3049) );
  OAI22_X1 U23003 ( .A1(n20115), .A2(n20637), .B1(n20114), .B2(n20632), .ZN(
        n20096) );
  INV_X1 U23004 ( .A(n20096), .ZN(n20098) );
  AOI22_X1 U23005 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20118), .B1(
        n20245), .B2(n20117), .ZN(n20097) );
  OAI211_X1 U23006 ( .C1(n20538), .C2(n20151), .A(n20098), .B(n20097), .ZN(
        P1_U3050) );
  OAI22_X1 U23007 ( .A1(n20151), .A2(n20543), .B1(n20114), .B2(n20639), .ZN(
        n20099) );
  INV_X1 U23008 ( .A(n20099), .ZN(n20101) );
  AOI22_X1 U23009 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20118), .B1(
        n20249), .B2(n20117), .ZN(n20100) );
  OAI211_X1 U23010 ( .C1(n20644), .C2(n20115), .A(n20101), .B(n20100), .ZN(
        P1_U3051) );
  OAI22_X1 U23011 ( .A1(n20151), .A2(n20548), .B1(n20114), .B2(n20646), .ZN(
        n20102) );
  INV_X1 U23012 ( .A(n20102), .ZN(n20104) );
  AOI22_X1 U23013 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20118), .B1(
        n20253), .B2(n20117), .ZN(n20103) );
  OAI211_X1 U23014 ( .C1(n20651), .C2(n20115), .A(n20104), .B(n20103), .ZN(
        P1_U3052) );
  OAI22_X1 U23015 ( .A1(n20115), .A2(n20256), .B1(n20114), .B2(n20414), .ZN(
        n20105) );
  INV_X1 U23016 ( .A(n20105), .ZN(n20107) );
  AOI22_X1 U23017 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20118), .B1(
        n20653), .B2(n20117), .ZN(n20106) );
  OAI211_X1 U23018 ( .C1(n20657), .C2(n20151), .A(n20107), .B(n20106), .ZN(
        P1_U3053) );
  OAI22_X1 U23019 ( .A1(n20115), .A2(n20667), .B1(n20114), .B2(n20418), .ZN(
        n20108) );
  INV_X1 U23020 ( .A(n20108), .ZN(n20110) );
  AOI22_X1 U23021 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20118), .B1(
        n20661), .B2(n20117), .ZN(n20109) );
  OAI211_X1 U23022 ( .C1(n20597), .C2(n20151), .A(n20110), .B(n20109), .ZN(
        P1_U3054) );
  OAI22_X1 U23023 ( .A1(n20151), .A2(n20674), .B1(n20114), .B2(n20669), .ZN(
        n20111) );
  INV_X1 U23024 ( .A(n20111), .ZN(n20113) );
  AOI22_X1 U23025 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20118), .B1(
        n20264), .B2(n20117), .ZN(n20112) );
  OAI211_X1 U23026 ( .C1(n20468), .C2(n20115), .A(n20113), .B(n20112), .ZN(
        P1_U3055) );
  OAI22_X1 U23027 ( .A1(n20115), .A2(n20610), .B1(n20114), .B2(n20678), .ZN(
        n20116) );
  INV_X1 U23028 ( .A(n20116), .ZN(n20120) );
  AOI22_X1 U23029 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20118), .B1(
        n20270), .B2(n20117), .ZN(n20119) );
  OAI211_X1 U23030 ( .C1(n20686), .C2(n20151), .A(n20120), .B(n20119), .ZN(
        P1_U3056) );
  NOR2_X1 U23031 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20434), .ZN(
        n20144) );
  INV_X1 U23032 ( .A(n20144), .ZN(n20150) );
  OAI22_X1 U23033 ( .A1(n20151), .A2(n20630), .B1(n20395), .B2(n20150), .ZN(
        n20122) );
  INV_X1 U23034 ( .A(n20122), .ZN(n20133) );
  AND2_X1 U23035 ( .A1(n20124), .A2(n20123), .ZN(n20611) );
  AOI21_X1 U23036 ( .B1(n20125), .B2(n20611), .A(n20144), .ZN(n20131) );
  AOI21_X1 U23037 ( .B1(n20126), .B2(n20625), .A(n20621), .ZN(n20130) );
  INV_X1 U23038 ( .A(n20130), .ZN(n20127) );
  AOI22_X1 U23039 ( .A1(n20131), .A2(n20127), .B1(n20567), .B2(n20129), .ZN(
        n20128) );
  NAND2_X1 U23040 ( .A1(n20624), .A2(n20128), .ZN(n20154) );
  OAI22_X1 U23041 ( .A1(n20131), .A2(n20130), .B1(n20689), .B2(n20129), .ZN(
        n20153) );
  AOI22_X1 U23042 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20154), .B1(
        n20618), .B2(n20153), .ZN(n20132) );
  OAI211_X1 U23043 ( .C1(n20232), .C2(n20187), .A(n20133), .B(n20132), .ZN(
        P1_U3057) );
  INV_X1 U23044 ( .A(n20538), .ZN(n20634) );
  INV_X1 U23045 ( .A(n20632), .ZN(n20492) );
  AOI22_X1 U23046 ( .A1(n20191), .A2(n20634), .B1(n20492), .B2(n20144), .ZN(
        n20135) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20154), .B1(
        n20245), .B2(n20153), .ZN(n20134) );
  OAI211_X1 U23048 ( .C1(n20637), .C2(n20151), .A(n20135), .B(n20134), .ZN(
        P1_U3058) );
  OAI22_X1 U23049 ( .A1(n20151), .A2(n20644), .B1(n20639), .B2(n20150), .ZN(
        n20136) );
  INV_X1 U23050 ( .A(n20136), .ZN(n20138) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20154), .B1(
        n20249), .B2(n20153), .ZN(n20137) );
  OAI211_X1 U23052 ( .C1(n20543), .C2(n20187), .A(n20138), .B(n20137), .ZN(
        P1_U3059) );
  INV_X1 U23053 ( .A(n20548), .ZN(n20648) );
  INV_X1 U23054 ( .A(n20646), .ZN(n20498) );
  AOI22_X1 U23055 ( .A1(n20191), .A2(n20648), .B1(n20498), .B2(n20144), .ZN(
        n20140) );
  AOI22_X1 U23056 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20154), .B1(
        n20253), .B2(n20153), .ZN(n20139) );
  OAI211_X1 U23057 ( .C1(n20651), .C2(n20151), .A(n20140), .B(n20139), .ZN(
        P1_U3060) );
  OAI22_X1 U23058 ( .A1(n20151), .A2(n20256), .B1(n20150), .B2(n20414), .ZN(
        n20141) );
  INV_X1 U23059 ( .A(n20141), .ZN(n20143) );
  AOI22_X1 U23060 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20154), .B1(
        n20653), .B2(n20153), .ZN(n20142) );
  OAI211_X1 U23061 ( .C1(n20657), .C2(n20187), .A(n20143), .B(n20142), .ZN(
        P1_U3061) );
  AOI22_X1 U23062 ( .A1(n20191), .A2(n20662), .B1(n20659), .B2(n20144), .ZN(
        n20146) );
  AOI22_X1 U23063 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20154), .B1(
        n20661), .B2(n20153), .ZN(n20145) );
  OAI211_X1 U23064 ( .C1(n20667), .C2(n20151), .A(n20146), .B(n20145), .ZN(
        P1_U3062) );
  OAI22_X1 U23065 ( .A1(n20151), .A2(n20468), .B1(n20669), .B2(n20150), .ZN(
        n20147) );
  INV_X1 U23066 ( .A(n20147), .ZN(n20149) );
  AOI22_X1 U23067 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20154), .B1(
        n20264), .B2(n20153), .ZN(n20148) );
  OAI211_X1 U23068 ( .C1(n20674), .C2(n20187), .A(n20149), .B(n20148), .ZN(
        P1_U3063) );
  OAI22_X1 U23069 ( .A1(n20151), .A2(n20610), .B1(n20150), .B2(n20678), .ZN(
        n20152) );
  INV_X1 U23070 ( .A(n20152), .ZN(n20156) );
  AOI22_X1 U23071 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20154), .B1(
        n20270), .B2(n20153), .ZN(n20155) );
  OAI211_X1 U23072 ( .C1(n20686), .C2(n20187), .A(n20156), .B(n20155), .ZN(
        P1_U3064) );
  NOR2_X1 U23073 ( .A1(n13583), .A2(n20157), .ZN(n20275) );
  NAND3_X1 U23074 ( .A1(n20275), .A2(n20625), .A3(n20315), .ZN(n20161) );
  INV_X1 U23075 ( .A(n20158), .ZN(n20159) );
  NAND2_X1 U23076 ( .A1(n20159), .A2(n20568), .ZN(n20160) );
  NAND2_X1 U23077 ( .A1(n20161), .A2(n20160), .ZN(n20181) );
  NAND3_X1 U23078 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20435), .A3(
        n20482), .ZN(n20196) );
  NOR2_X1 U23079 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20196), .ZN(
        n20180) );
  AOI22_X1 U23080 ( .A1(n20618), .A2(n20181), .B1(n20617), .B2(n20180), .ZN(
        n20168) );
  INV_X1 U23081 ( .A(n20275), .ZN(n20163) );
  OAI21_X1 U23082 ( .B1(n20191), .B2(n20214), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20162) );
  OAI21_X1 U23083 ( .B1(n20565), .B2(n20163), .A(n20162), .ZN(n20166) );
  INV_X1 U23084 ( .A(n20164), .ZN(n20393) );
  NOR2_X1 U23085 ( .A1(n20393), .A2(n20165), .ZN(n20577) );
  OAI221_X1 U23086 ( .B1(n20180), .B2(n20323), .C1(n20180), .C2(n20166), .A(
        n20577), .ZN(n20192) );
  INV_X1 U23087 ( .A(n20232), .ZN(n20627) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20192), .B1(
        n20214), .B2(n20627), .ZN(n20167) );
  OAI211_X1 U23089 ( .C1(n20630), .C2(n20187), .A(n20168), .B(n20167), .ZN(
        P1_U3065) );
  INV_X1 U23090 ( .A(n20180), .ZN(n20189) );
  INV_X1 U23091 ( .A(n20181), .ZN(n20188) );
  OAI22_X1 U23092 ( .A1(n20632), .A2(n20189), .B1(n20188), .B2(n20631), .ZN(
        n20169) );
  INV_X1 U23093 ( .A(n20169), .ZN(n20171) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20192), .B1(
        n20191), .B2(n20535), .ZN(n20170) );
  OAI211_X1 U23095 ( .C1(n20538), .C2(n20231), .A(n20171), .B(n20170), .ZN(
        P1_U3066) );
  OAI22_X1 U23096 ( .A1(n20639), .A2(n20189), .B1(n20188), .B2(n20638), .ZN(
        n20172) );
  INV_X1 U23097 ( .A(n20172), .ZN(n20174) );
  INV_X1 U23098 ( .A(n20543), .ZN(n20641) );
  AOI22_X1 U23099 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20192), .B1(
        n20214), .B2(n20641), .ZN(n20173) );
  OAI211_X1 U23100 ( .C1(n20644), .C2(n20187), .A(n20174), .B(n20173), .ZN(
        P1_U3067) );
  OAI22_X1 U23101 ( .A1(n20646), .A2(n20189), .B1(n20188), .B2(n20645), .ZN(
        n20175) );
  INV_X1 U23102 ( .A(n20175), .ZN(n20177) );
  AOI22_X1 U23103 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20192), .B1(
        n20214), .B2(n20648), .ZN(n20176) );
  OAI211_X1 U23104 ( .C1(n20651), .C2(n20187), .A(n20177), .B(n20176), .ZN(
        P1_U3068) );
  AOI22_X1 U23105 ( .A1(n20653), .A2(n20181), .B1(n20652), .B2(n20180), .ZN(
        n20179) );
  AOI22_X1 U23106 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20192), .B1(
        n20191), .B2(n20654), .ZN(n20178) );
  OAI211_X1 U23107 ( .C1(n20657), .C2(n20231), .A(n20179), .B(n20178), .ZN(
        P1_U3069) );
  AOI22_X1 U23108 ( .A1(n20661), .A2(n20181), .B1(n20659), .B2(n20180), .ZN(
        n20183) );
  INV_X1 U23109 ( .A(n20667), .ZN(n20594) );
  AOI22_X1 U23110 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20192), .B1(
        n20191), .B2(n20594), .ZN(n20182) );
  OAI211_X1 U23111 ( .C1(n20597), .C2(n20231), .A(n20183), .B(n20182), .ZN(
        P1_U3070) );
  OAI22_X1 U23112 ( .A1(n20669), .A2(n20189), .B1(n20188), .B2(n20668), .ZN(
        n20184) );
  INV_X1 U23113 ( .A(n20184), .ZN(n20186) );
  AOI22_X1 U23114 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20192), .B1(
        n20214), .B2(n20508), .ZN(n20185) );
  OAI211_X1 U23115 ( .C1(n20468), .C2(n20187), .A(n20186), .B(n20185), .ZN(
        P1_U3071) );
  OAI22_X1 U23116 ( .A1(n20678), .A2(n20189), .B1(n20188), .B2(n20675), .ZN(
        n20190) );
  INV_X1 U23117 ( .A(n20190), .ZN(n20194) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20192), .B1(
        n20191), .B2(n20680), .ZN(n20193) );
  OAI211_X1 U23119 ( .C1(n20686), .C2(n20231), .A(n20194), .B(n20193), .ZN(
        P1_U3072) );
  INV_X1 U23120 ( .A(n20522), .ZN(n20352) );
  NAND2_X1 U23121 ( .A1(n20275), .A2(n20352), .ZN(n20195) );
  NOR2_X1 U23122 ( .A1(n20521), .A2(n20196), .ZN(n20217) );
  INV_X1 U23123 ( .A(n20217), .ZN(n20225) );
  NAND2_X1 U23124 ( .A1(n20195), .A2(n20225), .ZN(n20199) );
  NAND2_X1 U23125 ( .A1(n20199), .A2(n20625), .ZN(n20198) );
  INV_X1 U23126 ( .A(n20196), .ZN(n20202) );
  NAND2_X1 U23127 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20202), .ZN(n20197) );
  NAND2_X1 U23128 ( .A1(n20198), .A2(n20197), .ZN(n20218) );
  AOI22_X1 U23129 ( .A1(n20618), .A2(n20218), .B1(n20617), .B2(n20217), .ZN(
        n20204) );
  INV_X1 U23130 ( .A(n20199), .ZN(n20200) );
  OAI211_X1 U23131 ( .C1(n20283), .C2(n20359), .A(n20625), .B(n20200), .ZN(
        n20201) );
  OAI211_X1 U23132 ( .C1(n20625), .C2(n20202), .A(n20624), .B(n20201), .ZN(
        n20228) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20228), .B1(
        n20214), .B2(n20530), .ZN(n20203) );
  OAI211_X1 U23134 ( .C1(n20232), .C2(n20274), .A(n20204), .B(n20203), .ZN(
        P1_U3073) );
  INV_X1 U23135 ( .A(n20218), .ZN(n20224) );
  OAI22_X1 U23136 ( .A1(n20632), .A2(n20225), .B1(n20224), .B2(n20631), .ZN(
        n20205) );
  INV_X1 U23137 ( .A(n20205), .ZN(n20207) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20228), .B1(
        n20214), .B2(n20535), .ZN(n20206) );
  OAI211_X1 U23139 ( .C1(n20538), .C2(n20274), .A(n20207), .B(n20206), .ZN(
        P1_U3074) );
  OAI22_X1 U23140 ( .A1(n20639), .A2(n20225), .B1(n20224), .B2(n20638), .ZN(
        n20208) );
  INV_X1 U23141 ( .A(n20208), .ZN(n20210) );
  AOI22_X1 U23142 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20228), .B1(
        n20214), .B2(n20540), .ZN(n20209) );
  OAI211_X1 U23143 ( .C1(n20543), .C2(n20274), .A(n20210), .B(n20209), .ZN(
        P1_U3075) );
  OAI22_X1 U23144 ( .A1(n20646), .A2(n20225), .B1(n20224), .B2(n20645), .ZN(
        n20211) );
  INV_X1 U23145 ( .A(n20211), .ZN(n20213) );
  INV_X1 U23146 ( .A(n20274), .ZN(n20227) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20228), .B1(
        n20227), .B2(n20648), .ZN(n20212) );
  OAI211_X1 U23148 ( .C1(n20651), .C2(n20231), .A(n20213), .B(n20212), .ZN(
        P1_U3076) );
  AOI22_X1 U23149 ( .A1(n20653), .A2(n20218), .B1(n20652), .B2(n20217), .ZN(
        n20216) );
  AOI22_X1 U23150 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20228), .B1(
        n20214), .B2(n20654), .ZN(n20215) );
  OAI211_X1 U23151 ( .C1(n20657), .C2(n20274), .A(n20216), .B(n20215), .ZN(
        P1_U3077) );
  AOI22_X1 U23152 ( .A1(n20661), .A2(n20218), .B1(n20659), .B2(n20217), .ZN(
        n20220) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20228), .B1(
        n20227), .B2(n20662), .ZN(n20219) );
  OAI211_X1 U23154 ( .C1(n20667), .C2(n20231), .A(n20220), .B(n20219), .ZN(
        P1_U3078) );
  OAI22_X1 U23155 ( .A1(n20669), .A2(n20225), .B1(n20224), .B2(n20668), .ZN(
        n20221) );
  INV_X1 U23156 ( .A(n20221), .ZN(n20223) );
  AOI22_X1 U23157 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20228), .B1(
        n20227), .B2(n20508), .ZN(n20222) );
  OAI211_X1 U23158 ( .C1(n20468), .C2(n20231), .A(n20223), .B(n20222), .ZN(
        P1_U3079) );
  OAI22_X1 U23159 ( .A1(n20678), .A2(n20225), .B1(n20224), .B2(n20675), .ZN(
        n20226) );
  INV_X1 U23160 ( .A(n20226), .ZN(n20230) );
  INV_X1 U23161 ( .A(n20686), .ZN(n20605) );
  AOI22_X1 U23162 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20228), .B1(
        n20227), .B2(n20605), .ZN(n20229) );
  OAI211_X1 U23163 ( .C1(n20610), .C2(n20231), .A(n20230), .B(n20229), .ZN(
        P1_U3080) );
  INV_X1 U23164 ( .A(n20285), .ZN(n20278) );
  OR2_X1 U23165 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20278), .ZN(
        n20267) );
  OAI22_X1 U23166 ( .A1(n20313), .A2(n20232), .B1(n20395), .B2(n20267), .ZN(
        n20233) );
  INV_X1 U23167 ( .A(n20233), .ZN(n20243) );
  NAND3_X1 U23168 ( .A1(n20313), .A2(n20274), .A3(n20625), .ZN(n20234) );
  NAND2_X1 U23169 ( .A1(n20234), .A2(n20479), .ZN(n20237) );
  NAND2_X1 U23170 ( .A1(n20275), .A2(n20565), .ZN(n20240) );
  AOI22_X1 U23171 ( .A1(n20237), .A2(n20240), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20267), .ZN(n20236) );
  NAND3_X1 U23172 ( .A1(n20577), .A2(n20236), .A3(n20235), .ZN(n20271) );
  INV_X1 U23173 ( .A(n20237), .ZN(n20241) );
  INV_X1 U23174 ( .A(n20568), .ZN(n20238) );
  OAI22_X1 U23175 ( .A1(n20241), .A2(n20240), .B1(n20239), .B2(n20238), .ZN(
        n20269) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20271), .B1(
        n20618), .B2(n20269), .ZN(n20242) );
  OAI211_X1 U23177 ( .C1(n20630), .C2(n20274), .A(n20243), .B(n20242), .ZN(
        P1_U3081) );
  OAI22_X1 U23178 ( .A1(n20313), .A2(n20538), .B1(n20632), .B2(n20267), .ZN(
        n20244) );
  INV_X1 U23179 ( .A(n20244), .ZN(n20247) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20271), .B1(
        n20245), .B2(n20269), .ZN(n20246) );
  OAI211_X1 U23181 ( .C1(n20637), .C2(n20274), .A(n20247), .B(n20246), .ZN(
        P1_U3082) );
  OAI22_X1 U23182 ( .A1(n20313), .A2(n20543), .B1(n20639), .B2(n20267), .ZN(
        n20248) );
  INV_X1 U23183 ( .A(n20248), .ZN(n20251) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20271), .B1(
        n20249), .B2(n20269), .ZN(n20250) );
  OAI211_X1 U23185 ( .C1(n20644), .C2(n20274), .A(n20251), .B(n20250), .ZN(
        P1_U3083) );
  OAI22_X1 U23186 ( .A1(n20274), .A2(n20651), .B1(n20646), .B2(n20267), .ZN(
        n20252) );
  INV_X1 U23187 ( .A(n20252), .ZN(n20255) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20271), .B1(
        n20253), .B2(n20269), .ZN(n20254) );
  OAI211_X1 U23189 ( .C1(n20548), .C2(n20313), .A(n20255), .B(n20254), .ZN(
        P1_U3084) );
  OAI22_X1 U23190 ( .A1(n20274), .A2(n20256), .B1(n20414), .B2(n20267), .ZN(
        n20257) );
  INV_X1 U23191 ( .A(n20257), .ZN(n20259) );
  AOI22_X1 U23192 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20271), .B1(
        n20653), .B2(n20269), .ZN(n20258) );
  OAI211_X1 U23193 ( .C1(n20657), .C2(n20313), .A(n20259), .B(n20258), .ZN(
        P1_U3085) );
  OAI22_X1 U23194 ( .A1(n20313), .A2(n20597), .B1(n20418), .B2(n20267), .ZN(
        n20260) );
  INV_X1 U23195 ( .A(n20260), .ZN(n20262) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20271), .B1(
        n20661), .B2(n20269), .ZN(n20261) );
  OAI211_X1 U23197 ( .C1(n20667), .C2(n20274), .A(n20262), .B(n20261), .ZN(
        P1_U3086) );
  OAI22_X1 U23198 ( .A1(n20274), .A2(n20468), .B1(n20669), .B2(n20267), .ZN(
        n20263) );
  INV_X1 U23199 ( .A(n20263), .ZN(n20266) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20271), .B1(
        n20264), .B2(n20269), .ZN(n20265) );
  OAI211_X1 U23201 ( .C1(n20674), .C2(n20313), .A(n20266), .B(n20265), .ZN(
        P1_U3087) );
  OAI22_X1 U23202 ( .A1(n20313), .A2(n20686), .B1(n20678), .B2(n20267), .ZN(
        n20268) );
  INV_X1 U23203 ( .A(n20268), .ZN(n20273) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20269), .ZN(n20272) );
  OAI211_X1 U23205 ( .C1(n20610), .C2(n20274), .A(n20273), .B(n20272), .ZN(
        P1_U3088) );
  NAND2_X1 U23206 ( .A1(n20275), .A2(n20611), .ZN(n20277) );
  INV_X1 U23207 ( .A(n20276), .ZN(n20300) );
  NAND2_X1 U23208 ( .A1(n20277), .A2(n20276), .ZN(n20281) );
  NAND2_X1 U23209 ( .A1(n20281), .A2(n20625), .ZN(n20280) );
  NAND2_X1 U23210 ( .A1(n20285), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20279) );
  NAND2_X1 U23211 ( .A1(n20280), .A2(n20279), .ZN(n20301) );
  AOI22_X1 U23212 ( .A1(n20618), .A2(n20301), .B1(n20617), .B2(n20300), .ZN(
        n20288) );
  INV_X1 U23213 ( .A(n20281), .ZN(n20282) );
  OAI211_X1 U23214 ( .C1(n20283), .C2(n20621), .A(n20625), .B(n20282), .ZN(
        n20284) );
  OAI211_X1 U23215 ( .C1(n20285), .C2(n20625), .A(n20624), .B(n20284), .ZN(
        n20310) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20310), .B1(
        n20348), .B2(n20627), .ZN(n20287) );
  OAI211_X1 U23217 ( .C1(n20630), .C2(n20313), .A(n20288), .B(n20287), .ZN(
        P1_U3089) );
  INV_X1 U23218 ( .A(n20301), .ZN(n20308) );
  OAI22_X1 U23219 ( .A1(n20632), .A2(n20276), .B1(n20308), .B2(n20631), .ZN(
        n20289) );
  INV_X1 U23220 ( .A(n20289), .ZN(n20291) );
  INV_X1 U23221 ( .A(n20313), .ZN(n20305) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20310), .B1(
        n20305), .B2(n20535), .ZN(n20290) );
  OAI211_X1 U23223 ( .C1(n20538), .C2(n20335), .A(n20291), .B(n20290), .ZN(
        P1_U3090) );
  OAI22_X1 U23224 ( .A1(n20639), .A2(n20276), .B1(n20308), .B2(n20638), .ZN(
        n20292) );
  INV_X1 U23225 ( .A(n20292), .ZN(n20294) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20310), .B1(
        n20305), .B2(n20540), .ZN(n20293) );
  OAI211_X1 U23227 ( .C1(n20543), .C2(n20335), .A(n20294), .B(n20293), .ZN(
        P1_U3091) );
  OAI22_X1 U23228 ( .A1(n20646), .A2(n20276), .B1(n20308), .B2(n20645), .ZN(
        n20295) );
  INV_X1 U23229 ( .A(n20295), .ZN(n20297) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20310), .B1(
        n20305), .B2(n20545), .ZN(n20296) );
  OAI211_X1 U23231 ( .C1(n20548), .C2(n20335), .A(n20297), .B(n20296), .ZN(
        P1_U3092) );
  AOI22_X1 U23232 ( .A1(n20653), .A2(n20301), .B1(n20652), .B2(n20300), .ZN(
        n20299) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20310), .B1(
        n20305), .B2(n20654), .ZN(n20298) );
  OAI211_X1 U23234 ( .C1(n20657), .C2(n20335), .A(n20299), .B(n20298), .ZN(
        P1_U3093) );
  AOI22_X1 U23235 ( .A1(n20661), .A2(n20301), .B1(n20659), .B2(n20300), .ZN(
        n20303) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20310), .B1(
        n20305), .B2(n20594), .ZN(n20302) );
  OAI211_X1 U23237 ( .C1(n20597), .C2(n20335), .A(n20303), .B(n20302), .ZN(
        P1_U3094) );
  OAI22_X1 U23238 ( .A1(n20669), .A2(n20276), .B1(n20308), .B2(n20668), .ZN(
        n20304) );
  INV_X1 U23239 ( .A(n20304), .ZN(n20307) );
  INV_X1 U23240 ( .A(n20468), .ZN(n20671) );
  AOI22_X1 U23241 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20310), .B1(
        n20305), .B2(n20671), .ZN(n20306) );
  OAI211_X1 U23242 ( .C1(n20674), .C2(n20335), .A(n20307), .B(n20306), .ZN(
        P1_U3095) );
  OAI22_X1 U23243 ( .A1(n20678), .A2(n20276), .B1(n20308), .B2(n20675), .ZN(
        n20309) );
  INV_X1 U23244 ( .A(n20309), .ZN(n20312) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20310), .B1(
        n20348), .B2(n20605), .ZN(n20311) );
  OAI211_X1 U23246 ( .C1(n20610), .C2(n20313), .A(n20312), .B(n20311), .ZN(
        P1_U3096) );
  AND2_X1 U23247 ( .A1(n20314), .A2(n13583), .ZN(n20433) );
  NAND3_X1 U23248 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20394), .A3(
        n20482), .ZN(n20354) );
  NOR2_X1 U23249 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20354), .ZN(
        n20338) );
  AOI21_X1 U23250 ( .B1(n20433), .B2(n20315), .A(n20338), .ZN(n20320) );
  OR2_X1 U23251 ( .A1(n20320), .A2(n20567), .ZN(n20318) );
  AND2_X1 U23252 ( .A1(n20316), .A2(n20392), .ZN(n20488) );
  NAND2_X1 U23253 ( .A1(n20488), .A2(n20393), .ZN(n20317) );
  NAND2_X1 U23254 ( .A1(n20318), .A2(n20317), .ZN(n20339) );
  AOI22_X1 U23255 ( .A1(n20618), .A2(n20339), .B1(n20617), .B2(n20338), .ZN(
        n20325) );
  NAND2_X1 U23256 ( .A1(n20446), .A2(n20319), .ZN(n20383) );
  OAI21_X1 U23257 ( .B1(n20387), .B2(n20348), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20321) );
  NAND2_X1 U23258 ( .A1(n20321), .A2(n20320), .ZN(n20322) );
  OAI211_X1 U23259 ( .C1(n20338), .C2(n20323), .A(n20402), .B(n20322), .ZN(
        n20349) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20349), .B1(
        n20387), .B2(n20627), .ZN(n20324) );
  OAI211_X1 U23261 ( .C1(n20630), .C2(n20335), .A(n20325), .B(n20324), .ZN(
        P1_U3097) );
  INV_X1 U23262 ( .A(n20338), .ZN(n20346) );
  INV_X1 U23263 ( .A(n20339), .ZN(n20345) );
  OAI22_X1 U23264 ( .A1(n20632), .A2(n20346), .B1(n20345), .B2(n20631), .ZN(
        n20326) );
  INV_X1 U23265 ( .A(n20326), .ZN(n20328) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20349), .B1(
        n20387), .B2(n20634), .ZN(n20327) );
  OAI211_X1 U23267 ( .C1(n20637), .C2(n20335), .A(n20328), .B(n20327), .ZN(
        P1_U3098) );
  OAI22_X1 U23268 ( .A1(n20639), .A2(n20346), .B1(n20345), .B2(n20638), .ZN(
        n20329) );
  INV_X1 U23269 ( .A(n20329), .ZN(n20331) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20349), .B1(
        n20387), .B2(n20641), .ZN(n20330) );
  OAI211_X1 U23271 ( .C1(n20644), .C2(n20335), .A(n20331), .B(n20330), .ZN(
        P1_U3099) );
  OAI22_X1 U23272 ( .A1(n20646), .A2(n20346), .B1(n20345), .B2(n20645), .ZN(
        n20332) );
  INV_X1 U23273 ( .A(n20332), .ZN(n20334) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20349), .B1(
        n20387), .B2(n20648), .ZN(n20333) );
  OAI211_X1 U23275 ( .C1(n20651), .C2(n20335), .A(n20334), .B(n20333), .ZN(
        P1_U3100) );
  AOI22_X1 U23276 ( .A1(n20653), .A2(n20339), .B1(n20652), .B2(n20338), .ZN(
        n20337) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20654), .ZN(n20336) );
  OAI211_X1 U23278 ( .C1(n20657), .C2(n20383), .A(n20337), .B(n20336), .ZN(
        P1_U3101) );
  AOI22_X1 U23279 ( .A1(n20661), .A2(n20339), .B1(n20659), .B2(n20338), .ZN(
        n20341) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20594), .ZN(n20340) );
  OAI211_X1 U23281 ( .C1(n20597), .C2(n20383), .A(n20341), .B(n20340), .ZN(
        P1_U3102) );
  OAI22_X1 U23282 ( .A1(n20669), .A2(n20346), .B1(n20345), .B2(n20668), .ZN(
        n20342) );
  INV_X1 U23283 ( .A(n20342), .ZN(n20344) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20671), .ZN(n20343) );
  OAI211_X1 U23285 ( .C1(n20674), .C2(n20383), .A(n20344), .B(n20343), .ZN(
        P1_U3103) );
  OAI22_X1 U23286 ( .A1(n20678), .A2(n20346), .B1(n20345), .B2(n20675), .ZN(
        n20347) );
  INV_X1 U23287 ( .A(n20347), .ZN(n20351) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20349), .B1(
        n20348), .B2(n20680), .ZN(n20350) );
  OAI211_X1 U23289 ( .C1(n20686), .C2(n20383), .A(n20351), .B(n20350), .ZN(
        P1_U3104) );
  NAND2_X1 U23290 ( .A1(n20433), .A2(n20352), .ZN(n20353) );
  NOR2_X1 U23291 ( .A1(n20521), .A2(n20354), .ZN(n20376) );
  INV_X1 U23292 ( .A(n20376), .ZN(n20385) );
  NAND2_X1 U23293 ( .A1(n20353), .A2(n20385), .ZN(n20357) );
  NAND2_X1 U23294 ( .A1(n20357), .A2(n20625), .ZN(n20356) );
  INV_X1 U23295 ( .A(n20354), .ZN(n20361) );
  NAND2_X1 U23296 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20361), .ZN(n20355) );
  NAND2_X1 U23297 ( .A1(n20356), .A2(n20355), .ZN(n20377) );
  AOI22_X1 U23298 ( .A1(n20618), .A2(n20377), .B1(n20617), .B2(n20376), .ZN(
        n20364) );
  INV_X1 U23299 ( .A(n20446), .ZN(n20442) );
  INV_X1 U23300 ( .A(n20357), .ZN(n20358) );
  OAI211_X1 U23301 ( .C1(n20442), .C2(n20359), .A(n20625), .B(n20358), .ZN(
        n20360) );
  OAI211_X1 U23302 ( .C1(n20625), .C2(n20361), .A(n20624), .B(n20360), .ZN(
        n20388) );
  NAND2_X1 U23303 ( .A1(n20446), .A2(n20362), .ZN(n20427) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20388), .B1(
        n20420), .B2(n20627), .ZN(n20363) );
  OAI211_X1 U23305 ( .C1(n20630), .C2(n20383), .A(n20364), .B(n20363), .ZN(
        P1_U3105) );
  INV_X1 U23306 ( .A(n20377), .ZN(n20384) );
  OAI22_X1 U23307 ( .A1(n20632), .A2(n20385), .B1(n20384), .B2(n20631), .ZN(
        n20365) );
  INV_X1 U23308 ( .A(n20365), .ZN(n20367) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20388), .B1(
        n20420), .B2(n20634), .ZN(n20366) );
  OAI211_X1 U23310 ( .C1(n20637), .C2(n20383), .A(n20367), .B(n20366), .ZN(
        P1_U3106) );
  OAI22_X1 U23311 ( .A1(n20639), .A2(n20385), .B1(n20384), .B2(n20638), .ZN(
        n20368) );
  INV_X1 U23312 ( .A(n20368), .ZN(n20370) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20388), .B1(
        n20420), .B2(n20641), .ZN(n20369) );
  OAI211_X1 U23314 ( .C1(n20644), .C2(n20383), .A(n20370), .B(n20369), .ZN(
        P1_U3107) );
  OAI22_X1 U23315 ( .A1(n20646), .A2(n20385), .B1(n20384), .B2(n20645), .ZN(
        n20371) );
  INV_X1 U23316 ( .A(n20371), .ZN(n20373) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20388), .B1(
        n20420), .B2(n20648), .ZN(n20372) );
  OAI211_X1 U23318 ( .C1(n20651), .C2(n20383), .A(n20373), .B(n20372), .ZN(
        P1_U3108) );
  AOI22_X1 U23319 ( .A1(n20653), .A2(n20377), .B1(n20652), .B2(n20376), .ZN(
        n20375) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20388), .B1(
        n20387), .B2(n20654), .ZN(n20374) );
  OAI211_X1 U23321 ( .C1(n20657), .C2(n20427), .A(n20375), .B(n20374), .ZN(
        P1_U3109) );
  AOI22_X1 U23322 ( .A1(n20661), .A2(n20377), .B1(n20659), .B2(n20376), .ZN(
        n20379) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20388), .B1(
        n20387), .B2(n20594), .ZN(n20378) );
  OAI211_X1 U23324 ( .C1(n20597), .C2(n20427), .A(n20379), .B(n20378), .ZN(
        P1_U3110) );
  OAI22_X1 U23325 ( .A1(n20669), .A2(n20385), .B1(n20384), .B2(n20668), .ZN(
        n20380) );
  INV_X1 U23326 ( .A(n20380), .ZN(n20382) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20388), .B1(
        n20420), .B2(n20508), .ZN(n20381) );
  OAI211_X1 U23328 ( .C1(n20468), .C2(n20383), .A(n20382), .B(n20381), .ZN(
        P1_U3111) );
  OAI22_X1 U23329 ( .A1(n20678), .A2(n20385), .B1(n20384), .B2(n20675), .ZN(
        n20386) );
  INV_X1 U23330 ( .A(n20386), .ZN(n20390) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20388), .B1(
        n20387), .B2(n20680), .ZN(n20389) );
  OAI211_X1 U23332 ( .C1(n20686), .C2(n20427), .A(n20390), .B(n20389), .ZN(
        P1_U3112) );
  NAND3_X1 U23333 ( .A1(n20467), .A2(n20427), .A3(n20625), .ZN(n20391) );
  NAND2_X1 U23334 ( .A1(n20391), .A2(n20479), .ZN(n20399) );
  AND2_X1 U23335 ( .A1(n20433), .A2(n20565), .ZN(n20397) );
  OR2_X1 U23336 ( .A1(n20392), .A2(n20435), .ZN(n20400) );
  INV_X1 U23337 ( .A(n20400), .ZN(n20569) );
  AOI22_X1 U23338 ( .A1(n20399), .A2(n20397), .B1(n20569), .B2(n20393), .ZN(
        n20432) );
  INV_X1 U23339 ( .A(n20618), .ZN(n20491) );
  NAND3_X1 U23340 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20394), .ZN(n20437) );
  OR2_X1 U23341 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20437), .ZN(
        n20426) );
  OAI22_X1 U23342 ( .A1(n20427), .A2(n20630), .B1(n20395), .B2(n20426), .ZN(
        n20396) );
  INV_X1 U23343 ( .A(n20396), .ZN(n20404) );
  INV_X1 U23344 ( .A(n20397), .ZN(n20398) );
  AOI22_X1 U23345 ( .A1(n20399), .A2(n20398), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20426), .ZN(n20401) );
  NAND2_X1 U23346 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20400), .ZN(n20576) );
  NAND3_X1 U23347 ( .A1(n20402), .A2(n20401), .A3(n20576), .ZN(n20429) );
  INV_X1 U23348 ( .A(n20467), .ZN(n20472) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20429), .B1(
        n20472), .B2(n20627), .ZN(n20403) );
  OAI211_X1 U23350 ( .C1(n20432), .C2(n20491), .A(n20404), .B(n20403), .ZN(
        P1_U3113) );
  OAI22_X1 U23351 ( .A1(n20467), .A2(n20538), .B1(n20632), .B2(n20426), .ZN(
        n20405) );
  INV_X1 U23352 ( .A(n20405), .ZN(n20407) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20429), .B1(
        n20420), .B2(n20535), .ZN(n20406) );
  OAI211_X1 U23354 ( .C1(n20432), .C2(n20631), .A(n20407), .B(n20406), .ZN(
        P1_U3114) );
  OAI22_X1 U23355 ( .A1(n20467), .A2(n20543), .B1(n20639), .B2(n20426), .ZN(
        n20408) );
  INV_X1 U23356 ( .A(n20408), .ZN(n20410) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20429), .B1(
        n20420), .B2(n20540), .ZN(n20409) );
  OAI211_X1 U23358 ( .C1(n20432), .C2(n20638), .A(n20410), .B(n20409), .ZN(
        P1_U3115) );
  OAI22_X1 U23359 ( .A1(n20467), .A2(n20548), .B1(n20646), .B2(n20426), .ZN(
        n20411) );
  INV_X1 U23360 ( .A(n20411), .ZN(n20413) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20429), .B1(
        n20420), .B2(n20545), .ZN(n20412) );
  OAI211_X1 U23362 ( .C1(n20432), .C2(n20645), .A(n20413), .B(n20412), .ZN(
        P1_U3116) );
  INV_X1 U23363 ( .A(n20653), .ZN(n20504) );
  OAI22_X1 U23364 ( .A1(n20467), .A2(n20657), .B1(n20414), .B2(n20426), .ZN(
        n20415) );
  INV_X1 U23365 ( .A(n20415), .ZN(n20417) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20429), .B1(
        n20420), .B2(n20654), .ZN(n20416) );
  OAI211_X1 U23367 ( .C1(n20432), .C2(n20504), .A(n20417), .B(n20416), .ZN(
        P1_U3117) );
  INV_X1 U23368 ( .A(n20661), .ZN(n20507) );
  OAI22_X1 U23369 ( .A1(n20467), .A2(n20597), .B1(n20418), .B2(n20426), .ZN(
        n20419) );
  INV_X1 U23370 ( .A(n20419), .ZN(n20422) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20429), .B1(
        n20420), .B2(n20594), .ZN(n20421) );
  OAI211_X1 U23372 ( .C1(n20432), .C2(n20507), .A(n20422), .B(n20421), .ZN(
        P1_U3118) );
  OAI22_X1 U23373 ( .A1(n20427), .A2(n20468), .B1(n20669), .B2(n20426), .ZN(
        n20423) );
  INV_X1 U23374 ( .A(n20423), .ZN(n20425) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20429), .B1(
        n20472), .B2(n20508), .ZN(n20424) );
  OAI211_X1 U23376 ( .C1(n20432), .C2(n20668), .A(n20425), .B(n20424), .ZN(
        P1_U3119) );
  OAI22_X1 U23377 ( .A1(n20427), .A2(n20610), .B1(n20678), .B2(n20426), .ZN(
        n20428) );
  INV_X1 U23378 ( .A(n20428), .ZN(n20431) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20429), .B1(
        n20472), .B2(n20605), .ZN(n20430) );
  OAI211_X1 U23380 ( .C1(n20432), .C2(n20675), .A(n20431), .B(n20430), .ZN(
        P1_U3120) );
  NAND2_X1 U23381 ( .A1(n20433), .A2(n20611), .ZN(n20436) );
  NOR2_X1 U23382 ( .A1(n20435), .A2(n20434), .ZN(n20460) );
  INV_X1 U23383 ( .A(n20460), .ZN(n20470) );
  NAND2_X1 U23384 ( .A1(n20436), .A2(n20470), .ZN(n20440) );
  NAND2_X1 U23385 ( .A1(n20440), .A2(n20625), .ZN(n20439) );
  INV_X1 U23386 ( .A(n20437), .ZN(n20444) );
  NAND2_X1 U23387 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20444), .ZN(n20438) );
  NAND2_X1 U23388 ( .A1(n20439), .A2(n20438), .ZN(n20461) );
  AOI22_X1 U23389 ( .A1(n20618), .A2(n20461), .B1(n20617), .B2(n20460), .ZN(
        n20448) );
  INV_X1 U23390 ( .A(n20440), .ZN(n20441) );
  OAI211_X1 U23391 ( .C1(n20442), .C2(n20621), .A(n20625), .B(n20441), .ZN(
        n20443) );
  OAI211_X1 U23392 ( .C1(n20625), .C2(n20444), .A(n20624), .B(n20443), .ZN(
        n20473) );
  NAND2_X1 U23393 ( .A1(n20446), .A2(n20445), .ZN(n20477) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20473), .B1(
        n20514), .B2(n20627), .ZN(n20447) );
  OAI211_X1 U23395 ( .C1(n20630), .C2(n20467), .A(n20448), .B(n20447), .ZN(
        P1_U3121) );
  INV_X1 U23396 ( .A(n20461), .ZN(n20469) );
  OAI22_X1 U23397 ( .A1(n20632), .A2(n20470), .B1(n20469), .B2(n20631), .ZN(
        n20449) );
  INV_X1 U23398 ( .A(n20449), .ZN(n20451) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20473), .B1(
        n20514), .B2(n20634), .ZN(n20450) );
  OAI211_X1 U23400 ( .C1(n20637), .C2(n20467), .A(n20451), .B(n20450), .ZN(
        P1_U3122) );
  OAI22_X1 U23401 ( .A1(n20639), .A2(n20470), .B1(n20469), .B2(n20638), .ZN(
        n20452) );
  INV_X1 U23402 ( .A(n20452), .ZN(n20454) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20473), .B1(
        n20514), .B2(n20641), .ZN(n20453) );
  OAI211_X1 U23404 ( .C1(n20644), .C2(n20467), .A(n20454), .B(n20453), .ZN(
        P1_U3123) );
  OAI22_X1 U23405 ( .A1(n20646), .A2(n20470), .B1(n20469), .B2(n20645), .ZN(
        n20455) );
  INV_X1 U23406 ( .A(n20455), .ZN(n20457) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20473), .B1(
        n20514), .B2(n20648), .ZN(n20456) );
  OAI211_X1 U23408 ( .C1(n20651), .C2(n20467), .A(n20457), .B(n20456), .ZN(
        P1_U3124) );
  AOI22_X1 U23409 ( .A1(n20653), .A2(n20461), .B1(n20652), .B2(n20460), .ZN(
        n20459) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20654), .ZN(n20458) );
  OAI211_X1 U23411 ( .C1(n20657), .C2(n20477), .A(n20459), .B(n20458), .ZN(
        P1_U3125) );
  AOI22_X1 U23412 ( .A1(n20661), .A2(n20461), .B1(n20659), .B2(n20460), .ZN(
        n20463) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20473), .B1(
        n20514), .B2(n20662), .ZN(n20462) );
  OAI211_X1 U23414 ( .C1(n20667), .C2(n20467), .A(n20463), .B(n20462), .ZN(
        P1_U3126) );
  OAI22_X1 U23415 ( .A1(n20669), .A2(n20470), .B1(n20469), .B2(n20668), .ZN(
        n20464) );
  INV_X1 U23416 ( .A(n20464), .ZN(n20466) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20473), .B1(
        n20514), .B2(n20508), .ZN(n20465) );
  OAI211_X1 U23418 ( .C1(n20468), .C2(n20467), .A(n20466), .B(n20465), .ZN(
        P1_U3127) );
  OAI22_X1 U23419 ( .A1(n20678), .A2(n20470), .B1(n20469), .B2(n20675), .ZN(
        n20471) );
  INV_X1 U23420 ( .A(n20471), .ZN(n20475) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20473), .B1(
        n20472), .B2(n20680), .ZN(n20474) );
  OAI211_X1 U23422 ( .C1(n20686), .C2(n20477), .A(n20475), .B(n20474), .ZN(
        P1_U3128) );
  NOR2_X2 U23423 ( .A1(n20622), .A2(n20476), .ZN(n20561) );
  INV_X1 U23424 ( .A(n20561), .ZN(n20478) );
  NAND3_X1 U23425 ( .A1(n20478), .A2(n20477), .A3(n20625), .ZN(n20480) );
  NAND2_X1 U23426 ( .A1(n20480), .A2(n20479), .ZN(n20486) );
  OR2_X1 U23427 ( .A1(n13583), .A2(n20481), .ZN(n20613) );
  NOR2_X1 U23428 ( .A1(n20613), .A2(n20565), .ZN(n20483) );
  AOI22_X1 U23429 ( .A1(n20486), .A2(n20483), .B1(n20488), .B2(n20568), .ZN(
        n20518) );
  NAND3_X1 U23430 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20482), .ZN(n20524) );
  NOR2_X1 U23431 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20524), .ZN(
        n20512) );
  AOI22_X1 U23432 ( .A1(n20617), .A2(n20512), .B1(n20561), .B2(n20627), .ZN(
        n20490) );
  INV_X1 U23433 ( .A(n20483), .ZN(n20485) );
  INV_X1 U23434 ( .A(n20512), .ZN(n20484) );
  AOI22_X1 U23435 ( .A1(n20486), .A2(n20485), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20484), .ZN(n20487) );
  OAI211_X1 U23436 ( .C1(n20488), .C2(n20689), .A(n20577), .B(n20487), .ZN(
        n20515) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20515), .B1(
        n20514), .B2(n20530), .ZN(n20489) );
  OAI211_X1 U23438 ( .C1(n20518), .C2(n20491), .A(n20490), .B(n20489), .ZN(
        P1_U3129) );
  AOI22_X1 U23439 ( .A1(n20492), .A2(n20512), .B1(n20561), .B2(n20634), .ZN(
        n20494) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20515), .B1(
        n20514), .B2(n20535), .ZN(n20493) );
  OAI211_X1 U23441 ( .C1(n20518), .C2(n20631), .A(n20494), .B(n20493), .ZN(
        P1_U3130) );
  INV_X1 U23442 ( .A(n20639), .ZN(n20495) );
  AOI22_X1 U23443 ( .A1(n20495), .A2(n20512), .B1(n20561), .B2(n20641), .ZN(
        n20497) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20515), .B1(
        n20514), .B2(n20540), .ZN(n20496) );
  OAI211_X1 U23445 ( .C1(n20518), .C2(n20638), .A(n20497), .B(n20496), .ZN(
        P1_U3131) );
  AOI22_X1 U23446 ( .A1(n20498), .A2(n20512), .B1(n20561), .B2(n20648), .ZN(
        n20500) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20515), .B1(
        n20514), .B2(n20545), .ZN(n20499) );
  OAI211_X1 U23448 ( .C1(n20518), .C2(n20645), .A(n20500), .B(n20499), .ZN(
        P1_U3132) );
  INV_X1 U23449 ( .A(n20657), .ZN(n20501) );
  AOI22_X1 U23450 ( .A1(n20652), .A2(n20512), .B1(n20561), .B2(n20501), .ZN(
        n20503) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20515), .B1(
        n20514), .B2(n20654), .ZN(n20502) );
  OAI211_X1 U23452 ( .C1(n20518), .C2(n20504), .A(n20503), .B(n20502), .ZN(
        P1_U3133) );
  AOI22_X1 U23453 ( .A1(n20659), .A2(n20512), .B1(n20561), .B2(n20662), .ZN(
        n20506) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20515), .B1(
        n20514), .B2(n20594), .ZN(n20505) );
  OAI211_X1 U23455 ( .C1(n20518), .C2(n20507), .A(n20506), .B(n20505), .ZN(
        P1_U3134) );
  INV_X1 U23456 ( .A(n20669), .ZN(n20509) );
  AOI22_X1 U23457 ( .A1(n20509), .A2(n20512), .B1(n20561), .B2(n20508), .ZN(
        n20511) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20515), .B1(
        n20514), .B2(n20671), .ZN(n20510) );
  OAI211_X1 U23459 ( .C1(n20518), .C2(n20668), .A(n20511), .B(n20510), .ZN(
        P1_U3135) );
  INV_X1 U23460 ( .A(n20678), .ZN(n20513) );
  AOI22_X1 U23461 ( .A1(n20513), .A2(n20512), .B1(n20561), .B2(n20605), .ZN(
        n20517) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20515), .B1(
        n20514), .B2(n20680), .ZN(n20516) );
  OAI211_X1 U23463 ( .C1(n20518), .C2(n20675), .A(n20517), .B(n20516), .ZN(
        P1_U3136) );
  AOI21_X1 U23464 ( .B1(n20524), .B2(n20520), .A(n20519), .ZN(n20534) );
  INV_X1 U23465 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20832) );
  NOR2_X1 U23466 ( .A1(n20521), .A2(n20524), .ZN(n20551) );
  INV_X1 U23467 ( .A(n20551), .ZN(n20559) );
  OAI21_X1 U23468 ( .B1(n20613), .B2(n20522), .A(n20559), .ZN(n20523) );
  NAND2_X1 U23469 ( .A1(n20523), .A2(n20625), .ZN(n20527) );
  INV_X1 U23470 ( .A(n20524), .ZN(n20525) );
  NAND2_X1 U23471 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20525), .ZN(n20526) );
  NAND2_X1 U23472 ( .A1(n20527), .A2(n20526), .ZN(n20552) );
  AOI22_X1 U23473 ( .A1(n20618), .A2(n20552), .B1(n20617), .B2(n20551), .ZN(
        n20532) );
  AOI22_X1 U23474 ( .A1(n20599), .A2(n20627), .B1(n20561), .B2(n20530), .ZN(
        n20531) );
  OAI211_X1 U23475 ( .C1(n20534), .C2(n20832), .A(n20532), .B(n20531), .ZN(
        P1_U3137) );
  INV_X1 U23476 ( .A(n20552), .ZN(n20558) );
  OAI22_X1 U23477 ( .A1(n20632), .A2(n20559), .B1(n20558), .B2(n20631), .ZN(
        n20533) );
  INV_X1 U23478 ( .A(n20533), .ZN(n20537) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20562), .B1(
        n20561), .B2(n20535), .ZN(n20536) );
  OAI211_X1 U23480 ( .C1(n20538), .C2(n20609), .A(n20537), .B(n20536), .ZN(
        P1_U3138) );
  OAI22_X1 U23481 ( .A1(n20639), .A2(n20559), .B1(n20558), .B2(n20638), .ZN(
        n20539) );
  INV_X1 U23482 ( .A(n20539), .ZN(n20542) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20562), .B1(
        n20561), .B2(n20540), .ZN(n20541) );
  OAI211_X1 U23484 ( .C1(n20543), .C2(n20609), .A(n20542), .B(n20541), .ZN(
        P1_U3139) );
  OAI22_X1 U23485 ( .A1(n20646), .A2(n20559), .B1(n20558), .B2(n20645), .ZN(
        n20544) );
  INV_X1 U23486 ( .A(n20544), .ZN(n20547) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20562), .B1(
        n20561), .B2(n20545), .ZN(n20546) );
  OAI211_X1 U23488 ( .C1(n20548), .C2(n20609), .A(n20547), .B(n20546), .ZN(
        P1_U3140) );
  AOI22_X1 U23489 ( .A1(n20653), .A2(n20552), .B1(n20652), .B2(n20551), .ZN(
        n20550) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20562), .B1(
        n20561), .B2(n20654), .ZN(n20549) );
  OAI211_X1 U23491 ( .C1(n20657), .C2(n20609), .A(n20550), .B(n20549), .ZN(
        P1_U3141) );
  AOI22_X1 U23492 ( .A1(n20661), .A2(n20552), .B1(n20659), .B2(n20551), .ZN(
        n20554) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20562), .B1(
        n20561), .B2(n20594), .ZN(n20553) );
  OAI211_X1 U23494 ( .C1(n20597), .C2(n20609), .A(n20554), .B(n20553), .ZN(
        P1_U3142) );
  OAI22_X1 U23495 ( .A1(n20669), .A2(n20559), .B1(n20558), .B2(n20668), .ZN(
        n20555) );
  INV_X1 U23496 ( .A(n20555), .ZN(n20557) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20562), .B1(
        n20561), .B2(n20671), .ZN(n20556) );
  OAI211_X1 U23498 ( .C1(n20674), .C2(n20609), .A(n20557), .B(n20556), .ZN(
        P1_U3143) );
  OAI22_X1 U23499 ( .A1(n20678), .A2(n20559), .B1(n20558), .B2(n20675), .ZN(
        n20560) );
  INV_X1 U23500 ( .A(n20560), .ZN(n20564) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20562), .B1(
        n20561), .B2(n20680), .ZN(n20563) );
  OAI211_X1 U23502 ( .C1(n20686), .C2(n20609), .A(n20564), .B(n20563), .ZN(
        P1_U3144) );
  INV_X1 U23503 ( .A(n20613), .ZN(n20566) );
  NAND2_X1 U23504 ( .A1(n20566), .A2(n20565), .ZN(n20574) );
  OR2_X1 U23505 ( .A1(n20574), .A2(n20567), .ZN(n20571) );
  NAND2_X1 U23506 ( .A1(n20569), .A2(n20568), .ZN(n20570) );
  NAND2_X1 U23507 ( .A1(n20571), .A2(n20570), .ZN(n20593) );
  NOR2_X1 U23508 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20614), .ZN(
        n20592) );
  AOI22_X1 U23509 ( .A1(n20618), .A2(n20593), .B1(n20617), .B2(n20592), .ZN(
        n20580) );
  NAND2_X1 U23510 ( .A1(n20573), .A2(n20572), .ZN(n20666) );
  OAI21_X1 U23511 ( .B1(n20599), .B2(n20681), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20575) );
  AOI21_X1 U23512 ( .B1(n20575), .B2(n20574), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20578) );
  OAI211_X1 U23513 ( .C1(n20592), .C2(n20578), .A(n20577), .B(n20576), .ZN(
        n20606) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20606), .B1(
        n20681), .B2(n20627), .ZN(n20579) );
  OAI211_X1 U23515 ( .C1(n20630), .C2(n20609), .A(n20580), .B(n20579), .ZN(
        P1_U3145) );
  INV_X1 U23516 ( .A(n20592), .ZN(n20603) );
  INV_X1 U23517 ( .A(n20593), .ZN(n20602) );
  OAI22_X1 U23518 ( .A1(n20632), .A2(n20603), .B1(n20602), .B2(n20631), .ZN(
        n20581) );
  INV_X1 U23519 ( .A(n20581), .ZN(n20583) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20606), .B1(
        n20681), .B2(n20634), .ZN(n20582) );
  OAI211_X1 U23521 ( .C1(n20637), .C2(n20609), .A(n20583), .B(n20582), .ZN(
        P1_U3146) );
  OAI22_X1 U23522 ( .A1(n20639), .A2(n20603), .B1(n20602), .B2(n20638), .ZN(
        n20584) );
  INV_X1 U23523 ( .A(n20584), .ZN(n20586) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20606), .B1(
        n20681), .B2(n20641), .ZN(n20585) );
  OAI211_X1 U23525 ( .C1(n20644), .C2(n20609), .A(n20586), .B(n20585), .ZN(
        P1_U3147) );
  OAI22_X1 U23526 ( .A1(n20646), .A2(n20603), .B1(n20602), .B2(n20645), .ZN(
        n20587) );
  INV_X1 U23527 ( .A(n20587), .ZN(n20589) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20606), .B1(
        n20681), .B2(n20648), .ZN(n20588) );
  OAI211_X1 U23529 ( .C1(n20651), .C2(n20609), .A(n20589), .B(n20588), .ZN(
        P1_U3148) );
  AOI22_X1 U23530 ( .A1(n20653), .A2(n20593), .B1(n20652), .B2(n20592), .ZN(
        n20591) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20606), .B1(
        n20599), .B2(n20654), .ZN(n20590) );
  OAI211_X1 U23532 ( .C1(n20657), .C2(n20666), .A(n20591), .B(n20590), .ZN(
        P1_U3149) );
  AOI22_X1 U23533 ( .A1(n20661), .A2(n20593), .B1(n20659), .B2(n20592), .ZN(
        n20596) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20606), .B1(
        n20599), .B2(n20594), .ZN(n20595) );
  OAI211_X1 U23535 ( .C1(n20597), .C2(n20666), .A(n20596), .B(n20595), .ZN(
        P1_U3150) );
  OAI22_X1 U23536 ( .A1(n20669), .A2(n20603), .B1(n20602), .B2(n20668), .ZN(
        n20598) );
  INV_X1 U23537 ( .A(n20598), .ZN(n20601) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20606), .B1(
        n20599), .B2(n20671), .ZN(n20600) );
  OAI211_X1 U23539 ( .C1(n20674), .C2(n20666), .A(n20601), .B(n20600), .ZN(
        P1_U3151) );
  OAI22_X1 U23540 ( .A1(n20678), .A2(n20603), .B1(n20602), .B2(n20675), .ZN(
        n20604) );
  INV_X1 U23541 ( .A(n20604), .ZN(n20608) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20606), .B1(
        n20681), .B2(n20605), .ZN(n20607) );
  OAI211_X1 U23543 ( .C1(n20610), .C2(n20609), .A(n20608), .B(n20607), .ZN(
        P1_U3152) );
  INV_X1 U23544 ( .A(n20611), .ZN(n20612) );
  INV_X1 U23545 ( .A(n20658), .ZN(n20677) );
  OAI21_X1 U23546 ( .B1(n20613), .B2(n20612), .A(n20677), .ZN(n20619) );
  NAND2_X1 U23547 ( .A1(n20619), .A2(n20625), .ZN(n20616) );
  INV_X1 U23548 ( .A(n20614), .ZN(n20626) );
  NAND2_X1 U23549 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20626), .ZN(n20615) );
  NAND2_X1 U23550 ( .A1(n20616), .A2(n20615), .ZN(n20660) );
  AOI22_X1 U23551 ( .A1(n20618), .A2(n20660), .B1(n20617), .B2(n20658), .ZN(
        n20629) );
  INV_X1 U23552 ( .A(n20619), .ZN(n20620) );
  OAI211_X1 U23553 ( .C1(n20622), .C2(n20621), .A(n20625), .B(n20620), .ZN(
        n20623) );
  OAI211_X1 U23554 ( .C1(n20626), .C2(n20625), .A(n20624), .B(n20623), .ZN(
        n20682) );
  INV_X1 U23555 ( .A(n20685), .ZN(n20663) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20682), .B1(
        n20663), .B2(n20627), .ZN(n20628) );
  OAI211_X1 U23557 ( .C1(n20630), .C2(n20666), .A(n20629), .B(n20628), .ZN(
        P1_U3153) );
  INV_X1 U23558 ( .A(n20660), .ZN(n20676) );
  OAI22_X1 U23559 ( .A1(n20632), .A2(n20677), .B1(n20676), .B2(n20631), .ZN(
        n20633) );
  INV_X1 U23560 ( .A(n20633), .ZN(n20636) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20682), .B1(
        n20663), .B2(n20634), .ZN(n20635) );
  OAI211_X1 U23562 ( .C1(n20637), .C2(n20666), .A(n20636), .B(n20635), .ZN(
        P1_U3154) );
  OAI22_X1 U23563 ( .A1(n20639), .A2(n20677), .B1(n20676), .B2(n20638), .ZN(
        n20640) );
  INV_X1 U23564 ( .A(n20640), .ZN(n20643) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20682), .B1(
        n20663), .B2(n20641), .ZN(n20642) );
  OAI211_X1 U23566 ( .C1(n20644), .C2(n20666), .A(n20643), .B(n20642), .ZN(
        P1_U3155) );
  OAI22_X1 U23567 ( .A1(n20646), .A2(n20677), .B1(n20676), .B2(n20645), .ZN(
        n20647) );
  INV_X1 U23568 ( .A(n20647), .ZN(n20650) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20682), .B1(
        n20663), .B2(n20648), .ZN(n20649) );
  OAI211_X1 U23570 ( .C1(n20651), .C2(n20666), .A(n20650), .B(n20649), .ZN(
        P1_U3156) );
  AOI22_X1 U23571 ( .A1(n20653), .A2(n20660), .B1(n20652), .B2(n20658), .ZN(
        n20656) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20682), .B1(
        n20681), .B2(n20654), .ZN(n20655) );
  OAI211_X1 U23573 ( .C1(n20657), .C2(n20685), .A(n20656), .B(n20655), .ZN(
        P1_U3157) );
  AOI22_X1 U23574 ( .A1(n20661), .A2(n20660), .B1(n20659), .B2(n20658), .ZN(
        n20665) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20682), .B1(
        n20663), .B2(n20662), .ZN(n20664) );
  OAI211_X1 U23576 ( .C1(n20667), .C2(n20666), .A(n20665), .B(n20664), .ZN(
        P1_U3158) );
  OAI22_X1 U23577 ( .A1(n20669), .A2(n20677), .B1(n20676), .B2(n20668), .ZN(
        n20670) );
  INV_X1 U23578 ( .A(n20670), .ZN(n20673) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20682), .B1(
        n20681), .B2(n20671), .ZN(n20672) );
  OAI211_X1 U23580 ( .C1(n20674), .C2(n20685), .A(n20673), .B(n20672), .ZN(
        P1_U3159) );
  OAI22_X1 U23581 ( .A1(n20678), .A2(n20677), .B1(n20676), .B2(n20675), .ZN(
        n20679) );
  INV_X1 U23582 ( .A(n20679), .ZN(n20684) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20682), .B1(
        n20681), .B2(n20680), .ZN(n20683) );
  OAI211_X1 U23584 ( .C1(n20686), .C2(n20685), .A(n20684), .B(n20683), .ZN(
        P1_U3160) );
  OAI211_X1 U23585 ( .C1(n20690), .C2(n20689), .A(n20688), .B(n20687), .ZN(
        P1_U3163) );
  INV_X1 U23586 ( .A(n20770), .ZN(n20766) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20766), .ZN(
        P1_U3164) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20766), .ZN(
        P1_U3165) );
  AND2_X1 U23589 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20766), .ZN(
        P1_U3166) );
  AND2_X1 U23590 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20766), .ZN(
        P1_U3167) );
  AND2_X1 U23591 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20766), .ZN(
        P1_U3168) );
  AND2_X1 U23592 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20766), .ZN(
        P1_U3169) );
  AND2_X1 U23593 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20766), .ZN(
        P1_U3170) );
  AND2_X1 U23594 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20766), .ZN(
        P1_U3171) );
  AND2_X1 U23595 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20766), .ZN(
        P1_U3172) );
  AND2_X1 U23596 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20766), .ZN(
        P1_U3173) );
  AND2_X1 U23597 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20766), .ZN(
        P1_U3174) );
  AND2_X1 U23598 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20766), .ZN(
        P1_U3175) );
  AND2_X1 U23599 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20766), .ZN(
        P1_U3176) );
  AND2_X1 U23600 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20766), .ZN(
        P1_U3177) );
  AND2_X1 U23601 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20766), .ZN(
        P1_U3178) );
  AND2_X1 U23602 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20766), .ZN(
        P1_U3179) );
  AND2_X1 U23603 ( .A1(n20766), .A2(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(
        P1_U3180) );
  AND2_X1 U23604 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20766), .ZN(
        P1_U3181) );
  AND2_X1 U23605 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20766), .ZN(
        P1_U3182) );
  AND2_X1 U23606 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20766), .ZN(
        P1_U3183) );
  AND2_X1 U23607 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20766), .ZN(
        P1_U3184) );
  AND2_X1 U23608 ( .A1(n20766), .A2(P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(
        P1_U3185) );
  AND2_X1 U23609 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20766), .ZN(P1_U3186) );
  AND2_X1 U23610 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20766), .ZN(P1_U3187) );
  AND2_X1 U23611 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20766), .ZN(P1_U3188) );
  AND2_X1 U23612 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20766), .ZN(P1_U3189) );
  AND2_X1 U23613 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20766), .ZN(P1_U3190) );
  AND2_X1 U23614 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20766), .ZN(P1_U3191) );
  AND2_X1 U23615 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20766), .ZN(P1_U3192) );
  AND2_X1 U23616 ( .A1(n20766), .A2(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(P1_U3193) );
  AOI21_X1 U23617 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20691), .A(n20701), 
        .ZN(n20703) );
  NOR2_X1 U23618 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20693) );
  NOR2_X1 U23619 ( .A1(n20693), .A2(n20692), .ZN(n20694) );
  INV_X1 U23620 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20699) );
  AOI211_X1 U23621 ( .C1(NA), .C2(n20701), .A(n20694), .B(n20699), .ZN(n20695)
         );
  OAI22_X1 U23622 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20703), .B1(n20794), 
        .B2(n20695), .ZN(P1_U3194) );
  NOR3_X1 U23623 ( .A1(NA), .A2(n20699), .A3(n20701), .ZN(n20697) );
  OAI22_X1 U23624 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20697), .B1(
        P1_STATE_REG_1__SCAN_IN), .B2(n20696), .ZN(n20702) );
  OAI211_X1 U23625 ( .C1(NA), .C2(n20797), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20704), .ZN(n20698) );
  OAI211_X1 U23626 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20699), .A(HOLD), .B(
        n20698), .ZN(n20700) );
  OAI22_X1 U23627 ( .A1(n20703), .A2(n20702), .B1(n20701), .B2(n20700), .ZN(
        P1_U3196) );
  NAND2_X1 U23628 ( .A1(n20794), .A2(n20704), .ZN(n20754) );
  INV_X1 U23629 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20707) );
  INV_X1 U23630 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20705) );
  AND2_X1 U23631 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20794), .ZN(n20751) );
  INV_X1 U23632 ( .A(n20751), .ZN(n20758) );
  OAI222_X1 U23633 ( .A1(n20754), .A2(n20707), .B1(n20705), .B2(n20794), .C1(
        n13525), .C2(n20758), .ZN(P1_U3197) );
  INV_X1 U23634 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20706) );
  OAI222_X1 U23635 ( .A1(n20758), .A2(n20707), .B1(n20706), .B2(n20794), .C1(
        n20709), .C2(n20754), .ZN(P1_U3198) );
  OAI222_X1 U23636 ( .A1(n20758), .A2(n20709), .B1(n20708), .B2(n20794), .C1(
        n20711), .C2(n20754), .ZN(P1_U3199) );
  INV_X1 U23637 ( .A(n20754), .ZN(n20748) );
  AOI22_X1 U23638 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20748), .ZN(n20710) );
  OAI21_X1 U23639 ( .B1(n20711), .B2(n20758), .A(n20710), .ZN(P1_U3200) );
  AOI22_X1 U23640 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20748), .ZN(n20712) );
  OAI21_X1 U23641 ( .B1(n15924), .B2(n20758), .A(n20712), .ZN(P1_U3201) );
  INV_X1 U23642 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20714) );
  AOI22_X1 U23643 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20748), .ZN(n20713) );
  OAI21_X1 U23644 ( .B1(n20714), .B2(n20758), .A(n20713), .ZN(P1_U3202) );
  AOI22_X1 U23645 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20751), .ZN(n20715) );
  OAI21_X1 U23646 ( .B1(n20717), .B2(n20754), .A(n20715), .ZN(P1_U3203) );
  AOI22_X1 U23647 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20748), .ZN(n20716) );
  OAI21_X1 U23648 ( .B1(n20717), .B2(n20758), .A(n20716), .ZN(P1_U3204) );
  AOI22_X1 U23649 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20751), .ZN(n20718) );
  OAI21_X1 U23650 ( .B1(n20720), .B2(n20754), .A(n20718), .ZN(P1_U3205) );
  AOI22_X1 U23651 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20748), .ZN(n20719) );
  OAI21_X1 U23652 ( .B1(n20720), .B2(n20758), .A(n20719), .ZN(P1_U3206) );
  AOI22_X1 U23653 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20751), .ZN(n20721) );
  OAI21_X1 U23654 ( .B1(n20723), .B2(n20754), .A(n20721), .ZN(P1_U3207) );
  INV_X1 U23655 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20722) );
  INV_X1 U23656 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20725) );
  OAI222_X1 U23657 ( .A1(n20758), .A2(n20723), .B1(n20722), .B2(n20794), .C1(
        n20725), .C2(n20754), .ZN(P1_U3208) );
  INV_X1 U23658 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20724) );
  OAI222_X1 U23659 ( .A1(n20758), .A2(n20725), .B1(n20724), .B2(n20794), .C1(
        n20726), .C2(n20754), .ZN(P1_U3209) );
  INV_X1 U23660 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20727) );
  OAI222_X1 U23661 ( .A1(n20754), .A2(n20729), .B1(n20727), .B2(n20794), .C1(
        n20726), .C2(n20758), .ZN(P1_U3210) );
  INV_X1 U23662 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20728) );
  OAI222_X1 U23663 ( .A1(n20758), .A2(n20729), .B1(n20728), .B2(n20794), .C1(
        n14773), .C2(n20754), .ZN(P1_U3211) );
  INV_X1 U23664 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20730) );
  OAI222_X1 U23665 ( .A1(n20758), .A2(n14773), .B1(n20730), .B2(n20794), .C1(
        n20732), .C2(n20754), .ZN(P1_U3212) );
  INV_X1 U23666 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20731) );
  OAI222_X1 U23667 ( .A1(n20758), .A2(n20732), .B1(n20731), .B2(n20794), .C1(
        n20734), .C2(n20754), .ZN(P1_U3213) );
  INV_X1 U23668 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20733) );
  OAI222_X1 U23669 ( .A1(n20758), .A2(n20734), .B1(n20733), .B2(n20794), .C1(
        n14744), .C2(n20754), .ZN(P1_U3214) );
  INV_X1 U23670 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20735) );
  OAI222_X1 U23671 ( .A1(n20754), .A2(n14728), .B1(n20735), .B2(n20794), .C1(
        n14744), .C2(n20758), .ZN(P1_U3215) );
  INV_X1 U23672 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20736) );
  OAI222_X1 U23673 ( .A1(n20758), .A2(n14728), .B1(n20736), .B2(n20794), .C1(
        n20738), .C2(n20754), .ZN(P1_U3216) );
  AOI22_X1 U23674 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20748), .ZN(n20737) );
  OAI21_X1 U23675 ( .B1(n20738), .B2(n20758), .A(n20737), .ZN(P1_U3217) );
  AOI22_X1 U23676 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20792), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20751), .ZN(n20739) );
  OAI21_X1 U23677 ( .B1(n20741), .B2(n20754), .A(n20739), .ZN(P1_U3218) );
  INV_X1 U23678 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20740) );
  OAI222_X1 U23679 ( .A1(n20758), .A2(n20741), .B1(n20740), .B2(n20794), .C1(
        n20743), .C2(n20754), .ZN(P1_U3219) );
  INV_X1 U23680 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20742) );
  OAI222_X1 U23681 ( .A1(n20758), .A2(n20743), .B1(n20742), .B2(n20794), .C1(
        n20745), .C2(n20754), .ZN(P1_U3220) );
  INV_X1 U23682 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20744) );
  OAI222_X1 U23683 ( .A1(n20758), .A2(n20745), .B1(n20744), .B2(n20794), .C1(
        n20747), .C2(n20754), .ZN(P1_U3221) );
  INV_X1 U23684 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20746) );
  OAI222_X1 U23685 ( .A1(n20758), .A2(n20747), .B1(n20746), .B2(n20794), .C1(
        n20750), .C2(n20754), .ZN(P1_U3222) );
  AOI22_X1 U23686 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20748), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20792), .ZN(n20749) );
  OAI21_X1 U23687 ( .B1(n20750), .B2(n20758), .A(n20749), .ZN(P1_U3223) );
  AOI22_X1 U23688 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20751), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20792), .ZN(n20752) );
  OAI21_X1 U23689 ( .B1(n20753), .B2(n20754), .A(n20752), .ZN(P1_U3224) );
  INV_X1 U23690 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20933) );
  OAI222_X1 U23691 ( .A1(n20754), .A2(n20757), .B1(n20933), .B2(n20794), .C1(
        n20753), .C2(n20758), .ZN(P1_U3225) );
  INV_X1 U23692 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20756) );
  OAI222_X1 U23693 ( .A1(n20758), .A2(n20757), .B1(n20756), .B2(n20794), .C1(
        n20755), .C2(n20754), .ZN(P1_U3226) );
  INV_X1 U23694 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20759) );
  AOI22_X1 U23695 ( .A1(n20794), .A2(n20760), .B1(n20759), .B2(n20792), .ZN(
        P1_U3458) );
  INV_X1 U23696 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20787) );
  INV_X1 U23697 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20761) );
  AOI22_X1 U23698 ( .A1(n20794), .A2(n20787), .B1(n20761), .B2(n20792), .ZN(
        P1_U3459) );
  INV_X1 U23699 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20762) );
  AOI22_X1 U23700 ( .A1(n20794), .A2(n20763), .B1(n20762), .B2(n20792), .ZN(
        P1_U3460) );
  INV_X1 U23701 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20790) );
  INV_X1 U23702 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20764) );
  AOI22_X1 U23703 ( .A1(n20794), .A2(n20790), .B1(n20764), .B2(n20792), .ZN(
        P1_U3461) );
  INV_X1 U23704 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20767) );
  INV_X1 U23705 ( .A(n20768), .ZN(n20765) );
  AOI21_X1 U23706 ( .B1(n20767), .B2(n20766), .A(n20765), .ZN(P1_U3464) );
  OAI21_X1 U23707 ( .B1(n20770), .B2(n20769), .A(n20768), .ZN(P1_U3465) );
  INV_X1 U23708 ( .A(n20771), .ZN(n20779) );
  OR2_X1 U23709 ( .A1(n20773), .A2(n20772), .ZN(n20778) );
  NAND3_X1 U23710 ( .A1(n20776), .A2(n20775), .A3(n20774), .ZN(n20777) );
  OAI211_X1 U23711 ( .C1(n20780), .C2(n20779), .A(n20778), .B(n20777), .ZN(
        n20782) );
  OAI22_X1 U23712 ( .A1(n20783), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n20782), .B2(n20781), .ZN(n20784) );
  INV_X1 U23713 ( .A(n20784), .ZN(P1_U3473) );
  AOI21_X1 U23714 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20785) );
  AOI22_X1 U23715 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20785), .B2(n13525), .ZN(n20788) );
  AOI22_X1 U23716 ( .A1(n20791), .A2(n20788), .B1(n20787), .B2(n20786), .ZN(
        P1_U3481) );
  OAI21_X1 U23717 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20791), .ZN(n20789) );
  OAI21_X1 U23718 ( .B1(n20791), .B2(n20790), .A(n20789), .ZN(P1_U3482) );
  AOI22_X1 U23719 ( .A1(n20794), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20793), 
        .B2(n20792), .ZN(P1_U3483) );
  AOI211_X1 U23720 ( .C1(n20798), .C2(n20797), .A(n20796), .B(n20795), .ZN(
        n20805) );
  OAI211_X1 U23721 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20800), .A(n20799), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20802) );
  AOI21_X1 U23722 ( .B1(n20802), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20801), 
        .ZN(n20804) );
  NAND2_X1 U23723 ( .A1(n20805), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20803) );
  OAI21_X1 U23724 ( .B1(n20805), .B2(n20804), .A(n20803), .ZN(P1_U3485) );
  MUX2_X1 U23725 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20794), .Z(P1_U3486) );
  OAI22_X1 U23726 ( .A1(n15307), .A2(keyinput47), .B1(n20807), .B2(keyinput10), 
        .ZN(n20806) );
  AOI221_X1 U23727 ( .B1(n15307), .B2(keyinput47), .C1(keyinput10), .C2(n20807), .A(n20806), .ZN(n20820) );
  INV_X1 U23728 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n20809) );
  OAI22_X1 U23729 ( .A1(n20810), .A2(keyinput63), .B1(n20809), .B2(keyinput28), 
        .ZN(n20808) );
  AOI221_X1 U23730 ( .B1(n20810), .B2(keyinput63), .C1(keyinput28), .C2(n20809), .A(n20808), .ZN(n20819) );
  OAI22_X1 U23731 ( .A1(n20813), .A2(keyinput37), .B1(n20812), .B2(keyinput16), 
        .ZN(n20811) );
  AOI221_X1 U23732 ( .B1(n20813), .B2(keyinput37), .C1(keyinput16), .C2(n20812), .A(n20811), .ZN(n20818) );
  OAI22_X1 U23733 ( .A1(n20816), .A2(keyinput55), .B1(n20815), .B2(keyinput24), 
        .ZN(n20814) );
  AOI221_X1 U23734 ( .B1(n20816), .B2(keyinput55), .C1(keyinput24), .C2(n20815), .A(n20814), .ZN(n20817) );
  NAND4_X1 U23735 ( .A1(n20820), .A2(n20819), .A3(n20818), .A4(n20817), .ZN(
        n20959) );
  INV_X1 U23736 ( .A(DATAI_25_), .ZN(n20822) );
  OAI22_X1 U23737 ( .A1(n20823), .A2(keyinput11), .B1(n20822), .B2(keyinput4), 
        .ZN(n20821) );
  AOI221_X1 U23738 ( .B1(n20823), .B2(keyinput11), .C1(keyinput4), .C2(n20822), 
        .A(n20821), .ZN(n20836) );
  INV_X1 U23739 ( .A(DATAI_16_), .ZN(n20826) );
  INV_X1 U23740 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n20825) );
  OAI22_X1 U23741 ( .A1(n20826), .A2(keyinput62), .B1(n20825), .B2(keyinput20), 
        .ZN(n20824) );
  AOI221_X1 U23742 ( .B1(n20826), .B2(keyinput62), .C1(keyinput20), .C2(n20825), .A(n20824), .ZN(n20835) );
  INV_X1 U23743 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n20828) );
  OAI22_X1 U23744 ( .A1(n20829), .A2(keyinput41), .B1(n20828), .B2(keyinput32), 
        .ZN(n20827) );
  AOI221_X1 U23745 ( .B1(n20829), .B2(keyinput41), .C1(keyinput32), .C2(n20828), .A(n20827), .ZN(n20834) );
  INV_X1 U23746 ( .A(keyinput5), .ZN(n20831) );
  OAI22_X1 U23747 ( .A1(n20832), .A2(keyinput3), .B1(n20831), .B2(
        P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20830) );
  AOI221_X1 U23748 ( .B1(n20832), .B2(keyinput3), .C1(
        P3_ADDRESS_REG_6__SCAN_IN), .C2(n20831), .A(n20830), .ZN(n20833) );
  NAND4_X1 U23749 ( .A1(n20836), .A2(n20835), .A3(n20834), .A4(n20833), .ZN(
        n20958) );
  INV_X1 U23750 ( .A(keyinput27), .ZN(n20838) );
  AOI22_X1 U23751 ( .A1(n20839), .A2(keyinput35), .B1(
        P2_DATAWIDTH_REG_27__SCAN_IN), .B2(n20838), .ZN(n20837) );
  OAI221_X1 U23752 ( .B1(n20839), .B2(keyinput35), .C1(n20838), .C2(
        P2_DATAWIDTH_REG_27__SCAN_IN), .A(n20837), .ZN(n20851) );
  AOI22_X1 U23753 ( .A1(n20842), .A2(keyinput9), .B1(n20841), .B2(keyinput60), 
        .ZN(n20840) );
  OAI221_X1 U23754 ( .B1(n20842), .B2(keyinput9), .C1(n20841), .C2(keyinput60), 
        .A(n20840), .ZN(n20850) );
  AOI22_X1 U23755 ( .A1(n20844), .A2(keyinput49), .B1(n13806), .B2(keyinput17), 
        .ZN(n20843) );
  OAI221_X1 U23756 ( .B1(n20844), .B2(keyinput49), .C1(n13806), .C2(keyinput17), .A(n20843), .ZN(n20849) );
  INV_X1 U23757 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n20846) );
  AOI22_X1 U23758 ( .A1(n20847), .A2(keyinput54), .B1(keyinput61), .B2(n20846), 
        .ZN(n20845) );
  OAI221_X1 U23759 ( .B1(n20847), .B2(keyinput54), .C1(n20846), .C2(keyinput61), .A(n20845), .ZN(n20848) );
  NOR4_X1 U23760 ( .A1(n20851), .A2(n20850), .A3(n20849), .A4(n20848), .ZN(
        n20900) );
  AOI22_X1 U23761 ( .A1(n20854), .A2(keyinput45), .B1(n20853), .B2(keyinput1), 
        .ZN(n20852) );
  OAI221_X1 U23762 ( .B1(n20854), .B2(keyinput45), .C1(n20853), .C2(keyinput1), 
        .A(n20852), .ZN(n20867) );
  INV_X1 U23763 ( .A(keyinput18), .ZN(n20857) );
  INV_X1 U23764 ( .A(keyinput22), .ZN(n20856) );
  AOI22_X1 U23765 ( .A1(n20857), .A2(P1_DATAWIDTH_REG_10__SCAN_IN), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n20856), .ZN(n20855) );
  OAI221_X1 U23766 ( .B1(n20857), .B2(P1_DATAWIDTH_REG_10__SCAN_IN), .C1(
        n20856), .C2(P3_ADDRESS_REG_2__SCAN_IN), .A(n20855), .ZN(n20866) );
  INV_X1 U23767 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20859) );
  AOI22_X1 U23768 ( .A1(n20860), .A2(keyinput39), .B1(n20859), .B2(keyinput51), 
        .ZN(n20858) );
  OAI221_X1 U23769 ( .B1(n20860), .B2(keyinput39), .C1(n20859), .C2(keyinput51), .A(n20858), .ZN(n20865) );
  INV_X1 U23770 ( .A(P3_LWORD_REG_1__SCAN_IN), .ZN(n20862) );
  AOI22_X1 U23771 ( .A1(n20863), .A2(keyinput23), .B1(keyinput31), .B2(n20862), 
        .ZN(n20861) );
  OAI221_X1 U23772 ( .B1(n20863), .B2(keyinput23), .C1(n20862), .C2(keyinput31), .A(n20861), .ZN(n20864) );
  NOR4_X1 U23773 ( .A1(n20867), .A2(n20866), .A3(n20865), .A4(n20864), .ZN(
        n20899) );
  INV_X1 U23774 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n20869) );
  AOI22_X1 U23775 ( .A1(n20870), .A2(keyinput33), .B1(n20869), .B2(keyinput34), 
        .ZN(n20868) );
  OAI221_X1 U23776 ( .B1(n20870), .B2(keyinput33), .C1(n20869), .C2(keyinput34), .A(n20868), .ZN(n20880) );
  INV_X1 U23777 ( .A(keyinput21), .ZN(n20872) );
  AOI22_X1 U23778 ( .A1(n12335), .A2(keyinput59), .B1(
        P1_DATAWIDTH_REG_2__SCAN_IN), .B2(n20872), .ZN(n20871) );
  OAI221_X1 U23779 ( .B1(n12335), .B2(keyinput59), .C1(n20872), .C2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A(n20871), .ZN(n20879) );
  INV_X1 U23780 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U23781 ( .A1(n20875), .A2(keyinput48), .B1(keyinput29), .B2(n20874), 
        .ZN(n20873) );
  OAI221_X1 U23782 ( .B1(n20875), .B2(keyinput48), .C1(n20874), .C2(keyinput29), .A(n20873), .ZN(n20878) );
  AOI22_X1 U23783 ( .A1(n12038), .A2(keyinput7), .B1(keyinput13), .B2(n12000), 
        .ZN(n20876) );
  OAI221_X1 U23784 ( .B1(n12038), .B2(keyinput7), .C1(n12000), .C2(keyinput13), 
        .A(n20876), .ZN(n20877) );
  NOR4_X1 U23785 ( .A1(n20880), .A2(n20879), .A3(n20878), .A4(n20877), .ZN(
        n20898) );
  INV_X1 U23786 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n20882) );
  AOI22_X1 U23787 ( .A1(n20883), .A2(keyinput46), .B1(keyinput38), .B2(n20882), 
        .ZN(n20881) );
  OAI221_X1 U23788 ( .B1(n20883), .B2(keyinput46), .C1(n20882), .C2(keyinput38), .A(n20881), .ZN(n20896) );
  AOI22_X1 U23789 ( .A1(n20886), .A2(keyinput57), .B1(keyinput50), .B2(n20885), 
        .ZN(n20884) );
  OAI221_X1 U23790 ( .B1(n20886), .B2(keyinput57), .C1(n20885), .C2(keyinput50), .A(n20884), .ZN(n20895) );
  AOI22_X1 U23791 ( .A1(n20889), .A2(keyinput52), .B1(n20888), .B2(keyinput53), 
        .ZN(n20887) );
  OAI221_X1 U23792 ( .B1(n20889), .B2(keyinput52), .C1(n20888), .C2(keyinput53), .A(n20887), .ZN(n20894) );
  INV_X1 U23793 ( .A(keyinput14), .ZN(n20891) );
  AOI22_X1 U23794 ( .A1(n20892), .A2(keyinput8), .B1(
        P1_DATAWIDTH_REG_15__SCAN_IN), .B2(n20891), .ZN(n20890) );
  OAI221_X1 U23795 ( .B1(n20892), .B2(keyinput8), .C1(n20891), .C2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A(n20890), .ZN(n20893) );
  NOR4_X1 U23796 ( .A1(n20896), .A2(n20895), .A3(n20894), .A4(n20893), .ZN(
        n20897) );
  NAND4_X1 U23797 ( .A1(n20900), .A2(n20899), .A3(n20898), .A4(n20897), .ZN(
        n20957) );
  NOR4_X1 U23798 ( .A1(keyinput62), .A2(keyinput47), .A3(keyinput42), .A4(
        keyinput30), .ZN(n20904) );
  NOR4_X1 U23799 ( .A1(keyinput26), .A2(keyinput19), .A3(keyinput15), .A4(
        keyinput11), .ZN(n20903) );
  NOR4_X1 U23800 ( .A1(keyinput6), .A2(keyinput3), .A3(keyinput2), .A4(
        keyinput37), .ZN(n20902) );
  NOR4_X1 U23801 ( .A1(keyinput25), .A2(keyinput40), .A3(keyinput56), .A4(
        keyinput20), .ZN(n20901) );
  NAND4_X1 U23802 ( .A1(n20904), .A2(n20903), .A3(n20902), .A4(n20901), .ZN(
        n20955) );
  NAND3_X1 U23803 ( .A1(keyinput27), .A2(keyinput9), .A3(keyinput60), .ZN(
        n20910) );
  NOR2_X1 U23804 ( .A1(keyinput54), .A2(keyinput17), .ZN(n20905) );
  NAND3_X1 U23805 ( .A1(keyinput49), .A2(keyinput61), .A3(n20905), .ZN(n20909)
         );
  NOR3_X1 U23806 ( .A1(keyinput45), .A2(keyinput1), .A3(keyinput22), .ZN(
        n20907) );
  NOR3_X1 U23807 ( .A1(keyinput39), .A2(keyinput51), .A3(keyinput31), .ZN(
        n20906) );
  NAND4_X1 U23808 ( .A1(keyinput18), .A2(n20907), .A3(keyinput23), .A4(n20906), 
        .ZN(n20908) );
  NOR4_X1 U23809 ( .A1(keyinput35), .A2(n20910), .A3(n20909), .A4(n20908), 
        .ZN(n20924) );
  INV_X1 U23810 ( .A(keyinput53), .ZN(n20911) );
  NOR4_X1 U23811 ( .A1(keyinput52), .A2(keyinput14), .A3(keyinput8), .A4(
        n20911), .ZN(n20923) );
  NOR2_X1 U23812 ( .A1(keyinput21), .A2(keyinput59), .ZN(n20912) );
  NAND3_X1 U23813 ( .A1(keyinput34), .A2(keyinput33), .A3(n20912), .ZN(n20916)
         );
  NAND3_X1 U23814 ( .A1(keyinput48), .A2(keyinput29), .A3(keyinput13), .ZN(
        n20915) );
  NOR2_X1 U23815 ( .A1(keyinput57), .A2(keyinput38), .ZN(n20913) );
  NAND3_X1 U23816 ( .A1(keyinput46), .A2(keyinput50), .A3(n20913), .ZN(n20914)
         );
  NOR4_X1 U23817 ( .A1(keyinput7), .A2(n20916), .A3(n20915), .A4(n20914), .ZN(
        n20922) );
  NAND4_X1 U23818 ( .A1(keyinput58), .A2(keyinput63), .A3(keyinput55), .A4(
        keyinput43), .ZN(n20920) );
  NAND4_X1 U23819 ( .A1(keyinput41), .A2(keyinput10), .A3(keyinput5), .A4(
        keyinput44), .ZN(n20919) );
  NAND4_X1 U23820 ( .A1(keyinput0), .A2(keyinput32), .A3(keyinput12), .A4(
        keyinput36), .ZN(n20918) );
  NAND4_X1 U23821 ( .A1(keyinput4), .A2(keyinput28), .A3(keyinput16), .A4(
        keyinput24), .ZN(n20917) );
  NOR4_X1 U23822 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20921) );
  NAND4_X1 U23823 ( .A1(n20924), .A2(n20923), .A3(n20922), .A4(n20921), .ZN(
        n20954) );
  AOI22_X1 U23824 ( .A1(n20927), .A2(keyinput26), .B1(n20926), .B2(keyinput0), 
        .ZN(n20925) );
  OAI221_X1 U23825 ( .B1(n20927), .B2(keyinput26), .C1(n20926), .C2(keyinput0), 
        .A(n20925), .ZN(n20937) );
  INV_X1 U23826 ( .A(keyinput42), .ZN(n20929) );
  AOI22_X1 U23827 ( .A1(n10651), .A2(keyinput44), .B1(
        P3_DATAWIDTH_REG_31__SCAN_IN), .B2(n20929), .ZN(n20928) );
  OAI221_X1 U23828 ( .B1(n10651), .B2(keyinput44), .C1(n20929), .C2(
        P3_DATAWIDTH_REG_31__SCAN_IN), .A(n20928), .ZN(n20936) );
  INV_X1 U23829 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20931) );
  AOI22_X1 U23830 ( .A1(n12257), .A2(keyinput19), .B1(keyinput25), .B2(n20931), 
        .ZN(n20930) );
  OAI221_X1 U23831 ( .B1(n12257), .B2(keyinput19), .C1(n20931), .C2(keyinput25), .A(n20930), .ZN(n20935) );
  AOI22_X1 U23832 ( .A1(n15008), .A2(keyinput58), .B1(n20933), .B2(keyinput43), 
        .ZN(n20932) );
  OAI221_X1 U23833 ( .B1(n15008), .B2(keyinput58), .C1(n20933), .C2(keyinput43), .A(n20932), .ZN(n20934) );
  NOR4_X1 U23834 ( .A1(n20937), .A2(n20936), .A3(n20935), .A4(n20934), .ZN(
        n20953) );
  INV_X1 U23835 ( .A(keyinput36), .ZN(n20939) );
  AOI22_X1 U23836 ( .A1(n20940), .A2(keyinput12), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n20939), .ZN(n20938) );
  OAI221_X1 U23837 ( .B1(n20940), .B2(keyinput12), .C1(n20939), .C2(
        P3_ADDRESS_REG_17__SCAN_IN), .A(n20938), .ZN(n20951) );
  AOI22_X1 U23838 ( .A1(n12236), .A2(keyinput2), .B1(keyinput40), .B2(n12983), 
        .ZN(n20941) );
  OAI221_X1 U23839 ( .B1(n12236), .B2(keyinput2), .C1(n12983), .C2(keyinput40), 
        .A(n20941), .ZN(n20950) );
  AOI22_X1 U23840 ( .A1(n20944), .A2(keyinput30), .B1(n20943), .B2(keyinput56), 
        .ZN(n20942) );
  OAI221_X1 U23841 ( .B1(n20944), .B2(keyinput30), .C1(n20943), .C2(keyinput56), .A(n20942), .ZN(n20949) );
  INV_X1 U23842 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20947) );
  INV_X1 U23843 ( .A(keyinput6), .ZN(n20946) );
  AOI22_X1 U23844 ( .A1(n20947), .A2(keyinput15), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n20946), .ZN(n20945) );
  OAI221_X1 U23845 ( .B1(n20947), .B2(keyinput15), .C1(n20946), .C2(
        P3_ADDRESS_REG_1__SCAN_IN), .A(n20945), .ZN(n20948) );
  NOR4_X1 U23846 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20952) );
  OAI211_X1 U23847 ( .C1(n20955), .C2(n20954), .A(n20953), .B(n20952), .ZN(
        n20956) );
  NOR4_X1 U23848 ( .A1(n20959), .A2(n20958), .A3(n20957), .A4(n20956), .ZN(
        n20963) );
  OAI21_X1 U23849 ( .B1(n20961), .B2(n19725), .A(n20960), .ZN(n20962) );
  XOR2_X1 U23850 ( .A(n20963), .B(n20962), .Z(P2_U2818) );
  CLKBUF_X2 U11369 ( .A(n9939), .Z(n10033) );
  AND2_X1 U12126 ( .A1(n11006), .A2(n13581), .ZN(n11035) );
  BUF_X1 U11157 ( .A(n10844), .Z(n16957) );
  NAND2_X1 U11407 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17222), .ZN(n17218) );
  CLKBUF_X1 U11068 ( .A(n11105), .Z(n11779) );
  CLKBUF_X2 U11085 ( .A(n11212), .Z(n11761) );
  CLKBUF_X1 U11109 ( .A(n11867), .Z(n11956) );
  CLKBUF_X1 U11160 ( .A(n10098), .Z(n13059) );
  OR2_X1 U11168 ( .A1(n11985), .A2(n11990), .ZN(n12196) );
  CLKBUF_X1 U11736 ( .A(n11121), .Z(n13671) );
  OR2_X1 U11838 ( .A1(n10658), .A2(n10666), .ZN(n9644) );
  CLKBUF_X1 U12010 ( .A(n17670), .Z(n9624) );
  CLKBUF_X1 U12029 ( .A(n14608), .Z(n14741) );
  CLKBUF_X1 U12084 ( .A(n19036), .Z(n19027) );
  INV_X2 U12165 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10651) );
  CLKBUF_X1 U12191 ( .A(n17388), .Z(n17396) );
endmodule

