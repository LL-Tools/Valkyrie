

module b17_C_SARLock_k_128_2 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9733, n9734, n9735, n9737, n9738, n9739, n9741, n9742, n9743, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21178;

  XNOR2_X1 U11178 ( .A(n14908), .B(n10053), .ZN(n14920) );
  INV_X1 U11179 ( .A(n20040), .ZN(n20054) );
  OR2_X1 U11180 ( .A1(n14245), .A2(n14244), .ZN(n14247) );
  INV_X2 U11181 ( .A(n12131), .ZN(n10051) );
  AND2_X1 U11182 ( .A1(n9869), .A2(n11870), .ZN(n10188) );
  AND4_X1 U11183 ( .A1(n17485), .A2(n15566), .A3(n18303), .A4(n15559), .ZN(
        n17523) );
  CLKBUF_X2 U11184 ( .A(n15602), .Z(n15595) );
  INV_X1 U11185 ( .A(n9735), .ZN(n9739) );
  NAND2_X1 U11187 ( .A1(n11822), .A2(n11823), .ZN(n11821) );
  INV_X1 U11188 ( .A(n20851), .ZN(n13138) );
  AND2_X1 U11189 ( .A1(n10452), .A2(n10438), .ZN(n10240) );
  AND2_X1 U11190 ( .A1(n11543), .A2(n12710), .ZN(n11586) );
  AND2_X1 U11191 ( .A1(n9749), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12414) );
  NAND2_X1 U11192 ( .A1(n20177), .A2(n13428), .ZN(n20851) );
  CLKBUF_X2 U11193 ( .A(n11723), .Z(n12901) );
  CLKBUF_X2 U11194 ( .A(n11672), .Z(n12870) );
  INV_X2 U11195 ( .A(n13626), .ZN(n20177) );
  INV_X1 U11196 ( .A(n13338), .ZN(n9873) );
  INV_X1 U11198 ( .A(n16993), .ZN(n17274) );
  INV_X1 U11199 ( .A(n9735), .ZN(n9738) );
  CLKBUF_X2 U11200 ( .A(n15481), .Z(n17272) );
  INV_X1 U11201 ( .A(n17288), .ZN(n17267) );
  CLKBUF_X2 U11202 ( .A(n15481), .Z(n17252) );
  CLKBUF_X1 U11203 ( .A(n15602), .Z(n17291) );
  OR2_X1 U11204 ( .A1(n15539), .A2(n17024), .ZN(n10254) );
  CLKBUF_X1 U11205 ( .A(n15624), .Z(n17196) );
  INV_X2 U11206 ( .A(n11013), .ZN(n10971) );
  INV_X1 U11207 ( .A(n10262), .ZN(n17285) );
  INV_X2 U11208 ( .A(n16993), .ZN(n15669) );
  NAND2_X1 U11209 ( .A1(n11776), .A2(n11750), .ZN(n11763) );
  AND4_X1 U11210 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11712) );
  AND2_X1 U11211 ( .A1(n10279), .A2(n10288), .ZN(n11068) );
  AND2_X4 U11212 ( .A1(n10279), .A2(n10284), .ZN(n10329) );
  AND2_X1 U11213 ( .A1(n10287), .A2(n14661), .ZN(n10746) );
  INV_X1 U11214 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11537) );
  CLKBUF_X1 U11215 ( .A(n15055), .Z(n9733) );
  NOR2_X1 U11216 ( .A1(n13092), .A2(n15585), .ZN(n15055) );
  AND2_X1 U11217 ( .A1(n11773), .A2(n12928), .ZN(n11752) );
  AND2_X2 U11218 ( .A1(n11542), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11551) );
  INV_X1 U11219 ( .A(n19290), .ZN(n12247) );
  OAI21_X1 U11220 ( .B1(n10560), .B2(n11427), .A(n10552), .ZN(n10578) );
  AND2_X1 U11221 ( .A1(n12710), .A2(n14000), .ZN(n11585) );
  AND2_X1 U11222 ( .A1(n11538), .A2(n11539), .ZN(n12735) );
  AOI21_X1 U11223 ( .B1(n9747), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11779), .ZN(n11796) );
  XNOR2_X1 U11225 ( .A(n10551), .B(n10550), .ZN(n10560) );
  AND3_X1 U11226 ( .A1(n11775), .A2(n11774), .A3(n11773), .ZN(n12260) );
  BUF_X1 U11227 ( .A(n11804), .Z(n12533) );
  AND2_X1 U11228 ( .A1(n14770), .A2(n12769), .ZN(n12746) );
  NAND2_X2 U11229 ( .A1(n11754), .A2(n12330), .ZN(n12450) );
  NAND2_X1 U11230 ( .A1(n9855), .A2(n11846), .ZN(n11934) );
  AND2_X1 U11231 ( .A1(n19290), .A2(n12255), .ZN(n11757) );
  INV_X1 U11232 ( .A(n9735), .ZN(n9737) );
  INV_X1 U11233 ( .A(n13428), .ZN(n20162) );
  INV_X1 U11234 ( .A(n10426), .ZN(n20214) );
  INV_X1 U11235 ( .A(n12587), .ZN(n11774) );
  NAND3_X1 U11236 ( .A1(n11757), .A2(n11730), .A3(n11754), .ZN(n12175) );
  INV_X1 U11237 ( .A(n17792), .ZN(n17856) );
  INV_X1 U11238 ( .A(n11286), .ZN(n14035) );
  NOR2_X1 U11239 ( .A1(n14886), .A2(n14897), .ZN(n14891) );
  OAI22_X1 U11240 ( .A1(n14910), .A2(n14909), .B1(n14920), .B2(n15134), .ZN(
        n14913) );
  INV_X1 U11241 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16435) );
  NAND2_X1 U11242 ( .A1(n18151), .A2(n18732), .ZN(n18168) );
  INV_X1 U11243 ( .A(n20031), .ZN(n15890) );
  NAND2_X1 U11245 ( .A1(n11821), .A2(n11824), .ZN(n13607) );
  NOR2_X1 U11247 ( .A1(n18929), .A2(n16657), .ZN(n17914) );
  AND2_X4 U11248 ( .A1(n10285), .A2(n10284), .ZN(n10681) );
  NOR2_X2 U11249 ( .A1(n17733), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17732) );
  INV_X1 U11250 ( .A(n12819), .ZN(n11718) );
  NOR3_X2 U11251 ( .A1(n12051), .A2(n12049), .A3(n11664), .ZN(n12066) );
  NOR2_X1 U11254 ( .A1(n15539), .A2(n15356), .ZN(n15494) );
  NAND2_X1 U11255 ( .A1(n14465), .A2(n14644), .ZN(n14487) );
  XNOR2_X2 U11256 ( .A(n11945), .B(n12001), .ZN(n12208) );
  AOI211_X2 U11257 ( .C1(n15100), .C2(n9733), .A(n14894), .B(n14893), .ZN(
        n14895) );
  OAI21_X2 U11258 ( .B1(n12086), .B2(n10051), .A(n15240), .ZN(n15016) );
  AND3_X4 U11259 ( .A1(n11795), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n16435), .ZN(n11722) );
  NOR2_X2 U11261 ( .A1(n15425), .A2(n15424), .ZN(n18303) );
  NOR2_X1 U11263 ( .A1(n14441), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15827) );
  NOR3_X2 U11264 ( .A1(n14454), .A2(n14501), .A3(n14609), .ZN(n15826) );
  AND2_X4 U11265 ( .A1(n12901), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11896) );
  XNOR2_X2 U11266 ( .A(n10488), .B(n10487), .ZN(n10570) );
  AND2_X1 U11267 ( .A1(n9860), .A2(n9859), .ZN(n14886) );
  NAND2_X1 U11268 ( .A1(n10197), .A2(n9848), .ZN(n14921) );
  INV_X1 U11269 ( .A(n14963), .ZN(n10197) );
  NOR2_X1 U11270 ( .A1(n14963), .A2(n10200), .ZN(n14947) );
  XNOR2_X1 U11271 ( .A(n12970), .B(n12926), .ZN(n16189) );
  NOR2_X1 U11272 ( .A1(n15705), .A2(n17691), .ZN(n17651) );
  XNOR2_X1 U11273 ( .A(n11968), .B(n16404), .ZN(n16333) );
  NOR2_X1 U11274 ( .A1(n17691), .A2(n17680), .ZN(n17722) );
  NAND2_X1 U11275 ( .A1(n11948), .A2(n13639), .ZN(n11968) );
  NAND2_X1 U11276 ( .A1(n18048), .A2(n17840), .ZN(n17755) );
  NAND2_X1 U11277 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  INV_X1 U11278 ( .A(n11847), .ZN(n9855) );
  MUX2_X1 U11279 ( .A(n10568), .B(n10567), .S(n10566), .Z(n20830) );
  INV_X2 U11280 ( .A(n18716), .ZN(n18722) );
  BUF_X2 U11281 ( .A(n16942), .Z(n16953) );
  XNOR2_X1 U11282 ( .A(n11798), .B(n11796), .ZN(n11825) );
  NOR2_X2 U11283 ( .A1(n20970), .A2(n17589), .ZN(n16680) );
  NOR2_X2 U11284 ( .A1(n11770), .A2(n11769), .ZN(n12464) );
  BUF_X2 U11285 ( .A(n11307), .Z(n9748) );
  AND2_X1 U11286 ( .A1(n14016), .A2(n14027), .ZN(n10438) );
  NOR2_X1 U11287 ( .A1(n10411), .A2(n14015), .ZN(n12992) );
  NAND2_X2 U11288 ( .A1(n12330), .A2(n12130), .ZN(n12281) );
  NAND2_X1 U11289 ( .A1(n20214), .A2(n14281), .ZN(n10437) );
  INV_X2 U11290 ( .A(n18929), .ZN(n9961) );
  NAND2_X1 U11291 ( .A1(n11764), .A2(n11743), .ZN(n11742) );
  BUF_X1 U11292 ( .A(n11764), .Z(n19307) );
  OR2_X1 U11293 ( .A1(n9950), .A2(n15640), .ZN(n15681) );
  BUF_X2 U11294 ( .A(n12293), .Z(n12458) );
  INV_X2 U11295 ( .A(n12973), .ZN(n11750) );
  INV_X2 U11296 ( .A(n12255), .ZN(n11751) );
  INV_X4 U11297 ( .A(n18316), .ZN(n17450) );
  BUF_X1 U11298 ( .A(n11744), .Z(n19297) );
  BUF_X1 U11299 ( .A(n11732), .Z(n12928) );
  NAND4_X1 U11300 ( .A1(n10377), .A2(n10376), .A3(n10375), .A4(n10374), .ZN(
        n14027) );
  AOI22_X1 U11301 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15366) );
  CLKBUF_X2 U11302 ( .A(n10746), .Z(n11206) );
  INV_X1 U11303 ( .A(n10382), .ZN(n11013) );
  BUF_X4 U11304 ( .A(n15418), .Z(n9741) );
  NOR2_X1 U11305 ( .A1(n15352), .A2(n15355), .ZN(n15481) );
  AND2_X1 U11306 ( .A1(n10279), .A2(n10287), .ZN(n10416) );
  INV_X2 U11307 ( .A(n11168), .ZN(n11205) );
  INV_X4 U11308 ( .A(n11010), .ZN(n9742) );
  INV_X2 U11309 ( .A(n11168), .ZN(n10970) );
  AND2_X1 U11310 ( .A1(n13353), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10285) );
  AND2_X1 U11311 ( .A1(n13370), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10279) );
  NOR2_X2 U11312 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11542) );
  NOR2_X1 U11313 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U11314 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15539) );
  OR2_X1 U11315 ( .A1(n12126), .A2(n12127), .ZN(n9860) );
  AND2_X1 U11316 ( .A1(n10184), .A2(n10187), .ZN(n13993) );
  NAND2_X1 U11317 ( .A1(n9864), .A2(n9863), .ZN(n9862) );
  INV_X1 U11318 ( .A(n9914), .ZN(n14916) );
  NAND2_X1 U11319 ( .A1(n9814), .A2(n9921), .ZN(n9920) );
  AOI21_X1 U11320 ( .B1(n15027), .B2(n10005), .A(n10004), .ZN(n10001) );
  OAI21_X1 U11321 ( .B1(n14424), .B2(n10026), .A(n10024), .ZN(n10023) );
  AOI211_X1 U11322 ( .C1(n15037), .C2(n10000), .A(n14975), .B(n10002), .ZN(
        n14990) );
  AOI21_X1 U11323 ( .B1(n14082), .B2(n14090), .A(n14081), .ZN(n14398) );
  NAND3_X1 U11324 ( .A1(n9809), .A2(n10063), .A3(n14595), .ZN(n14356) );
  NOR2_X1 U11325 ( .A1(n14389), .A2(n14515), .ZN(n14390) );
  NAND2_X1 U11326 ( .A1(n14416), .A2(n10025), .ZN(n10024) );
  NOR2_X1 U11327 ( .A1(n17593), .A2(n17592), .ZN(n17591) );
  NAND2_X1 U11328 ( .A1(n10014), .A2(n10017), .ZN(n15059) );
  NAND2_X1 U11329 ( .A1(n14409), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14389) );
  NOR2_X1 U11330 ( .A1(n10064), .A2(n14377), .ZN(n10063) );
  OR2_X1 U11331 ( .A1(n14104), .A2(n14069), .ZN(n14080) );
  OR2_X1 U11332 ( .A1(n14104), .A2(n14092), .ZN(n14090) );
  NOR2_X1 U11333 ( .A1(n14133), .A2(n14135), .ZN(n14134) );
  NOR2_X1 U11334 ( .A1(n14133), .A2(n10250), .ZN(n14116) );
  NAND2_X1 U11335 ( .A1(n14594), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11517) );
  OR2_X1 U11336 ( .A1(n14439), .A2(n11515), .ZN(n11516) );
  OR2_X1 U11337 ( .A1(n14733), .A2(n14732), .ZN(n15128) );
  NAND2_X1 U11338 ( .A1(n9947), .A2(n9945), .ZN(n16563) );
  NAND2_X1 U11339 ( .A1(n10091), .A2(n14499), .ZN(n10022) );
  NOR2_X1 U11340 ( .A1(n14752), .A2(n10134), .ZN(n14733) );
  NOR2_X1 U11341 ( .A1(n14752), .A2(n14744), .ZN(n14743) );
  NAND2_X1 U11342 ( .A1(n13963), .A2(n11501), .ZN(n14499) );
  AOI21_X1 U11343 ( .B1(n10193), .B2(n10195), .A(n10191), .ZN(n10190) );
  NAND2_X1 U11344 ( .A1(n15327), .A2(n12018), .ZN(n10196) );
  OR2_X1 U11345 ( .A1(n15327), .A2(n12018), .ZN(n10195) );
  OAI22_X1 U11346 ( .A1(n13844), .A2(n13843), .B1(n11967), .B2(n16405), .ZN(
        n16334) );
  OR2_X2 U11347 ( .A1(n14796), .A2(n10176), .ZN(n12745) );
  OAI21_X1 U11348 ( .B1(n12225), .B2(n12131), .A(n19089), .ZN(n12007) );
  NOR2_X1 U11349 ( .A1(n10090), .A2(n11502), .ZN(n10086) );
  NAND2_X1 U11350 ( .A1(n9887), .A2(n9922), .ZN(n16020) );
  OR2_X1 U11351 ( .A1(n12234), .A2(n10051), .ZN(n12236) );
  NOR2_X1 U11352 ( .A1(n9925), .A2(n9886), .ZN(n9885) );
  AOI21_X1 U11353 ( .B1(n16024), .B2(n9924), .A(n9923), .ZN(n9922) );
  AND2_X1 U11354 ( .A1(n17610), .A2(n16731), .ZN(n16738) );
  AND2_X1 U11355 ( .A1(n9974), .A2(n13711), .ZN(n9973) );
  NOR2_X1 U11356 ( .A1(n15701), .A2(n15700), .ZN(n17742) );
  NOR2_X1 U11357 ( .A1(n13849), .A2(n13848), .ZN(n13851) );
  NAND2_X1 U11358 ( .A1(n10617), .A2(n10616), .ZN(n13481) );
  XNOR2_X1 U11359 ( .A(n11477), .B(n10697), .ZN(n11486) );
  INV_X1 U11360 ( .A(n9734), .ZN(n17944) );
  NOR3_X1 U11361 ( .A1(n11886), .A2(n11885), .A3(n11884), .ZN(n11894) );
  OR2_X1 U11362 ( .A1(n10559), .A2(n10558), .ZN(n13376) );
  NOR2_X1 U11363 ( .A1(n12629), .A2(n10167), .ZN(n10166) );
  NAND2_X1 U11364 ( .A1(n18759), .A2(n9957), .ZN(n17943) );
  CLKBUF_X1 U11365 ( .A(n11436), .Z(n20431) );
  NAND2_X1 U11366 ( .A1(n9959), .A2(n9958), .ZN(n18759) );
  NAND2_X1 U11367 ( .A1(n13172), .A2(n12618), .ZN(n13118) );
  OR2_X1 U11368 ( .A1(n12628), .A2(n12625), .ZN(n12626) );
  OR2_X1 U11369 ( .A1(n13391), .A2(n13390), .ZN(n13397) );
  NAND2_X1 U11370 ( .A1(n9855), .A2(n10052), .ZN(n11917) );
  NAND3_X1 U11371 ( .A1(n10580), .A2(n10579), .A3(n10604), .ZN(n10636) );
  CLKBUF_X1 U11372 ( .A(n13014), .Z(n14343) );
  NAND2_X1 U11373 ( .A1(n11848), .A2(n11820), .ZN(n19602) );
  OR2_X1 U11374 ( .A1(n11836), .A2(n11827), .ZN(n19502) );
  NAND2_X1 U11375 ( .A1(n17866), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17865) );
  NOR2_X1 U11376 ( .A1(n11847), .A2(n13098), .ZN(n11848) );
  OR2_X1 U11377 ( .A1(n11843), .A2(n11842), .ZN(n19350) );
  OR2_X1 U11378 ( .A1(n11843), .A2(n11841), .ZN(n19275) );
  OR2_X1 U11379 ( .A1(n11836), .A2(n11842), .ZN(n19475) );
  OR2_X1 U11380 ( .A1(n11836), .A2(n11853), .ZN(n19444) );
  OR2_X1 U11381 ( .A1(n11836), .A2(n11841), .ZN(n19416) );
  OR2_X1 U11382 ( .A1(n11843), .A2(n11853), .ZN(n19325) );
  OR2_X1 U11383 ( .A1(n11843), .A2(n11827), .ZN(n19384) );
  INV_X2 U11384 ( .A(n13680), .ZN(n20119) );
  XNOR2_X1 U11385 ( .A(n12617), .B(n12615), .ZN(n13174) );
  NOR2_X1 U11386 ( .A1(n20328), .A2(n20193), .ZN(n20707) );
  NOR2_X1 U11387 ( .A1(n20328), .A2(n20200), .ZN(n20713) );
  NOR2_X1 U11388 ( .A1(n20328), .A2(n20208), .ZN(n20719) );
  NOR2_X1 U11389 ( .A1(n20328), .A2(n20185), .ZN(n20701) );
  NOR2_X1 U11390 ( .A1(n20328), .A2(n20227), .ZN(n20734) );
  NOR2_X1 U11391 ( .A1(n20328), .A2(n20163), .ZN(n20685) );
  NOR2_X1 U11392 ( .A1(n20328), .A2(n20215), .ZN(n20725) );
  NOR2_X1 U11393 ( .A1(n20328), .A2(n20179), .ZN(n20695) );
  NAND2_X1 U11394 ( .A1(n12604), .A2(n12603), .ZN(n12617) );
  NAND2_X1 U11395 ( .A1(n13089), .A2(n15585), .ZN(n19259) );
  NAND2_X1 U11396 ( .A1(n12611), .A2(n12610), .ZN(n13612) );
  AND2_X1 U11397 ( .A1(n10141), .A2(n10140), .ZN(n10139) );
  OR2_X1 U11398 ( .A1(n13607), .A2(n16471), .ZN(n12611) );
  NOR2_X1 U11399 ( .A1(n13512), .A2(n10142), .ZN(n10141) );
  NAND2_X1 U11400 ( .A1(n10526), .A2(n10525), .ZN(n10551) );
  OAI21_X4 U11401 ( .B1(n13989), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12937), 
        .ZN(n12939) );
  OAI211_X1 U11402 ( .C1(n20164), .C2(n11520), .A(n10465), .B(n10464), .ZN(
        n10466) );
  XNOR2_X1 U11403 ( .A(n12936), .B(n14684), .ZN(n13989) );
  AND2_X1 U11404 ( .A1(n12011), .A2(n12010), .ZN(n12022) );
  NOR2_X1 U11405 ( .A1(n13504), .A2(n13505), .ZN(n13579) );
  NAND2_X1 U11406 ( .A1(n13054), .A2(n13053), .ZN(n13052) );
  CLKBUF_X1 U11407 ( .A(n11825), .Z(n11830) );
  NAND2_X1 U11408 ( .A1(n17896), .A2(n15689), .ZN(n15692) );
  NOR2_X1 U11409 ( .A1(n12004), .A2(n12003), .ZN(n12015) );
  NAND2_X1 U11410 ( .A1(n12200), .A2(n12198), .ZN(n16449) );
  OAI21_X1 U11411 ( .B1(n11801), .B2(n16435), .A(n11802), .ZN(n11818) );
  XOR2_X1 U11412 ( .A(n16689), .B(n16486), .Z(n16942) );
  OR2_X1 U11413 ( .A1(n13609), .A2(n12245), .ZN(n12595) );
  NAND3_X2 U11414 ( .A1(n9961), .A2(n17523), .A3(n17522), .ZN(n17586) );
  OAI211_X1 U11415 ( .C1(n11804), .C2(n13085), .A(n11782), .B(n11781), .ZN(
        n11783) );
  NOR2_X1 U11416 ( .A1(n12964), .A2(n16227), .ZN(n12965) );
  NAND2_X1 U11417 ( .A1(n10395), .A2(n10394), .ZN(n10241) );
  CLKBUF_X1 U11418 ( .A(n12992), .Z(n13412) );
  AND2_X1 U11419 ( .A1(n10446), .A2(n10436), .ZN(n13342) );
  OR2_X1 U11420 ( .A1(n13348), .A2(n10427), .ZN(n13436) );
  AND3_X1 U11421 ( .A1(n13429), .A2(n10433), .A3(n10432), .ZN(n10445) );
  NAND2_X1 U11422 ( .A1(n11307), .A2(n11286), .ZN(n13501) );
  NAND2_X1 U11423 ( .A1(n10438), .A2(n13326), .ZN(n13366) );
  NAND2_X1 U11424 ( .A1(n12260), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11804) );
  OAI211_X1 U11425 ( .C1(n12249), .C2(n11760), .A(n11759), .B(n11758), .ZN(
        n11771) );
  INV_X1 U11426 ( .A(n12175), .ZN(n12162) );
  AND2_X1 U11427 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11773), .ZN(n9745) );
  AND2_X1 U11428 ( .A1(n13741), .A2(n20851), .ZN(n14033) );
  CLKBUF_X1 U11429 ( .A(n12159), .Z(n16456) );
  INV_X1 U11430 ( .A(n12627), .ZN(n10167) );
  NAND2_X1 U11431 ( .A1(n11424), .A2(n9873), .ZN(n14015) );
  NOR2_X1 U11432 ( .A1(n9773), .A2(n15006), .ZN(n12955) );
  AND2_X1 U11433 ( .A1(n11777), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U11434 ( .A1(n11763), .A2(n12587), .ZN(n12246) );
  OR2_X1 U11435 ( .A1(n11620), .A2(n11619), .ZN(n11869) );
  NAND2_X2 U11436 ( .A1(n13428), .A2(n13626), .ZN(n11302) );
  OR2_X1 U11437 ( .A1(n11603), .A2(n11602), .ZN(n12216) );
  AND2_X1 U11438 ( .A1(n12169), .A2(n12929), .ZN(n9746) );
  AND2_X1 U11439 ( .A1(n11703), .A2(n11739), .ZN(n11735) );
  OR2_X1 U11440 ( .A1(n11550), .A2(n11549), .ZN(n11912) );
  NOR2_X4 U11441 ( .A1(n13428), .A2(n13626), .ZN(n10451) );
  INV_X1 U11442 ( .A(n11732), .ZN(n11764) );
  NAND2_X1 U11443 ( .A1(n12951), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12950) );
  NAND2_X1 U11444 ( .A1(n12283), .A2(n12973), .ZN(n12587) );
  NAND2_X2 U11445 ( .A1(n11679), .A2(n11678), .ZN(n12929) );
  INV_X4 U11446 ( .A(n12283), .ZN(n11776) );
  MUX2_X1 U11447 ( .A(n11729), .B(n11728), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12255) );
  AND4_X2 U11448 ( .A1(n9788), .A2(n10355), .A3(n10354), .A4(n9890), .ZN(
        n20199) );
  AND4_X1 U11449 ( .A1(n10413), .A2(n10417), .A3(n9970), .A4(n9969), .ZN(n9968) );
  AND2_X1 U11450 ( .A1(n12947), .A2(n9758), .ZN(n12951) );
  AND4_X1 U11451 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n11713) );
  NOR2_X1 U11452 ( .A1(n9791), .A2(n9971), .ZN(n9970) );
  AND3_X1 U11453 ( .A1(n9891), .A2(n10339), .A3(n10338), .ZN(n9890) );
  NOR2_X2 U11454 ( .A1(n12944), .A2(n16315), .ZN(n12947) );
  AND4_X1 U11455 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n10355) );
  AND4_X1 U11456 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n10293) );
  AND4_X1 U11457 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10375) );
  AND4_X1 U11458 ( .A1(n10300), .A2(n10299), .A3(n10298), .A4(n10297), .ZN(
        n10319) );
  AND4_X1 U11459 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10376) );
  AOI22_X1 U11460 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15365) );
  NAND2_X1 U11461 ( .A1(n20158), .A2(n20156), .ZN(n20220) );
  NAND2_X2 U11462 ( .A1(n18872), .A2(n18807), .ZN(n18868) );
  BUF_X2 U11463 ( .A(n15460), .Z(n15430) );
  CLKBUF_X3 U11464 ( .A(n11721), .Z(n12900) );
  AND2_X2 U11465 ( .A1(n11718), .A2(n11537), .ZN(n12729) );
  NOR2_X1 U11466 ( .A1(n12943), .A2(n16325), .ZN(n12945) );
  CLKBUF_X2 U11467 ( .A(n15460), .Z(n17273) );
  AND2_X2 U11468 ( .A1(n16569), .A2(n19913), .ZN(n16642) );
  NAND2_X2 U11469 ( .A1(n19969), .A2(n19866), .ZN(n19915) );
  OAI21_X2 U11470 ( .B1(n12925), .B2(n12924), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n19268) );
  INV_X2 U11471 ( .A(n20845), .ZN(n20799) );
  NAND2_X1 U11472 ( .A1(n10279), .A2(n13359), .ZN(n11199) );
  AND2_X2 U11473 ( .A1(n11540), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11721) );
  AND2_X1 U11474 ( .A1(n10285), .A2(n10288), .ZN(n10415) );
  CLKBUF_X1 U11475 ( .A(n11551), .Z(n12802) );
  OR2_X1 U11476 ( .A1(n15357), .A2(n18741), .ZN(n16993) );
  BUF_X4 U11477 ( .A(n15495), .Z(n9743) );
  OR2_X1 U11478 ( .A1(n15355), .A2(n18741), .ZN(n9779) );
  NAND2_X1 U11479 ( .A1(n11542), .A2(n11532), .ZN(n12829) );
  NAND2_X1 U11480 ( .A1(n18896), .A2(n18886), .ZN(n15355) );
  NAND2_X1 U11481 ( .A1(n18903), .A2(n18910), .ZN(n17024) );
  NAND2_X1 U11482 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18896), .ZN(
        n15354) );
  NOR3_X2 U11483 ( .A1(n16976), .A2(n16978), .A3(n16485), .ZN(n17872) );
  AND2_X1 U11484 ( .A1(n14661), .A2(n10288), .ZN(n10419) );
  NAND2_X1 U11485 ( .A1(n14661), .A2(n10284), .ZN(n11168) );
  AND2_X1 U11486 ( .A1(n9966), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10287) );
  INV_X1 U11487 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18903) );
  INV_X2 U11488 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18896) );
  INV_X1 U11489 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18886) );
  NAND2_X2 U11490 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18741) );
  INV_X1 U11491 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13353) );
  NOR2_X2 U11492 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14661) );
  AND2_X2 U11493 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10286) );
  OAI211_X1 U11494 ( .C1(n12465), .C2(n11750), .A(n12251), .B(n11741), .ZN(
        n11784) );
  NAND2_X1 U11495 ( .A1(n9745), .A2(n12464), .ZN(n11789) );
  NAND2_X1 U11496 ( .A1(n11771), .A2(n12587), .ZN(n11772) );
  NOR2_X2 U11497 ( .A1(n9966), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13359) );
  NAND2_X1 U11498 ( .A1(n11753), .A2(n11752), .ZN(n12249) );
  XNOR2_X1 U11499 ( .A(n15681), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17932) );
  OR2_X2 U11500 ( .A1(n14247), .A2(n10073), .ZN(n9774) );
  XNOR2_X2 U11501 ( .A(n11391), .B(n11390), .ZN(n14525) );
  AOI21_X2 U11502 ( .B1(n16942), .B2(n17708), .A(n16849), .ZN(n16817) );
  NOR2_X2 U11503 ( .A1(n17849), .A2(n17767), .ZN(n17782) );
  NAND2_X2 U11504 ( .A1(n20599), .A2(n10548), .ZN(n14182) );
  INV_X2 U11505 ( .A(n11199), .ZN(n11125) );
  NAND2_X1 U11506 ( .A1(n11789), .A2(n11772), .ZN(n11803) );
  INV_X2 U11507 ( .A(n13935), .ZN(n14876) );
  NOR2_X2 U11508 ( .A1(n13570), .A2(n13571), .ZN(n13803) );
  NOR2_X2 U11509 ( .A1(n13217), .A2(n13218), .ZN(n13216) );
  NAND2_X1 U11510 ( .A1(n12246), .A2(n9746), .ZN(n11770) );
  INV_X1 U11511 ( .A(n11744), .ZN(n12169) );
  OR2_X1 U11512 ( .A1(n12794), .A2(n12793), .ZN(n10265) );
  NAND2_X1 U11513 ( .A1(n13119), .A2(n13118), .ZN(n10168) );
  AOI21_X1 U11514 ( .B1(n11803), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11807), .ZN(n11817) );
  NAND2_X1 U11515 ( .A1(n11789), .A2(n11772), .ZN(n9747) );
  NAND2_X1 U11516 ( .A1(n10168), .A2(n10166), .ZN(n12630) );
  NAND2_X1 U11517 ( .A1(n14952), .A2(n14948), .ZN(n9864) );
  NAND2_X1 U11518 ( .A1(n20192), .A2(n13428), .ZN(n11307) );
  NAND2_X1 U11519 ( .A1(n10054), .A2(n10267), .ZN(n14908) );
  NOR2_X2 U11520 ( .A1(n12842), .A2(n12841), .ZN(n12861) );
  NOR2_X2 U11521 ( .A1(n14739), .A2(n12818), .ZN(n12842) );
  NOR2_X2 U11522 ( .A1(n15017), .A2(n14999), .ZN(n15000) );
  XNOR2_X2 U11523 ( .A(n12794), .B(n12790), .ZN(n14749) );
  AND2_X1 U11524 ( .A1(n11538), .A2(n11795), .ZN(n9749) );
  AND2_X1 U11525 ( .A1(n11538), .A2(n11795), .ZN(n9750) );
  XNOR2_X2 U11526 ( .A(n12210), .B(n12318), .ZN(n13835) );
  NAND2_X2 U11527 ( .A1(n10189), .A2(n10188), .ZN(n12210) );
  INV_X1 U11528 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16978) );
  NAND2_X1 U11529 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16976) );
  NAND2_X2 U11530 ( .A1(n12009), .A2(n12008), .ZN(n15076) );
  NOR4_X2 U11531 ( .A1(n16700), .A2(n16699), .A3(n17006), .A4(n18787), .ZN(
        n16691) );
  INV_X2 U11532 ( .A(n12829), .ZN(n11672) );
  AOI21_X2 U11533 ( .B1(n9778), .B2(n14970), .A(n14969), .ZN(n15039) );
  AND2_X2 U11534 ( .A1(n10008), .A2(n10009), .ZN(n9778) );
  XOR2_X1 U11535 ( .A(n16689), .B(n16486), .Z(n9751) );
  NAND2_X1 U11536 ( .A1(n11820), .A2(n11826), .ZN(n11843) );
  NOR2_X4 U11537 ( .A1(n14225), .A2(n10243), .ZN(n14144) );
  NAND2_X2 U11538 ( .A1(n14239), .A2(n14236), .ZN(n14225) );
  NAND2_X2 U11540 ( .A1(n18944), .A2(n18933), .ZN(n18148) );
  AOI21_X1 U11541 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19933), .A(
        n11610), .ZN(n12138) );
  AND3_X1 U11542 ( .A1(n10286), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n10581), .ZN(n10382) );
  NOR2_X1 U11543 ( .A1(n10517), .A2(n10516), .ZN(n11428) );
  AND2_X1 U11544 ( .A1(n11608), .A2(n11607), .ZN(n11610) );
  NAND2_X1 U11545 ( .A1(n11944), .A2(n11943), .ZN(n11999) );
  OAI22_X1 U11546 ( .A1(n11917), .A2(n11890), .B1(n19733), .B2(n11889), .ZN(
        n11891) );
  NOR2_X1 U11547 ( .A1(n9806), .A2(n9980), .ZN(n9979) );
  INV_X1 U11548 ( .A(n9981), .ZN(n9980) );
  OR2_X1 U11549 ( .A1(n14070), .A2(n14069), .ZN(n11162) );
  NOR2_X1 U11550 ( .A1(n14203), .A2(n9982), .ZN(n9981) );
  INV_X1 U11551 ( .A(n14209), .ZN(n9982) );
  OR2_X1 U11552 ( .A1(n14027), .A2(n20260), .ZN(n11186) );
  NOR2_X1 U11553 ( .A1(n10090), .A2(n9929), .ZN(n9927) );
  INV_X1 U11554 ( .A(n11501), .ZN(n9929) );
  NOR2_X1 U11555 ( .A1(n14271), .A2(n10071), .ZN(n10070) );
  INV_X1 U11556 ( .A(n13956), .ZN(n10071) );
  AOI21_X1 U11557 ( .B1(n11426), .B2(n11469), .A(n9916), .ZN(n9915) );
  NAND2_X1 U11558 ( .A1(n20830), .A2(n11426), .ZN(n9917) );
  NAND2_X1 U11559 ( .A1(n10520), .A2(n13428), .ZN(n11260) );
  NAND2_X1 U11560 ( .A1(n10019), .A2(n9879), .ZN(n9877) );
  NAND2_X1 U11561 ( .A1(n10020), .A2(n9879), .ZN(n9878) );
  AOI221_X1 U11562 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11233), 
        .C1(n16169), .C2(n11233), .A(n11232), .ZN(n11275) );
  NAND2_X1 U11563 ( .A1(n10019), .A2(n9883), .ZN(n9881) );
  NOR2_X1 U11564 ( .A1(n11954), .A2(n11957), .ZN(n11953) );
  NOR2_X1 U11565 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U11566 ( .A1(n12624), .A2(n12623), .ZN(n12628) );
  AND2_X1 U11567 ( .A1(n12131), .A2(n12130), .ZN(n12331) );
  NOR2_X1 U11568 ( .A1(n10137), .A2(n14744), .ZN(n10136) );
  INV_X1 U11569 ( .A(n14731), .ZN(n10137) );
  NAND2_X1 U11570 ( .A1(n10059), .A2(n12042), .ZN(n10057) );
  NOR2_X1 U11571 ( .A1(n14973), .A2(n10006), .ZN(n10005) );
  INV_X1 U11572 ( .A(n15025), .ZN(n10006) );
  NOR2_X1 U11573 ( .A1(n14973), .A2(n10007), .ZN(n10004) );
  NOR2_X1 U11574 ( .A1(n16282), .A2(n10061), .ZN(n10060) );
  INV_X1 U11575 ( .A(n15058), .ZN(n10061) );
  NOR2_X1 U11576 ( .A1(n10013), .A2(n12042), .ZN(n10012) );
  INV_X1 U11577 ( .A(n10017), .ZN(n10013) );
  INV_X1 U11578 ( .A(n13557), .ZN(n10142) );
  INV_X1 U11579 ( .A(n10195), .ZN(n10194) );
  INV_X1 U11580 ( .A(n10196), .ZN(n10193) );
  AND4_X1 U11581 ( .A1(n11655), .A2(n11654), .A3(n11653), .A4(n11652), .ZN(
        n11656) );
  OR2_X1 U11582 ( .A1(n12197), .A2(n12194), .ZN(n12195) );
  OR2_X1 U11583 ( .A1(n17024), .A2(n15357), .ZN(n15493) );
  NOR2_X1 U11584 ( .A1(n15352), .A2(n15357), .ZN(n15495) );
  NOR2_X1 U11585 ( .A1(n15354), .A2(n17024), .ZN(n15418) );
  NOR2_X1 U11586 ( .A1(n15352), .A2(n15354), .ZN(n15602) );
  NOR2_X1 U11587 ( .A1(n17458), .A2(n15666), .ZN(n15664) );
  NOR2_X1 U11588 ( .A1(n18316), .A2(n18294), .ZN(n15566) );
  NAND2_X1 U11589 ( .A1(n17920), .A2(n15683), .ZN(n15686) );
  INV_X1 U11590 ( .A(n15715), .ZN(n15577) );
  AOI21_X1 U11591 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21010), .A(
        n15440), .ZN(n15576) );
  OR2_X1 U11592 ( .A1(n14032), .A2(n13299), .ZN(n13332) );
  NOR2_X1 U11593 ( .A1(n14057), .A2(n14044), .ZN(n14043) );
  NAND2_X1 U11594 ( .A1(n16020), .A2(n11494), .ZN(n10080) );
  AND2_X1 U11595 ( .A1(n14032), .A2(n13422), .ZN(n15805) );
  NAND2_X1 U11596 ( .A1(n14356), .A2(n14501), .ZN(n9921) );
  AND2_X2 U11597 ( .A1(n14125), .A2(n10065), .ZN(n14068) );
  AND2_X1 U11598 ( .A1(n9768), .A2(n14066), .ZN(n10065) );
  NAND2_X1 U11599 ( .A1(n14575), .A2(n16064), .ZN(n14522) );
  INV_X1 U11600 ( .A(n11423), .ZN(n14417) );
  NAND2_X1 U11601 ( .A1(n19975), .A2(n9880), .ZN(n11520) );
  AND2_X1 U11602 ( .A1(n13421), .A2(n13420), .ZN(n13438) );
  OR2_X1 U11603 ( .A1(n16445), .A2(n16443), .ZN(n13200) );
  AND2_X1 U11604 ( .A1(n12114), .A2(n9781), .ZN(n12109) );
  NAND2_X1 U11605 ( .A1(n12092), .A2(n12114), .ZN(n12048) );
  NAND2_X1 U11606 ( .A1(n12968), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12967) );
  NAND2_X1 U11607 ( .A1(n12221), .A2(n13834), .ZN(n12224) );
  NAND2_X1 U11608 ( .A1(n13672), .A2(n13647), .ZN(n10046) );
  AND2_X1 U11609 ( .A1(n19565), .A2(n19953), .ZN(n19471) );
  INV_X1 U11610 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19509) );
  INV_X1 U11611 ( .A(n17451), .ZN(n16545) );
  OR2_X1 U11612 ( .A1(n16484), .A2(n18757), .ZN(n9958) );
  NAND2_X1 U11613 ( .A1(n18750), .A2(n9960), .ZN(n9959) );
  NOR2_X1 U11614 ( .A1(n13200), .A2(n16479), .ZN(n18951) );
  NOR2_X1 U11615 ( .A1(n11256), .A2(n11240), .ZN(n11247) );
  INV_X1 U11616 ( .A(n10635), .ZN(n10634) );
  NAND2_X1 U11617 ( .A1(n19940), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11529) );
  AND2_X1 U11618 ( .A1(n13342), .A2(n11519), .ZN(n13324) );
  INV_X1 U11619 ( .A(n10566), .ZN(n9978) );
  OR2_X1 U11620 ( .A1(n13428), .A2(n9880), .ZN(n10586) );
  OR2_X1 U11621 ( .A1(n13435), .A2(n9880), .ZN(n11243) );
  OR2_X1 U11622 ( .A1(n20851), .A2(n20199), .ZN(n10432) );
  NAND2_X1 U11623 ( .A1(n9901), .A2(n9898), .ZN(n9897) );
  AOI21_X1 U11624 ( .B1(n11248), .B2(n9903), .A(n9902), .ZN(n9901) );
  OAI21_X1 U11625 ( .B1(n11248), .B2(n9903), .A(n9899), .ZN(n9898) );
  NOR2_X1 U11626 ( .A1(n11241), .A2(n9792), .ZN(n9903) );
  INV_X1 U11627 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U11628 ( .A1(n11243), .A2(n10586), .ZN(n11256) );
  NAND2_X1 U11629 ( .A1(n11742), .A2(n12169), .ZN(n12167) );
  XNOR2_X1 U11630 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11607) );
  AND2_X1 U11631 ( .A1(n9831), .A2(n10163), .ZN(n10162) );
  INV_X1 U11632 ( .A(n14826), .ZN(n10163) );
  OAI211_X1 U11633 ( .C1(n11804), .C2(n13764), .A(n11778), .B(n10043), .ZN(
        n11779) );
  NOR2_X1 U11634 ( .A1(n12929), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12282) );
  AND2_X1 U11635 ( .A1(n11744), .A2(n11732), .ZN(n11739) );
  AND4_X1 U11636 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n11684) );
  NOR2_X1 U11637 ( .A1(n17466), .A2(n15668), .ZN(n15667) );
  NAND2_X1 U11638 ( .A1(n17450), .A2(n18277), .ZN(n15556) );
  AOI21_X1 U11639 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18725), .A(
        n15437), .ZN(n15446) );
  AND2_X1 U11640 ( .A1(n15575), .A2(n15574), .ZN(n15437) );
  AOI22_X1 U11641 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18746), .B2(n18896), .ZN(
        n15445) );
  NAND2_X1 U11642 ( .A1(n20214), .A2(n20199), .ZN(n14016) );
  INV_X1 U11643 ( .A(n14101), .ZN(n10067) );
  NAND2_X1 U11644 ( .A1(n10247), .A2(n10910), .ZN(n10246) );
  INV_X1 U11645 ( .A(n14220), .ZN(n10247) );
  NAND2_X1 U11646 ( .A1(n14656), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11221) );
  INV_X1 U11647 ( .A(n11221), .ZN(n11188) );
  INV_X1 U11648 ( .A(n11279), .ZN(n11224) );
  INV_X1 U11649 ( .A(n11490), .ZN(n11496) );
  OR2_X1 U11650 ( .A1(n12998), .A2(n20260), .ZN(n10816) );
  INV_X1 U11651 ( .A(n13563), .ZN(n9974) );
  NOR2_X2 U11652 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11279) );
  NAND2_X1 U11653 ( .A1(n10077), .A2(n14229), .ZN(n10076) );
  INV_X1 U11654 ( .A(n14242), .ZN(n10077) );
  INV_X1 U11655 ( .A(n14233), .ZN(n10078) );
  INV_X1 U11656 ( .A(n14266), .ZN(n10069) );
  NAND2_X1 U11657 ( .A1(n13303), .A2(n11383), .ZN(n11381) );
  OAI21_X1 U11658 ( .B1(n11427), .B2(n20177), .A(n11431), .ZN(n11433) );
  AND2_X1 U11659 ( .A1(n13435), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U11660 ( .A1(n10286), .A2(n10284), .ZN(n10507) );
  NAND2_X1 U11661 ( .A1(n10580), .A2(n10579), .ZN(n10605) );
  NOR2_X1 U11662 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10224), .ZN(n10223) );
  NAND2_X1 U11663 ( .A1(n12512), .A2(n12516), .ZN(n10224) );
  NAND2_X1 U11664 ( .A1(n10179), .A2(n10177), .ZN(n10176) );
  INV_X1 U11665 ( .A(n14771), .ZN(n10177) );
  NOR2_X1 U11666 ( .A1(n9817), .A2(n10180), .ZN(n10179) );
  INV_X1 U11667 ( .A(n14780), .ZN(n10180) );
  NOR2_X1 U11668 ( .A1(n16308), .A2(n10123), .ZN(n10122) );
  INV_X1 U11669 ( .A(n13312), .ZN(n10131) );
  INV_X1 U11670 ( .A(n11999), .ZN(n11945) );
  AOI21_X1 U11671 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11815), .ZN(n12498) );
  INV_X1 U11672 ( .A(n10165), .ZN(n9853) );
  NAND2_X1 U11673 ( .A1(n9864), .A2(n9805), .ZN(n12122) );
  AND2_X1 U11674 ( .A1(n12116), .A2(n14929), .ZN(n10225) );
  NOR2_X1 U11675 ( .A1(n10235), .A2(n10237), .ZN(n10227) );
  NAND2_X1 U11676 ( .A1(n10236), .A2(n10266), .ZN(n10235) );
  INV_X1 U11677 ( .A(n14961), .ZN(n10236) );
  AND2_X1 U11678 ( .A1(n12075), .A2(n10060), .ZN(n10059) );
  AND2_X1 U11679 ( .A1(n12074), .A2(n12073), .ZN(n12075) );
  AND2_X1 U11680 ( .A1(n10005), .A2(n14998), .ZN(n10003) );
  NAND2_X1 U11681 ( .A1(n10160), .A2(n10159), .ZN(n10158) );
  INV_X1 U11682 ( .A(n13509), .ZN(n10159) );
  INV_X1 U11683 ( .A(n13584), .ZN(n10140) );
  NAND2_X1 U11684 ( .A1(n9868), .A2(n9866), .ZN(n10014) );
  AND2_X1 U11685 ( .A1(n10015), .A2(n9867), .ZN(n9866) );
  INV_X1 U11686 ( .A(n15313), .ZN(n9868) );
  INV_X1 U11687 ( .A(n15310), .ZN(n9867) );
  NOR2_X1 U11688 ( .A1(n10018), .A2(n9833), .ZN(n10017) );
  INV_X1 U11689 ( .A(n16298), .ZN(n10018) );
  NOR2_X1 U11690 ( .A1(n11644), .A2(n11643), .ZN(n12326) );
  INV_X1 U11691 ( .A(n13167), .ZN(n10127) );
  NAND2_X1 U11692 ( .A1(n10049), .A2(n10050), .ZN(n10047) );
  NAND2_X1 U11693 ( .A1(n11817), .A2(n11810), .ZN(n11811) );
  INV_X1 U11694 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11795) );
  AND2_X1 U11695 ( .A1(n11785), .A2(n11774), .ZN(n11749) );
  INV_X1 U11696 ( .A(n12450), .ZN(n12459) );
  OR2_X1 U11697 ( .A1(n12812), .A2(n12606), .ZN(n12615) );
  AND2_X1 U11698 ( .A1(n21158), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12619) );
  OR3_X1 U11699 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18903), .A3(
        n15539), .ZN(n17288) );
  NOR2_X1 U11700 ( .A1(n9954), .A2(n9952), .ZN(n9951) );
  INV_X1 U11701 ( .A(n15638), .ZN(n9954) );
  NOR2_X1 U11702 ( .A1(n15732), .A2(n17845), .ZN(n15700) );
  INV_X1 U11703 ( .A(n18287), .ZN(n15551) );
  NAND2_X1 U11704 ( .A1(n15735), .A2(n18171), .ZN(n9949) );
  NAND2_X1 U11705 ( .A1(n17873), .A2(n15694), .ZN(n15695) );
  NOR4_X1 U11706 ( .A1(n15548), .A2(n15712), .A3(n15556), .A4(n15711), .ZN(
        n15565) );
  AND2_X1 U11707 ( .A1(n15565), .A2(n15551), .ZN(n15567) );
  AOI21_X1 U11708 ( .B1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B2(n15595), .A(
        n9992), .ZN(n9991) );
  INV_X1 U11709 ( .A(n15413), .ZN(n9992) );
  INV_X1 U11710 ( .A(n15411), .ZN(n9993) );
  NOR2_X1 U11711 ( .A1(n15564), .A2(n15550), .ZN(n15724) );
  AND2_X1 U11712 ( .A1(n18310), .A2(n15712), .ZN(n15572) );
  NAND2_X1 U11713 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n9965) );
  NOR2_X1 U11714 ( .A1(n15727), .A2(n18752), .ZN(n15580) );
  NAND2_X1 U11715 ( .A1(n18928), .A2(n15573), .ZN(n17483) );
  NOR2_X1 U11716 ( .A1(n10361), .A2(n10360), .ZN(n10377) );
  INV_X1 U11717 ( .A(n11186), .ZN(n11226) );
  NAND2_X1 U11718 ( .A1(n14144), .A2(n9793), .ZN(n14057) );
  OR2_X1 U11719 ( .A1(n11139), .A2(n11138), .ZN(n11163) );
  INV_X1 U11720 ( .A(n10252), .ZN(n10250) );
  NAND2_X1 U11721 ( .A1(n10944), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10987) );
  AND2_X1 U11722 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10641), .ZN(
        n10668) );
  NAND2_X1 U11723 ( .A1(n9928), .A2(n16009), .ZN(n14594) );
  AOI211_X1 U11724 ( .C1(n11513), .C2(n11512), .A(n10086), .B(n10085), .ZN(
        n10084) );
  NAND2_X1 U11725 ( .A1(n14455), .A2(n10087), .ZN(n10085) );
  AND2_X1 U11726 ( .A1(n9906), .A2(n9905), .ZN(n14513) );
  NAND2_X1 U11727 ( .A1(n14626), .A2(n9916), .ZN(n9906) );
  INV_X1 U11728 ( .A(n10083), .ZN(n10091) );
  NAND2_X1 U11729 ( .A1(n10083), .A2(n11512), .ZN(n10088) );
  NOR2_X1 U11730 ( .A1(n14489), .A2(n9893), .ZN(n15994) );
  NAND2_X1 U11731 ( .A1(n14487), .A2(n14484), .ZN(n9893) );
  NAND2_X1 U11732 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15995) );
  NAND2_X1 U11733 ( .A1(n16031), .A2(n9885), .ZN(n9887) );
  INV_X1 U11734 ( .A(n11476), .ZN(n9924) );
  INV_X1 U11735 ( .A(n16131), .ZN(n16113) );
  OR2_X1 U11736 ( .A1(n13438), .A2(n20135), .ZN(n9905) );
  NAND2_X1 U11737 ( .A1(n10585), .A2(n10584), .ZN(n20322) );
  NAND2_X1 U11738 ( .A1(n9907), .A2(n11268), .ZN(n14032) );
  OAI21_X1 U11739 ( .B1(n11265), .B2(n11264), .A(n9908), .ZN(n9907) );
  NAND2_X1 U11740 ( .A1(n20815), .A2(n20812), .ZN(n20294) );
  NAND2_X1 U11741 ( .A1(n10547), .A2(n10546), .ZN(n20599) );
  NOR2_X1 U11742 ( .A1(n20489), .A2(n20328), .ZN(n20651) );
  OR2_X1 U11743 ( .A1(n20688), .A2(n20609), .ZN(n20645) );
  NAND2_X1 U11744 ( .A1(n20431), .A2(n10604), .ZN(n20688) );
  AOI21_X1 U11745 ( .B1(n20834), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20328), 
        .ZN(n20689) );
  NAND2_X1 U11746 ( .A1(n9880), .A2(n20161), .ZN(n20328) );
  AND2_X1 U11747 ( .A1(n11284), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15819) );
  AOI221_X1 U11748 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12138), 
        .C1(n15589), .C2(n12138), .A(n12137), .ZN(n12197) );
  NAND2_X1 U11749 ( .A1(n12015), .A2(n12331), .ZN(n12114) );
  NOR2_X1 U11750 ( .A1(n12096), .A2(n10222), .ZN(n10221) );
  INV_X1 U11751 ( .A(n11665), .ZN(n10222) );
  NAND2_X1 U11752 ( .A1(n10214), .A2(n9766), .ZN(n12092) );
  INV_X1 U11753 ( .A(n12051), .ZN(n10214) );
  NOR2_X1 U11754 ( .A1(n10211), .A2(n12059), .ZN(n10210) );
  INV_X1 U11755 ( .A(n10212), .ZN(n10211) );
  AND2_X1 U11756 ( .A1(n13548), .A2(n13546), .ZN(n13547) );
  OR2_X1 U11757 ( .A1(n13511), .A2(n12633), .ZN(n13523) );
  NAND2_X1 U11758 ( .A1(n10257), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10174) );
  AND2_X1 U11759 ( .A1(n12839), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13163) );
  NAND2_X1 U11760 ( .A1(n9834), .A2(n10136), .ZN(n10135) );
  INV_X1 U11761 ( .A(n12979), .ZN(n10138) );
  OR2_X1 U11762 ( .A1(n16209), .A2(n10051), .ZN(n14909) );
  NAND2_X1 U11763 ( .A1(n10197), .A2(n10198), .ZN(n14933) );
  NOR2_X1 U11764 ( .A1(n14963), .A2(n13976), .ZN(n14945) );
  NOR2_X1 U11765 ( .A1(n14961), .A2(n14959), .ZN(n10232) );
  NAND2_X1 U11766 ( .A1(n12090), .A2(n10234), .ZN(n10233) );
  INV_X1 U11767 ( .A(n10235), .ZN(n10234) );
  NAND2_X1 U11768 ( .A1(n10062), .A2(n10059), .ZN(n12090) );
  INV_X1 U11769 ( .A(n10001), .ZN(n15017) );
  NAND2_X1 U11770 ( .A1(n10010), .A2(n10060), .ZN(n10009) );
  INV_X1 U11771 ( .A(n10012), .ZN(n10010) );
  NAND2_X1 U11772 ( .A1(n10014), .A2(n10012), .ZN(n10062) );
  NOR2_X1 U11773 ( .A1(n13373), .A2(n10161), .ZN(n10160) );
  INV_X1 U11774 ( .A(n15300), .ZN(n10161) );
  NAND2_X1 U11775 ( .A1(n13216), .A2(n13262), .ZN(n13372) );
  NAND2_X1 U11776 ( .A1(n10192), .A2(n10195), .ZN(n15084) );
  NAND2_X1 U11777 ( .A1(n15329), .A2(n10196), .ZN(n10192) );
  AOI21_X1 U11778 ( .B1(n13647), .B2(n12131), .A(n12264), .ZN(n10049) );
  INV_X1 U11779 ( .A(n10189), .ZN(n11950) );
  INV_X1 U11780 ( .A(n10188), .ZN(n11949) );
  AND4_X1 U11781 ( .A1(n11648), .A2(n11647), .A3(n11646), .A4(n11645), .ZN(
        n11659) );
  OAI21_X1 U11782 ( .B1(n11801), .B2(n11795), .A(n11794), .ZN(n11823) );
  NOR2_X1 U11783 ( .A1(n11793), .A2(n11792), .ZN(n11794) );
  NAND2_X1 U11784 ( .A1(n11804), .A2(n11791), .ZN(n11792) );
  INV_X1 U11785 ( .A(n11789), .ZN(n11793) );
  NAND2_X1 U11786 ( .A1(n12600), .A2(n19509), .ZN(n12622) );
  INV_X1 U11787 ( .A(n12939), .ZN(n19108) );
  AND2_X1 U11788 ( .A1(n13078), .A2(n12614), .ZN(n13173) );
  NAND2_X1 U11789 ( .A1(n13174), .A2(n13173), .ZN(n13172) );
  AND2_X1 U11790 ( .A1(n19936), .A2(n19925), .ZN(n19923) );
  NOR2_X1 U11791 ( .A1(n13098), .A2(n11820), .ZN(n10239) );
  BUF_X1 U11792 ( .A(n11765), .Z(n19302) );
  INV_X1 U11793 ( .A(n19782), .ZN(n19723) );
  NOR2_X1 U11794 ( .A1(n19936), .A2(n19943), .ZN(n19782) );
  AOI22_X2 U11795 ( .A1(n21158), .A2(n16474), .B1(n15857), .B2(n15856), .ZN(
        n19778) );
  NAND2_X1 U11796 ( .A1(n18277), .A2(n18929), .ZN(n15726) );
  NOR2_X1 U11797 ( .A1(n17479), .A2(n9995), .ZN(n9994) );
  NOR2_X1 U11798 ( .A1(n17555), .A2(n9997), .ZN(n9996) );
  NOR2_X1 U11799 ( .A1(n18736), .A2(n9988), .ZN(n15859) );
  AND2_X1 U11800 ( .A1(n17523), .A2(n18929), .ZN(n9988) );
  OAI21_X1 U11801 ( .B1(n15578), .B2(n15577), .A(n15576), .ZN(n18749) );
  INV_X1 U11802 ( .A(n18277), .ZN(n17485) );
  AND2_X1 U11803 ( .A1(n17638), .A2(n10093), .ZN(n10095) );
  NOR2_X1 U11804 ( .A1(n10094), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10093) );
  INV_X1 U11805 ( .A(n9832), .ZN(n10094) );
  NAND2_X1 U11806 ( .A1(n15707), .A2(n17856), .ZN(n15708) );
  NOR2_X1 U11807 ( .A1(n18090), .A2(n17615), .ZN(n17946) );
  NAND2_X1 U11808 ( .A1(n10096), .A2(n10095), .ZN(n17619) );
  OR2_X1 U11809 ( .A1(n17639), .A2(n17626), .ZN(n10096) );
  INV_X1 U11810 ( .A(n18135), .ZN(n17808) );
  NAND2_X1 U11811 ( .A1(n18739), .A2(n18722), .ZN(n15734) );
  NOR2_X1 U11812 ( .A1(n15548), .A2(n15551), .ZN(n15730) );
  INV_X1 U11813 ( .A(n18168), .ZN(n9962) );
  XNOR2_X1 U11814 ( .A(n15686), .B(n15685), .ZN(n17912) );
  NAND2_X1 U11815 ( .A1(n15724), .A2(n15723), .ZN(n18757) );
  AND2_X1 U11816 ( .A1(n18730), .A2(n9989), .ZN(n18736) );
  INV_X1 U11817 ( .A(n15728), .ZN(n9989) );
  NAND2_X1 U11818 ( .A1(n13625), .A2(n13046), .ZN(n20846) );
  INV_X1 U11819 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20814) );
  INV_X1 U11820 ( .A(n14182), .ZN(n20647) );
  AND2_X1 U11821 ( .A1(n16037), .A2(n20131), .ZN(n16033) );
  AND2_X2 U11822 ( .A1(n11420), .A2(n20813), .ZN(n20158) );
  XNOR2_X1 U11823 ( .A(n9888), .B(n20899), .ZN(n9896) );
  NAND2_X1 U11824 ( .A1(n9889), .A2(n9919), .ZN(n9888) );
  NAND2_X1 U11825 ( .A1(n9920), .A2(n9824), .ZN(n9889) );
  OR2_X1 U11826 ( .A1(n14068), .A2(n14067), .ZN(n14561) );
  XNOR2_X1 U11827 ( .A(n14382), .B(n14381), .ZN(n14562) );
  NAND2_X1 U11828 ( .A1(n16054), .A2(n14531), .ZN(n14518) );
  OAI21_X1 U11829 ( .B1(n20830), .B2(n11469), .A(n11426), .ZN(n20128) );
  AND2_X1 U11830 ( .A1(n13438), .A2(n13437), .ZN(n20145) );
  INV_X1 U11831 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20834) );
  CLKBUF_X1 U11832 ( .A(n13445), .Z(n13446) );
  OR2_X1 U11833 ( .A1(n13045), .A2(n13044), .ZN(n13092) );
  OAI21_X1 U11834 ( .B1(n12990), .B2(n19090), .A(n10147), .ZN(n10146) );
  INV_X1 U11835 ( .A(n12989), .ZN(n10147) );
  OR2_X1 U11836 ( .A1(n15112), .A2(n19105), .ZN(n10148) );
  NAND2_X1 U11837 ( .A1(n10113), .A2(n16195), .ZN(n10109) );
  OR2_X1 U11838 ( .A1(n10110), .A2(n10108), .ZN(n10107) );
  INV_X1 U11839 ( .A(n16195), .ZN(n10108) );
  NAND2_X1 U11840 ( .A1(n12913), .A2(n19838), .ZN(n12914) );
  NAND2_X1 U11841 ( .A1(n10183), .A2(n10182), .ZN(n13992) );
  NAND2_X1 U11842 ( .A1(n9914), .A2(n9851), .ZN(n10183) );
  OAI21_X1 U11843 ( .B1(n14916), .B2(n10185), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10182) );
  XNOR2_X1 U11844 ( .A(n9857), .B(n9815), .ZN(n13994) );
  NAND2_X1 U11845 ( .A1(n9858), .A2(n9813), .ZN(n9857) );
  AND2_X1 U11846 ( .A1(n12598), .A2(n19962), .ZN(n16400) );
  AND2_X1 U11847 ( .A1(n12598), .A2(n19963), .ZN(n16423) );
  NAND2_X1 U11848 ( .A1(n12598), .A2(n12597), .ZN(n16388) );
  NAND2_X1 U11849 ( .A1(n13084), .A2(n13083), .ZN(n19953) );
  INV_X1 U11850 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19933) );
  NAND2_X1 U11851 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17308), .ZN(n17302) );
  NOR2_X1 U11852 ( .A1(n15601), .A2(n15600), .ZN(n17451) );
  NAND2_X1 U11853 ( .A1(n16530), .A2(n10104), .ZN(n10103) );
  OR2_X1 U11854 ( .A1(n16554), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10104) );
  INV_X1 U11855 ( .A(n10106), .ZN(n10105) );
  AOI21_X1 U11856 ( .B1(n16558), .B2(n16531), .A(n16532), .ZN(n10106) );
  NAND3_X1 U11857 ( .A1(n16675), .A2(n17940), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n17786) );
  NOR2_X2 U11858 ( .A1(n17451), .A2(n17943), .ZN(n17857) );
  NAND2_X1 U11859 ( .A1(n9934), .A2(n9930), .ZN(n16541) );
  NAND2_X1 U11860 ( .A1(n9935), .A2(n16496), .ZN(n9934) );
  NAND2_X1 U11861 ( .A1(n9932), .A2(n9931), .ZN(n9930) );
  NAND2_X1 U11862 ( .A1(n9937), .A2(n9936), .ZN(n9935) );
  XNOR2_X1 U11863 ( .A(n15710), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16529) );
  INV_X1 U11864 ( .A(n18258), .ZN(n18251) );
  NOR2_X1 U11865 ( .A1(n18117), .A2(n18217), .ZN(n18258) );
  INV_X1 U11866 ( .A(n10636), .ZN(n10021) );
  NOR2_X1 U11867 ( .A1(n9797), .A2(n9900), .ZN(n9899) );
  INV_X1 U11868 ( .A(n11270), .ZN(n9900) );
  INV_X1 U11869 ( .A(n11254), .ZN(n9902) );
  OAI21_X1 U11870 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18896), .A(
        n15438), .ZN(n15439) );
  OR2_X1 U11871 ( .A1(n15445), .A2(n15446), .ZN(n15438) );
  AND2_X1 U11872 ( .A1(n10633), .A2(n10632), .ZN(n10635) );
  NAND2_X1 U11873 ( .A1(n10021), .A2(n10634), .ZN(n10666) );
  INV_X1 U11874 ( .A(n11512), .ZN(n10090) );
  NOR2_X1 U11875 ( .A1(n10481), .A2(n10480), .ZN(n11440) );
  NOR2_X1 U11876 ( .A1(n13370), .A2(n9880), .ZN(n9879) );
  OR2_X1 U11877 ( .A1(n10601), .A2(n10600), .ZN(n11457) );
  NOR2_X1 U11878 ( .A1(n13353), .A2(n9880), .ZN(n9883) );
  NAND2_X1 U11879 ( .A1(n10020), .A2(n9883), .ZN(n9882) );
  NOR2_X1 U11880 ( .A1(n14029), .A2(n10425), .ZN(n10429) );
  INV_X1 U11881 ( .A(n13436), .ZN(n10428) );
  NAND2_X1 U11882 ( .A1(n10019), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10457) );
  INV_X1 U11883 ( .A(n14755), .ZN(n10171) );
  INV_X1 U11884 ( .A(n14833), .ZN(n10164) );
  NOR2_X1 U11885 ( .A1(n16300), .A2(n10016), .ZN(n10015) );
  INV_X1 U11886 ( .A(n15069), .ZN(n10016) );
  INV_X1 U11887 ( .A(n15083), .ZN(n10191) );
  NAND2_X1 U11888 ( .A1(n11746), .A2(n11751), .ZN(n11747) );
  NAND2_X1 U11889 ( .A1(n12605), .A2(n15585), .ZN(n12812) );
  INV_X1 U11890 ( .A(n11763), .ZN(n11753) );
  AND2_X1 U11891 ( .A1(n11529), .A2(n11528), .ZN(n11605) );
  NAND2_X1 U11892 ( .A1(n17285), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n9953) );
  NAND2_X1 U11893 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18903), .ZN(
        n15356) );
  NOR2_X1 U11894 ( .A1(n17462), .A2(n15749), .ZN(n15739) );
  OR2_X1 U11895 ( .A1(n15551), .A2(n15572), .ZN(n15558) );
  INV_X1 U11896 ( .A(n11225), .ZN(n10886) );
  OAI22_X1 U11897 ( .A1(n9742), .A2(n10414), .B1(n9972), .B2(n11013), .ZN(
        n9967) );
  INV_X1 U11898 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10414) );
  INV_X1 U11899 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n9972) );
  NAND2_X1 U11900 ( .A1(n14105), .A2(n10252), .ZN(n10251) );
  NOR2_X1 U11901 ( .A1(n10253), .A2(n14135), .ZN(n10252) );
  AND2_X1 U11902 ( .A1(n10248), .A2(n13954), .ZN(n9983) );
  AND2_X1 U11903 ( .A1(n10818), .A2(n10249), .ZN(n10248) );
  OR2_X1 U11904 ( .A1(n14153), .A2(n14275), .ZN(n10249) );
  AND2_X1 U11905 ( .A1(n14261), .A2(n14157), .ZN(n10818) );
  INV_X1 U11906 ( .A(n14087), .ZN(n10066) );
  INV_X1 U11907 ( .A(n11517), .ZN(n10064) );
  NAND2_X1 U11908 ( .A1(n11517), .A2(n16009), .ZN(n14409) );
  INV_X1 U11909 ( .A(n14527), .ZN(n10087) );
  NAND2_X1 U11910 ( .A1(n14461), .A2(n9798), .ZN(n11513) );
  NAND2_X1 U11911 ( .A1(n14465), .A2(n11503), .ZN(n14484) );
  OR2_X1 U11912 ( .A1(n10502), .A2(n10501), .ZN(n11490) );
  INV_X1 U11913 ( .A(n16024), .ZN(n9925) );
  INV_X1 U11914 ( .A(n16030), .ZN(n9886) );
  INV_X1 U11915 ( .A(n16023), .ZN(n9923) );
  OR2_X1 U11916 ( .A1(n10540), .A2(n10539), .ZN(n11437) );
  AOI21_X1 U11917 ( .B1(n10568), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9978), 
        .ZN(n9977) );
  OAI21_X1 U11918 ( .B1(n10020), .B2(n10019), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n9884) );
  INV_X1 U11919 ( .A(n11260), .ZN(n11263) );
  AOI21_X1 U11920 ( .B1(n9897), .B2(n11259), .A(n9825), .ZN(n11261) );
  INV_X1 U11921 ( .A(n9909), .ZN(n9908) );
  OAI211_X1 U11922 ( .C1(n11273), .C2(n11266), .A(n11267), .B(n9910), .ZN(
        n9909) );
  NAND2_X1 U11923 ( .A1(n9880), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9910) );
  INV_X1 U11924 ( .A(n10604), .ZN(n20321) );
  INV_X1 U11925 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10352) );
  NOR2_X1 U11926 ( .A1(n10349), .A2(n9892), .ZN(n9891) );
  OR2_X1 U11927 ( .A1(n11610), .A2(n11609), .ZN(n12139) );
  NAND2_X1 U11928 ( .A1(n12135), .A2(n12110), .ZN(n12119) );
  NOR2_X1 U11929 ( .A1(n10220), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10219) );
  INV_X1 U11930 ( .A(n10221), .ZN(n10220) );
  OR2_X1 U11931 ( .A1(n11664), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U11932 ( .A1(n12043), .A2(n10213), .ZN(n10212) );
  INV_X1 U11933 ( .A(n12039), .ZN(n10213) );
  OR2_X1 U11934 ( .A1(n11632), .A2(n11631), .ZN(n11942) );
  NAND2_X1 U11935 ( .A1(n10207), .A2(n9799), .ZN(n11954) );
  NAND2_X1 U11936 ( .A1(n12152), .A2(n12130), .ZN(n10207) );
  AND2_X1 U11937 ( .A1(n12447), .A2(n12446), .ZN(n14826) );
  INV_X1 U11938 ( .A(n14784), .ZN(n10181) );
  NAND2_X1 U11939 ( .A1(n10117), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10116) );
  NOR2_X1 U11940 ( .A1(n19025), .A2(n14705), .ZN(n10117) );
  XNOR2_X1 U11941 ( .A(n14683), .B(n9842), .ZN(n12132) );
  NAND2_X1 U11942 ( .A1(n9865), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12125) );
  AND2_X1 U11943 ( .A1(n15182), .A2(n10162), .ZN(n14825) );
  NOR2_X1 U11944 ( .A1(n10200), .A2(n10199), .ZN(n10198) );
  NAND2_X1 U11945 ( .A1(n15182), .A2(n9831), .ZN(n14835) );
  OR2_X1 U11946 ( .A1(n16228), .A2(n10051), .ZN(n12123) );
  INV_X1 U11947 ( .A(n14949), .ZN(n9863) );
  NAND2_X1 U11948 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U11949 ( .A1(n10204), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10203) );
  INV_X1 U11950 ( .A(n10205), .ZN(n10204) );
  NAND2_X1 U11951 ( .A1(n12472), .A2(n15218), .ZN(n10205) );
  NOR2_X1 U11952 ( .A1(n13929), .A2(n13928), .ZN(n10144) );
  AND2_X1 U11953 ( .A1(n10060), .A2(n10015), .ZN(n10011) );
  AND2_X1 U11954 ( .A1(n12311), .A2(n10151), .ZN(n10150) );
  AND2_X1 U11955 ( .A1(n13531), .A2(n13535), .ZN(n10151) );
  INV_X1 U11956 ( .A(n12500), .ZN(n9854) );
  OR2_X1 U11957 ( .A1(n11798), .A2(n11797), .ZN(n11799) );
  NAND2_X1 U11958 ( .A1(n11790), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11791) );
  OR2_X1 U11959 ( .A1(n12812), .A2(n12612), .ZN(n12613) );
  AND2_X1 U11960 ( .A1(n13176), .A2(n13098), .ZN(n10052) );
  NAND2_X1 U11961 ( .A1(n10258), .A2(n10259), .ZN(n11689) );
  NAND3_X1 U11962 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19928), .A3(n19731), 
        .ZN(n19269) );
  NAND2_X1 U11963 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18910), .ZN(
        n15352) );
  OR2_X1 U11964 ( .A1(n15539), .A2(n18741), .ZN(n9775) );
  NAND2_X1 U11965 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .ZN(n9997) );
  NOR2_X1 U11966 ( .A1(n18910), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n15574) );
  NOR2_X1 U11967 ( .A1(n17333), .A2(n15558), .ZN(n15559) );
  NAND2_X1 U11968 ( .A1(n9943), .A2(n17792), .ZN(n9942) );
  INV_X1 U11969 ( .A(n16494), .ZN(n9943) );
  NAND2_X1 U11970 ( .A1(n9948), .A2(n17792), .ZN(n15699) );
  NAND2_X1 U11971 ( .A1(n17775), .A2(n10255), .ZN(n9948) );
  AND2_X1 U11972 ( .A1(n10100), .A2(n17841), .ZN(n10099) );
  AND2_X1 U11973 ( .A1(n17819), .A2(n10101), .ZN(n10100) );
  INV_X1 U11974 ( .A(n15726), .ZN(n9955) );
  NOR2_X1 U11975 ( .A1(n15755), .A2(n17886), .ZN(n15757) );
  AND2_X1 U11976 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15753), .ZN(
        n15755) );
  OAI22_X1 U11977 ( .A1(n18903), .A2(n18725), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15575) );
  AOI21_X1 U11978 ( .B1(n15446), .B2(n15445), .A(n15444), .ZN(n15715) );
  NAND2_X1 U11979 ( .A1(n18886), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15357) );
  NOR2_X1 U11980 ( .A1(n10943), .A2(n14450), .ZN(n10944) );
  OR2_X1 U11981 ( .A1(n20021), .A2(n14161), .ZN(n15944) );
  INV_X1 U11982 ( .A(n15944), .ZN(n15952) );
  NAND2_X1 U11983 ( .A1(n10724), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10741) );
  INV_X1 U11984 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20001) );
  NAND2_X1 U11985 ( .A1(n14125), .A2(n9830), .ZN(n14099) );
  AND2_X1 U11986 ( .A1(n14205), .A2(n14132), .ZN(n14130) );
  AND2_X1 U11987 ( .A1(n11368), .A2(n11367), .ZN(n14204) );
  NOR2_X1 U11988 ( .A1(n14214), .A2(n14204), .ZN(n14205) );
  AND2_X1 U11989 ( .A1(n11347), .A2(n11346), .ZN(n14242) );
  NAND2_X1 U11990 ( .A1(n12997), .A2(n12996), .ZN(n13322) );
  AND2_X1 U11991 ( .A1(n14032), .A2(n13142), .ZN(n20072) );
  OR2_X1 U11992 ( .A1(n11163), .A2(n20944), .ZN(n11282) );
  OR2_X1 U11993 ( .A1(n11142), .A2(n11141), .ZN(n14070) );
  NAND2_X1 U11994 ( .A1(n11137), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11159) );
  INV_X1 U11995 ( .A(n11157), .ZN(n11137) );
  NAND2_X1 U11996 ( .A1(n11049), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11078) );
  INV_X1 U11997 ( .A(n11051), .ZN(n11049) );
  NAND2_X1 U11998 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n11025), .ZN(
        n11051) );
  INV_X1 U11999 ( .A(n11024), .ZN(n11025) );
  NOR2_X1 U12000 ( .A1(n10987), .A2(n15984), .ZN(n10988) );
  AND2_X1 U12001 ( .A1(n10965), .A2(n10964), .ZN(n14209) );
  NAND2_X1 U12002 ( .A1(n10244), .A2(n14146), .ZN(n10243) );
  INV_X1 U12003 ( .A(n10246), .ZN(n10244) );
  NOR2_X1 U12004 ( .A1(n10906), .A2(n15908), .ZN(n10907) );
  NAND2_X1 U12005 ( .A1(n10245), .A2(n10910), .ZN(n14228) );
  INV_X1 U12006 ( .A(n14225), .ZN(n10245) );
  NOR2_X2 U12007 ( .A1(n14249), .A2(n14238), .ZN(n14239) );
  NOR2_X1 U12008 ( .A1(n10870), .A2(n14478), .ZN(n10871) );
  NAND2_X1 U12009 ( .A1(n10871), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10906) );
  NAND2_X1 U12010 ( .A1(n10835), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10870) );
  NOR2_X1 U12011 ( .A1(n10819), .A2(n14164), .ZN(n10835) );
  NAND2_X1 U12012 ( .A1(n10812), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10819) );
  INV_X1 U12013 ( .A(n10811), .ZN(n10812) );
  AND2_X1 U12014 ( .A1(n10762), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10763) );
  NOR2_X1 U12015 ( .A1(n13944), .A2(n13856), .ZN(n10242) );
  NOR2_X1 U12016 ( .A1(n20883), .A2(n10698), .ZN(n10724) );
  NAND2_X1 U12017 ( .A1(n10688), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10698) );
  NOR2_X1 U12018 ( .A1(n13595), .A2(n13563), .ZN(n13712) );
  AND2_X1 U12019 ( .A1(n10668), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10688) );
  NOR2_X1 U12020 ( .A1(n10609), .A2(n10608), .ZN(n10641) );
  NAND2_X1 U12021 ( .A1(n13378), .A2(n10577), .ZN(n13482) );
  NAND2_X1 U12022 ( .A1(n10607), .A2(n10848), .ZN(n10617) );
  CLKBUF_X1 U12023 ( .A(n13480), .Z(n13596) );
  AND2_X1 U12024 ( .A1(n11376), .A2(n11375), .ZN(n14111) );
  NAND2_X1 U12025 ( .A1(n14125), .A2(n14111), .ZN(n14110) );
  AND2_X1 U12026 ( .A1(n14130), .A2(n14123), .ZN(n14125) );
  NAND2_X1 U12027 ( .A1(n10075), .A2(n10074), .ZN(n10073) );
  INV_X1 U12028 ( .A(n10076), .ZN(n10075) );
  NOR2_X1 U12029 ( .A1(n10078), .A2(n14221), .ZN(n10074) );
  NOR3_X1 U12030 ( .A1(n14247), .A2(n10078), .A3(n14242), .ZN(n14235) );
  NOR2_X1 U12031 ( .A1(n14247), .A2(n14242), .ZN(n14241) );
  OR2_X1 U12032 ( .A1(n16009), .A2(n11509), .ZN(n14472) );
  OR2_X1 U12033 ( .A1(n11423), .A2(n16079), .ZN(n14471) );
  NAND2_X1 U12034 ( .A1(n15995), .A2(n9756), .ZN(n14489) );
  AND2_X1 U12035 ( .A1(n13957), .A2(n9826), .ZN(n14256) );
  INV_X1 U12036 ( .A(n9844), .ZN(n10068) );
  AND2_X1 U12037 ( .A1(n11336), .A2(n11335), .ZN(n14266) );
  NAND2_X1 U12038 ( .A1(n13957), .A2(n10070), .ZN(n14274) );
  NAND2_X1 U12039 ( .A1(n13957), .A2(n13956), .ZN(n14272) );
  NAND2_X1 U12040 ( .A1(n14499), .A2(n11502), .ZN(n14496) );
  NAND2_X1 U12041 ( .A1(n10080), .A2(n10079), .ZN(n11500) );
  AND2_X1 U12042 ( .A1(n9796), .A2(n11495), .ZN(n10079) );
  AND2_X1 U12043 ( .A1(n11327), .A2(n11326), .ZN(n13945) );
  AND2_X1 U12044 ( .A1(n13946), .A2(n13945), .ZN(n13957) );
  OR2_X1 U12045 ( .A1(n13787), .A2(n11318), .ZN(n13858) );
  OR2_X1 U12046 ( .A1(n13577), .A2(n13565), .ZN(n13787) );
  NAND2_X1 U12047 ( .A1(n13579), .A2(n13578), .ZN(n13577) );
  OR2_X1 U12048 ( .A1(n13402), .A2(n13401), .ZN(n13504) );
  AND2_X1 U12049 ( .A1(n13416), .A2(n13341), .ZN(n14022) );
  XNOR2_X1 U12050 ( .A(n11432), .B(n11433), .ZN(n13317) );
  INV_X1 U12051 ( .A(n10466), .ZN(n9876) );
  INV_X1 U12052 ( .A(n13366), .ZN(n14656) );
  NAND2_X1 U12053 ( .A1(n10286), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13448) );
  NAND2_X1 U12054 ( .A1(n20158), .A2(n20157), .ZN(n20222) );
  NOR2_X1 U12055 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20682) );
  AND2_X1 U12056 ( .A1(n12242), .A2(n12241), .ZN(n16441) );
  AND2_X1 U12057 ( .A1(n10209), .A2(n10208), .ZN(n12152) );
  INV_X1 U12058 ( .A(n12189), .ZN(n10208) );
  NAND2_X1 U12059 ( .A1(n12216), .A2(n11774), .ZN(n10209) );
  NOR2_X1 U12060 ( .A1(n12140), .A2(n12139), .ZN(n12192) );
  NAND2_X1 U12061 ( .A1(n10218), .A2(n10217), .ZN(n14683) );
  INV_X1 U12062 ( .A(n12128), .ZN(n10217) );
  INV_X1 U12063 ( .A(n12132), .ZN(n16187) );
  INV_X1 U12064 ( .A(n16222), .ZN(n10114) );
  INV_X1 U12065 ( .A(n10111), .ZN(n10110) );
  OAI21_X1 U12066 ( .B1(n12939), .B2(n10112), .A(n12939), .ZN(n10111) );
  NOR3_X1 U12067 ( .A1(n12051), .A2(n10215), .A3(n12049), .ZN(n12063) );
  NAND2_X1 U12068 ( .A1(n12033), .A2(n9765), .ZN(n12058) );
  NAND2_X1 U12069 ( .A1(n12033), .A2(n10212), .ZN(n12060) );
  NAND2_X1 U12070 ( .A1(n12033), .A2(n12039), .ZN(n12044) );
  NAND2_X1 U12071 ( .A1(n12022), .A2(n12512), .ZN(n12025) );
  AND2_X1 U12072 ( .A1(n12015), .A2(n12013), .ZN(n12011) );
  NOR2_X1 U12073 ( .A1(n11964), .A2(n11966), .ZN(n11947) );
  NAND2_X1 U12074 ( .A1(n15182), .A2(n14843), .ZN(n14845) );
  NAND2_X1 U12075 ( .A1(n14876), .A2(n9763), .ZN(n14870) );
  NAND2_X1 U12076 ( .A1(n14876), .A2(n14877), .ZN(n14879) );
  NOR2_X1 U12077 ( .A1(n14796), .A2(n14797), .ZN(n14795) );
  NAND2_X1 U12078 ( .A1(n12637), .A2(n10173), .ZN(n10172) );
  INV_X1 U12079 ( .A(n10174), .ZN(n10173) );
  OR2_X1 U12080 ( .A1(n12647), .A2(n12646), .ZN(n13800) );
  OR2_X2 U12081 ( .A1(n13372), .A2(n10155), .ZN(n13570) );
  NAND2_X1 U12082 ( .A1(n10156), .A2(n13528), .ZN(n10155) );
  INV_X1 U12083 ( .A(n10158), .ZN(n10156) );
  AND2_X1 U12084 ( .A1(n14836), .A2(n12930), .ZN(n13126) );
  AND2_X1 U12085 ( .A1(n19186), .A2(n19850), .ZN(n19218) );
  INV_X1 U12086 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14902) );
  AND2_X1 U12087 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12934), .ZN(
        n12968) );
  AND2_X1 U12088 ( .A1(n12955), .A2(n9764), .ZN(n12963) );
  NAND2_X1 U12089 ( .A1(n12963), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12964) );
  NAND2_X1 U12090 ( .A1(n12955), .A2(n9762), .ZN(n12938) );
  AND2_X1 U12091 ( .A1(n12955), .A2(n9820), .ZN(n12960) );
  NAND2_X1 U12092 ( .A1(n10144), .A2(n10143), .ZN(n14794) );
  INV_X1 U12093 ( .A(n14791), .ZN(n10143) );
  AND2_X1 U12094 ( .A1(n12955), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12962) );
  INV_X1 U12095 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15006) );
  NOR2_X1 U12096 ( .A1(n12950), .A2(n10116), .ZN(n12954) );
  NAND2_X1 U12097 ( .A1(n12947), .A2(n9755), .ZN(n12948) );
  AND2_X1 U12098 ( .A1(n12947), .A2(n10122), .ZN(n12949) );
  NAND2_X1 U12099 ( .A1(n12947), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12946) );
  NAND2_X1 U12100 ( .A1(n13558), .A2(n13557), .ZN(n13560) );
  NAND2_X1 U12101 ( .A1(n10126), .A2(n9804), .ZN(n13391) );
  NOR2_X1 U12102 ( .A1(n13266), .A2(n10131), .ZN(n10130) );
  NOR2_X1 U12103 ( .A1(n16339), .A2(n10120), .ZN(n10119) );
  NOR2_X1 U12104 ( .A1(n12940), .A2(n13673), .ZN(n12942) );
  NOR2_X1 U12105 ( .A1(n13168), .A2(n13167), .ZN(n13211) );
  NOR2_X1 U12106 ( .A1(n15092), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10186) );
  NAND2_X1 U12107 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10185) );
  INV_X1 U12108 ( .A(n12109), .ZN(n12135) );
  NAND2_X1 U12109 ( .A1(n9860), .A2(n9856), .ZN(n9858) );
  AND2_X1 U12110 ( .A1(n9859), .A2(n14888), .ZN(n9856) );
  INV_X1 U12111 ( .A(n10136), .ZN(n10134) );
  NAND2_X1 U12112 ( .A1(n14733), .A2(n14726), .ZN(n14728) );
  OR2_X1 U12113 ( .A1(n16198), .A2(n10051), .ZN(n14911) );
  INV_X1 U12114 ( .A(n14909), .ZN(n10053) );
  OR2_X1 U12115 ( .A1(n12123), .A2(n15158), .ZN(n14938) );
  NAND2_X1 U12116 ( .A1(n10058), .A2(n10056), .ZN(n10228) );
  AND2_X1 U12117 ( .A1(n10227), .A2(n10057), .ZN(n10056) );
  NAND2_X1 U12118 ( .A1(n15059), .A2(n10059), .ZN(n10058) );
  NOR2_X1 U12119 ( .A1(n13974), .A2(n10232), .ZN(n10230) );
  NAND2_X1 U12120 ( .A1(n10202), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10201) );
  INV_X1 U12121 ( .A(n10203), .ZN(n10202) );
  OR2_X1 U12122 ( .A1(n15018), .A2(n10203), .ZN(n14984) );
  OR2_X1 U12123 ( .A1(n18978), .A2(n12088), .ZN(n14977) );
  NOR2_X1 U12124 ( .A1(n15018), .A2(n10205), .ZN(n14991) );
  AND2_X1 U12125 ( .A1(n10004), .A2(n14998), .ZN(n10002) );
  AND2_X1 U12126 ( .A1(n10003), .A2(n14972), .ZN(n10000) );
  OR2_X1 U12127 ( .A1(n15018), .A2(n15215), .ZN(n15002) );
  INV_X1 U12128 ( .A(n10144), .ZN(n14792) );
  NAND2_X1 U12129 ( .A1(n13558), .A2(n9794), .ZN(n13544) );
  NAND2_X1 U12130 ( .A1(n13558), .A2(n10141), .ZN(n13585) );
  AND2_X1 U12131 ( .A1(n13558), .A2(n10139), .ZN(n13587) );
  NOR2_X1 U12132 ( .A1(n12470), .A2(n16383), .ZN(n15295) );
  NAND2_X1 U12133 ( .A1(n15067), .A2(n15069), .ZN(n16299) );
  INV_X1 U12134 ( .A(n15295), .ZN(n16368) );
  OR2_X1 U12135 ( .A1(n15077), .A2(n15324), .ZN(n10238) );
  NAND2_X1 U12136 ( .A1(n13919), .A2(n12233), .ZN(n15329) );
  NAND2_X1 U12137 ( .A1(n13635), .A2(n12327), .ZN(n15343) );
  NOR2_X1 U12138 ( .A1(n10128), .A2(n13168), .ZN(n13311) );
  NAND2_X1 U12139 ( .A1(n10132), .A2(n10129), .ZN(n10128) );
  INV_X1 U12140 ( .A(n13266), .ZN(n10129) );
  OR2_X1 U12141 ( .A1(n13168), .A2(n10133), .ZN(n13265) );
  INV_X1 U12142 ( .A(n10132), .ZN(n10133) );
  AOI22_X1 U12143 ( .A1(n9818), .A2(n10048), .B1(n12131), .B2(n9759), .ZN(
        n10045) );
  INV_X1 U12144 ( .A(n10049), .ZN(n10048) );
  NAND2_X1 U12145 ( .A1(n12292), .A2(n12291), .ZN(n12295) );
  AND2_X1 U12146 ( .A1(n16451), .A2(n12463), .ZN(n16443) );
  AOI21_X1 U12147 ( .B1(n14005), .B2(n12619), .A(n12609), .ZN(n13075) );
  CLKBUF_X1 U12148 ( .A(n11542), .Z(n11543) );
  AND2_X1 U12149 ( .A1(n19565), .A2(n19534), .ZN(n19513) );
  INV_X1 U12150 ( .A(n19329), .ZN(n19566) );
  INV_X1 U12151 ( .A(n19697), .ZN(n19687) );
  INV_X1 U12152 ( .A(n19311), .ZN(n19313) );
  INV_X1 U12153 ( .A(n19312), .ZN(n19314) );
  NOR2_X2 U12154 ( .A1(n19270), .A2(n19269), .ZN(n19311) );
  NOR2_X2 U12155 ( .A1(n19268), .A2(n19269), .ZN(n19312) );
  OR2_X1 U12156 ( .A1(n19565), .A2(n19953), .ZN(n19688) );
  OR2_X1 U12157 ( .A1(n19565), .A2(n19534), .ZN(n19724) );
  NAND2_X1 U12158 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19731), .ZN(n19315) );
  NAND2_X1 U12159 ( .A1(n12144), .A2(n12143), .ZN(n16445) );
  OR2_X1 U12160 ( .A1(n15567), .A2(n17523), .ZN(n9956) );
  NOR3_X1 U12161 ( .A1(n17523), .A2(n16673), .A3(n18736), .ZN(n18754) );
  NOR2_X1 U12162 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16896), .ZN(n16889) );
  NOR2_X1 U12163 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16903), .ZN(n16902) );
  INV_X1 U12164 ( .A(n16942), .ZN(n17006) );
  NOR2_X1 U12165 ( .A1(n17450), .A2(n10034), .ZN(n10033) );
  INV_X1 U12166 ( .A(n10035), .ZN(n10034) );
  NOR2_X1 U12167 ( .A1(n20879), .A2(n10036), .ZN(n10035) );
  INV_X1 U12168 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10036) );
  NOR2_X1 U12169 ( .A1(n17311), .A2(n10028), .ZN(n10027) );
  INV_X1 U12170 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n10028) );
  NOR2_X1 U12171 ( .A1(n17543), .A2(n9999), .ZN(n9998) );
  AOI211_X1 U12172 ( .C1(n17298), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n15631), .B(n15630), .ZN(n15632) );
  NAND2_X1 U12173 ( .A1(n9789), .A2(n9951), .ZN(n9950) );
  NOR2_X1 U12174 ( .A1(n17484), .A2(n17483), .ZN(n17503) );
  NOR2_X1 U12175 ( .A1(n18925), .A2(n18749), .ZN(n17522) );
  NOR2_X1 U12176 ( .A1(n17633), .A2(n17634), .ZN(n16487) );
  NAND2_X1 U12177 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16487), .ZN(
        n17589) );
  NAND2_X1 U12178 ( .A1(n17658), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17633) );
  NAND2_X1 U12179 ( .A1(n17695), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17672) );
  NOR2_X1 U12180 ( .A1(n17711), .A2(n17713), .ZN(n17695) );
  NOR2_X1 U12181 ( .A1(n17744), .A2(n17748), .ZN(n17735) );
  INV_X1 U12182 ( .A(n17940), .ZN(n17889) );
  NAND2_X1 U12183 ( .A1(n9942), .A2(n9938), .ZN(n9937) );
  NOR2_X1 U12184 ( .A1(n16495), .A2(n9939), .ZN(n9938) );
  AND2_X1 U12185 ( .A1(n18890), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9939) );
  INV_X1 U12186 ( .A(n16539), .ZN(n9936) );
  NAND2_X1 U12187 ( .A1(n9933), .A2(n9942), .ZN(n9932) );
  OAI21_X1 U12188 ( .B1(n16495), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9933) );
  INV_X1 U12189 ( .A(n16496), .ZN(n9931) );
  NOR2_X1 U12190 ( .A1(n15833), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16494) );
  AND2_X1 U12191 ( .A1(n9941), .A2(n9940), .ZN(n16495) );
  NOR2_X1 U12192 ( .A1(n16548), .A2(n16531), .ZN(n9940) );
  INV_X1 U12193 ( .A(n16552), .ZN(n9941) );
  INV_X1 U12194 ( .A(n16513), .ZN(n17615) );
  AND2_X1 U12195 ( .A1(n15704), .A2(n15703), .ZN(n15705) );
  OR2_X1 U12196 ( .A1(n17742), .A2(n17959), .ZN(n15704) );
  NOR2_X1 U12197 ( .A1(n17722), .A2(n9845), .ZN(n17655) );
  NOR2_X1 U12198 ( .A1(n18098), .A2(n17773), .ZN(n17772) );
  NAND2_X1 U12199 ( .A1(n17831), .A2(n10099), .ZN(n17802) );
  NAND2_X1 U12200 ( .A1(n17831), .A2(n17841), .ZN(n17821) );
  NOR2_X1 U12201 ( .A1(n15767), .A2(n17854), .ZN(n18135) );
  INV_X1 U12202 ( .A(n9949), .ZN(n17831) );
  NAND2_X1 U12203 ( .A1(n17865), .A2(n15697), .ZN(n17846) );
  NAND2_X1 U12204 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17846), .ZN(
        n17845) );
  NOR2_X1 U12205 ( .A1(n17855), .A2(n18171), .ZN(n17854) );
  XNOR2_X1 U12206 ( .A(n15695), .B(n10098), .ZN(n17866) );
  INV_X1 U12207 ( .A(n15696), .ZN(n10098) );
  NOR2_X1 U12208 ( .A1(n17879), .A2(n18195), .ZN(n17878) );
  NAND2_X1 U12209 ( .A1(n17912), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17911) );
  NOR2_X1 U12210 ( .A1(n18942), .A2(n15727), .ZN(n18751) );
  NAND2_X1 U12211 ( .A1(n17333), .A2(n17336), .ZN(n15711) );
  OR2_X1 U12212 ( .A1(n9990), .A2(n15410), .ZN(n15712) );
  INV_X1 U12213 ( .A(n18750), .ZN(n18117) );
  INV_X1 U12214 ( .A(n18730), .ZN(n18733) );
  INV_X1 U12215 ( .A(n18751), .ZN(n18739) );
  AND2_X1 U12216 ( .A1(n9963), .A2(n9801), .ZN(n18277) );
  NOR2_X1 U12217 ( .A1(n15372), .A2(n9964), .ZN(n9963) );
  NOR2_X1 U12218 ( .A1(n15436), .A2(n15435), .ZN(n18287) );
  NOR2_X1 U12219 ( .A1(n15394), .A2(n15393), .ZN(n18294) );
  INV_X1 U12220 ( .A(n15712), .ZN(n18298) );
  NAND2_X1 U12221 ( .A1(n18933), .A2(n18275), .ZN(n18367) );
  NOR3_X1 U12222 ( .A1(n15580), .A2(n15719), .A3(n15579), .ZN(n18761) );
  INV_X1 U12223 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20883) );
  INV_X1 U12224 ( .A(n20059), .ZN(n20044) );
  AND2_X1 U12225 ( .A1(n14158), .A2(n13745), .ZN(n20040) );
  AND2_X1 U12226 ( .A1(n11412), .A2(n11411), .ZN(n20046) );
  AND2_X1 U12227 ( .A1(n14158), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20059) );
  NAND2_X1 U12228 ( .A1(n11412), .A2(n11410), .ZN(n20021) );
  AND2_X1 U12229 ( .A1(n11412), .A2(n11392), .ZN(n20027) );
  INV_X1 U12230 ( .A(n14280), .ZN(n14268) );
  INV_X1 U12231 ( .A(n14278), .ZN(n14267) );
  INV_X1 U12232 ( .A(n14270), .ZN(n13782) );
  NAND2_X2 U12233 ( .A1(n13302), .A2(n13301), .ZN(n14278) );
  OR2_X1 U12234 ( .A1(n13332), .A2(n19976), .ZN(n13302) );
  INV_X1 U12235 ( .A(n13782), .ZN(n14277) );
  INV_X1 U12236 ( .A(n14398), .ZN(n14303) );
  INV_X1 U12237 ( .A(n15972), .ZN(n14348) );
  NOR2_X1 U12238 ( .A1(n14348), .A2(n13289), .ZN(n15969) );
  INV_X1 U12239 ( .A(n15969), .ZN(n14353) );
  AND2_X1 U12241 ( .A1(n20851), .A2(n16173), .ZN(n13624) );
  INV_X1 U12242 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14450) );
  INV_X1 U12243 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14478) );
  NAND2_X1 U12244 ( .A1(n10080), .A2(n11495), .ZN(n13911) );
  OR2_X1 U12245 ( .A1(n20134), .A2(n11521), .ZN(n16037) );
  OR3_X1 U12246 ( .A1(n14549), .A2(n14521), .A3(n14540), .ZN(n14542) );
  INV_X1 U12247 ( .A(n9920), .ZN(n14373) );
  NAND2_X1 U12248 ( .A1(n14517), .A2(n14522), .ZN(n16054) );
  XNOR2_X1 U12249 ( .A(n9894), .B(n20932), .ZN(n15979) );
  OAI211_X1 U12250 ( .C1(n16113), .C2(n14601), .A(n14513), .B(n14512), .ZN(
        n15846) );
  NAND2_X1 U12251 ( .A1(n10022), .A2(n11512), .ZN(n14456) );
  NAND2_X1 U12252 ( .A1(n9926), .A2(n11476), .ZN(n16026) );
  NAND2_X1 U12253 ( .A1(n16031), .A2(n16030), .ZN(n9926) );
  OAI21_X1 U12254 ( .B1(n14509), .B2(n14642), .A(n16132), .ZN(n16156) );
  NAND2_X1 U12255 ( .A1(n13438), .A2(n14022), .ZN(n14642) );
  INV_X1 U12256 ( .A(n16089), .ZN(n20143) );
  INV_X1 U12257 ( .A(n9905), .ZN(n20142) );
  NAND2_X1 U12258 ( .A1(n9976), .A2(n10568), .ZN(n10567) );
  INV_X1 U12259 ( .A(n20682), .ZN(n20829) );
  INV_X1 U12260 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20825) );
  NAND2_X1 U12261 ( .A1(n14032), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14671) );
  INV_X1 U12262 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16169) );
  NOR2_X1 U12263 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n19975) );
  OAI21_X1 U12264 ( .B1(n20264), .B2(n20263), .A(n20262), .ZN(n20285) );
  INV_X1 U12265 ( .A(n20300), .ZN(n20317) );
  OAI21_X1 U12266 ( .B1(n20345), .B2(n20329), .A(n20651), .ZN(n20347) );
  INV_X1 U12267 ( .A(n20436), .ZN(n20457) );
  INV_X1 U12268 ( .A(n20496), .ZN(n20520) );
  INV_X1 U12269 ( .A(n20513), .ZN(n20518) );
  INV_X1 U12270 ( .A(n20641), .ZN(n20591) );
  AOI22_X1 U12271 ( .A1(n20566), .A2(n20563), .B1(n20561), .B2(n20560), .ZN(
        n20597) );
  OAI211_X1 U12272 ( .C1(n20670), .C2(n20652), .A(n20651), .B(n20650), .ZN(
        n20673) );
  NOR2_X1 U12273 ( .A1(n20260), .A2(n11284), .ZN(n16179) );
  NAND2_X1 U12274 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20848) );
  OAI21_X1 U12275 ( .B1(n16233), .B2(n10112), .A(n10110), .ZN(n16196) );
  NAND2_X1 U12276 ( .A1(n16221), .A2(n16222), .ZN(n16220) );
  NAND2_X1 U12277 ( .A1(n16233), .A2(n12939), .ZN(n16221) );
  AND2_X1 U12278 ( .A1(n12109), .A2(n12105), .ZN(n16217) );
  NAND2_X1 U12279 ( .A1(n16234), .A2(n16235), .ZN(n16233) );
  NAND2_X1 U12280 ( .A1(n16247), .A2(n12939), .ZN(n16234) );
  NAND2_X1 U12281 ( .A1(n16257), .A2(n12939), .ZN(n16248) );
  NAND2_X1 U12282 ( .A1(n16248), .A2(n16249), .ZN(n16247) );
  NAND2_X1 U12283 ( .A1(n12048), .A2(n10221), .ZN(n12098) );
  NAND2_X1 U12284 ( .A1(n14691), .A2(n12939), .ZN(n15783) );
  NAND2_X1 U12285 ( .A1(n18992), .A2(n12939), .ZN(n18981) );
  NAND2_X1 U12286 ( .A1(n18981), .A2(n18982), .ZN(n18980) );
  NAND2_X1 U12287 ( .A1(n14711), .A2(n12939), .ZN(n19004) );
  INV_X1 U12288 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14705) );
  OR2_X1 U12289 ( .A1(n12953), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10125) );
  OR2_X1 U12290 ( .A1(n12953), .A2(n12937), .ZN(n10124) );
  OR2_X1 U12291 ( .A1(n15028), .A2(n14702), .ZN(n14711) );
  NAND2_X1 U12292 ( .A1(n14685), .A2(n12987), .ZN(n19117) );
  OR2_X1 U12293 ( .A1(n18951), .A2(n12985), .ZN(n19059) );
  NAND2_X1 U12294 ( .A1(n19059), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19024) );
  OR3_X1 U12295 ( .A1(n12981), .A2(n12978), .A3(n12977), .ZN(n19090) );
  INV_X1 U12296 ( .A(n19024), .ZN(n19130) );
  INV_X1 U12297 ( .A(n14992), .ZN(n18976) );
  OR2_X1 U12298 ( .A1(n12280), .A2(n12279), .ZN(n13589) );
  OR2_X1 U12299 ( .A1(n13270), .A2(n10175), .ZN(n13310) );
  INV_X1 U12300 ( .A(n14785), .ZN(n14798) );
  OR2_X1 U12301 ( .A1(n14799), .A2(n19316), .ZN(n14785) );
  NOR2_X1 U12302 ( .A1(n9786), .A2(n12746), .ZN(n14756) );
  AND2_X1 U12303 ( .A1(n13126), .A2(n19268), .ZN(n19134) );
  AND2_X1 U12304 ( .A1(n14836), .A2(n11754), .ZN(n16265) );
  NOR2_X1 U12305 ( .A1(n19175), .A2(n19173), .ZN(n19138) );
  NAND2_X1 U12306 ( .A1(n10168), .A2(n12627), .ZN(n13165) );
  INV_X1 U12307 ( .A(n19953), .ZN(n19534) );
  INV_X1 U12308 ( .A(n16267), .ZN(n19173) );
  INV_X1 U12309 ( .A(n14836), .ZN(n19172) );
  NOR2_X1 U12310 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15857), .ZN(n19244) );
  CLKBUF_X1 U12311 ( .A(n13259), .Z(n13282) );
  INV_X1 U12312 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19025) );
  INV_X1 U12313 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16308) );
  INV_X1 U12314 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16315) );
  INV_X1 U12315 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16325) );
  INV_X1 U12316 ( .A(n16327), .ZN(n19267) );
  AND2_X1 U12317 ( .A1(n16338), .A2(n19942), .ZN(n19263) );
  INV_X1 U12318 ( .A(n19259), .ZN(n16335) );
  NAND2_X1 U12319 ( .A1(n13092), .A2(n13087), .ZN(n16338) );
  INV_X1 U12320 ( .A(n9733), .ZN(n19257) );
  AND2_X1 U12321 ( .A1(n16338), .A2(n13104), .ZN(n16327) );
  INV_X1 U12322 ( .A(n19263), .ZN(n16287) );
  NAND2_X1 U12323 ( .A1(n15090), .A2(n16417), .ZN(n15098) );
  INV_X1 U12324 ( .A(n15095), .ZN(n15096) );
  NAND2_X1 U12325 ( .A1(n10233), .A2(n10231), .ZN(n13975) );
  INV_X1 U12326 ( .A(n10232), .ZN(n10231) );
  AOI21_X1 U12327 ( .B1(n15027), .B2(n15025), .A(n15024), .ZN(n15015) );
  NAND2_X1 U12328 ( .A1(n10062), .A2(n15058), .ZN(n16284) );
  OR2_X1 U12329 ( .A1(n13372), .A2(n10157), .ZN(n13508) );
  INV_X1 U12330 ( .A(n10160), .ZN(n10157) );
  BUF_X1 U12331 ( .A(n19255), .Z(n19103) );
  INV_X1 U12332 ( .A(n16388), .ZN(n16417) );
  OAI21_X1 U12333 ( .B1(n13672), .B2(n12131), .A(n9759), .ZN(n13668) );
  NAND2_X1 U12334 ( .A1(n10046), .A2(n10049), .ZN(n13667) );
  AND2_X1 U12335 ( .A1(n13028), .A2(n13027), .ZN(n19165) );
  OR2_X1 U12336 ( .A1(n11823), .A2(n11822), .ZN(n11824) );
  INV_X1 U12337 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19958) );
  INV_X1 U12338 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19940) );
  INV_X1 U12339 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15858) );
  NAND2_X1 U12340 ( .A1(n13172), .A2(n13175), .ZN(n19936) );
  OAI21_X1 U12341 ( .B1(n19284), .B2(n19283), .A(n19282), .ZN(n19319) );
  OAI21_X1 U12342 ( .B1(n19284), .B2(n19279), .A(n19278), .ZN(n19320) );
  INV_X1 U12343 ( .A(n19470), .ZN(n19459) );
  AND2_X1 U12344 ( .A1(n19513), .A2(n19697), .ZN(n19497) );
  NOR2_X1 U12345 ( .A1(n19723), .A2(n19472), .ZN(n19522) );
  OAI21_X1 U12346 ( .B1(n19542), .B2(n19541), .A(n19540), .ZN(n19559) );
  OR2_X1 U12347 ( .A1(n19724), .A2(n19566), .ZN(n19596) );
  NOR2_X1 U12348 ( .A1(n19724), .A2(n19635), .ZN(n19654) );
  NOR2_X1 U12349 ( .A1(n19662), .A2(n19660), .ZN(n19682) );
  OAI22_X1 U12350 ( .A1(n20169), .A2(n19314), .B1(n19271), .B2(n19313), .ZN(
        n19725) );
  INV_X1 U12351 ( .A(n19805), .ZN(n19747) );
  OR2_X1 U12352 ( .A1(n19688), .A2(n19687), .ZN(n19760) );
  OAI22_X1 U12353 ( .A1(n21037), .A2(n19314), .B1(n19306), .B2(n19313), .ZN(
        n19757) );
  OAI21_X1 U12354 ( .B1(n19737), .B2(n19736), .A(n19735), .ZN(n19765) );
  INV_X1 U12355 ( .A(n19740), .ZN(n19784) );
  INV_X1 U12356 ( .A(n19704), .ZN(n19790) );
  INV_X1 U12357 ( .A(n19835), .ZN(n19821) );
  INV_X1 U12358 ( .A(n19757), .ZN(n19825) );
  OR2_X1 U12359 ( .A1(n19724), .A2(n19723), .ZN(n19835) );
  INV_X1 U12360 ( .A(n19824), .ZN(n19831) );
  INV_X1 U12361 ( .A(n19769), .ZN(n19830) );
  INV_X1 U12362 ( .A(n19764), .ZN(n19836) );
  OAI21_X1 U12363 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n21158), .ZN(n16473) );
  AND2_X1 U12364 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12206), .ZN(n19838) );
  INV_X1 U12365 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n21158) );
  NOR2_X1 U12366 ( .A1(n18754), .A2(n17484), .ZN(n18947) );
  NAND2_X1 U12367 ( .A1(n18947), .A2(n17485), .ZN(n18945) );
  INV_X1 U12368 ( .A(n18947), .ZN(n18943) );
  INV_X1 U12369 ( .A(n9956), .ZN(n16656) );
  NAND2_X1 U12370 ( .A1(n18759), .A2(n18771), .ZN(n16657) );
  NOR2_X1 U12371 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16872), .ZN(n16858) );
  INV_X1 U12372 ( .A(n17036), .ZN(n17026) );
  NOR2_X2 U12373 ( .A1(n18945), .A2(n18773), .ZN(n17018) );
  NOR2_X2 U12374 ( .A1(n18880), .A2(n16974), .ZN(n17021) );
  NOR2_X1 U12375 ( .A1(n17050), .A2(n17049), .ZN(n17077) );
  NAND2_X1 U12376 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17096), .ZN(n17087) );
  NOR2_X1 U12377 ( .A1(n21154), .A2(n17091), .ZN(n17096) );
  AND2_X1 U12378 ( .A1(n17156), .A2(n10030), .ZN(n17104) );
  NOR2_X1 U12379 ( .A1(n10032), .A2(n10031), .ZN(n10030) );
  NAND2_X1 U12380 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .ZN(n10031) );
  INV_X1 U12381 ( .A(n10033), .ZN(n10032) );
  NAND2_X1 U12382 ( .A1(n17156), .A2(n10033), .ZN(n17105) );
  NAND2_X1 U12383 ( .A1(n17156), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17142) );
  AND2_X1 U12384 ( .A1(n17251), .A2(n9753), .ZN(n17144) );
  NOR2_X1 U12385 ( .A1(n16812), .A2(n17157), .ZN(n17156) );
  NAND2_X1 U12386 ( .A1(n17251), .A2(n9752), .ZN(n17195) );
  AND2_X1 U12387 ( .A1(n17251), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n15537) );
  NOR2_X1 U12388 ( .A1(n17236), .A2(n17263), .ZN(n17251) );
  NAND2_X1 U12389 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17283), .ZN(n17263) );
  NOR2_X1 U12390 ( .A1(n17265), .A2(n17302), .ZN(n17283) );
  AND2_X1 U12391 ( .A1(n17320), .A2(n9843), .ZN(n17308) );
  NAND2_X1 U12392 ( .A1(n17320), .A2(n9770), .ZN(n17309) );
  NAND2_X1 U12393 ( .A1(n17320), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n17314) );
  NOR2_X1 U12394 ( .A1(n17316), .A2(n17321), .ZN(n17320) );
  NAND2_X1 U12395 ( .A1(n9821), .A2(P3_EBX_REG_2__SCAN_IN), .ZN(n17321) );
  NOR2_X1 U12396 ( .A1(n15860), .A2(n10037), .ZN(n17324) );
  NAND2_X1 U12397 ( .A1(n18929), .A2(n10038), .ZN(n10037) );
  NOR2_X1 U12398 ( .A1(n18277), .A2(n18925), .ZN(n10038) );
  NAND2_X1 U12399 ( .A1(n17324), .A2(P3_EBX_REG_0__SCAN_IN), .ZN(n17328) );
  INV_X1 U12400 ( .A(n17342), .ZN(n17338) );
  AND2_X1 U12401 ( .A1(n17363), .A2(n9772), .ZN(n17346) );
  NAND2_X1 U12402 ( .A1(n17363), .A2(n9771), .ZN(n17354) );
  INV_X1 U12403 ( .A(n17367), .ZN(n17363) );
  NAND2_X1 U12404 ( .A1(n17363), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17362) );
  NOR2_X1 U12405 ( .A1(n17372), .A2(n17450), .ZN(n17368) );
  NOR2_X1 U12406 ( .A1(n17408), .A2(n9986), .ZN(n17373) );
  NAND2_X1 U12407 ( .A1(n9847), .A2(n9987), .ZN(n9986) );
  INV_X1 U12408 ( .A(n17377), .ZN(n9987) );
  NAND2_X1 U12409 ( .A1(n17373), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17372) );
  NAND2_X1 U12410 ( .A1(n17412), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17408) );
  INV_X1 U12411 ( .A(n17378), .ZN(n17406) );
  NOR2_X2 U12412 ( .A1(n17336), .A2(n17465), .ZN(n17407) );
  NOR2_X1 U12413 ( .A1(n17587), .A2(n17418), .ZN(n17412) );
  NAND4_X1 U12414 ( .A1(n17417), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_9__SCAN_IN), .A4(n9754), .ZN(n17418) );
  NOR2_X1 U12415 ( .A1(n15863), .A2(n17479), .ZN(n17447) );
  INV_X1 U12416 ( .A(n9994), .ZN(n17445) );
  NOR2_X1 U12417 ( .A1(n15612), .A2(n15611), .ZN(n17458) );
  NOR2_X1 U12418 ( .A1(n15622), .A2(n15621), .ZN(n17466) );
  NAND2_X1 U12419 ( .A1(n17450), .A2(n17332), .ZN(n17465) );
  NOR2_X1 U12420 ( .A1(n17557), .A2(n17469), .ZN(n17475) );
  INV_X1 U12421 ( .A(n17478), .ZN(n17476) );
  NOR2_X1 U12422 ( .A1(n15679), .A2(n15678), .ZN(n17939) );
  OAI21_X1 U12423 ( .B1(n15862), .B2(n15861), .A(n18771), .ZN(n17479) );
  NOR3_X1 U12424 ( .A1(n15860), .A2(n17485), .A3(n18929), .ZN(n15861) );
  NOR3_X1 U12425 ( .A1(n18931), .A2(n15859), .A3(n18749), .ZN(n15862) );
  INV_X1 U12426 ( .A(n17479), .ZN(n17332) );
  NOR2_X1 U12427 ( .A1(n15864), .A2(n17479), .ZN(n17478) );
  NOR2_X1 U12428 ( .A1(n9961), .A2(n17583), .ZN(n17544) );
  OAI211_X1 U12429 ( .C1(n9961), .C2(n18796), .A(n17523), .B(n17522), .ZN(
        n17578) );
  BUF_X1 U12430 ( .A(n17578), .Z(n17583) );
  NOR2_X1 U12432 ( .A1(n16500), .A2(n16499), .ZN(n16501) );
  NOR2_X1 U12433 ( .A1(n17672), .A2(n17673), .ZN(n17658) );
  NOR2_X1 U12434 ( .A1(n18020), .A2(n17755), .ZN(n17719) );
  NAND2_X1 U12435 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17772), .ZN(
        n18079) );
  INV_X1 U12436 ( .A(n17777), .ZN(n16499) );
  NOR2_X2 U12437 ( .A1(n18620), .A2(n18367), .ZN(n18662) );
  INV_X1 U12438 ( .A(n18662), .ZN(n18365) );
  OAI21_X1 U12439 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18267), .A(n16657), 
        .ZN(n17940) );
  NOR2_X1 U12440 ( .A1(n9961), .A2(n18925), .ZN(n9957) );
  INV_X1 U12441 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18889) );
  INV_X1 U12442 ( .A(n16553), .ZN(n16549) );
  NAND2_X1 U12443 ( .A1(n16560), .A2(n16559), .ZN(n16561) );
  NAND2_X1 U12444 ( .A1(n10096), .A2(n9946), .ZN(n9945) );
  OR2_X1 U12445 ( .A1(n15708), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9947) );
  AND2_X1 U12446 ( .A1(n10095), .A2(n17953), .ZN(n9946) );
  AND2_X1 U12447 ( .A1(n17638), .A2(n9832), .ZN(n10097) );
  INV_X1 U12448 ( .A(n18226), .ZN(n18164) );
  INV_X1 U12449 ( .A(n18245), .ZN(n18189) );
  NAND2_X1 U12450 ( .A1(n18254), .A2(n16551), .ZN(n18162) );
  INV_X1 U12451 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18171) );
  OR2_X1 U12452 ( .A1(n18180), .A2(n18197), .ZN(n18196) );
  NAND2_X1 U12453 ( .A1(n18730), .A2(n15728), .ZN(n18716) );
  NOR2_X1 U12454 ( .A1(n18217), .A2(n18757), .ZN(n18260) );
  INV_X1 U12455 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18725) );
  INV_X1 U12456 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18746) );
  INV_X1 U12457 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21010) );
  AOI211_X1 U12458 ( .C1(n18771), .C2(n18744), .A(n18276), .B(n15581), .ZN(
        n18911) );
  INV_X1 U12459 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18282) );
  INV_X1 U12460 ( .A(n16929), .ZN(n18787) );
  NAND2_X1 U12461 ( .A1(n18889), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18783) );
  NAND2_X1 U12462 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18796) );
  NOR3_X1 U12463 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18812), .A3(n18793), 
        .ZN(n18928) );
  INV_X1 U12464 ( .A(n19268), .ZN(n19270) );
  NOR3_X1 U12465 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(n13024), .ZN(n16569) );
  INV_X1 U12466 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19913) );
  OAI21_X1 U12467 ( .B1(n14536), .B2(n19981), .A(n9985), .ZN(P1_U2968) );
  AOI21_X1 U12468 ( .B1(n13003), .B2(n20158), .A(n11524), .ZN(n9985) );
  INV_X1 U12469 ( .A(n9896), .ZN(n14536) );
  NAND2_X1 U12470 ( .A1(n9896), .A2(n20140), .ZN(n9895) );
  OAI21_X1 U12471 ( .B1(n14562), .B2(n16160), .A(n10081), .ZN(P1_U3003) );
  NOR2_X1 U12472 ( .A1(n14563), .A2(n10082), .ZN(n10081) );
  AND2_X1 U12473 ( .A1(n14571), .A2(n14564), .ZN(n10082) );
  OR2_X1 U12474 ( .A1(n12991), .A2(n9802), .ZN(P2_U2826) );
  AOI21_X1 U12475 ( .B1(n15109), .B2(n19121), .A(n10146), .ZN(n10145) );
  OAI21_X1 U12476 ( .B1(n13994), .B2(n16393), .A(n9911), .ZN(P2_U3015) );
  NAND2_X1 U12477 ( .A1(n10153), .A2(n9913), .ZN(n9912) );
  OAI21_X1 U12478 ( .B1(n16529), .B2(n17844), .A(n9795), .ZN(P3_U2801) );
  AND2_X1 U12479 ( .A1(n10103), .A2(n16528), .ZN(n10102) );
  OR2_X1 U12480 ( .A1(n16544), .A2(n18251), .ZN(n9944) );
  INV_X1 U12481 ( .A(n10475), .ZN(n11087) );
  XNOR2_X1 U12482 ( .A(n11816), .B(n11819), .ZN(n11845) );
  AND2_X2 U12483 ( .A1(n12710), .A2(n11541), .ZN(n11904) );
  INV_X2 U12484 ( .A(n9779), .ZN(n17290) );
  INV_X2 U12485 ( .A(n9779), .ZN(n15653) );
  NAND4_X2 U12486 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n12131) );
  INV_X1 U12487 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13673) );
  NAND2_X1 U12488 ( .A1(n10178), .A2(n10179), .ZN(n14769) );
  AND2_X1 U12489 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .ZN(n9752) );
  AND3_X1 U12490 ( .A1(n9850), .A2(n9752), .A3(P3_EBX_REG_18__SCAN_IN), .ZN(
        n9753) );
  AND2_X1 U12492 ( .A1(n12900), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11897) );
  CLKBUF_X3 U12493 ( .A(n11897), .Z(n12383) );
  INV_X2 U12494 ( .A(n14035), .ZN(n11383) );
  INV_X1 U12495 ( .A(n11423), .ZN(n14501) );
  INV_X2 U12496 ( .A(n14417), .ZN(n16009) );
  AND2_X1 U12497 ( .A1(n9994), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U12498 ( .A1(n14144), .A2(n14209), .ZN(n14201) );
  AND2_X1 U12499 ( .A1(n10122), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9755) );
  OR2_X1 U12500 ( .A1(n14417), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9756) );
  XNOR2_X1 U12501 ( .A(n12462), .B(n12461), .ZN(n19133) );
  INV_X1 U12502 ( .A(n19133), .ZN(n10154) );
  AND2_X1 U12503 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10284) );
  AND2_X1 U12504 ( .A1(n11512), .A2(n9849), .ZN(n9757) );
  AND2_X1 U12505 ( .A1(n9755), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9758) );
  AND2_X1 U12506 ( .A1(n13647), .A2(n12264), .ZN(n9759) );
  NOR2_X1 U12507 ( .A1(n14796), .A2(n9817), .ZN(n14779) );
  AND2_X1 U12508 ( .A1(n17156), .A2(n10035), .ZN(n9760) );
  INV_X1 U12509 ( .A(n12940), .ZN(n10121) );
  AND4_X1 U12510 ( .A1(n10121), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9761) );
  AND2_X1 U12511 ( .A1(n9820), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9762) );
  AND2_X1 U12512 ( .A1(n9837), .A2(n10152), .ZN(n13532) );
  AND2_X1 U12513 ( .A1(n12436), .A2(n14877), .ZN(n9763) );
  AND2_X1 U12514 ( .A1(n9762), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9764) );
  AND2_X1 U12515 ( .A1(n10210), .A2(n12056), .ZN(n9765) );
  NOR3_X1 U12516 ( .A1(n10215), .A2(n12049), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n9766) );
  AND2_X1 U12517 ( .A1(n17320), .A2(n10027), .ZN(n9767) );
  AND2_X1 U12518 ( .A1(n9830), .A2(n10066), .ZN(n9768) );
  AND2_X1 U12519 ( .A1(n10219), .A2(n12564), .ZN(n9769) );
  AND2_X1 U12520 ( .A1(n10027), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n9770) );
  AND2_X1 U12521 ( .A1(n9998), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9771) );
  AND2_X1 U12522 ( .A1(n9771), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9772) );
  OR3_X1 U12523 ( .A1(n12950), .A2(n10116), .A3(n10115), .ZN(n9773) );
  NOR2_X1 U12524 ( .A1(n15357), .A2(n15356), .ZN(n15419) );
  BUF_X1 U12525 ( .A(n15419), .Z(n15625) );
  AND4_X1 U12526 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n9776) );
  OR2_X1 U12527 ( .A1(n15354), .A2(n15356), .ZN(n9777) );
  INV_X2 U12528 ( .A(n15493), .ZN(n17060) );
  NAND2_X1 U12529 ( .A1(n15049), .A2(n12266), .ZN(n15018) );
  AND2_X1 U12530 ( .A1(n14144), .A2(n9979), .ZN(n14056) );
  INV_X1 U12531 ( .A(n9862), .ZN(n14928) );
  OR2_X1 U12532 ( .A1(n14752), .A2(n10135), .ZN(n9780) );
  NAND2_X1 U12533 ( .A1(n13953), .A2(n14153), .ZN(n14152) );
  OR2_X1 U12534 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n12104), .ZN(n9781) );
  AND2_X1 U12535 ( .A1(n14125), .A2(n9768), .ZN(n9782) );
  NOR2_X1 U12536 ( .A1(n14225), .A2(n10246), .ZN(n14143) );
  OR2_X1 U12537 ( .A1(n14794), .A2(n14786), .ZN(n9783) );
  AND2_X1 U12538 ( .A1(n17363), .A2(n9998), .ZN(n9784) );
  AND2_X1 U12539 ( .A1(n12048), .A2(n10219), .ZN(n9785) );
  AND2_X1 U12540 ( .A1(n13943), .A2(n13954), .ZN(n13953) );
  NAND2_X1 U12541 ( .A1(n12090), .A2(n10266), .ZN(n14958) );
  INV_X1 U12542 ( .A(n10218), .ZN(n12129) );
  NOR2_X1 U12543 ( .A1(n12119), .A2(n12118), .ZN(n10218) );
  AND2_X1 U12544 ( .A1(n14765), .A2(n14764), .ZN(n9786) );
  NAND4_X1 U12545 ( .A1(n10296), .A2(n10295), .A3(n10294), .A4(n10293), .ZN(
        n10426) );
  AND2_X1 U12546 ( .A1(n12297), .A2(n10149), .ZN(n9787) );
  NAND2_X1 U12547 ( .A1(n15082), .A2(n12237), .ZN(n15049) );
  AND4_X1 U12548 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n9788) );
  AND3_X1 U12549 ( .A1(n15637), .A2(n15642), .A3(n15636), .ZN(n9789) );
  AND2_X1 U12550 ( .A1(n11777), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n9790) );
  AND2_X1 U12551 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n9791) );
  AND2_X1 U12552 ( .A1(n11263), .A2(n11270), .ZN(n9792) );
  INV_X1 U12553 ( .A(n20199), .ZN(n13435) );
  AND2_X1 U12554 ( .A1(n9979), .A2(n14058), .ZN(n9793) );
  AND2_X1 U12555 ( .A1(n10139), .A2(n13525), .ZN(n9794) );
  AND3_X1 U12556 ( .A1(n16527), .A2(n10105), .A3(n10102), .ZN(n9795) );
  NAND2_X1 U12557 ( .A1(n13909), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9796) );
  AND2_X1 U12558 ( .A1(n11247), .A2(n13626), .ZN(n9797) );
  OR2_X1 U12559 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9798) );
  OR2_X1 U12560 ( .A1(n12130), .A2(n10206), .ZN(n9799) );
  AND2_X1 U12561 ( .A1(n15730), .A2(n15572), .ZN(n9800) );
  AND4_X1 U12562 ( .A1(n15371), .A2(n15370), .A3(n15369), .A4(n15368), .ZN(
        n9801) );
  NAND2_X1 U12563 ( .A1(n10148), .A2(n10145), .ZN(n9802) );
  NOR2_X1 U12564 ( .A1(n14756), .A2(n14755), .ZN(n9803) );
  AND2_X1 U12565 ( .A1(n10132), .A2(n10130), .ZN(n9804) );
  AND2_X1 U12566 ( .A1(n10225), .A2(n9863), .ZN(n9805) );
  NOR2_X1 U12567 ( .A1(n14809), .A2(n14811), .ZN(n12453) );
  INV_X1 U12568 ( .A(n11502), .ZN(n10092) );
  OR2_X1 U12569 ( .A1(n11162), .A2(n10251), .ZN(n9806) );
  AND2_X1 U12570 ( .A1(n12599), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9807) );
  NAND2_X1 U12571 ( .A1(n14144), .A2(n9981), .ZN(n14133) );
  INV_X1 U12572 ( .A(n10216), .ZN(n12069) );
  NOR2_X1 U12573 ( .A1(n12051), .A2(n12049), .ZN(n10216) );
  AND2_X1 U12574 ( .A1(n12095), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10237) );
  AND2_X1 U12575 ( .A1(n14595), .A2(n10063), .ZN(n9808) );
  INV_X1 U12576 ( .A(n10229), .ZN(n15176) );
  NAND2_X1 U12577 ( .A1(n10233), .A2(n10230), .ZN(n10229) );
  AND2_X1 U12578 ( .A1(n14389), .A2(n14557), .ZN(n9809) );
  OR2_X1 U12579 ( .A1(n12477), .A2(n10260), .ZN(n9810) );
  INV_X1 U12580 ( .A(n15568), .ZN(n16673) );
  NAND2_X1 U12581 ( .A1(n9956), .A2(n9955), .ZN(n15568) );
  AND2_X1 U12582 ( .A1(n14409), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14416) );
  AND2_X1 U12583 ( .A1(n12033), .A2(n10210), .ZN(n9811) );
  INV_X1 U12584 ( .A(n18310), .ZN(n17333) );
  NOR2_X1 U12585 ( .A1(n15404), .A2(n15403), .ZN(n18310) );
  AND2_X1 U12586 ( .A1(n9876), .A2(n10460), .ZN(n9812) );
  NOR2_X1 U12587 ( .A1(n14897), .A2(n14887), .ZN(n9813) );
  NAND2_X1 U12588 ( .A1(n14390), .A2(n14556), .ZN(n9814) );
  INV_X1 U12589 ( .A(n10416), .ZN(n10992) );
  INV_X1 U12590 ( .A(n10419), .ZN(n11193) );
  AND2_X1 U12592 ( .A1(n13438), .A2(n13425), .ZN(n20140) );
  NOR2_X1 U12593 ( .A1(n13270), .A2(n10174), .ZN(n13393) );
  INV_X1 U12595 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19949) );
  XOR2_X1 U12596 ( .A(n12136), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(
        n9815) );
  NOR2_X1 U12597 ( .A1(n13372), .A2(n13373), .ZN(n9816) );
  AND3_X1 U12598 ( .A1(n10703), .A2(n10704), .A3(n10242), .ZN(n13943) );
  NAND2_X1 U12599 ( .A1(n13943), .A2(n9983), .ZN(n14156) );
  OR2_X1 U12600 ( .A1(n14797), .A2(n10181), .ZN(n9817) );
  INV_X1 U12601 ( .A(n11469), .ZN(n9918) );
  AND2_X1 U12602 ( .A1(n13670), .A2(n10047), .ZN(n9818) );
  AND2_X1 U12603 ( .A1(n10070), .A2(n10069), .ZN(n9819) );
  AND2_X1 U12604 ( .A1(n13803), .A2(n13804), .ZN(n13802) );
  NAND2_X1 U12605 ( .A1(n10703), .A2(n10704), .ZN(n13769) );
  NOR2_X1 U12606 ( .A1(n13729), .A2(n13730), .ZN(n13123) );
  NOR2_X1 U12607 ( .A1(n13372), .A2(n10158), .ZN(n13507) );
  AND2_X1 U12608 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9820) );
  INV_X1 U12609 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U12610 ( .A1(n17328), .A2(n17325), .ZN(n9821) );
  OR3_X1 U12611 ( .A1(n14247), .A2(n10076), .A3(n10078), .ZN(n9822) );
  OR3_X1 U12612 ( .A1(n12950), .A2(n10118), .A3(n19025), .ZN(n9823) );
  NOR2_X1 U12613 ( .A1(n14370), .A2(n14540), .ZN(n9824) );
  AND2_X1 U12614 ( .A1(n11260), .A2(n11272), .ZN(n9825) );
  INV_X1 U12615 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13980) );
  INV_X1 U12616 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9880) );
  NAND3_X2 U12617 ( .A1(n15366), .A2(n15365), .A3(n15364), .ZN(n18929) );
  INV_X1 U12618 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10206) );
  AND2_X1 U12619 ( .A1(n12123), .A2(n15158), .ZN(n14937) );
  INV_X1 U12620 ( .A(n14937), .ZN(n10055) );
  AND2_X1 U12621 ( .A1(n9819), .A2(n10068), .ZN(n9826) );
  AND2_X1 U12622 ( .A1(n10634), .A2(n10664), .ZN(n9827) );
  AND2_X1 U12623 ( .A1(n9983), .A2(n10834), .ZN(n9828) );
  OR2_X1 U12624 ( .A1(n9818), .A2(n9759), .ZN(n9829) );
  INV_X1 U12625 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16339) );
  INV_X2 U12626 ( .A(n12897), .ZN(n11531) );
  AND2_X1 U12627 ( .A1(n10127), .A2(n13212), .ZN(n10132) );
  NAND2_X1 U12628 ( .A1(n12598), .A2(n12467), .ZN(n16413) );
  INV_X1 U12629 ( .A(n16413), .ZN(n16396) );
  INV_X1 U12630 ( .A(n15024), .ZN(n10007) );
  AND2_X1 U12631 ( .A1(n10067), .A2(n14111), .ZN(n9830) );
  INV_X1 U12632 ( .A(n14115), .ZN(n10253) );
  AND2_X1 U12633 ( .A1(n10164), .A2(n14843), .ZN(n9831) );
  OR2_X1 U12634 ( .A1(n17792), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9832) );
  NOR2_X1 U12635 ( .A1(n12967), .A2(n14902), .ZN(n12935) );
  NAND2_X1 U12636 ( .A1(n10636), .A2(n10606), .ZN(n20812) );
  NAND2_X1 U12637 ( .A1(n13957), .A2(n9819), .ZN(n10072) );
  AND2_X1 U12638 ( .A1(n13717), .A2(n12037), .ZN(n9833) );
  AND2_X1 U12639 ( .A1(n14726), .A2(n10138), .ZN(n9834) );
  NAND2_X1 U12640 ( .A1(n10099), .A2(n18095), .ZN(n9835) );
  INV_X1 U12641 ( .A(n10113), .ZN(n10112) );
  NOR2_X1 U12642 ( .A1(n16207), .A2(n10114), .ZN(n10113) );
  AND2_X1 U12643 ( .A1(n10171), .A2(n14764), .ZN(n9836) );
  AND2_X1 U12644 ( .A1(n12311), .A2(n13531), .ZN(n9837) );
  AND2_X1 U12645 ( .A1(n10152), .A2(n12311), .ZN(n9838) );
  AND2_X1 U12646 ( .A1(n10162), .A2(n14819), .ZN(n9839) );
  AND2_X1 U12647 ( .A1(n9763), .A2(n12439), .ZN(n9840) );
  AND2_X1 U12648 ( .A1(n12769), .A2(n12768), .ZN(n12770) );
  INV_X1 U12649 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n9916) );
  AND2_X1 U12650 ( .A1(n17324), .A2(n17450), .ZN(n17323) );
  INV_X1 U12651 ( .A(n17323), .ZN(n17318) );
  AND2_X1 U12652 ( .A1(n9742), .A2(n9904), .ZN(n9841) );
  INV_X1 U12653 ( .A(n18752), .ZN(n9960) );
  NOR2_X2 U12654 ( .A1(n15384), .A2(n15383), .ZN(n18316) );
  INV_X1 U12655 ( .A(n10834), .ZN(n9984) );
  NAND2_X2 U12656 ( .A1(n16545), .A2(n16549), .ZN(n17792) );
  OR2_X1 U12657 ( .A1(n12130), .A2(n12585), .ZN(n9842) );
  NOR2_X1 U12658 ( .A1(n18930), .A2(n18783), .ZN(n18771) );
  INV_X1 U12659 ( .A(n18771), .ZN(n18925) );
  INV_X1 U12660 ( .A(n11551), .ZN(n12819) );
  AND2_X1 U12661 ( .A1(n9770), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U12662 ( .A1(n11338), .A2(n11337), .ZN(n9844) );
  OR2_X1 U12663 ( .A1(n17594), .A2(n21129), .ZN(n9845) );
  AND4_X1 U12664 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n9846) );
  INV_X1 U12665 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10581) );
  INV_X2 U12666 ( .A(n10254), .ZN(n17298) );
  AND4_X1 U12667 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_22__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n9847)
         );
  AND2_X1 U12668 ( .A1(n10198), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9848) );
  NOR2_X1 U12669 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n9849) );
  INV_X1 U12670 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n9999) );
  AND4_X1 U12671 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(P3_EBX_REG_15__SCAN_IN), .A4(P3_EBX_REG_14__SCAN_IN), .ZN(n9850)
         );
  INV_X1 U12672 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10115) );
  INV_X1 U12673 ( .A(n15140), .ZN(n10199) );
  AND2_X1 U12674 ( .A1(n10186), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9851) );
  INV_X1 U12675 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10123) );
  INV_X1 U12676 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n10029) );
  NOR3_X2 U12677 ( .A1(n18781), .A2(n18725), .A3(n18409), .ZN(n18383) );
  NOR3_X2 U12678 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18781), .A3(
        n18503), .ZN(n18472) );
  NOR3_X2 U12679 ( .A1(n18781), .A2(n18574), .A3(n18550), .ZN(n18543) );
  AOI221_X2 U12680 ( .B1(n18621), .B2(n18622), .C1(n18620), .C2(n18622), .A(
        n18619), .ZN(n18656) );
  CLKBUF_X1 U12681 ( .A(n19794), .Z(n9852) );
  NOR2_X2 U12682 ( .A1(n20225), .A2(n9873), .ZN(n20702) );
  NAND2_X1 U12683 ( .A1(n12497), .A2(n9853), .ZN(n12502) );
  XNOR2_X2 U12684 ( .A(n12498), .B(n9854), .ZN(n10165) );
  NAND2_X1 U12685 ( .A1(n10239), .A2(n9855), .ZN(n19733) );
  INV_X1 U12686 ( .A(n9860), .ZN(n14898) );
  INV_X1 U12687 ( .A(n14896), .ZN(n9859) );
  AND2_X4 U12688 ( .A1(n12162), .A2(n11777), .ZN(n12574) );
  NAND2_X1 U12689 ( .A1(n12162), .A2(n9790), .ZN(n11805) );
  NAND2_X1 U12690 ( .A1(n12162), .A2(n9861), .ZN(n11781) );
  INV_X1 U12691 ( .A(n12122), .ZN(n9865) );
  NOR2_X2 U12692 ( .A1(n15313), .A2(n15310), .ZN(n15067) );
  NAND3_X2 U12693 ( .A1(n10189), .A2(n10188), .A3(n11912), .ZN(n12001) );
  NAND4_X1 U12694 ( .A1(n11868), .A2(n11866), .A3(n11865), .A4(n11867), .ZN(
        n9869) );
  AND2_X2 U12695 ( .A1(n9870), .A2(n11911), .ZN(n10189) );
  NAND4_X1 U12696 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11895), .ZN(
        n9870) );
  NAND2_X1 U12697 ( .A1(n9873), .A2(n14281), .ZN(n11429) );
  NAND2_X1 U12698 ( .A1(n10393), .A2(n9873), .ZN(n10394) );
  NAND2_X1 U12699 ( .A1(n9872), .A2(n9871), .ZN(n13419) );
  NAND2_X1 U12700 ( .A1(n13414), .A2(n13338), .ZN(n9871) );
  NAND2_X1 U12701 ( .A1(n13413), .A2(n9873), .ZN(n9872) );
  NAND2_X1 U12702 ( .A1(n13485), .A2(n9874), .ZN(n11448) );
  XNOR2_X1 U12703 ( .A(n13485), .B(n9874), .ZN(n13500) );
  NAND2_X1 U12704 ( .A1(n11445), .A2(n11444), .ZN(n9874) );
  NAND2_X1 U12705 ( .A1(n10548), .A2(n10460), .ZN(n9875) );
  NAND2_X2 U12706 ( .A1(n9875), .A2(n10466), .ZN(n13462) );
  NAND2_X1 U12707 ( .A1(n9812), .A2(n10548), .ZN(n10467) );
  NAND3_X1 U12708 ( .A1(n9878), .A2(n10444), .A3(n9877), .ZN(n10488) );
  NAND3_X1 U12709 ( .A1(n9882), .A2(n10442), .A3(n9881), .ZN(n10443) );
  OR2_X1 U12710 ( .A1(n9884), .A2(n9966), .ZN(n10465) );
  OR2_X1 U12711 ( .A1(n9884), .A2(n10581), .ZN(n10585) );
  NAND2_X1 U12712 ( .A1(n10337), .A2(n10336), .ZN(n9892) );
  NAND4_X4 U12713 ( .A1(n10318), .A2(n10319), .A3(n10316), .A4(n10317), .ZN(
        n14281) );
  INV_X2 U12715 ( .A(n10435), .ZN(n13136) );
  OAI22_X1 U12716 ( .A1(n15979), .A2(n19981), .B1(n20137), .B2(n15978), .ZN(
        n15980) );
  AOI22_X1 U12717 ( .A1(n15827), .A2(n14501), .B1(n15826), .B2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9894) );
  OR2_X2 U12718 ( .A1(n11513), .A2(n10092), .ZN(n10083) );
  AOI21_X2 U12719 ( .B1(n14473), .B2(n14463), .A(n11507), .ZN(n14461) );
  AND2_X4 U12720 ( .A1(n10287), .A2(n10286), .ZN(n10896) );
  NAND2_X1 U12721 ( .A1(n14535), .A2(n9895), .ZN(P1_U3000) );
  NAND2_X1 U12722 ( .A1(n13448), .A2(n10581), .ZN(n9904) );
  AOI211_X2 U12723 ( .C1(n13992), .C2(n16400), .A(n9810), .B(n9912), .ZN(n9911) );
  AOI21_X1 U12724 ( .B1(n10154), .B2(n16396), .A(n9807), .ZN(n9913) );
  OAI21_X2 U12725 ( .B1(n13672), .B2(n13671), .A(n12220), .ZN(n13834) );
  NAND2_X2 U12726 ( .A1(n11951), .A2(n12210), .ZN(n13672) );
  NOR2_X2 U12727 ( .A1(n14921), .A2(n15117), .ZN(n9914) );
  OR2_X2 U12728 ( .A1(n15018), .A2(n10201), .ZN(n14963) );
  NAND2_X1 U12729 ( .A1(n9917), .A2(n9915), .ZN(n11432) );
  NAND2_X1 U12730 ( .A1(n13317), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11435) );
  NAND3_X1 U12731 ( .A1(n9814), .A2(n9921), .A3(n11518), .ZN(n9919) );
  NAND2_X1 U12732 ( .A1(n10084), .A2(n10089), .ZN(n9928) );
  NAND2_X1 U12733 ( .A1(n13963), .A2(n9927), .ZN(n10089) );
  NAND2_X1 U12734 ( .A1(n17874), .A2(n17875), .ZN(n17873) );
  INV_X2 U12735 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18910) );
  NAND3_X1 U12736 ( .A1(n16542), .A2(n16543), .A3(n9944), .ZN(P3_U2831) );
  NOR2_X2 U12737 ( .A1(n9949), .A2(n9835), .ZN(n17775) );
  NAND3_X1 U12738 ( .A1(n15639), .A2(n15641), .A3(n9953), .ZN(n9952) );
  NOR2_X2 U12739 ( .A1(n17732), .A2(n17856), .ZN(n17691) );
  AOI21_X2 U12740 ( .B1(n18730), .B2(n15730), .A(n15729), .ZN(n18732) );
  AOI21_X2 U12741 ( .B1(n18731), .B2(n18303), .A(n16673), .ZN(n18730) );
  NOR2_X2 U12742 ( .A1(n15729), .A2(n9800), .ZN(n18731) );
  AND2_X2 U12743 ( .A1(n9962), .A2(n9961), .ZN(n18750) );
  NAND3_X1 U12744 ( .A1(n15374), .A2(n15373), .A3(n9965), .ZN(n9964) );
  AND2_X4 U12745 ( .A1(n13359), .A2(n14661), .ZN(n10412) );
  INV_X1 U12746 ( .A(n9967), .ZN(n9969) );
  INV_X1 U12747 ( .A(n10418), .ZN(n9971) );
  NAND2_X4 U12748 ( .A1(n9968), .A2(n9776), .ZN(n13626) );
  INV_X1 U12749 ( .A(n13595), .ZN(n9975) );
  NAND2_X1 U12750 ( .A1(n9975), .A2(n9973), .ZN(n13710) );
  OAI21_X1 U12751 ( .B1(n10570), .B2(n10518), .A(n9977), .ZN(n10526) );
  NAND2_X1 U12752 ( .A1(n10570), .A2(n9880), .ZN(n9976) );
  NAND2_X1 U12753 ( .A1(n13943), .A2(n9828), .ZN(n14248) );
  NAND3_X1 U12754 ( .A1(n9993), .A2(n9991), .A3(n15412), .ZN(n9990) );
  NAND3_X1 U12755 ( .A1(n9996), .A2(n9846), .A3(P3_EAX_REG_0__SCAN_IN), .ZN(
        n9995) );
  AND2_X1 U12756 ( .A1(n15037), .A2(n14972), .ZN(n15027) );
  NAND2_X1 U12757 ( .A1(n15067), .A2(n10011), .ZN(n10008) );
  NAND2_X1 U12758 ( .A1(n10440), .A2(n10445), .ZN(n10020) );
  NAND2_X1 U12759 ( .A1(n10430), .A2(n13424), .ZN(n10019) );
  INV_X2 U12760 ( .A(n14417), .ZN(n14465) );
  NAND2_X1 U12761 ( .A1(n10021), .A2(n9827), .ZN(n10694) );
  NAND2_X1 U12762 ( .A1(n10022), .A2(n9757), .ZN(n14439) );
  INV_X1 U12763 ( .A(n16050), .ZN(n16047) );
  XNOR2_X1 U12764 ( .A(n10023), .B(n16053), .ZN(n16050) );
  NOR2_X1 U12765 ( .A1(n14501), .A2(n14530), .ZN(n10025) );
  NAND2_X1 U12766 ( .A1(n14429), .A2(n14530), .ZN(n10026) );
  NAND2_X1 U12767 ( .A1(n14408), .A2(n14501), .ZN(n14424) );
  INV_X1 U12768 ( .A(n15537), .ZN(n17234) );
  INV_X2 U12769 ( .A(n11743), .ZN(n11765) );
  NAND2_X2 U12770 ( .A1(n10040), .A2(n10039), .ZN(n11743) );
  NAND2_X1 U12771 ( .A1(n10042), .A2(n11537), .ZN(n10039) );
  NAND2_X1 U12772 ( .A1(n10041), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10040) );
  NAND4_X1 U12773 ( .A1(n11575), .A2(n11574), .A3(n11572), .A4(n11573), .ZN(
        n10041) );
  NAND4_X1 U12774 ( .A1(n11577), .A2(n11579), .A3(n11578), .A4(n11576), .ZN(
        n10042) );
  NAND3_X1 U12775 ( .A1(n12162), .A2(n11777), .A3(P2_REIP_REG_1__SCAN_IN), 
        .ZN(n10043) );
  NAND2_X1 U12776 ( .A1(n13672), .A2(n9829), .ZN(n10044) );
  NAND2_X1 U12777 ( .A1(n10044), .A2(n10045), .ZN(n13844) );
  INV_X1 U12778 ( .A(n13647), .ZN(n10050) );
  NAND3_X1 U12779 ( .A1(n14928), .A2(n14929), .A3(n10055), .ZN(n10054) );
  NAND2_X2 U12780 ( .A1(n11477), .A2(n11422), .ZN(n11423) );
  OR2_X2 U12781 ( .A1(n10694), .A2(n10695), .ZN(n11477) );
  NAND2_X1 U12782 ( .A1(n14595), .A2(n11517), .ZN(n14425) );
  INV_X1 U12783 ( .A(n10072), .ZN(n14265) );
  NAND3_X1 U12784 ( .A1(n10089), .A2(n14455), .A3(n10088), .ZN(n14454) );
  NAND2_X1 U12785 ( .A1(n17921), .A2(n17922), .ZN(n17920) );
  AND2_X1 U12786 ( .A1(n17619), .A2(n15708), .ZN(n15709) );
  NAND2_X1 U12787 ( .A1(n10096), .A2(n10097), .ZN(n17621) );
  INV_X1 U12788 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10101) );
  OAI21_X1 U12789 ( .B1(n16233), .B2(n10109), .A(n10107), .ZN(n16205) );
  NOR2_X1 U12790 ( .A1(n12950), .A2(n19025), .ZN(n12952) );
  INV_X1 U12791 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U12792 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10120) );
  NAND3_X1 U12793 ( .A1(n10121), .A2(n10119), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12943) );
  NAND3_X1 U12794 ( .A1(n10121), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12941) );
  OAI21_X1 U12795 ( .B1(n13989), .B2(n10125), .A(n10124), .ZN(n14702) );
  AND2_X2 U12796 ( .A1(n12929), .A2(n11765), .ZN(n11754) );
  INV_X1 U12797 ( .A(n13168), .ZN(n10126) );
  NOR2_X2 U12798 ( .A1(n14693), .A2(n9783), .ZN(n14773) );
  NAND3_X1 U12799 ( .A1(n11754), .A2(n12330), .A3(P2_REIP_REG_1__SCAN_IN), 
        .ZN(n10149) );
  AND2_X2 U12800 ( .A1(n14876), .A2(n9840), .ZN(n14853) );
  NAND2_X1 U12801 ( .A1(n13052), .A2(n10150), .ZN(n13536) );
  CLKBUF_X1 U12802 ( .A(n13052), .Z(n10152) );
  OR2_X1 U12803 ( .A1(n14714), .A2(n16388), .ZN(n10153) );
  NAND2_X1 U12805 ( .A1(n15182), .A2(n9839), .ZN(n14809) );
  NAND2_X1 U12806 ( .A1(n11854), .A2(n13120), .ZN(n11858) );
  OR2_X1 U12807 ( .A1(n11826), .A2(n19118), .ZN(n11847) );
  NAND2_X1 U12808 ( .A1(n13120), .A2(n11855), .ZN(n11859) );
  INV_X2 U12809 ( .A(n11826), .ZN(n13120) );
  NAND2_X1 U12810 ( .A1(n11845), .A2(n11826), .ZN(n11836) );
  XNOR2_X2 U12811 ( .A(n12497), .B(n10165), .ZN(n11826) );
  AND2_X2 U12812 ( .A1(n12626), .A2(n13162), .ZN(n13119) );
  NAND2_X1 U12813 ( .A1(n14765), .A2(n9836), .ZN(n10169) );
  AOI21_X1 U12814 ( .B1(n12746), .B2(n10171), .A(n12770), .ZN(n10170) );
  AND2_X2 U12815 ( .A1(n10169), .A2(n10170), .ZN(n12794) );
  NOR2_X2 U12816 ( .A1(n13270), .A2(n10172), .ZN(n13801) );
  INV_X1 U12817 ( .A(n10257), .ZN(n10175) );
  INV_X1 U12818 ( .A(n14796), .ZN(n10178) );
  INV_X1 U12819 ( .A(n12208), .ZN(n12209) );
  NAND2_X1 U12820 ( .A1(n12208), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16329) );
  NOR2_X1 U12821 ( .A1(n14916), .A2(n14901), .ZN(n14900) );
  NAND2_X1 U12822 ( .A1(n13992), .A2(n9733), .ZN(n10184) );
  NOR2_X1 U12823 ( .A1(n13991), .A2(n13990), .ZN(n10187) );
  OAI21_X1 U12824 ( .B1(n15329), .B2(n10194), .A(n10190), .ZN(n15082) );
  NAND2_X1 U12825 ( .A1(n11947), .A2(n11946), .ZN(n12004) );
  NAND2_X1 U12826 ( .A1(n12048), .A2(n9769), .ZN(n12104) );
  NAND2_X1 U12827 ( .A1(n12048), .A2(n11665), .ZN(n12097) );
  NAND2_X1 U12828 ( .A1(n12022), .A2(n10223), .ZN(n11661) );
  INV_X1 U12829 ( .A(n11661), .ZN(n12038) );
  NAND2_X1 U12830 ( .A1(n12002), .A2(n12234), .ZN(n12225) );
  NAND2_X1 U12831 ( .A1(n10226), .A2(n12000), .ZN(n12234) );
  INV_X1 U12832 ( .A(n12001), .ZN(n10226) );
  OAI21_X2 U12833 ( .B1(n10230), .B2(n10237), .A(n10228), .ZN(n14952) );
  OAI21_X2 U12834 ( .B1(n15076), .B2(n10238), .A(n12020), .ZN(n15313) );
  NAND2_X2 U12835 ( .A1(n10241), .A2(n10240), .ZN(n13344) );
  NAND3_X1 U12836 ( .A1(n10241), .A2(n10240), .A3(n10410), .ZN(n11276) );
  NAND3_X1 U12837 ( .A1(n10703), .A2(n10704), .A3(n10723), .ZN(n13854) );
  OR2_X2 U12838 ( .A1(n14133), .A2(n10251), .ZN(n14104) );
  XNOR2_X2 U12839 ( .A(n10443), .B(n10457), .ZN(n20289) );
  OR2_X2 U12840 ( .A1(n17024), .A2(n15355), .ZN(n10262) );
  XNOR2_X1 U12841 ( .A(n15692), .B(n15691), .ZN(n17885) );
  AOI21_X2 U12842 ( .B1(n14070), .B2(n14080), .A(n14056), .ZN(n14387) );
  NAND2_X1 U12843 ( .A1(n14761), .A2(n14760), .ZN(n14759) );
  CLKBUF_X1 U12844 ( .A(n11544), .Z(n14000) );
  INV_X1 U12845 ( .A(n11719), .ZN(n13185) );
  NAND2_X1 U12846 ( .A1(n11677), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11678) );
  OR2_X2 U12847 ( .A1(n11858), .A2(n13176), .ZN(n11921) );
  NOR2_X1 U12848 ( .A1(n13176), .A2(n14005), .ZN(n11846) );
  NAND2_X1 U12849 ( .A1(n12230), .A2(n10256), .ZN(n12228) );
  XNOR2_X1 U12850 ( .A(n13119), .B(n13118), .ZN(n19565) );
  INV_X1 U12851 ( .A(n12745), .ZN(n14770) );
  CLKBUF_X1 U12852 ( .A(n13799), .Z(n13830) );
  NOR2_X1 U12853 ( .A1(n19290), .A2(n19315), .ZN(n19794) );
  XNOR2_X1 U12854 ( .A(n11764), .B(n11743), .ZN(n12166) );
  AND2_X1 U12855 ( .A1(n11743), .A2(n12929), .ZN(n11703) );
  XNOR2_X1 U12856 ( .A(n10580), .B(n10578), .ZN(n11436) );
  NAND2_X1 U12857 ( .A1(n10647), .A2(n10646), .ZN(n13595) );
  INV_X1 U12858 ( .A(n13597), .ZN(n10646) );
  INV_X1 U12859 ( .A(n13480), .ZN(n10647) );
  CLKBUF_X1 U12860 ( .A(n14248), .Z(n14252) );
  INV_X1 U12861 ( .A(n13799), .ZN(n12659) );
  AOI21_X1 U12862 ( .B1(n12122), .B2(n12121), .A(n14911), .ZN(n12127) );
  NAND2_X1 U12863 ( .A1(n11740), .A2(n11750), .ZN(n11741) );
  NOR2_X2 U12864 ( .A1(n14741), .A2(n14740), .ZN(n14739) );
  INV_X1 U12865 ( .A(n10437), .ZN(n13326) );
  NAND2_X1 U12866 ( .A1(n10437), .A2(n14281), .ZN(n10393) );
  AND2_X1 U12867 ( .A1(n10488), .A2(n10486), .ZN(n10545) );
  NOR2_X1 U12868 ( .A1(n13344), .A2(n13137), .ZN(n15789) );
  NOR2_X1 U12869 ( .A1(n13344), .A2(n12995), .ZN(n13464) );
  OR2_X1 U12870 ( .A1(n20606), .A2(n20830), .ZN(n20609) );
  OR2_X1 U12871 ( .A1(n20606), .A2(n20151), .ZN(n20555) );
  AOI21_X1 U12872 ( .B1(n10673), .B2(n10848), .A(n10672), .ZN(n13563) );
  INV_X1 U12874 ( .A(n14354), .ZN(n15970) );
  NAND2_X2 U12875 ( .A1(n15972), .A2(n13289), .ZN(n14354) );
  NAND2_X1 U12876 ( .A1(n14278), .A2(n20224), .ZN(n14280) );
  INV_X1 U12877 ( .A(n20134), .ZN(n19981) );
  INV_X2 U12878 ( .A(n13681), .ZN(n20118) );
  AND3_X1 U12879 ( .A1(n18098), .A2(n18132), .A3(n15698), .ZN(n10255) );
  INV_X1 U12880 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15589) );
  INV_X1 U12881 ( .A(n10816), .ZN(n10848) );
  INV_X2 U12882 ( .A(n18940), .ZN(n18872) );
  AND2_X1 U12883 ( .A1(n16329), .A2(n12231), .ZN(n10256) );
  AND2_X1 U12884 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10257) );
  AND3_X1 U12885 ( .A1(n11686), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11685), .ZN(n10258) );
  AND2_X1 U12886 ( .A1(n11688), .A2(n11687), .ZN(n10259) );
  INV_X1 U12887 ( .A(n13377), .ZN(n10576) );
  INV_X1 U12888 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15698) );
  INV_X1 U12889 ( .A(n14679), .ZN(n11790) );
  INV_X1 U12890 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12512) );
  AND4_X1 U12891 ( .A1(n15105), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n12476), .ZN(n10260) );
  CLKBUF_X1 U12892 ( .A(n16648), .Z(n16649) );
  OR2_X1 U12893 ( .A1(n13501), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10261) );
  NOR2_X1 U12894 ( .A1(n15355), .A2(n15356), .ZN(n15624) );
  CLKBUF_X3 U12895 ( .A(n15624), .Z(n17284) );
  NOR2_X1 U12896 ( .A1(n20487), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10263) );
  INV_X1 U12897 ( .A(n19841), .ZN(n19080) );
  AND2_X1 U12898 ( .A1(n13080), .A2(n19838), .ZN(n14790) );
  INV_X2 U12899 ( .A(n14790), .ZN(n14799) );
  INV_X1 U12900 ( .A(n11068), .ZN(n11172) );
  INV_X2 U12901 ( .A(n17447), .ZN(n17473) );
  AND2_X1 U12902 ( .A1(n12814), .A2(n12838), .ZN(n10264) );
  AND3_X1 U12903 ( .A1(n12089), .A2(n15013), .A3(n14977), .ZN(n10266) );
  AND2_X1 U12904 ( .A1(n14938), .A2(n12124), .ZN(n10267) );
  INV_X1 U12905 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16467) );
  NAND2_X1 U12906 ( .A1(n11877), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11878) );
  AND3_X1 U12907 ( .A1(n10455), .A2(n13298), .A3(n10439), .ZN(n10440) );
  OR2_X1 U12908 ( .A1(n10661), .A2(n10660), .ZN(n11479) );
  AND2_X1 U12909 ( .A1(n12167), .A2(n12929), .ZN(n11745) );
  INV_X1 U12910 ( .A(n11242), .ZN(n11238) );
  INV_X1 U12911 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10305) );
  OR2_X1 U12912 ( .A1(n10551), .A2(n10550), .ZN(n10552) );
  INV_X1 U12913 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11532) );
  INV_X1 U12914 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11530) );
  AND2_X1 U12915 ( .A1(n11236), .A2(n11237), .ZN(n11234) );
  OR2_X1 U12916 ( .A1(n10687), .A2(n10686), .ZN(n11488) );
  NOR2_X1 U12917 ( .A1(n11013), .A2(n10348), .ZN(n10349) );
  INV_X1 U12918 ( .A(n12892), .ZN(n12871) );
  AND2_X1 U12919 ( .A1(n12817), .A2(n10264), .ZN(n12818) );
  AND2_X1 U12920 ( .A1(n14976), .A2(n14974), .ZN(n12073) );
  OR2_X1 U12921 ( .A1(n12236), .A2(n20961), .ZN(n12237) );
  AOI21_X1 U12922 ( .B1(n20825), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11234), .ZN(n11233) );
  AND2_X1 U12923 ( .A1(n11358), .A2(n11357), .ZN(n14211) );
  AND4_X1 U12924 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10317) );
  AND2_X1 U12925 ( .A1(n12998), .A2(n14027), .ZN(n13337) );
  OR2_X1 U12926 ( .A1(n11159), .A2(n14396), .ZN(n11139) );
  INV_X1 U12927 ( .A(n11078), .ZN(n11077) );
  INV_X1 U12928 ( .A(n13856), .ZN(n10723) );
  INV_X1 U12929 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10608) );
  AND3_X1 U12930 ( .A1(n11421), .A2(n9918), .A3(n11490), .ZN(n11422) );
  OR2_X1 U12931 ( .A1(n10631), .A2(n10630), .ZN(n11461) );
  AND2_X1 U12932 ( .A1(n13298), .A2(n13297), .ZN(n13341) );
  AND4_X1 U12933 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10294) );
  AND3_X1 U12934 ( .A1(n15589), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n12138), .ZN(n12140) );
  AND2_X1 U12935 ( .A1(n12728), .A2(n12727), .ZN(n12763) );
  INV_X1 U12936 ( .A(n12894), .ZN(n12887) );
  AOI21_X1 U12937 ( .B1(n14909), .B2(n15134), .A(n14937), .ZN(n12116) );
  AND3_X1 U12938 ( .A1(n11651), .A2(n11650), .A3(n11649), .ZN(n11658) );
  INV_X1 U12939 ( .A(n12282), .ZN(n12296) );
  NOR2_X1 U12940 ( .A1(n17455), .A2(n15756), .ZN(n15760) );
  OR2_X1 U12941 ( .A1(n15740), .A2(n17466), .ZN(n15749) );
  INV_X1 U12942 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20977) );
  NOR2_X1 U12943 ( .A1(n11260), .A2(n11469), .ZN(n11262) );
  INV_X1 U12944 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n11284) );
  INV_X1 U12945 ( .A(n20846), .ZN(n13742) );
  INV_X1 U12946 ( .A(n13501), .ZN(n11374) );
  INV_X1 U12947 ( .A(n10671), .ZN(n10672) );
  AND2_X1 U12948 ( .A1(n13337), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10615) );
  NOR2_X1 U12949 ( .A1(n11282), .A2(n14045), .ZN(n11283) );
  OR2_X1 U12950 ( .A1(n14082), .A2(n14092), .ZN(n14069) );
  NAND2_X1 U12951 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11157) );
  INV_X1 U12952 ( .A(n14226), .ZN(n10910) );
  AND2_X1 U12953 ( .A1(n20260), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11225) );
  AND2_X1 U12954 ( .A1(n13324), .A2(n13136), .ZN(n13422) );
  OR2_X1 U12955 ( .A1(n14465), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14371) );
  NAND2_X1 U12956 ( .A1(n14281), .A2(n13626), .ZN(n11469) );
  NOR2_X1 U12957 ( .A1(n16113), .A2(n13492), .ZN(n14643) );
  INV_X1 U12958 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20490) );
  OR2_X1 U12959 ( .A1(n19961), .A2(n16469), .ZN(n12157) );
  AND2_X1 U12960 ( .A1(n12788), .A2(n12787), .ZN(n12791) );
  AND2_X1 U12961 ( .A1(n12839), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12625) );
  OR2_X1 U12962 ( .A1(n12813), .A2(n12815), .ZN(n12838) );
  INV_X1 U12963 ( .A(n12812), .ZN(n12839) );
  INV_X1 U12964 ( .A(n13831), .ZN(n12658) );
  AND2_X1 U12965 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n12474), .ZN(
        n15153) );
  NOR2_X1 U12966 ( .A1(n16368), .A2(n12471), .ZN(n15286) );
  INV_X1 U12967 ( .A(n15265), .ZN(n15330) );
  AND3_X1 U12968 ( .A1(n12259), .A2(n12258), .A3(n12257), .ZN(n13606) );
  OR2_X1 U12969 ( .A1(n13174), .A2(n13173), .ZN(n13175) );
  NOR2_X1 U12970 ( .A1(n18791), .A2(n17889), .ZN(n16488) );
  NAND2_X1 U12971 ( .A1(n16556), .A2(n16555), .ZN(n16557) );
  NOR2_X1 U12972 ( .A1(n17846), .A2(n17856), .ZN(n15735) );
  AOI211_X1 U12973 ( .C1(n15711), .C2(n15564), .A(n15563), .B(n15562), .ZN(
        n15571) );
  OR2_X1 U12974 ( .A1(n18904), .A2(n18788), .ZN(n18275) );
  NAND2_X1 U12975 ( .A1(n12992), .A2(n13428), .ZN(n14029) );
  AND2_X1 U12976 ( .A1(n14023), .A2(n11277), .ZN(n14030) );
  OR3_X1 U12977 ( .A1(n14096), .A2(n21109), .A3(n16045), .ZN(n14074) );
  OR3_X1 U12978 ( .A1(n20021), .A2(n11405), .A3(n11404), .ZN(n14138) );
  NAND2_X1 U12979 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n10907), .ZN(
        n10943) );
  INV_X1 U12980 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14164) );
  INV_X1 U12981 ( .A(n20046), .ZN(n20060) );
  OR3_X1 U12982 ( .A1(n20846), .A2(n20135), .A3(n11281), .ZN(n14158) );
  INV_X1 U12983 ( .A(n11302), .ZN(n13303) );
  OR2_X1 U12984 ( .A1(n11161), .A2(n11160), .ZN(n14092) );
  INV_X1 U12985 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15908) );
  NOR2_X1 U12986 ( .A1(n10741), .A2(n20001), .ZN(n10762) );
  INV_X1 U12987 ( .A(n19976), .ZN(n13420) );
  INV_X1 U12988 ( .A(n16133), .ZN(n16064) );
  INV_X1 U12989 ( .A(n20145), .ZN(n16135) );
  OAI21_X1 U12990 ( .B1(n20852), .B2(n16179), .A(n14671), .ZN(n20161) );
  AND3_X1 U12991 ( .A1(n13335), .A2(n13334), .A3(n13333), .ZN(n15792) );
  INV_X1 U12992 ( .A(n20431), .ZN(n20815) );
  OR2_X1 U12993 ( .A1(n20534), .A2(n20609), .ZN(n20513) );
  INV_X1 U12994 ( .A(n20829), .ZN(n20813) );
  AND2_X1 U12995 ( .A1(n20524), .A2(n10463), .ZN(n20164) );
  NAND3_X1 U12996 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n9880), .A3(n20161), 
        .ZN(n20225) );
  INV_X1 U12997 ( .A(n19117), .ZN(n19101) );
  XNOR2_X1 U12998 ( .A(n12817), .B(n10264), .ZN(n14741) );
  AND2_X1 U12999 ( .A1(n12636), .A2(n13547), .ZN(n12637) );
  NAND2_X1 U13000 ( .A1(n14836), .A2(n19316), .ZN(n16267) );
  INV_X1 U13001 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16227) );
  OR2_X1 U13002 ( .A1(n15018), .A2(n15291), .ZN(n15042) );
  OR2_X1 U13003 ( .A1(n15091), .A2(n15092), .ZN(n15097) );
  OR2_X1 U13004 ( .A1(n15331), .A2(n16403), .ZN(n16383) );
  INV_X1 U13005 ( .A(n11912), .ZN(n12318) );
  AND3_X1 U13006 ( .A1(n13207), .A2(n13206), .A3(n13205), .ZN(n16458) );
  INV_X1 U13007 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19951) );
  INV_X1 U13008 ( .A(n19923), .ZN(n19635) );
  INV_X1 U13009 ( .A(n19943), .ZN(n19925) );
  INV_X1 U13010 ( .A(n12253), .ZN(n16469) );
  INV_X1 U13011 ( .A(n18791), .ZN(n17709) );
  OR2_X1 U13012 ( .A1(n16711), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n16701) );
  OR3_X1 U13013 ( .A1(n17029), .A2(n16759), .A3(n18853), .ZN(n16749) );
  INV_X1 U13014 ( .A(n17035), .ZN(n17028) );
  AND4_X1 U13015 ( .A1(n18316), .A2(n18298), .A3(n15552), .A4(n15730), .ZN(
        n15449) );
  NOR2_X1 U13016 ( .A1(n16720), .A2(n16525), .ZN(n16524) );
  NOR2_X1 U13017 ( .A1(n17615), .A2(n18079), .ZN(n17945) );
  INV_X1 U13018 ( .A(n18005), .ZN(n18010) );
  INV_X1 U13019 ( .A(n18090), .ZN(n18001) );
  INV_X1 U13020 ( .A(n16859), .ZN(n17780) );
  NOR2_X1 U13021 ( .A1(n15735), .A2(n18171), .ZN(n17809) );
  INV_X1 U13022 ( .A(n16488), .ZN(n17694) );
  NAND2_X1 U13023 ( .A1(n17651), .A2(n17986), .ZN(n17650) );
  NOR2_X1 U13024 ( .A1(n17742), .A2(n18054), .ZN(n17680) );
  INV_X1 U13025 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18098) );
  INV_X1 U13026 ( .A(n15690), .ZN(n15691) );
  INV_X1 U13027 ( .A(n15684), .ZN(n15685) );
  NAND2_X1 U13028 ( .A1(n15819), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19976) );
  AND2_X1 U13029 ( .A1(n14158), .A2(n11285), .ZN(n20031) );
  INV_X1 U13030 ( .A(n20021), .ZN(n20019) );
  INV_X1 U13031 ( .A(n14027), .ZN(n20224) );
  INV_X1 U13032 ( .A(n14306), .ZN(n14340) );
  NAND2_X1 U13033 ( .A1(n13322), .A2(n13420), .ZN(n13001) );
  NOR2_X2 U13034 ( .A1(n20118), .A2(n20177), .ZN(n20110) );
  AND2_X1 U13035 ( .A1(n11282), .A2(n11164), .ZN(n14369) );
  NAND2_X1 U13036 ( .A1(n10988), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11024) );
  NAND2_X1 U13037 ( .A1(n10763), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10811) );
  INV_X1 U13038 ( .A(n16037), .ZN(n20132) );
  AND2_X1 U13039 ( .A1(n15805), .A2(n13420), .ZN(n20134) );
  OAI21_X1 U13040 ( .B1(n16094), .B2(n14613), .A(n14576), .ZN(n16082) );
  OR2_X1 U13041 ( .A1(n20139), .A2(n20143), .ZN(n16133) );
  OAI22_X1 U13042 ( .A1(n20167), .A2(n20166), .B1(n20435), .B2(n20324), .ZN(
        n20228) );
  INV_X1 U13043 ( .A(n20232), .ZN(n20253) );
  INV_X1 U13044 ( .A(n20279), .ZN(n20284) );
  OAI211_X1 U13045 ( .C1(n20396), .C2(n20568), .A(n20651), .B(n20381), .ZN(
        n20398) );
  NOR2_X2 U13046 ( .A1(n20819), .A2(n20609), .ZN(n20397) );
  NAND2_X1 U13047 ( .A1(n20431), .A2(n20321), .ZN(n20819) );
  INV_X1 U13048 ( .A(n20534), .ZN(n20528) );
  INV_X1 U13049 ( .A(n20554), .ZN(n20519) );
  OR2_X1 U13050 ( .A1(n20812), .A2(n20431), .ZN(n20534) );
  INV_X1 U13051 ( .A(n20556), .ZN(n20592) );
  OAI21_X1 U13052 ( .B1(n20608), .B2(n20607), .A(n20689), .ZN(n20638) );
  INV_X1 U13053 ( .A(n20645), .ZN(n20672) );
  INV_X1 U13054 ( .A(n20731), .ZN(n20738) );
  INV_X1 U13055 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19972) );
  OR2_X1 U13056 ( .A1(n16451), .A2(n16479), .ZN(n19181) );
  NAND2_X1 U13057 ( .A1(n14692), .A2(n14983), .ZN(n14691) );
  NAND2_X1 U13058 ( .A1(n19004), .A2(n19005), .ZN(n19003) );
  AND2_X1 U13059 ( .A1(n13258), .A2(n12976), .ZN(n19121) );
  INV_X1 U13060 ( .A(n19059), .ZN(n19122) );
  INV_X1 U13061 ( .A(n19105), .ZN(n19119) );
  OR2_X1 U13062 ( .A1(n12393), .A2(n12392), .ZN(n13524) );
  OR2_X1 U13063 ( .A1(n12341), .A2(n12340), .ZN(n13394) );
  INV_X1 U13064 ( .A(n13612), .ZN(n13084) );
  AND2_X1 U13065 ( .A1(n13126), .A2(n19270), .ZN(n19135) );
  AND2_X1 U13066 ( .A1(n12429), .A2(n12428), .ZN(n13571) );
  INV_X1 U13067 ( .A(n19168), .ZN(n19175) );
  INV_X1 U13068 ( .A(n12196), .ZN(n19187) );
  OAI21_X1 U13069 ( .B1(n11776), .B2(n15853), .A(n13180), .ZN(n13259) );
  AND2_X1 U13070 ( .A1(n14752), .A2(n14751), .ZN(n16232) );
  INV_X1 U13071 ( .A(n16338), .ZN(n19256) );
  AND2_X1 U13072 ( .A1(n12124), .A2(n12108), .ZN(n14929) );
  AND2_X1 U13073 ( .A1(n11790), .A2(n19928), .ZN(n19255) );
  AND2_X1 U13074 ( .A1(n12207), .A2(n19838), .ZN(n12598) );
  NOR2_X2 U13075 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19928) );
  INV_X1 U13076 ( .A(n19778), .ZN(n19731) );
  AND2_X1 U13077 ( .A1(n16449), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16474) );
  AND2_X1 U13078 ( .A1(n19936), .A2(n19943), .ZN(n19329) );
  INV_X1 U13079 ( .A(n19354), .ZN(n19376) );
  INV_X1 U13080 ( .A(n19441), .ZN(n19431) );
  OAI21_X1 U13081 ( .B1(n19420), .B2(n19419), .A(n19418), .ZN(n19437) );
  NOR2_X1 U13082 ( .A1(n19936), .A2(n19925), .ZN(n19697) );
  INV_X1 U13083 ( .A(n19563), .ZN(n19555) );
  INV_X1 U13084 ( .A(n19596), .ZN(n19588) );
  INV_X1 U13085 ( .A(n19591), .ZN(n19622) );
  OAI21_X1 U13086 ( .B1(n19666), .B2(n19665), .A(n19664), .ZN(n19683) );
  INV_X1 U13087 ( .A(n19799), .ZN(n19743) );
  INV_X1 U13088 ( .A(n19760), .ZN(n19763) );
  OAI22_X1 U13089 ( .A1(n20221), .A2(n19314), .B1(n20992), .B2(n19313), .ZN(
        n19764) );
  NAND2_X1 U13090 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n15857) );
  INV_X1 U13091 ( .A(n15853), .ZN(n19857) );
  INV_X1 U13092 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19866) );
  INV_X1 U13093 ( .A(n17522), .ZN(n17484) );
  NOR3_X1 U13094 ( .A1(n18857), .A2(n18855), .A3(n16749), .ZN(n16733) );
  NOR2_X1 U13095 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16831), .ZN(n16815) );
  NOR2_X1 U13096 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16854), .ZN(n16836) );
  INV_X1 U13097 ( .A(n17018), .ZN(n17029) );
  INV_X1 U13098 ( .A(n17039), .ZN(n16974) );
  NOR2_X1 U13099 ( .A1(n18255), .A2(n16929), .ZN(n16967) );
  INV_X1 U13100 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20879) );
  INV_X1 U13101 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17265) );
  NOR2_X1 U13102 ( .A1(n15580), .A2(n15449), .ZN(n15860) );
  NOR3_X1 U13103 ( .A1(n17450), .A2(n17408), .A3(n17377), .ZN(n17396) );
  INV_X1 U13104 ( .A(n15732), .ZN(n18048) );
  INV_X1 U13105 ( .A(n17786), .ZN(n17801) );
  NAND2_X1 U13106 ( .A1(n17808), .A2(n18048), .ZN(n18090) );
  INV_X1 U13107 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18095) );
  INV_X1 U13108 ( .A(n18162), .ZN(n18175) );
  INV_X1 U13109 ( .A(n18254), .ZN(n18217) );
  XNOR2_X1 U13110 ( .A(n15682), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17922) );
  INV_X1 U13111 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18930) );
  NOR2_X1 U13112 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18880), .ZN(
        n18904) );
  NOR2_X1 U13113 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18906) );
  INV_X1 U13114 ( .A(n18713), .ZN(n18360) );
  CLKBUF_X1 U13115 ( .A(n18356), .Z(n18384) );
  INV_X1 U13116 ( .A(n18364), .ZN(n18426) );
  INV_X1 U13117 ( .A(n18480), .ZN(n18520) );
  INV_X1 U13118 ( .A(n18547), .ZN(n18614) );
  AND2_X1 U13119 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18662), .ZN(n18681) );
  INV_X1 U13120 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18933) );
  INV_X1 U13121 ( .A(n18796), .ZN(n18931) );
  AND2_X1 U13122 ( .A1(n18872), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18812) );
  NAND2_X1 U13123 ( .A1(n14032), .A2(n11269), .ZN(n13625) );
  INV_X1 U13124 ( .A(n11417), .ZN(n11418) );
  INV_X1 U13125 ( .A(n20027), .ZN(n20062) );
  INV_X1 U13126 ( .A(n20067), .ZN(n14190) );
  NAND2_X1 U13127 ( .A1(n14278), .A2(n14027), .ZN(n14270) );
  NOR2_X1 U13128 ( .A1(n13018), .A2(n13017), .ZN(n13019) );
  AND2_X1 U13129 ( .A1(n13690), .A2(n13689), .ZN(n20227) );
  NAND2_X1 U13130 ( .A1(n13001), .A2(n13000), .ZN(n15972) );
  INV_X1 U13131 ( .A(n20072), .ZN(n20095) );
  NOR2_X1 U13132 ( .A1(n13625), .A2(n13624), .ZN(n13681) );
  OR2_X1 U13133 ( .A1(n20118), .A2(n13626), .ZN(n13680) );
  INV_X1 U13134 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15984) );
  INV_X1 U13135 ( .A(n16033), .ZN(n16029) );
  INV_X1 U13136 ( .A(n20140), .ZN(n16160) );
  INV_X1 U13137 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20562) );
  AOI21_X1 U13138 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n9880), .A(n16166), 
        .ZN(n16165) );
  OR2_X1 U13139 ( .A1(n20294), .A2(n20555), .ZN(n20232) );
  OR2_X1 U13140 ( .A1(n20294), .A2(n20609), .ZN(n20279) );
  AOI22_X1 U13141 ( .A1(n20259), .A2(n20263), .B1(n10263), .B2(n20489), .ZN(
        n20288) );
  INV_X1 U13142 ( .A(n20293), .ZN(n20320) );
  OR2_X1 U13143 ( .A1(n20819), .A2(n20555), .ZN(n20373) );
  AOI22_X1 U13144 ( .A1(n20380), .A2(n20377), .B1(n20561), .B2(n10263), .ZN(
        n20401) );
  OR2_X1 U13145 ( .A1(n20819), .A2(n20533), .ZN(n20436) );
  NAND2_X1 U13146 ( .A1(n20528), .A2(n20432), .ZN(n20485) );
  AOI22_X1 U13147 ( .A1(n20495), .A2(n20491), .B1(n20489), .B2(n20488), .ZN(
        n20523) );
  OR2_X1 U13148 ( .A1(n20534), .A2(n20642), .ZN(n20554) );
  INV_X1 U13149 ( .A(n20685), .ZN(n20571) );
  INV_X1 U13150 ( .A(n20719), .ZN(n20586) );
  OR2_X1 U13151 ( .A1(n20688), .A2(n20555), .ZN(n20641) );
  INV_X1 U13152 ( .A(n20737), .ZN(n20676) );
  OR2_X1 U13153 ( .A1(n20688), .A2(n20533), .ZN(n20731) );
  OR2_X1 U13154 ( .A1(n20688), .A2(n20642), .ZN(n20742) );
  INV_X1 U13155 ( .A(n20811), .ZN(n20747) );
  OR2_X1 U13156 ( .A1(n16445), .A2(n12975), .ZN(n13179) );
  INV_X1 U13157 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19661) );
  OR3_X1 U13158 ( .A1(n12981), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19857), 
        .ZN(n19105) );
  INV_X1 U13159 ( .A(n19121), .ZN(n19100) );
  AND2_X1 U13160 ( .A1(n13078), .A2(n13077), .ZN(n19943) );
  NAND2_X1 U13161 ( .A1(n12915), .A2(n12914), .ZN(n14836) );
  NAND2_X1 U13162 ( .A1(n14836), .A2(n12916), .ZN(n19168) );
  NOR2_X2 U13163 ( .A1(n16265), .A2(n13126), .ZN(n19180) );
  NAND2_X1 U13164 ( .A1(n19218), .A2(n19187), .ZN(n19216) );
  INV_X1 U13165 ( .A(n19218), .ZN(n19253) );
  OR2_X1 U13166 ( .A1(n13179), .A2(n15585), .ZN(n19185) );
  INV_X1 U13167 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16291) );
  INV_X1 U13168 ( .A(n16423), .ZN(n16393) );
  INV_X1 U13169 ( .A(n16400), .ZN(n16420) );
  AND2_X1 U13170 ( .A1(n15259), .A2(n15264), .ZN(n15265) );
  INV_X1 U13171 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14010) );
  NAND2_X1 U13172 ( .A1(n19329), .A2(n19471), .ZN(n19349) );
  NAND2_X1 U13173 ( .A1(n19471), .A2(n19923), .ZN(n19409) );
  NAND2_X1 U13174 ( .A1(n19513), .A2(n19923), .ZN(n19441) );
  NAND2_X1 U13175 ( .A1(n19471), .A2(n19697), .ZN(n19470) );
  INV_X1 U13176 ( .A(n19522), .ZN(n19533) );
  NAND2_X1 U13177 ( .A1(n19513), .A2(n19782), .ZN(n19563) );
  OR2_X1 U13178 ( .A1(n19688), .A2(n19566), .ZN(n19591) );
  INV_X1 U13179 ( .A(n19654), .ZN(n19626) );
  NAND2_X1 U13180 ( .A1(n19627), .A2(n19923), .ZN(n19686) );
  INV_X1 U13181 ( .A(n19725), .ZN(n19787) );
  OR2_X1 U13182 ( .A1(n19688), .A2(n19723), .ZN(n19824) );
  AOI211_X1 U13183 ( .C1(n16472), .C2(n16471), .A(n11790), .B(n16470), .ZN(
        n19843) );
  INV_X1 U13184 ( .A(n19922), .ZN(n19844) );
  NAND2_X1 U13185 ( .A1(n19845), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19970) );
  INV_X1 U13186 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16675) );
  NAND2_X1 U13187 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18805), .ZN(n18940) );
  INV_X1 U13188 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16720) );
  INV_X1 U13189 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17236) );
  INV_X1 U13190 ( .A(n17021), .ZN(n17014) );
  OAI211_X1 U13191 ( .C1(n18783), .C2(n18777), .A(n18943), .B(n16967), .ZN(
        n17039) );
  AND3_X1 U13192 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17209), .ZN(n17208) );
  INV_X1 U13193 ( .A(n17323), .ZN(n17331) );
  OR3_X1 U13194 ( .A1(n17535), .A2(n17533), .A3(n17392), .ZN(n17383) );
  INV_X1 U13195 ( .A(n17465), .ZN(n17470) );
  NOR2_X1 U13196 ( .A1(n17561), .A2(n17461), .ZN(n17464) );
  INV_X1 U13197 ( .A(n17503), .ZN(n17521) );
  INV_X1 U13198 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17553) );
  AOI21_X1 U13199 ( .B1(n16541), .B2(n17857), .A(n16501), .ZN(n16502) );
  INV_X1 U13200 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17986) );
  INV_X1 U13201 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17819) );
  INV_X1 U13202 ( .A(n17857), .ZN(n17844) );
  INV_X1 U13203 ( .A(n17934), .ZN(n17919) );
  NAND2_X1 U13204 ( .A1(n16561), .A2(n18148), .ZN(n16565) );
  INV_X1 U13205 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17998) );
  NAND2_X1 U13206 ( .A1(n18148), .A2(n18217), .ZN(n18245) );
  INV_X1 U13207 ( .A(n18260), .ZN(n18247) );
  INV_X1 U13208 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18273) );
  INV_X1 U13209 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18285) );
  INV_X1 U13210 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18313) );
  INV_X1 U13211 ( .A(n18449), .ZN(n18432) );
  INV_X1 U13212 ( .A(n18471), .ZN(n18431) );
  INV_X1 U13213 ( .A(n18542), .ZN(n18476) );
  INV_X1 U13214 ( .A(n18566), .ZN(n18500) );
  INV_X1 U13215 ( .A(n18623), .ZN(n18666) );
  INV_X1 U13216 ( .A(n18626), .ZN(n18672) );
  INV_X1 U13217 ( .A(n18645), .ZN(n18702) );
  INV_X1 U13218 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18880) );
  INV_X1 U13219 ( .A(n18792), .ZN(n18876) );
  INV_X1 U13220 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18805) );
  AND2_X2 U13221 ( .A1(n13013), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20156)
         );
  INV_X1 U13222 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19871) );
  NAND2_X1 U13223 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10271) );
  AND2_X4 U13224 ( .A1(n13359), .A2(n10285), .ZN(n10475) );
  NAND2_X1 U13225 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10270) );
  NAND2_X1 U13226 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10269) );
  NAND2_X1 U13227 ( .A1(n11205), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10268) );
  NAND4_X1 U13228 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n10274) );
  INV_X2 U13229 ( .A(n10507), .ZN(n11010) );
  INV_X1 U13230 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10272) );
  NOR2_X1 U13231 ( .A1(n9742), .A2(n10272), .ZN(n10273) );
  NOR2_X1 U13232 ( .A1(n10274), .A2(n10273), .ZN(n10296) );
  INV_X1 U13233 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U13234 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10276) );
  NAND2_X1 U13235 ( .A1(n10419), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10275) );
  OAI211_X1 U13236 ( .C1(n11013), .C2(n10277), .A(n10276), .B(n10275), .ZN(
        n10278) );
  INV_X1 U13237 ( .A(n10278), .ZN(n10295) );
  NAND2_X1 U13238 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10283) );
  NAND2_X1 U13239 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10282) );
  NAND2_X1 U13240 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10281) );
  NAND2_X1 U13241 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10280) );
  NAND2_X1 U13242 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10292) );
  NAND2_X1 U13243 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10291) );
  NAND2_X1 U13244 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10290) );
  AND2_X4 U13245 ( .A1(n10288), .A2(n10286), .ZN(n11207) );
  NAND2_X1 U13246 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10289) );
  NAND2_X1 U13247 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10300) );
  NAND2_X1 U13248 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10299) );
  NAND2_X1 U13249 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10298) );
  NAND2_X1 U13250 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U13251 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10304) );
  NAND2_X1 U13252 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10303) );
  NAND2_X1 U13253 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U13254 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10301) );
  NAND4_X1 U13255 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10307) );
  NOR2_X1 U13256 ( .A1(n9742), .A2(n10305), .ZN(n10306) );
  NOR2_X1 U13257 ( .A1(n10307), .A2(n10306), .ZN(n10318) );
  NAND2_X1 U13258 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10311) );
  NAND2_X1 U13259 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10310) );
  NAND2_X1 U13260 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10309) );
  NAND2_X1 U13261 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10308) );
  INV_X1 U13262 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U13263 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U13264 ( .A1(n10419), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10312) );
  OAI211_X1 U13265 ( .C1(n11013), .C2(n10314), .A(n10313), .B(n10312), .ZN(
        n10315) );
  INV_X1 U13266 ( .A(n10315), .ZN(n10316) );
  INV_X1 U13267 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U13268 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10321) );
  NAND2_X1 U13269 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10320) );
  OAI211_X1 U13270 ( .C1(n9742), .C2(n10322), .A(n10321), .B(n10320), .ZN(
        n10323) );
  INV_X1 U13271 ( .A(n10323), .ZN(n10328) );
  INV_X1 U13272 ( .A(n10415), .ZN(n10324) );
  AOI22_X1 U13273 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10415), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13274 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10326) );
  NAND2_X1 U13275 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10325) );
  NAND4_X1 U13276 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10335) );
  INV_X2 U13277 ( .A(n11199), .ZN(n10976) );
  AOI22_X1 U13278 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13279 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10332) );
  INV_X4 U13280 ( .A(n11195), .ZN(n11126) );
  AOI22_X1 U13281 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10419), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13282 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10330) );
  NAND4_X1 U13283 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10334) );
  OR2_X2 U13284 ( .A1(n10335), .A2(n10334), .ZN(n11424) );
  NAND2_X1 U13285 ( .A1(n10437), .A2(n11424), .ZN(n10452) );
  NAND2_X1 U13286 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10339) );
  NAND2_X1 U13287 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10338) );
  NAND2_X1 U13288 ( .A1(n10419), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10337) );
  NAND2_X1 U13289 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10336) );
  NAND2_X1 U13290 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10343) );
  NAND2_X1 U13291 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10342) );
  NAND2_X1 U13292 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10341) );
  NAND2_X1 U13293 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10340) );
  NAND2_X1 U13294 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10347) );
  NAND2_X1 U13295 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10346) );
  NAND2_X1 U13296 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10345) );
  NAND2_X1 U13297 ( .A1(n11205), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10344) );
  NAND2_X1 U13298 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10351) );
  NAND2_X1 U13299 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10350) );
  OAI211_X1 U13300 ( .C1(n9742), .C2(n10352), .A(n10351), .B(n10350), .ZN(
        n10353) );
  INV_X1 U13301 ( .A(n10353), .ZN(n10354) );
  NAND2_X1 U13302 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10359) );
  NAND2_X1 U13303 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10358) );
  NAND2_X1 U13304 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10357) );
  NAND2_X1 U13305 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10356) );
  NAND4_X1 U13306 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10361) );
  NOR2_X1 U13307 ( .A1(n11013), .A2(n20977), .ZN(n10360) );
  NAND2_X1 U13308 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10365) );
  NAND2_X1 U13309 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10364) );
  NAND2_X1 U13310 ( .A1(n10746), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10363) );
  NAND2_X1 U13311 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10362) );
  NAND2_X1 U13312 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10369) );
  NAND2_X1 U13313 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10368) );
  NAND2_X1 U13314 ( .A1(n10419), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10367) );
  NAND2_X1 U13315 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10366) );
  INV_X1 U13316 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10372) );
  NAND2_X1 U13317 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10371) );
  NAND2_X1 U13318 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10370) );
  OAI211_X1 U13319 ( .C1(n9742), .C2(n10372), .A(n10371), .B(n10370), .ZN(
        n10373) );
  INV_X1 U13320 ( .A(n10373), .ZN(n10374) );
  INV_X1 U13321 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U13322 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10379) );
  NAND2_X1 U13323 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10378) );
  OAI211_X1 U13324 ( .C1(n9742), .C2(n10380), .A(n10379), .B(n10378), .ZN(
        n10381) );
  INV_X1 U13325 ( .A(n10381), .ZN(n10386) );
  AOI22_X1 U13326 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10415), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13327 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U13328 ( .A1(n10382), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10383) );
  NAND4_X1 U13329 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10392) );
  AOI22_X1 U13330 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13331 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13332 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10419), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13333 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10387) );
  NAND4_X1 U13334 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10391) );
  OR2_X2 U13335 ( .A1(n10392), .A2(n10391), .ZN(n13338) );
  NAND2_X1 U13336 ( .A1(n13136), .A2(n13338), .ZN(n10395) );
  INV_X1 U13337 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U13338 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10397) );
  NAND2_X1 U13339 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10396) );
  OAI211_X1 U13340 ( .C1(n9742), .C2(n10398), .A(n10397), .B(n10396), .ZN(
        n10399) );
  INV_X1 U13341 ( .A(n10399), .ZN(n10403) );
  AOI22_X1 U13342 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10415), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13343 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10401) );
  NAND2_X1 U13344 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10400) );
  NAND4_X1 U13345 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10409) );
  AOI22_X1 U13346 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13347 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13348 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10419), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U13349 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10404) );
  NAND4_X1 U13350 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10408) );
  OR2_X4 U13351 ( .A1(n10409), .A2(n10408), .ZN(n13428) );
  NOR2_X1 U13352 ( .A1(n10435), .A2(n13428), .ZN(n10410) );
  NAND4_X1 U13353 ( .A1(n20207), .A2(n20214), .A3(n20199), .A4(n14027), .ZN(
        n10411) );
  NAND2_X1 U13354 ( .A1(n11276), .A2(n14029), .ZN(n10424) );
  NAND2_X1 U13355 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10413) );
  AOI22_X1 U13356 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10415), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U13357 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10746), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13358 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10423) );
  AOI22_X1 U13359 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U13360 ( .A1(n10419), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U13361 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U13362 ( .A1(n20162), .A2(n13626), .ZN(n13741) );
  NAND2_X1 U13363 ( .A1(n10424), .A2(n14033), .ZN(n13424) );
  XNOR2_X1 U13364 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n10425) );
  NOR2_X2 U13365 ( .A1(n11424), .A2(n13338), .ZN(n13450) );
  NAND2_X1 U13366 ( .A1(n13450), .A2(n20207), .ZN(n13348) );
  NAND2_X1 U13367 ( .A1(n10451), .A2(n13337), .ZN(n10427) );
  NOR2_X1 U13368 ( .A1(n10429), .A2(n10428), .ZN(n10430) );
  NAND2_X2 U13369 ( .A1(n11424), .A2(n13626), .ZN(n11286) );
  NAND2_X1 U13370 ( .A1(n13136), .A2(n14035), .ZN(n13429) );
  NAND2_X1 U13371 ( .A1(n13428), .A2(n13338), .ZN(n10431) );
  AND2_X1 U13372 ( .A1(n13741), .A2(n10431), .ZN(n10433) );
  NAND2_X1 U13373 ( .A1(n20207), .A2(n12998), .ZN(n10434) );
  AND2_X1 U13374 ( .A1(n10434), .A2(n14027), .ZN(n10446) );
  OR2_X1 U13375 ( .A1(n10435), .A2(n12998), .ZN(n10436) );
  NAND2_X1 U13376 ( .A1(n13342), .A2(n20199), .ZN(n13328) );
  NAND2_X1 U13377 ( .A1(n13328), .A2(n13366), .ZN(n10455) );
  INV_X1 U13378 ( .A(n11424), .ZN(n20192) );
  NAND2_X1 U13379 ( .A1(n13501), .A2(n14015), .ZN(n13298) );
  OAI21_X1 U13380 ( .B1(n13344), .B2(n13450), .A(n20162), .ZN(n10439) );
  NAND2_X1 U13381 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10462) );
  OAI21_X1 U13382 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n10462), .ZN(n20487) );
  OR2_X1 U13383 ( .A1(n15819), .A2(n20490), .ZN(n10456) );
  OAI21_X1 U13384 ( .B1(n11520), .B2(n20487), .A(n10456), .ZN(n10441) );
  INV_X1 U13385 ( .A(n10441), .ZN(n10442) );
  MUX2_X1 U13386 ( .A(n11520), .B(n15819), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10444) );
  INV_X1 U13387 ( .A(n10445), .ZN(n10450) );
  INV_X1 U13388 ( .A(n10446), .ZN(n10447) );
  NAND2_X1 U13389 ( .A1(n10447), .A2(n13138), .ZN(n10448) );
  NAND2_X1 U13390 ( .A1(n13450), .A2(n20214), .ZN(n13426) );
  NAND4_X1 U13391 ( .A1(n10448), .A2(n13426), .A3(n19975), .A4(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n10449) );
  NOR2_X1 U13392 ( .A1(n10450), .A2(n10449), .ZN(n10454) );
  OAI21_X1 U13393 ( .B1(n10451), .B2(n10452), .A(n13344), .ZN(n10453) );
  OAI211_X1 U13394 ( .C1(n10455), .C2(n20177), .A(n10454), .B(n10453), .ZN(
        n10486) );
  NAND2_X1 U13395 ( .A1(n20289), .A2(n10545), .ZN(n10548) );
  INV_X1 U13396 ( .A(n10456), .ZN(n10459) );
  INV_X1 U13397 ( .A(n10457), .ZN(n10458) );
  OAI21_X1 U13398 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n10459), .A(
        n10458), .ZN(n10460) );
  INV_X1 U13399 ( .A(n10462), .ZN(n10461) );
  NAND2_X1 U13400 ( .A1(n10461), .A2(n20562), .ZN(n20524) );
  NAND2_X1 U13401 ( .A1(n10462), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10463) );
  INV_X1 U13402 ( .A(n15819), .ZN(n15812) );
  NAND2_X1 U13403 ( .A1(n15812), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13404 ( .A1(n13462), .A2(n10467), .ZN(n13445) );
  INV_X1 U13405 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U13406 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10469) );
  NAND2_X1 U13407 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10468) );
  OAI211_X1 U13408 ( .C1(n9742), .C2(n10482), .A(n10469), .B(n10468), .ZN(
        n10470) );
  INV_X1 U13409 ( .A(n10470), .ZN(n10474) );
  AOI22_X1 U13410 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10473) );
  INV_X2 U13411 ( .A(n10992), .ZN(n11094) );
  AOI22_X1 U13412 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10472) );
  NAND2_X1 U13413 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10471) );
  NAND4_X1 U13414 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10481) );
  AOI22_X1 U13415 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13416 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10478) );
  INV_X2 U13417 ( .A(n11193), .ZN(n10595) );
  AOI22_X1 U13418 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U13419 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10476) );
  NAND4_X1 U13420 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10480) );
  OAI22_X2 U13421 ( .A1(n13445), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11440), 
        .B2(n11243), .ZN(n10485) );
  OAI22_X1 U13422 ( .A1(n11260), .A2(n10482), .B1(n10586), .B2(n11440), .ZN(
        n10483) );
  INV_X1 U13423 ( .A(n10483), .ZN(n10484) );
  XNOR2_X2 U13424 ( .A(n10485), .B(n10484), .ZN(n10580) );
  INV_X1 U13425 ( .A(n10486), .ZN(n10487) );
  INV_X1 U13426 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10491) );
  NAND2_X1 U13427 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10490) );
  NAND2_X1 U13428 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10489) );
  OAI211_X1 U13429 ( .C1(n9742), .C2(n10491), .A(n10490), .B(n10489), .ZN(
        n10492) );
  INV_X1 U13430 ( .A(n10492), .ZN(n10496) );
  AOI22_X1 U13431 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13432 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10494) );
  NAND2_X1 U13433 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10493) );
  NAND4_X1 U13434 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .ZN(
        n10502) );
  AOI22_X1 U13435 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13436 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13437 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13438 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10497) );
  NAND4_X1 U13439 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10501) );
  NOR2_X1 U13440 ( .A1(n11243), .A2(n11490), .ZN(n10519) );
  NOR2_X1 U13441 ( .A1(n11243), .A2(n11496), .ZN(n10524) );
  NAND2_X1 U13442 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10506) );
  NAND2_X1 U13443 ( .A1(n11196), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10505) );
  NAND2_X1 U13444 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U13445 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10503) );
  AND4_X1 U13446 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10511) );
  AOI22_X1 U13447 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10510) );
  NAND2_X1 U13448 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10509) );
  NAND2_X1 U13449 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10508) );
  NAND4_X1 U13450 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10517) );
  AOI22_X1 U13451 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13452 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13453 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13454 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10512) );
  NAND4_X1 U13455 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10516) );
  MUX2_X1 U13456 ( .A(n10519), .B(n10524), .S(n11428), .Z(n10518) );
  INV_X1 U13457 ( .A(n10518), .ZN(n10568) );
  INV_X1 U13458 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20172) );
  INV_X1 U13459 ( .A(n10519), .ZN(n10543) );
  INV_X1 U13460 ( .A(n10520), .ZN(n10521) );
  NAND2_X1 U13461 ( .A1(n10543), .A2(n10521), .ZN(n10523) );
  INV_X1 U13462 ( .A(n11428), .ZN(n11438) );
  NAND2_X1 U13463 ( .A1(n20162), .A2(n11438), .ZN(n10522) );
  OAI211_X1 U13464 ( .C1(n11260), .C2(n20172), .A(n10523), .B(n10522), .ZN(
        n10566) );
  INV_X1 U13465 ( .A(n10524), .ZN(n10525) );
  INV_X1 U13466 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10544) );
  INV_X1 U13467 ( .A(n10586), .ZN(n10541) );
  NAND2_X1 U13468 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13469 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10529) );
  NAND2_X1 U13470 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10528) );
  NAND2_X1 U13471 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10527) );
  AND4_X1 U13472 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10534) );
  AOI22_X1 U13473 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13474 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10532) );
  NAND2_X1 U13475 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10531) );
  NAND4_X1 U13476 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n10540) );
  AOI22_X1 U13477 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13478 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13479 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13480 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10535) );
  NAND4_X1 U13481 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10539) );
  NAND2_X1 U13482 ( .A1(n10541), .A2(n11437), .ZN(n10542) );
  OAI211_X1 U13483 ( .C1(n11260), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        n10550) );
  INV_X1 U13484 ( .A(n20289), .ZN(n10547) );
  INV_X1 U13485 ( .A(n10545), .ZN(n10546) );
  INV_X1 U13486 ( .A(n11243), .ZN(n11421) );
  NAND2_X1 U13487 ( .A1(n11421), .A2(n11437), .ZN(n10549) );
  OAI21_X2 U13488 ( .B1(n14182), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10549), 
        .ZN(n11427) );
  AND2_X1 U13489 ( .A1(n11436), .A2(n10848), .ZN(n10559) );
  INV_X2 U13490 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20260) );
  NAND2_X1 U13491 ( .A1(n11225), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10577) );
  INV_X1 U13492 ( .A(n10577), .ZN(n10557) );
  INV_X1 U13493 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n10554) );
  XNOR2_X1 U13494 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13746) );
  AOI21_X1 U13495 ( .B1(n11279), .B2(n13746), .A(n11225), .ZN(n10553) );
  OAI21_X1 U13496 ( .B1(n11186), .B2(n10554), .A(n10553), .ZN(n10555) );
  AOI21_X1 U13497 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n10615), .A(
        n10555), .ZN(n10556) );
  NOR2_X1 U13498 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  XNOR2_X2 U13499 ( .A(n10560), .B(n11427), .ZN(n20606) );
  NAND2_X1 U13500 ( .A1(n20606), .A2(n10848), .ZN(n10565) );
  INV_X1 U13501 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n10562) );
  INV_X1 U13502 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10561) );
  OAI22_X1 U13503 ( .A1(n11186), .A2(n10562), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n10561), .ZN(n10563) );
  AOI21_X1 U13504 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n10615), .A(
        n10563), .ZN(n10564) );
  NAND2_X1 U13505 ( .A1(n10565), .A2(n10564), .ZN(n13293) );
  NAND2_X1 U13506 ( .A1(n20830), .A2(n20214), .ZN(n10569) );
  NAND2_X1 U13507 ( .A1(n10569), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13285) );
  INV_X1 U13508 ( .A(n10615), .ZN(n10640) );
  NAND2_X1 U13509 ( .A1(n20260), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10572) );
  NAND2_X1 U13510 ( .A1(n11226), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10571) );
  OAI211_X1 U13511 ( .C1(n10640), .C2(n13370), .A(n10572), .B(n10571), .ZN(
        n10573) );
  AOI21_X1 U13512 ( .B1(n10570), .B2(n10848), .A(n10573), .ZN(n10574) );
  OR2_X1 U13513 ( .A1(n13285), .A2(n10574), .ZN(n13286) );
  INV_X1 U13514 ( .A(n10574), .ZN(n13287) );
  OR2_X1 U13515 ( .A1(n13287), .A2(n11224), .ZN(n10575) );
  NAND2_X1 U13516 ( .A1(n13286), .A2(n10575), .ZN(n13292) );
  NAND2_X1 U13517 ( .A1(n13293), .A2(n13292), .ZN(n13377) );
  NAND2_X1 U13518 ( .A1(n13376), .A2(n10576), .ZN(n13378) );
  INV_X1 U13519 ( .A(n10578), .ZN(n10579) );
  NAND3_X1 U13520 ( .A1(n20825), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20376) );
  INV_X1 U13521 ( .A(n20376), .ZN(n20410) );
  NAND2_X1 U13522 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20410), .ZN(
        n20402) );
  NAND2_X1 U13523 ( .A1(n20825), .A2(n20402), .ZN(n10582) );
  NAND3_X1 U13524 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20687) );
  INV_X1 U13525 ( .A(n20687), .ZN(n20681) );
  NAND2_X1 U13526 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20681), .ZN(
        n20677) );
  NAND2_X1 U13527 ( .A1(n10582), .A2(n20677), .ZN(n20433) );
  OAI22_X1 U13528 ( .A1(n11520), .A2(n20433), .B1(n15819), .B2(n20825), .ZN(
        n10583) );
  INV_X1 U13529 ( .A(n10583), .ZN(n10584) );
  XNOR2_X2 U13530 ( .A(n13462), .B(n20322), .ZN(n20817) );
  NAND2_X1 U13531 ( .A1(n20817), .A2(n9880), .ZN(n10603) );
  INV_X1 U13532 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U13533 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10588) );
  NAND2_X1 U13534 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10587) );
  OAI211_X1 U13535 ( .C1(n9742), .C2(n10589), .A(n10588), .B(n10587), .ZN(
        n10590) );
  INV_X1 U13536 ( .A(n10590), .ZN(n10594) );
  INV_X2 U13537 ( .A(n11172), .ZN(n11093) );
  INV_X2 U13538 ( .A(n10324), .ZN(n11196) );
  AOI22_X1 U13539 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13540 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U13541 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10591) );
  NAND4_X1 U13542 ( .A1(n10594), .A2(n10593), .A3(n10592), .A4(n10591), .ZN(
        n10601) );
  AOI22_X1 U13543 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13544 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13545 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13546 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10596) );
  NAND4_X1 U13547 ( .A1(n10599), .A2(n10598), .A3(n10597), .A4(n10596), .ZN(
        n10600) );
  AOI22_X1 U13548 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11263), .B1(
        n11256), .B2(n11457), .ZN(n10602) );
  NAND2_X1 U13549 ( .A1(n10605), .A2(n20321), .ZN(n10606) );
  INV_X1 U13550 ( .A(n20812), .ZN(n10607) );
  INV_X1 U13551 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n10613) );
  NAND2_X1 U13552 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10609) );
  INV_X1 U13553 ( .A(n10609), .ZN(n10611) );
  INV_X1 U13554 ( .A(n10641), .ZN(n10610) );
  OAI21_X1 U13555 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10611), .A(
        n10610), .ZN(n14173) );
  AOI22_X1 U13556 ( .A1(n11279), .A2(n14173), .B1(n11225), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10612) );
  OAI21_X1 U13557 ( .B1(n11186), .B2(n10613), .A(n10612), .ZN(n10614) );
  AOI21_X1 U13558 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n10615), .A(
        n10614), .ZN(n10616) );
  NAND2_X1 U13559 ( .A1(n13482), .A2(n13481), .ZN(n13480) );
  NAND2_X1 U13560 ( .A1(n11263), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10633) );
  NAND2_X1 U13561 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10621) );
  NAND2_X1 U13562 ( .A1(n11196), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10620) );
  NAND2_X1 U13563 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10619) );
  NAND2_X1 U13564 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10618) );
  AND4_X1 U13565 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10625) );
  AOI22_X1 U13566 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10624) );
  NAND2_X1 U13567 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10623) );
  NAND2_X1 U13568 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10622) );
  NAND4_X1 U13569 ( .A1(n10625), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10631) );
  AOI22_X1 U13570 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13571 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10628) );
  INV_X1 U13572 ( .A(n11207), .ZN(n11059) );
  AOI22_X1 U13573 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10412), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13574 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11093), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10626) );
  NAND4_X1 U13575 ( .A1(n10629), .A2(n10628), .A3(n10627), .A4(n10626), .ZN(
        n10630) );
  NAND2_X1 U13576 ( .A1(n11256), .A2(n11461), .ZN(n10632) );
  NAND2_X1 U13577 ( .A1(n10636), .A2(n10635), .ZN(n10637) );
  AND2_X1 U13578 ( .A1(n10666), .A2(n10637), .ZN(n11456) );
  OAI21_X1 U13579 ( .B1(n20814), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20260), .ZN(n10639) );
  NAND2_X1 U13580 ( .A1(n11226), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10638) );
  OAI211_X1 U13581 ( .C1(n10640), .C2(n16169), .A(n10639), .B(n10638), .ZN(
        n10644) );
  NOR2_X1 U13582 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10641), .ZN(
        n10642) );
  NOR2_X1 U13583 ( .A1(n10668), .A2(n10642), .ZN(n13598) );
  NAND2_X1 U13584 ( .A1(n13598), .A2(n11279), .ZN(n10643) );
  AND2_X1 U13585 ( .A1(n10644), .A2(n10643), .ZN(n10645) );
  AOI21_X1 U13586 ( .B1(n11456), .B2(n10848), .A(n10645), .ZN(n13597) );
  INV_X1 U13587 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10650) );
  NAND2_X1 U13588 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10649) );
  NAND2_X1 U13589 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10648) );
  OAI211_X1 U13590 ( .C1(n9742), .C2(n10650), .A(n10649), .B(n10648), .ZN(
        n10651) );
  INV_X1 U13591 ( .A(n10651), .ZN(n10655) );
  AOI22_X1 U13592 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13593 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10653) );
  NAND2_X1 U13594 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10652) );
  NAND4_X1 U13595 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(
        n10661) );
  AOI22_X1 U13596 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13597 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13598 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13599 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10656) );
  NAND4_X1 U13600 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n10660) );
  NAND2_X1 U13601 ( .A1(n11256), .A2(n11479), .ZN(n10663) );
  OR2_X1 U13602 ( .A1(n11260), .A2(n10650), .ZN(n10662) );
  NAND2_X1 U13603 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  INV_X1 U13604 ( .A(n10664), .ZN(n10665) );
  NAND2_X1 U13605 ( .A1(n10666), .A2(n10665), .ZN(n10667) );
  NAND2_X1 U13606 ( .A1(n10694), .A2(n10667), .ZN(n11470) );
  INV_X1 U13607 ( .A(n11470), .ZN(n10673) );
  NOR2_X1 U13608 ( .A1(n10668), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10669) );
  NOR2_X1 U13609 ( .A1(n10688), .A2(n10669), .ZN(n20039) );
  INV_X1 U13610 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20043) );
  OAI22_X1 U13611 ( .A1(n20039), .A2(n11224), .B1(n10886), .B2(n20043), .ZN(
        n10670) );
  AOI21_X1 U13612 ( .B1(n11226), .B2(P1_EAX_REG_5__SCAN_IN), .A(n10670), .ZN(
        n10671) );
  INV_X1 U13613 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11167) );
  NAND2_X1 U13614 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10675) );
  NAND2_X1 U13615 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10674) );
  OAI211_X1 U13616 ( .C1(n9742), .C2(n11167), .A(n10675), .B(n10674), .ZN(
        n10676) );
  INV_X1 U13617 ( .A(n10676), .ZN(n10680) );
  AOI22_X1 U13618 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13619 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U13620 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10677) );
  NAND4_X1 U13621 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(
        n10687) );
  AOI22_X1 U13622 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13623 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13624 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13625 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10682) );
  NAND4_X1 U13626 ( .A1(n10685), .A2(n10684), .A3(n10683), .A4(n10682), .ZN(
        n10686) );
  NAND2_X1 U13627 ( .A1(n11256), .A2(n11488), .ZN(n10695) );
  OAI211_X1 U13628 ( .C1(n11167), .C2(n11260), .A(n10694), .B(n10695), .ZN(
        n11478) );
  NAND2_X1 U13629 ( .A1(n11478), .A2(n10848), .ZN(n10693) );
  INV_X1 U13630 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10690) );
  OAI21_X1 U13631 ( .B1(n10688), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n10698), .ZN(n20025) );
  AOI22_X1 U13632 ( .A1(n20025), .A2(n11279), .B1(n11225), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10689) );
  OAI21_X1 U13633 ( .B1(n11186), .B2(n10690), .A(n10689), .ZN(n10691) );
  INV_X1 U13634 ( .A(n10691), .ZN(n10692) );
  NAND2_X1 U13635 ( .A1(n10693), .A2(n10692), .ZN(n13711) );
  INV_X1 U13636 ( .A(n13710), .ZN(n10704) );
  NAND2_X1 U13637 ( .A1(n11256), .A2(n11490), .ZN(n10696) );
  OAI21_X1 U13638 ( .B1(n10491), .B2(n11260), .A(n10696), .ZN(n10697) );
  INV_X1 U13639 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13772) );
  NAND2_X1 U13640 ( .A1(n10698), .A2(n20883), .ZN(n10700) );
  INV_X1 U13641 ( .A(n10724), .ZN(n10699) );
  NAND2_X1 U13642 ( .A1(n10700), .A2(n10699), .ZN(n20010) );
  AOI22_X1 U13643 ( .A1(n20010), .A2(n11279), .B1(n11225), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10701) );
  OAI21_X1 U13644 ( .B1(n11186), .B2(n13772), .A(n10701), .ZN(n10702) );
  AOI21_X1 U13645 ( .B1(n11486), .B2(n10848), .A(n10702), .ZN(n13770) );
  INV_X1 U13646 ( .A(n13770), .ZN(n10703) );
  INV_X1 U13647 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13887) );
  XNOR2_X1 U13648 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10724), .ZN(
        n13913) );
  AOI22_X1 U13649 ( .A1(n11279), .A2(n13913), .B1(n11225), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10705) );
  OAI21_X1 U13650 ( .B1(n11186), .B2(n13887), .A(n10705), .ZN(n10722) );
  INV_X1 U13651 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10708) );
  NAND2_X1 U13652 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10707) );
  NAND2_X1 U13653 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10706) );
  OAI211_X1 U13654 ( .C1(n9742), .C2(n10708), .A(n10707), .B(n10706), .ZN(
        n10709) );
  INV_X1 U13655 ( .A(n10709), .ZN(n10713) );
  AOI22_X1 U13656 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13657 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10711) );
  NAND2_X1 U13658 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10710) );
  NAND4_X1 U13659 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10719) );
  AOI22_X1 U13660 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13661 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13662 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13663 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10714) );
  NAND4_X1 U13664 ( .A1(n10717), .A2(n10716), .A3(n10715), .A4(n10714), .ZN(
        n10718) );
  NOR2_X1 U13665 ( .A1(n10719), .A2(n10718), .ZN(n10720) );
  NOR2_X1 U13666 ( .A1(n10816), .A2(n10720), .ZN(n10721) );
  NOR2_X1 U13667 ( .A1(n10722), .A2(n10721), .ZN(n13856) );
  XOR2_X1 U13668 ( .A(n20001), .B(n10741), .Z(n20004) );
  INV_X1 U13669 ( .A(n20004), .ZN(n13965) );
  AOI22_X1 U13670 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13671 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13672 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13673 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10725) );
  NAND4_X1 U13674 ( .A1(n10728), .A2(n10727), .A3(n10726), .A4(n10725), .ZN(
        n10736) );
  AOI22_X1 U13675 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13676 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10729) );
  AND2_X1 U13677 ( .A1(n10730), .A2(n10729), .ZN(n10734) );
  AOI22_X1 U13678 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13679 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10732) );
  NAND2_X1 U13680 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10731) );
  NAND4_X1 U13681 ( .A1(n10734), .A2(n10733), .A3(n10732), .A4(n10731), .ZN(
        n10735) );
  OAI21_X1 U13682 ( .B1(n10736), .B2(n10735), .A(n10848), .ZN(n10739) );
  NAND2_X1 U13683 ( .A1(n11226), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10738) );
  NAND2_X1 U13684 ( .A1(n11225), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10737) );
  NAND3_X1 U13685 ( .A1(n10739), .A2(n10738), .A3(n10737), .ZN(n10740) );
  AOI21_X1 U13686 ( .B1(n13965), .B2(n11279), .A(n10740), .ZN(n13944) );
  INV_X1 U13687 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14504) );
  XNOR2_X1 U13688 ( .A(n10762), .B(n14504), .ZN(n15959) );
  OR2_X1 U13689 ( .A1(n15959), .A2(n11224), .ZN(n10761) );
  INV_X1 U13690 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U13691 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10743) );
  NAND2_X1 U13692 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10742) );
  OAI211_X1 U13693 ( .C1(n9742), .C2(n10744), .A(n10743), .B(n10742), .ZN(
        n10745) );
  INV_X1 U13694 ( .A(n10745), .ZN(n10750) );
  AOI22_X1 U13695 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13696 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U13697 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10747) );
  NAND4_X1 U13698 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10756) );
  AOI22_X1 U13699 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13700 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13701 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13702 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10751) );
  NAND4_X1 U13703 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10755) );
  NOR2_X1 U13704 ( .A1(n10756), .A2(n10755), .ZN(n10757) );
  OAI22_X1 U13705 ( .A1(n10816), .A2(n10757), .B1(n10886), .B2(n14504), .ZN(
        n10759) );
  INV_X1 U13706 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13972) );
  NOR2_X1 U13707 ( .A1(n11186), .A2(n13972), .ZN(n10758) );
  NOR2_X1 U13708 ( .A1(n10759), .A2(n10758), .ZN(n10760) );
  NAND2_X1 U13709 ( .A1(n10761), .A2(n10760), .ZN(n13954) );
  INV_X1 U13710 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14351) );
  OAI21_X1 U13711 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10763), .A(
        n10811), .ZN(n16017) );
  AOI22_X1 U13712 ( .A1(n11279), .A2(n16017), .B1(n11225), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10764) );
  OAI21_X1 U13713 ( .B1(n11186), .B2(n14351), .A(n10764), .ZN(n14153) );
  INV_X1 U13714 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U13715 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10766) );
  NAND2_X1 U13716 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10765) );
  OAI211_X1 U13717 ( .C1(n9742), .C2(n10767), .A(n10766), .B(n10765), .ZN(
        n10768) );
  INV_X1 U13718 ( .A(n10768), .ZN(n10772) );
  AOI22_X1 U13719 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11094), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13720 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U13721 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10769) );
  NAND4_X1 U13722 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10778) );
  AOI22_X1 U13723 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13724 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13725 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13726 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10773) );
  NAND4_X1 U13727 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        n10777) );
  NOR2_X1 U13728 ( .A1(n10778), .A2(n10777), .ZN(n10779) );
  NOR2_X1 U13729 ( .A1(n10816), .A2(n10779), .ZN(n14275) );
  AOI22_X1 U13730 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10329), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13731 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10780) );
  AND2_X1 U13732 ( .A1(n10781), .A2(n10780), .ZN(n10785) );
  AOI22_X1 U13733 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11093), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13734 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10783) );
  NAND2_X1 U13735 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10782) );
  NAND4_X1 U13736 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n10791) );
  AOI22_X1 U13737 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10412), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13738 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13739 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13740 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11094), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10786) );
  NAND4_X1 U13741 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10790) );
  NOR2_X1 U13742 ( .A1(n10791), .A2(n10790), .ZN(n10796) );
  NAND2_X1 U13743 ( .A1(n11226), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10795) );
  XNOR2_X1 U13744 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10811), .ZN(
        n16005) );
  INV_X1 U13745 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10792) );
  OAI22_X1 U13746 ( .A1(n16005), .A2(n11224), .B1(n10886), .B2(n10792), .ZN(
        n10793) );
  INV_X1 U13747 ( .A(n10793), .ZN(n10794) );
  OAI211_X1 U13748 ( .C1(n10796), .C2(n10816), .A(n10795), .B(n10794), .ZN(
        n14261) );
  INV_X1 U13749 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U13750 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10798) );
  NAND2_X1 U13751 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10797) );
  OAI211_X1 U13752 ( .C1(n9742), .C2(n10799), .A(n10798), .B(n10797), .ZN(
        n10800) );
  INV_X1 U13753 ( .A(n10800), .ZN(n10804) );
  AOI22_X1 U13754 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13755 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10802) );
  NAND2_X1 U13756 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10801) );
  NAND4_X1 U13757 ( .A1(n10804), .A2(n10803), .A3(n10802), .A4(n10801), .ZN(
        n10810) );
  AOI22_X1 U13758 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13759 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13760 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13761 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10805) );
  NAND4_X1 U13762 ( .A1(n10808), .A2(n10807), .A3(n10806), .A4(n10805), .ZN(
        n10809) );
  NOR2_X1 U13763 ( .A1(n10810), .A2(n10809), .ZN(n10817) );
  NAND2_X1 U13764 ( .A1(n11226), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10815) );
  INV_X1 U13765 ( .A(n10819), .ZN(n10813) );
  XNOR2_X1 U13766 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10813), .ZN(
        n14491) );
  AOI22_X1 U13767 ( .A1(n11279), .A2(n14491), .B1(n11225), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10814) );
  OAI211_X1 U13768 ( .C1(n10817), .C2(n10816), .A(n10815), .B(n10814), .ZN(
        n14157) );
  XOR2_X1 U13769 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n10835), .Z(
        n16000) );
  AOI22_X1 U13770 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13771 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13772 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13773 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10820) );
  AND4_X1 U13774 ( .A1(n10823), .A2(n10822), .A3(n10821), .A4(n10820), .ZN(
        n10830) );
  AOI22_X1 U13775 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13776 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13777 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U13778 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10824) );
  AND3_X1 U13779 ( .A1(n10826), .A2(n10825), .A3(n10824), .ZN(n10828) );
  NAND2_X1 U13780 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10827) );
  NAND4_X1 U13781 ( .A1(n10830), .A2(n10829), .A3(n10828), .A4(n10827), .ZN(
        n10831) );
  AOI22_X1 U13782 ( .A1(n10848), .A2(n10831), .B1(n11225), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10833) );
  NAND2_X1 U13783 ( .A1(n11226), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10832) );
  OAI211_X1 U13784 ( .C1(n16000), .C2(n11224), .A(n10833), .B(n10832), .ZN(
        n10834) );
  XNOR2_X1 U13785 ( .A(n10870), .B(n14478), .ZN(n15928) );
  NAND2_X1 U13786 ( .A1(n11226), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13787 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13788 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U13789 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10836) );
  AND3_X1 U13790 ( .A1(n10838), .A2(n10837), .A3(n10836), .ZN(n10846) );
  AOI22_X1 U13791 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13792 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13793 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13794 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10839) );
  AND4_X1 U13795 ( .A1(n10842), .A2(n10841), .A3(n10840), .A4(n10839), .ZN(
        n10845) );
  AOI22_X1 U13796 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U13797 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10843) );
  NAND4_X1 U13798 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10847) );
  NAND2_X1 U13799 ( .A1(n10848), .A2(n10847), .ZN(n10849) );
  OAI211_X1 U13800 ( .C1(n10886), .C2(n14478), .A(n10850), .B(n10849), .ZN(
        n10851) );
  AOI21_X1 U13801 ( .B1(n15928), .B2(n11279), .A(n10851), .ZN(n14251) );
  OR2_X2 U13802 ( .A1(n14248), .A2(n14251), .ZN(n14249) );
  INV_X1 U13803 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10854) );
  NAND2_X1 U13804 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10853) );
  NAND2_X1 U13805 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10852) );
  OAI211_X1 U13806 ( .C1(n9742), .C2(n10854), .A(n10853), .B(n10852), .ZN(
        n10855) );
  INV_X1 U13807 ( .A(n10855), .ZN(n10859) );
  AOI22_X1 U13808 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13809 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10857) );
  NAND2_X1 U13810 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10856) );
  NAND4_X1 U13811 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10865) );
  AOI22_X1 U13812 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13813 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11094), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13814 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13815 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10860) );
  NAND4_X1 U13816 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n10864) );
  NOR2_X1 U13817 ( .A1(n10865), .A2(n10864), .ZN(n10869) );
  NAND2_X1 U13818 ( .A1(n20260), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10866) );
  NAND2_X1 U13819 ( .A1(n11224), .A2(n10866), .ZN(n10867) );
  AOI21_X1 U13820 ( .B1(n11226), .B2(P1_EAX_REG_16__SCAN_IN), .A(n10867), .ZN(
        n10868) );
  OAI21_X1 U13821 ( .B1(n11221), .B2(n10869), .A(n10868), .ZN(n10873) );
  OAI21_X1 U13822 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10871), .A(
        n10906), .ZN(n15993) );
  OR2_X1 U13823 ( .A1(n11224), .A2(n15993), .ZN(n10872) );
  NAND2_X1 U13824 ( .A1(n10873), .A2(n10872), .ZN(n14238) );
  AOI22_X1 U13825 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13826 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13827 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13828 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10874) );
  AND4_X1 U13829 ( .A1(n10877), .A2(n10876), .A3(n10875), .A4(n10874), .ZN(
        n10884) );
  AOI22_X1 U13830 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U13831 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13832 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10879) );
  NAND2_X1 U13833 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10878) );
  AND3_X1 U13834 ( .A1(n10880), .A2(n10879), .A3(n10878), .ZN(n10882) );
  NAND2_X1 U13835 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10881) );
  NAND4_X1 U13836 ( .A1(n10884), .A2(n10883), .A3(n10882), .A4(n10881), .ZN(
        n10885) );
  NAND2_X1 U13837 ( .A1(n11188), .A2(n10885), .ZN(n10889) );
  XNOR2_X1 U13838 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10906), .ZN(
        n15910) );
  OAI22_X1 U13839 ( .A1(n11224), .A2(n15910), .B1(n10886), .B2(n15908), .ZN(
        n10887) );
  AOI21_X1 U13840 ( .B1(n11226), .B2(P1_EAX_REG_17__SCAN_IN), .A(n10887), .ZN(
        n10888) );
  NAND2_X1 U13841 ( .A1(n10889), .A2(n10888), .ZN(n14236) );
  AOI22_X1 U13842 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U13843 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10890) );
  AND2_X1 U13844 ( .A1(n10891), .A2(n10890), .ZN(n10895) );
  AOI22_X1 U13845 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13846 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U13847 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10892) );
  NAND4_X1 U13848 ( .A1(n10895), .A2(n10894), .A3(n10893), .A4(n10892), .ZN(
        n10902) );
  AOI22_X1 U13849 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13850 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13851 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13852 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10897) );
  NAND4_X1 U13853 ( .A1(n10900), .A2(n10899), .A3(n10898), .A4(n10897), .ZN(
        n10901) );
  NOR2_X1 U13854 ( .A1(n10902), .A2(n10901), .ZN(n10905) );
  OAI21_X1 U13855 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20814), .A(
        n20260), .ZN(n10904) );
  NAND2_X1 U13856 ( .A1(n11226), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n10903) );
  OAI211_X1 U13857 ( .C1(n11221), .C2(n10905), .A(n10904), .B(n10903), .ZN(
        n10909) );
  OAI21_X1 U13858 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10907), .A(
        n10943), .ZN(n15897) );
  OR2_X1 U13859 ( .A1(n11224), .A2(n15897), .ZN(n10908) );
  NAND2_X1 U13860 ( .A1(n10909), .A2(n10908), .ZN(n14226) );
  AOI22_X1 U13861 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13862 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U13863 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10911) );
  AND3_X1 U13864 ( .A1(n10913), .A2(n10912), .A3(n10911), .ZN(n10921) );
  AOI22_X1 U13865 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13866 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13867 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13868 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10914) );
  AND4_X1 U13869 ( .A1(n10917), .A2(n10916), .A3(n10915), .A4(n10914), .ZN(
        n10920) );
  AOI22_X1 U13870 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10919) );
  NAND2_X1 U13871 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10918) );
  NAND4_X1 U13872 ( .A1(n10921), .A2(n10920), .A3(n10919), .A4(n10918), .ZN(
        n10922) );
  NAND2_X1 U13873 ( .A1(n11188), .A2(n10922), .ZN(n10925) );
  OAI21_X1 U13874 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14450), .A(n11224), 
        .ZN(n10923) );
  AOI21_X1 U13875 ( .B1(n11226), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10923), .ZN(
        n10924) );
  NAND2_X1 U13876 ( .A1(n10925), .A2(n10924), .ZN(n10927) );
  XNOR2_X1 U13877 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n10943), .ZN(
        n15894) );
  NAND2_X1 U13878 ( .A1(n15894), .A2(n11279), .ZN(n10926) );
  NAND2_X1 U13879 ( .A1(n10927), .A2(n10926), .ZN(n14220) );
  AOI22_X1 U13880 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10929) );
  NAND2_X1 U13881 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10928) );
  AND2_X1 U13882 ( .A1(n10929), .A2(n10928), .ZN(n10933) );
  AOI22_X1 U13883 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11093), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13884 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11094), .B1(
        n11126), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10931) );
  NAND2_X1 U13885 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10930) );
  NAND4_X1 U13886 ( .A1(n10933), .A2(n10932), .A3(n10931), .A4(n10930), .ZN(
        n10939) );
  AOI22_X1 U13887 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10475), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13888 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13889 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U13890 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10934) );
  NAND4_X1 U13891 ( .A1(n10937), .A2(n10936), .A3(n10935), .A4(n10934), .ZN(
        n10938) );
  NOR2_X1 U13892 ( .A1(n10939), .A2(n10938), .ZN(n10940) );
  OR2_X1 U13893 ( .A1(n11221), .A2(n10940), .ZN(n10947) );
  NAND2_X1 U13894 ( .A1(n20260), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10941) );
  NAND2_X1 U13895 ( .A1(n11224), .A2(n10941), .ZN(n10942) );
  AOI21_X1 U13896 ( .B1(n11226), .B2(P1_EAX_REG_20__SCAN_IN), .A(n10942), .ZN(
        n10946) );
  OAI21_X1 U13897 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10944), .A(
        n10987), .ZN(n14442) );
  NOR2_X1 U13898 ( .A1(n14442), .A2(n11224), .ZN(n10945) );
  AOI21_X1 U13899 ( .B1(n10947), .B2(n10946), .A(n10945), .ZN(n14146) );
  INV_X1 U13900 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U13901 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10949) );
  NAND2_X1 U13902 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10948) );
  OAI211_X1 U13903 ( .C1(n11193), .C2(n11119), .A(n10949), .B(n10948), .ZN(
        n10950) );
  INV_X1 U13904 ( .A(n10950), .ZN(n10954) );
  AOI22_X1 U13905 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U13906 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10952) );
  NAND2_X1 U13907 ( .A1(n11010), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10951) );
  NAND4_X1 U13908 ( .A1(n10954), .A2(n10953), .A3(n10952), .A4(n10951), .ZN(
        n10960) );
  AOI22_X1 U13909 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13910 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13911 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13912 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10955) );
  NAND4_X1 U13913 ( .A1(n10958), .A2(n10957), .A3(n10956), .A4(n10955), .ZN(
        n10959) );
  NOR2_X1 U13914 ( .A1(n10960), .A2(n10959), .ZN(n10963) );
  AOI21_X1 U13915 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15984), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10961) );
  AOI21_X1 U13916 ( .B1(n11226), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10961), .ZN(
        n10962) );
  OAI21_X1 U13917 ( .B1(n11221), .B2(n10963), .A(n10962), .ZN(n10965) );
  XNOR2_X1 U13918 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n10987), .ZN(
        n15981) );
  NAND2_X1 U13919 ( .A1(n15981), .A2(n11279), .ZN(n10964) );
  INV_X1 U13920 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U13921 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10967) );
  NAND2_X1 U13922 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10966) );
  OAI211_X1 U13923 ( .C1(n9742), .C2(n10968), .A(n10967), .B(n10966), .ZN(
        n10969) );
  INV_X1 U13924 ( .A(n10969), .ZN(n10975) );
  AOI22_X1 U13925 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13926 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10973) );
  NAND2_X1 U13927 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10972) );
  NAND4_X1 U13928 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10982) );
  AOI22_X1 U13929 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U13930 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U13931 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13932 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10977) );
  NAND4_X1 U13933 ( .A1(n10980), .A2(n10979), .A3(n10978), .A4(n10977), .ZN(
        n10981) );
  NOR2_X1 U13934 ( .A1(n10982), .A2(n10981), .ZN(n10986) );
  NAND2_X1 U13935 ( .A1(n20260), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10983) );
  NAND2_X1 U13936 ( .A1(n11224), .A2(n10983), .ZN(n10984) );
  AOI21_X1 U13937 ( .B1(n11226), .B2(P1_EAX_REG_22__SCAN_IN), .A(n10984), .ZN(
        n10985) );
  OAI21_X1 U13938 ( .B1(n11221), .B2(n10986), .A(n10985), .ZN(n10990) );
  OAI21_X1 U13939 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10988), .A(
        n11024), .ZN(n15977) );
  OR2_X1 U13940 ( .A1(n11224), .A2(n15977), .ZN(n10989) );
  NAND2_X1 U13941 ( .A1(n10990), .A2(n10989), .ZN(n14203) );
  INV_X1 U13942 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10999) );
  INV_X1 U13943 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10991) );
  OAI22_X1 U13944 ( .A1(n10992), .A2(n10991), .B1(n11168), .B2(n20172), .ZN(
        n10996) );
  INV_X1 U13945 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10994) );
  INV_X1 U13946 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10993) );
  OAI22_X1 U13947 ( .A1(n11172), .A2(n10994), .B1(n10324), .B2(n10993), .ZN(
        n10995) );
  AOI211_X1 U13948 ( .C1(n10971), .C2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n10996), .B(n10995), .ZN(n10998) );
  AOI22_X1 U13949 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10997) );
  OAI211_X1 U13950 ( .C1(n9742), .C2(n10999), .A(n10998), .B(n10997), .ZN(
        n11005) );
  AOI22_X1 U13951 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U13952 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U13953 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13954 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11000) );
  NAND4_X1 U13955 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11004) );
  NOR2_X1 U13956 ( .A1(n11005), .A2(n11004), .ZN(n11030) );
  INV_X1 U13957 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11198) );
  INV_X1 U13958 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11194) );
  INV_X1 U13959 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11192) );
  OAI22_X1 U13960 ( .A1(n10992), .A2(n11194), .B1(n10324), .B2(n11192), .ZN(
        n11009) );
  INV_X1 U13961 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11007) );
  INV_X1 U13962 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11006) );
  OAI22_X1 U13963 ( .A1(n11199), .A2(n11007), .B1(n11087), .B2(n11006), .ZN(
        n11008) );
  AOI211_X1 U13964 ( .C1(n11010), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11009), .B(n11008), .ZN(n11012) );
  AOI22_X1 U13965 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11011) );
  OAI211_X1 U13966 ( .C1(n11013), .C2(n11198), .A(n11012), .B(n11011), .ZN(
        n11019) );
  AOI22_X1 U13967 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U13968 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U13969 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U13970 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11014) );
  NAND4_X1 U13971 ( .A1(n11017), .A2(n11016), .A3(n11015), .A4(n11014), .ZN(
        n11018) );
  NOR2_X1 U13972 ( .A1(n11019), .A2(n11018), .ZN(n11029) );
  XOR2_X1 U13973 ( .A(n11030), .B(n11029), .Z(n11020) );
  NAND2_X1 U13974 ( .A1(n11020), .A2(n11188), .ZN(n11023) );
  INV_X1 U13975 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20941) );
  OAI21_X1 U13976 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20941), .A(n11224), 
        .ZN(n11021) );
  AOI21_X1 U13977 ( .B1(n11226), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11021), .ZN(
        n11022) );
  NAND2_X1 U13978 ( .A1(n11023), .A2(n11022), .ZN(n11028) );
  NAND2_X1 U13979 ( .A1(n20941), .A2(n11024), .ZN(n11026) );
  AND2_X1 U13980 ( .A1(n11026), .A2(n11051), .ZN(n14434) );
  NAND2_X1 U13981 ( .A1(n14434), .A2(n11279), .ZN(n11027) );
  NAND2_X1 U13982 ( .A1(n11028), .A2(n11027), .ZN(n14135) );
  NOR2_X1 U13983 ( .A1(n11030), .A2(n11029), .ZN(n11057) );
  INV_X1 U13984 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11033) );
  NAND2_X1 U13985 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11032) );
  NAND2_X1 U13986 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11031) );
  OAI211_X1 U13987 ( .C1(n9742), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        n11034) );
  INV_X1 U13988 ( .A(n11034), .ZN(n11038) );
  AOI22_X1 U13989 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U13990 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U13991 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11035) );
  NAND4_X1 U13992 ( .A1(n11038), .A2(n11037), .A3(n11036), .A4(n11035), .ZN(
        n11044) );
  AOI22_X1 U13993 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U13994 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11041) );
  INV_X1 U13995 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U13996 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U13997 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11039) );
  NAND4_X1 U13998 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(
        n11043) );
  OR2_X1 U13999 ( .A1(n11044), .A2(n11043), .ZN(n11056) );
  INV_X1 U14000 ( .A(n11056), .ZN(n11045) );
  XNOR2_X1 U14001 ( .A(n11057), .B(n11045), .ZN(n11046) );
  NAND2_X1 U14002 ( .A1(n11046), .A2(n11188), .ZN(n11055) );
  NAND2_X1 U14003 ( .A1(n20260), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11047) );
  NAND2_X1 U14004 ( .A1(n11224), .A2(n11047), .ZN(n11048) );
  AOI21_X1 U14005 ( .B1(n11226), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11048), .ZN(
        n11054) );
  INV_X1 U14006 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11050) );
  NAND2_X1 U14007 ( .A1(n11051), .A2(n11050), .ZN(n11052) );
  NAND2_X1 U14008 ( .A1(n11078), .A2(n11052), .ZN(n14420) );
  NOR2_X1 U14009 ( .A1(n14420), .A2(n11224), .ZN(n11053) );
  AOI21_X1 U14010 ( .B1(n11055), .B2(n11054), .A(n11053), .ZN(n14115) );
  NAND2_X1 U14011 ( .A1(n11057), .A2(n11056), .ZN(n11101) );
  INV_X1 U14012 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11067) );
  INV_X1 U14013 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11060) );
  INV_X1 U14014 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11058) );
  OAI22_X1 U14015 ( .A1(n11087), .A2(n11060), .B1(n11059), .B2(n11058), .ZN(
        n11064) );
  INV_X1 U14016 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11062) );
  INV_X1 U14017 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11061) );
  OAI22_X1 U14018 ( .A1(n11199), .A2(n11062), .B1(n10992), .B2(n11061), .ZN(
        n11063) );
  AOI211_X1 U14019 ( .C1(n10971), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n11064), .B(n11063), .ZN(n11066) );
  AOI22_X1 U14020 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11065) );
  OAI211_X1 U14021 ( .C1(n9742), .C2(n11067), .A(n11066), .B(n11065), .ZN(
        n11074) );
  AOI22_X1 U14022 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14023 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14024 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14025 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11069) );
  NAND4_X1 U14026 ( .A1(n11072), .A2(n11071), .A3(n11070), .A4(n11069), .ZN(
        n11073) );
  NOR2_X1 U14027 ( .A1(n11074), .A2(n11073), .ZN(n11102) );
  XOR2_X1 U14028 ( .A(n11101), .B(n11102), .Z(n11075) );
  NAND2_X1 U14029 ( .A1(n11075), .A2(n11188), .ZN(n11082) );
  INV_X1 U14030 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n20911) );
  OAI21_X1 U14031 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20911), .A(n11224), 
        .ZN(n11076) );
  AOI21_X1 U14032 ( .B1(n11226), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11076), .ZN(
        n11081) );
  NAND2_X1 U14033 ( .A1(n11078), .A2(n20911), .ZN(n11079) );
  NAND2_X1 U14034 ( .A1(n11157), .A2(n11079), .ZN(n14412) );
  NOR2_X1 U14035 ( .A1(n14412), .A2(n11224), .ZN(n11080) );
  AOI21_X1 U14036 ( .B1(n11082), .B2(n11081), .A(n11080), .ZN(n14105) );
  INV_X1 U14037 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11092) );
  INV_X1 U14038 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11084) );
  INV_X1 U14039 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11083) );
  OAI22_X1 U14040 ( .A1(n11199), .A2(n11084), .B1(n11168), .B2(n11083), .ZN(
        n11089) );
  INV_X1 U14041 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11086) );
  INV_X1 U14042 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11085) );
  OAI22_X1 U14043 ( .A1(n11087), .A2(n11086), .B1(n11195), .B2(n11085), .ZN(
        n11088) );
  AOI211_X1 U14044 ( .C1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .C2(n10971), .A(
        n11089), .B(n11088), .ZN(n11091) );
  AOI22_X1 U14045 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10412), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11090) );
  OAI211_X1 U14046 ( .C1(n11092), .C2(n9742), .A(n11091), .B(n11090), .ZN(
        n11100) );
  AOI22_X1 U14047 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11093), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14048 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11094), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14049 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U14050 ( .A1(n10681), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11095) );
  NAND4_X1 U14051 ( .A1(n11098), .A2(n11097), .A3(n11096), .A4(n11095), .ZN(
        n11099) );
  NOR2_X1 U14052 ( .A1(n11100), .A2(n11099), .ZN(n11143) );
  NOR2_X1 U14053 ( .A1(n11102), .A2(n11101), .ZN(n11153) );
  INV_X1 U14054 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14055 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11104) );
  NAND2_X1 U14056 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11103) );
  OAI211_X1 U14057 ( .C1(n9742), .C2(n11105), .A(n11104), .B(n11103), .ZN(
        n11106) );
  INV_X1 U14058 ( .A(n11106), .ZN(n11110) );
  AOI22_X1 U14059 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14060 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11108) );
  NAND2_X1 U14061 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11107) );
  NAND4_X1 U14062 ( .A1(n11110), .A2(n11109), .A3(n11108), .A4(n11107), .ZN(
        n11116) );
  AOI22_X1 U14063 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14064 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14065 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14066 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11111) );
  NAND4_X1 U14067 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(
        n11115) );
  OR2_X1 U14068 ( .A1(n11116), .A2(n11115), .ZN(n11151) );
  NAND2_X1 U14069 ( .A1(n11153), .A2(n11151), .ZN(n11144) );
  NOR2_X1 U14070 ( .A1(n11143), .A2(n11144), .ZN(n11166) );
  NAND2_X1 U14071 ( .A1(n10896), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11118) );
  NAND2_X1 U14072 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11117) );
  OAI211_X1 U14073 ( .C1(n9742), .C2(n11119), .A(n11118), .B(n11117), .ZN(
        n11120) );
  INV_X1 U14074 ( .A(n11120), .ZN(n11124) );
  AOI22_X1 U14075 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U14076 ( .A1(n11094), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U14077 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11121) );
  NAND4_X1 U14078 ( .A1(n11124), .A2(n11123), .A3(n11122), .A4(n11121), .ZN(
        n11132) );
  AOI22_X1 U14079 ( .A1(n11125), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11206), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11130) );
  INV_X1 U14080 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n20939) );
  AOI22_X1 U14081 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14082 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10595), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14083 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11127) );
  NAND4_X1 U14084 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11131) );
  OR2_X1 U14085 ( .A1(n11132), .A2(n11131), .ZN(n11165) );
  INV_X1 U14086 ( .A(n11165), .ZN(n11133) );
  XNOR2_X1 U14087 ( .A(n11166), .B(n11133), .ZN(n11136) );
  INV_X1 U14088 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14291) );
  NAND2_X1 U14089 ( .A1(n20260), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11134) );
  OAI211_X1 U14090 ( .C1(n11186), .C2(n14291), .A(n11224), .B(n11134), .ZN(
        n11135) );
  AOI21_X1 U14091 ( .B1(n11136), .B2(n11188), .A(n11135), .ZN(n11142) );
  INV_X1 U14092 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14396) );
  INV_X1 U14093 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U14094 ( .A1(n11139), .A2(n11138), .ZN(n11140) );
  NAND2_X1 U14095 ( .A1(n11163), .A2(n11140), .ZN(n14385) );
  NOR2_X1 U14096 ( .A1(n14385), .A2(n11224), .ZN(n11141) );
  XOR2_X1 U14097 ( .A(n11144), .B(n11143), .Z(n11145) );
  NAND2_X1 U14098 ( .A1(n11145), .A2(n11188), .ZN(n11148) );
  AOI21_X1 U14099 ( .B1(n14396), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11146) );
  AOI21_X1 U14100 ( .B1(n11226), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11146), .ZN(
        n11147) );
  NAND2_X1 U14101 ( .A1(n11148), .A2(n11147), .ZN(n11150) );
  XNOR2_X1 U14102 ( .A(n11159), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14394) );
  NAND2_X1 U14103 ( .A1(n14394), .A2(n11279), .ZN(n11149) );
  NAND2_X1 U14104 ( .A1(n11150), .A2(n11149), .ZN(n14082) );
  INV_X1 U14105 ( .A(n11151), .ZN(n11152) );
  XNOR2_X1 U14106 ( .A(n11153), .B(n11152), .ZN(n11156) );
  INV_X1 U14107 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14304) );
  NAND2_X1 U14108 ( .A1(n20260), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11154) );
  OAI211_X1 U14109 ( .C1(n11186), .C2(n14304), .A(n11224), .B(n11154), .ZN(
        n11155) );
  AOI21_X1 U14110 ( .B1(n11156), .B2(n11188), .A(n11155), .ZN(n11161) );
  INV_X1 U14111 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U14112 ( .A1(n11157), .A2(n14093), .ZN(n11158) );
  NAND2_X1 U14113 ( .A1(n11159), .A2(n11158), .ZN(n14403) );
  NOR2_X1 U14114 ( .A1(n14403), .A2(n11224), .ZN(n11160) );
  INV_X1 U14115 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20944) );
  NAND2_X1 U14116 ( .A1(n11163), .A2(n20944), .ZN(n11164) );
  NAND2_X1 U14117 ( .A1(n11166), .A2(n11165), .ZN(n11215) );
  INV_X1 U14118 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11177) );
  INV_X1 U14119 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11169) );
  OAI22_X1 U14120 ( .A1(n11199), .A2(n11169), .B1(n11168), .B2(n11167), .ZN(
        n11174) );
  INV_X1 U14121 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11171) );
  INV_X1 U14122 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11170) );
  OAI22_X1 U14123 ( .A1(n11172), .A2(n11171), .B1(n10992), .B2(n11170), .ZN(
        n11173) );
  AOI211_X1 U14124 ( .C1(n10971), .C2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n11174), .B(n11173), .ZN(n11176) );
  AOI22_X1 U14125 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U14126 ( .C1(n9742), .C2(n11177), .A(n11176), .B(n11175), .ZN(
        n11183) );
  AOI22_X1 U14127 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11196), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14128 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10412), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14129 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14130 ( .A1(n10595), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11178) );
  NAND4_X1 U14131 ( .A1(n11181), .A2(n11180), .A3(n11179), .A4(n11178), .ZN(
        n11182) );
  NOR2_X1 U14132 ( .A1(n11183), .A2(n11182), .ZN(n11216) );
  XOR2_X1 U14133 ( .A(n11215), .B(n11216), .Z(n11189) );
  INV_X1 U14134 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n11185) );
  NOR2_X1 U14135 ( .A1(n20814), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11184) );
  OAI22_X1 U14136 ( .A1(n11186), .A2(n11185), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11184), .ZN(n11187) );
  AOI21_X1 U14137 ( .B1(n11189), .B2(n11188), .A(n11187), .ZN(n11190) );
  AOI21_X1 U14138 ( .B1(n11279), .B2(n14369), .A(n11190), .ZN(n14058) );
  INV_X1 U14139 ( .A(n11282), .ZN(n11191) );
  XNOR2_X1 U14140 ( .A(n11191), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14363) );
  INV_X1 U14141 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11204) );
  OAI22_X1 U14142 ( .A1(n11195), .A2(n11194), .B1(n11193), .B2(n11192), .ZN(
        n11201) );
  INV_X1 U14143 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11197) );
  OAI22_X1 U14144 ( .A1(n11199), .A2(n11198), .B1(n10324), .B2(n11197), .ZN(
        n11200) );
  AOI211_X1 U14145 ( .C1(n10971), .C2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n11201), .B(n11200), .ZN(n11203) );
  AOI22_X1 U14146 ( .A1(n10412), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10896), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11202) );
  OAI211_X1 U14147 ( .C1(n9742), .C2(n11204), .A(n11203), .B(n11202), .ZN(
        n11214) );
  AOI22_X1 U14148 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11094), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14149 ( .A1(n10475), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10681), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14150 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11205), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14151 ( .A1(n10329), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11209) );
  NAND4_X1 U14152 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11213) );
  NOR2_X1 U14153 ( .A1(n11214), .A2(n11213), .ZN(n11218) );
  NOR2_X1 U14154 ( .A1(n11216), .A2(n11215), .ZN(n11217) );
  XOR2_X1 U14155 ( .A(n11218), .B(n11217), .Z(n11222) );
  AOI21_X1 U14156 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20260), .A(
        n11279), .ZN(n11220) );
  NAND2_X1 U14157 ( .A1(n11226), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11219) );
  OAI211_X1 U14158 ( .C1(n11222), .C2(n11221), .A(n11220), .B(n11219), .ZN(
        n11223) );
  OAI21_X1 U14159 ( .B1(n11224), .B2(n14363), .A(n11223), .ZN(n14044) );
  AOI22_X1 U14160 ( .A1(n11226), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11225), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11227) );
  XNOR2_X1 U14161 ( .A(n14043), .B(n11227), .ZN(n13003) );
  XNOR2_X1 U14162 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U14163 ( .A1(n20834), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11242) );
  NAND2_X1 U14164 ( .A1(n11239), .A2(n11238), .ZN(n11229) );
  NAND2_X1 U14165 ( .A1(n20490), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11228) );
  NAND2_X1 U14166 ( .A1(n11229), .A2(n11228), .ZN(n11250) );
  MUX2_X1 U14167 ( .A(n20562), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11249) );
  NAND2_X1 U14168 ( .A1(n11250), .A2(n11249), .ZN(n11231) );
  NAND2_X1 U14169 ( .A1(n20562), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11230) );
  NAND2_X1 U14170 ( .A1(n11231), .A2(n11230), .ZN(n11236) );
  XNOR2_X1 U14171 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11237) );
  INV_X1 U14172 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20150) );
  NOR2_X1 U14173 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20150), .ZN(
        n11232) );
  NAND2_X1 U14174 ( .A1(n11275), .A2(n11262), .ZN(n11268) );
  NAND2_X1 U14175 ( .A1(n11275), .A2(n11256), .ZN(n11267) );
  NAND3_X1 U14176 ( .A1(n16169), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11233), .ZN(n11273) );
  INV_X1 U14177 ( .A(n11262), .ZN(n11266) );
  INV_X1 U14178 ( .A(n11234), .ZN(n11235) );
  OAI21_X1 U14179 ( .B1(n11237), .B2(n11236), .A(n11235), .ZN(n11272) );
  XNOR2_X1 U14180 ( .A(n11239), .B(n11238), .ZN(n11270) );
  NOR2_X1 U14181 ( .A1(n14281), .A2(n9880), .ZN(n11240) );
  AOI21_X1 U14182 ( .B1(n20177), .B2(n14281), .A(n11247), .ZN(n11241) );
  INV_X1 U14183 ( .A(n11256), .ZN(n11253) );
  OAI21_X1 U14184 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20834), .A(
        n11242), .ZN(n11245) );
  NOR2_X1 U14185 ( .A1(n11253), .A2(n11245), .ZN(n11246) );
  AND2_X1 U14186 ( .A1(n20207), .A2(n13428), .ZN(n14017) );
  INV_X1 U14187 ( .A(n13741), .ZN(n13296) );
  AOI211_X1 U14188 ( .C1(n11243), .C2(n13626), .A(n14017), .B(n13296), .ZN(
        n11244) );
  OAI22_X1 U14189 ( .A1(n11262), .A2(n11246), .B1(n11245), .B2(n11244), .ZN(
        n11248) );
  XNOR2_X1 U14190 ( .A(n11250), .B(n11249), .ZN(n11271) );
  INV_X1 U14191 ( .A(n14017), .ZN(n11251) );
  NAND2_X1 U14192 ( .A1(n11251), .A2(n20177), .ZN(n11255) );
  NAND2_X1 U14193 ( .A1(n11263), .A2(n11271), .ZN(n11252) );
  OAI211_X1 U14194 ( .C1(n11253), .C2(n11271), .A(n11255), .B(n11252), .ZN(
        n11254) );
  INV_X1 U14195 ( .A(n11271), .ZN(n11258) );
  INV_X1 U14196 ( .A(n11255), .ZN(n11257) );
  NAND3_X1 U14197 ( .A1(n11258), .A2(n11257), .A3(n11256), .ZN(n11259) );
  AOI21_X1 U14198 ( .B1(n11262), .B2(n11272), .A(n11261), .ZN(n11265) );
  NOR2_X1 U14199 ( .A1(n11263), .A2(n11273), .ZN(n11264) );
  NOR2_X1 U14200 ( .A1(n14029), .A2(n19976), .ZN(n11269) );
  NOR3_X1 U14201 ( .A1(n11272), .A2(n11271), .A3(n11270), .ZN(n11274) );
  OAI21_X1 U14202 ( .B1(n11275), .B2(n11274), .A(n11273), .ZN(n14023) );
  INV_X1 U14203 ( .A(n11276), .ZN(n11277) );
  NAND2_X1 U14204 ( .A1(n14030), .A2(n13420), .ZN(n13046) );
  OR2_X2 U14205 ( .A1(n11520), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20042) );
  INV_X2 U14206 ( .A(n20042), .ZN(n20135) );
  NOR2_X1 U14207 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20852) );
  NAND2_X1 U14208 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20852), .ZN(n16174) );
  AND2_X1 U14209 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n9880), .ZN(n11278) );
  NAND2_X1 U14210 ( .A1(n11279), .A2(n11278), .ZN(n11280) );
  OAI21_X1 U14211 ( .B1(n16174), .B2(n9880), .A(n11280), .ZN(n11281) );
  INV_X1 U14212 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14045) );
  XNOR2_X1 U14213 ( .A(n11283), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13744) );
  NOR2_X1 U14214 ( .A1(n13744), .A2(n11284), .ZN(n11285) );
  NAND2_X1 U14215 ( .A1(n13003), .A2(n20031), .ZN(n11419) );
  AOI22_X1 U14216 ( .A1(n13501), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n11302), .ZN(n14040) );
  NOR2_X1 U14217 ( .A1(n11286), .A2(n11302), .ZN(n11287) );
  CLKBUF_X3 U14218 ( .A(n11287), .Z(n11387) );
  INV_X1 U14219 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13307) );
  NAND2_X1 U14220 ( .A1(n11387), .A2(n13307), .ZN(n11291) );
  INV_X1 U14221 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U14222 ( .A1(n9748), .A2(n11288), .ZN(n11289) );
  OAI211_X1 U14223 ( .C1(n11302), .C2(P1_EBX_REG_1__SCAN_IN), .A(n11289), .B(
        n11383), .ZN(n11290) );
  NAND2_X1 U14224 ( .A1(n11291), .A2(n11290), .ZN(n11295) );
  NAND2_X1 U14225 ( .A1(n9748), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11294) );
  INV_X1 U14226 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11292) );
  NAND2_X1 U14227 ( .A1(n11383), .A2(n11292), .ZN(n11293) );
  NAND2_X1 U14228 ( .A1(n11294), .A2(n11293), .ZN(n13502) );
  XNOR2_X1 U14229 ( .A(n11295), .B(n13502), .ZN(n13304) );
  NAND2_X1 U14230 ( .A1(n13304), .A2(n13303), .ZN(n13306) );
  NAND2_X1 U14231 ( .A1(n13306), .A2(n11295), .ZN(n13402) );
  INV_X1 U14232 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13404) );
  NAND2_X1 U14233 ( .A1(n11387), .A2(n13404), .ZN(n11298) );
  INV_X1 U14234 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U14235 ( .A1(n9748), .A2(n13493), .ZN(n11296) );
  OAI211_X1 U14236 ( .C1(n11302), .C2(P1_EBX_REG_2__SCAN_IN), .A(n11296), .B(
        n11383), .ZN(n11297) );
  AND2_X1 U14237 ( .A1(n11298), .A2(n11297), .ZN(n13401) );
  MUX2_X1 U14238 ( .A(n11381), .B(n11383), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11300) );
  INV_X1 U14239 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13616) );
  NAND2_X1 U14240 ( .A1(n11374), .A2(n13616), .ZN(n11299) );
  NAND2_X1 U14241 ( .A1(n11300), .A2(n11299), .ZN(n13505) );
  INV_X1 U14242 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n11301) );
  NAND2_X1 U14243 ( .A1(n11387), .A2(n11301), .ZN(n11306) );
  NAND2_X1 U14244 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11303) );
  NAND2_X1 U14245 ( .A1(n9748), .A2(n11303), .ZN(n11304) );
  OAI21_X1 U14246 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n11302), .A(n11304), .ZN(
        n11305) );
  NAND2_X1 U14247 ( .A1(n11306), .A2(n11305), .ZN(n13578) );
  NAND2_X1 U14248 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11308) );
  OAI211_X1 U14249 ( .C1(n11302), .C2(P1_EBX_REG_5__SCAN_IN), .A(n9748), .B(
        n11308), .ZN(n11309) );
  OAI21_X1 U14250 ( .B1(n11381), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11309), .ZN(
        n13565) );
  INV_X1 U14251 ( .A(n11381), .ZN(n11355) );
  INV_X1 U14252 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20011) );
  NAND2_X1 U14253 ( .A1(n11355), .A2(n20011), .ZN(n11312) );
  NAND2_X1 U14254 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11310) );
  OAI211_X1 U14255 ( .C1(n11302), .C2(P1_EBX_REG_7__SCAN_IN), .A(n9748), .B(
        n11310), .ZN(n11311) );
  AND2_X1 U14256 ( .A1(n11312), .A2(n11311), .ZN(n13784) );
  INV_X1 U14257 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U14258 ( .A1(n11387), .A2(n11313), .ZN(n11317) );
  NAND2_X1 U14259 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11314) );
  NAND2_X1 U14260 ( .A1(n9748), .A2(n11314), .ZN(n11315) );
  OAI21_X1 U14261 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n11302), .A(n11315), .ZN(
        n11316) );
  NAND2_X1 U14262 ( .A1(n11317), .A2(n11316), .ZN(n13783) );
  NAND2_X1 U14263 ( .A1(n13784), .A2(n13783), .ZN(n11318) );
  INV_X1 U14264 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n11319) );
  NAND2_X1 U14265 ( .A1(n11387), .A2(n11319), .ZN(n11323) );
  NAND2_X1 U14266 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11320) );
  NAND2_X1 U14267 ( .A1(n9748), .A2(n11320), .ZN(n11321) );
  OAI21_X1 U14268 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n11302), .A(n11321), .ZN(
        n11322) );
  AND2_X1 U14269 ( .A1(n11323), .A2(n11322), .ZN(n13857) );
  NOR2_X2 U14270 ( .A1(n13858), .A2(n13857), .ZN(n13946) );
  INV_X1 U14271 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14272 ( .A1(n11355), .A2(n11324), .ZN(n11327) );
  NAND2_X1 U14273 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11325) );
  OAI211_X1 U14274 ( .C1(n11302), .C2(P1_EBX_REG_9__SCAN_IN), .A(n9748), .B(
        n11325), .ZN(n11326) );
  INV_X1 U14275 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13959) );
  NAND2_X1 U14276 ( .A1(n11387), .A2(n13959), .ZN(n11330) );
  INV_X1 U14277 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14500) );
  NAND2_X1 U14278 ( .A1(n9748), .A2(n14500), .ZN(n11328) );
  OAI211_X1 U14279 ( .C1(n11302), .C2(P1_EBX_REG_10__SCAN_IN), .A(n11328), .B(
        n11383), .ZN(n11329) );
  NAND2_X1 U14280 ( .A1(n11330), .A2(n11329), .ZN(n13956) );
  MUX2_X1 U14281 ( .A(n11381), .B(n11383), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11331) );
  NAND2_X1 U14282 ( .A1(n11331), .A2(n10261), .ZN(n14271) );
  INV_X1 U14283 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14284 ( .A1(n11387), .A2(n11332), .ZN(n11336) );
  NAND2_X1 U14285 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14286 ( .A1(n9748), .A2(n11333), .ZN(n11334) );
  OAI21_X1 U14287 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(n11302), .A(n11334), .ZN(
        n11335) );
  INV_X1 U14288 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16094) );
  NAND2_X1 U14289 ( .A1(n11374), .A2(n16094), .ZN(n11338) );
  MUX2_X1 U14290 ( .A(n11381), .B(n11383), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11337) );
  INV_X1 U14291 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U14292 ( .A1(n11387), .A2(n11339), .ZN(n11342) );
  INV_X1 U14293 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11508) );
  NAND2_X1 U14294 ( .A1(n9748), .A2(n11508), .ZN(n11340) );
  OAI211_X1 U14295 ( .C1(n11302), .C2(P1_EBX_REG_14__SCAN_IN), .A(n11340), .B(
        n11383), .ZN(n11341) );
  NAND2_X1 U14296 ( .A1(n11342), .A2(n11341), .ZN(n14254) );
  NAND2_X1 U14297 ( .A1(n14256), .A2(n14254), .ZN(n14245) );
  MUX2_X1 U14298 ( .A(n11381), .B(n11383), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11344) );
  INV_X1 U14299 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U14300 ( .A1(n11374), .A2(n16079), .ZN(n11343) );
  NAND2_X1 U14301 ( .A1(n11344), .A2(n11343), .ZN(n14244) );
  INV_X1 U14302 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n20912) );
  NAND2_X1 U14303 ( .A1(n11387), .A2(n20912), .ZN(n11347) );
  INV_X1 U14304 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16072) );
  NAND2_X1 U14305 ( .A1(n9748), .A2(n16072), .ZN(n11345) );
  OAI211_X1 U14306 ( .C1(n11302), .C2(P1_EBX_REG_16__SCAN_IN), .A(n11345), .B(
        n11383), .ZN(n11346) );
  INV_X1 U14307 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14627) );
  NAND2_X1 U14308 ( .A1(n11374), .A2(n14627), .ZN(n11349) );
  MUX2_X1 U14309 ( .A(n11381), .B(n11383), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11348) );
  AND2_X1 U14310 ( .A1(n11349), .A2(n11348), .ZN(n14233) );
  INV_X1 U14311 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15898) );
  NAND2_X1 U14312 ( .A1(n11387), .A2(n15898), .ZN(n11352) );
  INV_X1 U14313 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16059) );
  NAND2_X1 U14314 ( .A1(n9748), .A2(n16059), .ZN(n11350) );
  OAI211_X1 U14315 ( .C1(n11302), .C2(P1_EBX_REG_18__SCAN_IN), .A(n11350), .B(
        n11383), .ZN(n11351) );
  NAND2_X1 U14316 ( .A1(n11352), .A2(n11351), .ZN(n14229) );
  NAND2_X1 U14317 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11353) );
  OAI211_X1 U14318 ( .C1(n11302), .C2(P1_EBX_REG_19__SCAN_IN), .A(n9748), .B(
        n11353), .ZN(n11354) );
  OAI21_X1 U14319 ( .B1(n11381), .B2(P1_EBX_REG_19__SCAN_IN), .A(n11354), .ZN(
        n14221) );
  INV_X1 U14320 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14216) );
  NAND2_X1 U14321 ( .A1(n11355), .A2(n14216), .ZN(n11358) );
  NAND2_X1 U14322 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11356) );
  OAI211_X1 U14323 ( .C1(n11302), .C2(P1_EBX_REG_21__SCAN_IN), .A(n9748), .B(
        n11356), .ZN(n11357) );
  INV_X1 U14324 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n11359) );
  NAND2_X1 U14325 ( .A1(n11387), .A2(n11359), .ZN(n11363) );
  NAND2_X1 U14326 ( .A1(n11383), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11360) );
  NAND2_X1 U14327 ( .A1(n9748), .A2(n11360), .ZN(n11361) );
  OAI21_X1 U14328 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n11302), .A(n11361), .ZN(
        n11362) );
  NAND2_X1 U14329 ( .A1(n11363), .A2(n11362), .ZN(n14210) );
  NAND2_X1 U14330 ( .A1(n14211), .A2(n14210), .ZN(n11364) );
  OR2_X2 U14331 ( .A1(n9774), .A2(n11364), .ZN(n14214) );
  INV_X1 U14332 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15869) );
  NAND2_X1 U14333 ( .A1(n11387), .A2(n15869), .ZN(n11368) );
  INV_X1 U14334 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11365) );
  NAND2_X1 U14335 ( .A1(n9748), .A2(n11365), .ZN(n11366) );
  OAI211_X1 U14336 ( .C1(n11302), .C2(P1_EBX_REG_22__SCAN_IN), .A(n11366), .B(
        n11286), .ZN(n11367) );
  MUX2_X1 U14337 ( .A(n11381), .B(n11286), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11370) );
  NAND2_X1 U14338 ( .A1(n11374), .A2(n14429), .ZN(n11369) );
  AND2_X1 U14339 ( .A1(n11370), .A2(n11369), .ZN(n14132) );
  INV_X1 U14340 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U14341 ( .A1(n11387), .A2(n14199), .ZN(n11373) );
  NAND2_X1 U14342 ( .A1(n9748), .A2(n14530), .ZN(n11371) );
  OAI211_X1 U14343 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n11302), .A(n11371), .B(
        n11286), .ZN(n11372) );
  NAND2_X1 U14344 ( .A1(n11373), .A2(n11372), .ZN(n14123) );
  MUX2_X1 U14345 ( .A(n11381), .B(n11286), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11376) );
  INV_X1 U14346 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16053) );
  NAND2_X1 U14347 ( .A1(n11374), .A2(n16053), .ZN(n11375) );
  INV_X1 U14348 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n11377) );
  NAND2_X1 U14349 ( .A1(n11387), .A2(n11377), .ZN(n11380) );
  INV_X1 U14350 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16042) );
  NAND2_X1 U14351 ( .A1(n9748), .A2(n16042), .ZN(n11378) );
  OAI211_X1 U14352 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n11302), .A(n11378), .B(
        n11286), .ZN(n11379) );
  AND2_X1 U14353 ( .A1(n11380), .A2(n11379), .ZN(n14101) );
  MUX2_X1 U14354 ( .A(n11381), .B(n11286), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11382) );
  OAI21_X1 U14355 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13501), .A(
        n11382), .ZN(n14087) );
  INV_X1 U14356 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14195) );
  NAND2_X1 U14357 ( .A1(n11387), .A2(n14195), .ZN(n11386) );
  INV_X1 U14358 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14381) );
  NAND2_X1 U14359 ( .A1(n9748), .A2(n14381), .ZN(n11384) );
  OAI211_X1 U14360 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n11302), .A(n11384), .B(
        n11383), .ZN(n11385) );
  NAND2_X1 U14361 ( .A1(n11386), .A2(n11385), .ZN(n14066) );
  OAI22_X1 U14362 ( .A1(n13501), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n11302), .ZN(n14036) );
  OR2_X1 U14363 ( .A1(n14036), .A2(n14035), .ZN(n11389) );
  INV_X1 U14364 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14194) );
  NAND2_X1 U14365 ( .A1(n11387), .A2(n14194), .ZN(n11388) );
  NAND2_X1 U14366 ( .A1(n11389), .A2(n11388), .ZN(n14053) );
  NAND2_X1 U14367 ( .A1(n14068), .A2(n14053), .ZN(n14055) );
  MUX2_X1 U14368 ( .A(n14040), .B(n11286), .S(n14055), .Z(n11391) );
  AOI22_X1 U14369 ( .A1(n13501), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11302), .ZN(n11390) );
  NOR2_X1 U14370 ( .A1(n13742), .A2(n20162), .ZN(n11412) );
  NAND2_X1 U14371 ( .A1(n13626), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n11408) );
  AND2_X1 U14372 ( .A1(n20848), .A2(n20814), .ZN(n11395) );
  NOR2_X1 U14373 ( .A1(n11408), .A2(n11395), .ZN(n11392) );
  AND2_X1 U14374 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n11403) );
  INV_X1 U14375 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20762) );
  NAND2_X1 U14376 ( .A1(n19972), .A2(n20762), .ZN(n20749) );
  INV_X1 U14377 ( .A(n20749), .ZN(n11393) );
  NOR2_X1 U14378 ( .A1(n11393), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20757) );
  NAND2_X1 U14379 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n11394) );
  NAND2_X1 U14380 ( .A1(n20757), .A2(n11394), .ZN(n15842) );
  INV_X1 U14381 ( .A(n11395), .ZN(n11396) );
  AOI21_X1 U14382 ( .B1(n20177), .B2(n15842), .A(n11396), .ZN(n11410) );
  NAND2_X1 U14383 ( .A1(n20021), .A2(n14158), .ZN(n15951) );
  INV_X1 U14384 ( .A(n15951), .ZN(n13778) );
  INV_X1 U14385 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15896) );
  INV_X1 U14386 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n16063) );
  INV_X1 U14387 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20775) );
  INV_X1 U14388 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20773) );
  NAND4_X1 U14389 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20018)
         );
  NAND3_X1 U14390 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n13860) );
  NOR3_X1 U14391 ( .A1(n20773), .A2(n20018), .A3(n13860), .ZN(n20000) );
  NAND2_X1 U14392 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20000), .ZN(n15961) );
  NOR2_X1 U14393 ( .A1(n20775), .A2(n15961), .ZN(n14160) );
  INV_X1 U14394 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20785) );
  NAND4_X1 U14395 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n15919) );
  NAND2_X1 U14396 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15917) );
  NOR3_X1 U14397 ( .A1(n20785), .A2(n15919), .A3(n15917), .ZN(n15885) );
  NAND2_X1 U14398 ( .A1(n14160), .A2(n15885), .ZN(n15884) );
  NOR3_X1 U14399 ( .A1(n15896), .A2(n16063), .A3(n15884), .ZN(n14148) );
  AND4_X1 U14400 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .A4(P1_REIP_REG_21__SCAN_IN), .ZN(n11397) );
  NAND3_X1 U14401 ( .A1(n14158), .A2(n14148), .A3(n11397), .ZN(n11398) );
  NAND2_X1 U14402 ( .A1(n15951), .A2(n11398), .ZN(n14137) );
  AND2_X1 U14403 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n11406) );
  INV_X1 U14404 ( .A(n11406), .ZN(n14106) );
  INV_X1 U14405 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n16045) );
  NOR2_X1 U14406 ( .A1(n14106), .A2(n16045), .ZN(n11399) );
  OR2_X1 U14407 ( .A1(n20021), .A2(n11399), .ZN(n11400) );
  NAND2_X1 U14408 ( .A1(n14137), .A2(n11400), .ZN(n14094) );
  AND2_X1 U14409 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n11401) );
  NOR2_X1 U14410 ( .A1(n20021), .A2(n11401), .ZN(n11402) );
  NOR2_X1 U14411 ( .A1(n14094), .A2(n11402), .ZN(n14075) );
  OAI21_X1 U14412 ( .B1(n11403), .B2(n13778), .A(n14075), .ZN(n14046) );
  INV_X1 U14413 ( .A(n14148), .ZN(n11405) );
  NAND3_X1 U14414 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_21__SCAN_IN), .ZN(n11404) );
  INV_X1 U14415 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14432) );
  NOR2_X1 U14416 ( .A1(n14138), .A2(n14432), .ZN(n14119) );
  NAND2_X1 U14417 ( .A1(n14119), .A2(n11406), .ZN(n14096) );
  INV_X1 U14418 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21109) );
  INV_X1 U14419 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14383) );
  NOR2_X1 U14420 ( .A1(n14074), .A2(n14383), .ZN(n14063) );
  INV_X1 U14421 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n11407) );
  NAND4_X1 U14422 ( .A1(n14063), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .A4(n11407), .ZN(n11414) );
  INV_X1 U14423 ( .A(n11408), .ZN(n11409) );
  NOR2_X1 U14424 ( .A1(n11410), .A2(n11409), .ZN(n11411) );
  AOI22_X1 U14425 ( .A1(n20046), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20059), .ZN(n11413) );
  NAND2_X1 U14426 ( .A1(n11414), .A2(n11413), .ZN(n11415) );
  AOI21_X1 U14427 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(n14046), .A(n11415), 
        .ZN(n11416) );
  OAI21_X1 U14428 ( .B1(n14525), .B2(n20062), .A(n11416), .ZN(n11417) );
  NAND2_X1 U14429 ( .A1(n11419), .A2(n11418), .ZN(P1_U2809) );
  NAND3_X1 U14430 ( .A1(n9880), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16172) );
  INV_X1 U14431 ( .A(n16172), .ZN(n11420) );
  NAND2_X1 U14432 ( .A1(n14465), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14370) );
  INV_X1 U14433 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14540) );
  NOR2_X1 U14434 ( .A1(n14371), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11518) );
  NAND2_X1 U14435 ( .A1(n20162), .A2(n11424), .ZN(n11441) );
  OAI21_X1 U14436 ( .B1(n11438), .B2(n20851), .A(n11441), .ZN(n11425) );
  INV_X1 U14437 ( .A(n11425), .ZN(n11426) );
  XNOR2_X1 U14438 ( .A(n11428), .B(n11437), .ZN(n11430) );
  AOI21_X1 U14439 ( .B1(n11430), .B2(n13138), .A(n11429), .ZN(n11431) );
  INV_X1 U14440 ( .A(n11432), .ZN(n20129) );
  NAND2_X1 U14441 ( .A1(n20129), .A2(n11433), .ZN(n11434) );
  NAND2_X1 U14442 ( .A1(n11435), .A2(n11434), .ZN(n11446) );
  XNOR2_X1 U14443 ( .A(n11446), .B(n13493), .ZN(n13485) );
  NAND2_X1 U14444 ( .A1(n11436), .A2(n9918), .ZN(n11445) );
  NAND2_X1 U14445 ( .A1(n11438), .A2(n11437), .ZN(n11439) );
  NAND2_X1 U14446 ( .A1(n11439), .A2(n11440), .ZN(n11458) );
  OAI21_X1 U14447 ( .B1(n11440), .B2(n11439), .A(n11458), .ZN(n11443) );
  INV_X1 U14448 ( .A(n11441), .ZN(n11442) );
  AOI21_X1 U14449 ( .B1(n11443), .B2(n13138), .A(n11442), .ZN(n11444) );
  NAND2_X1 U14450 ( .A1(n11446), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11447) );
  NAND2_X1 U14451 ( .A1(n11448), .A2(n11447), .ZN(n11453) );
  XNOR2_X1 U14452 ( .A(n11453), .B(n13616), .ZN(n13518) );
  OR2_X1 U14453 ( .A1(n20812), .A2(n11469), .ZN(n11452) );
  INV_X1 U14454 ( .A(n11457), .ZN(n11449) );
  XNOR2_X1 U14455 ( .A(n11458), .B(n11449), .ZN(n11450) );
  NAND2_X1 U14456 ( .A1(n11450), .A2(n13138), .ZN(n11451) );
  NAND2_X1 U14457 ( .A1(n11452), .A2(n11451), .ZN(n13517) );
  NAND2_X1 U14458 ( .A1(n13518), .A2(n13517), .ZN(n11455) );
  NAND2_X1 U14459 ( .A1(n11453), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11454) );
  NAND2_X1 U14460 ( .A1(n11455), .A2(n11454), .ZN(n13574) );
  NAND2_X1 U14461 ( .A1(n11456), .A2(n9918), .ZN(n11464) );
  NAND2_X1 U14462 ( .A1(n11458), .A2(n11457), .ZN(n11460) );
  INV_X1 U14463 ( .A(n11460), .ZN(n11462) );
  INV_X1 U14464 ( .A(n11461), .ZN(n11459) );
  OR2_X1 U14465 ( .A1(n11460), .A2(n11459), .ZN(n11481) );
  OAI211_X1 U14466 ( .C1(n11462), .C2(n11461), .A(n13138), .B(n11481), .ZN(
        n11463) );
  NAND2_X1 U14467 ( .A1(n11464), .A2(n11463), .ZN(n11466) );
  INV_X1 U14468 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11465) );
  XNOR2_X1 U14469 ( .A(n11466), .B(n11465), .ZN(n13573) );
  NAND2_X1 U14470 ( .A1(n13574), .A2(n13573), .ZN(n11468) );
  NAND2_X1 U14471 ( .A1(n11466), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11467) );
  NAND2_X1 U14472 ( .A1(n11468), .A2(n11467), .ZN(n16031) );
  OR2_X1 U14473 ( .A1(n11470), .A2(n11469), .ZN(n11473) );
  XNOR2_X1 U14474 ( .A(n11481), .B(n11479), .ZN(n11471) );
  NAND2_X1 U14475 ( .A1(n11471), .A2(n13138), .ZN(n11472) );
  NAND2_X1 U14476 ( .A1(n11473), .A2(n11472), .ZN(n11475) );
  INV_X1 U14477 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11474) );
  XNOR2_X1 U14478 ( .A(n11475), .B(n11474), .ZN(n16030) );
  NAND2_X1 U14479 ( .A1(n11475), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11476) );
  NAND3_X1 U14480 ( .A1(n11478), .A2(n11477), .A3(n9918), .ZN(n11484) );
  INV_X1 U14481 ( .A(n11479), .ZN(n11480) );
  OR2_X1 U14482 ( .A1(n11481), .A2(n11480), .ZN(n11487) );
  XNOR2_X1 U14483 ( .A(n11487), .B(n11488), .ZN(n11482) );
  NAND2_X1 U14484 ( .A1(n11482), .A2(n13138), .ZN(n11483) );
  NAND2_X1 U14485 ( .A1(n11484), .A2(n11483), .ZN(n11485) );
  OR2_X1 U14486 ( .A1(n11485), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16024) );
  NAND2_X1 U14487 ( .A1(n11485), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16023) );
  NAND2_X1 U14488 ( .A1(n11486), .A2(n9918), .ZN(n11493) );
  INV_X1 U14489 ( .A(n11487), .ZN(n11489) );
  NAND2_X1 U14490 ( .A1(n11489), .A2(n11488), .ZN(n11497) );
  XNOR2_X1 U14491 ( .A(n11497), .B(n11490), .ZN(n11491) );
  NAND2_X1 U14492 ( .A1(n11491), .A2(n13138), .ZN(n11492) );
  NAND2_X1 U14493 ( .A1(n11493), .A2(n11492), .ZN(n16018) );
  OR2_X1 U14494 ( .A1(n16018), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11494) );
  NAND2_X1 U14495 ( .A1(n16018), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11495) );
  OR3_X1 U14496 ( .A1(n11497), .A2(n11496), .A3(n20851), .ZN(n11498) );
  NAND2_X1 U14497 ( .A1(n14465), .A2(n11498), .ZN(n13909) );
  OR2_X1 U14498 ( .A1(n13909), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U14499 ( .A1(n11500), .A2(n11499), .ZN(n13963) );
  INV_X1 U14500 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16126) );
  OR2_X1 U14501 ( .A1(n16009), .A2(n16126), .ZN(n11501) );
  NAND2_X1 U14502 ( .A1(n14465), .A2(n16126), .ZN(n11502) );
  INV_X1 U14503 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14644) );
  NAND2_X1 U14504 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14505 ( .A1(n14465), .A2(n11508), .ZN(n11504) );
  NAND2_X1 U14506 ( .A1(n15994), .A2(n11504), .ZN(n14473) );
  NOR2_X1 U14507 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11505) );
  OR2_X1 U14508 ( .A1(n16009), .A2(n11505), .ZN(n11506) );
  AND2_X1 U14509 ( .A1(n14471), .A2(n11506), .ZN(n14463) );
  XNOR2_X1 U14510 ( .A(n16009), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15988) );
  NAND2_X1 U14511 ( .A1(n14465), .A2(n16079), .ZN(n15985) );
  NAND2_X1 U14512 ( .A1(n15988), .A2(n15985), .ZN(n11507) );
  NOR2_X1 U14513 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14460) );
  AND4_X1 U14514 ( .A1(n14460), .A2(n11508), .A3(n16094), .A4(n14644), .ZN(
        n11509) );
  NAND2_X1 U14515 ( .A1(n14471), .A2(n14472), .ZN(n15986) );
  NOR2_X1 U14516 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11510) );
  NOR2_X1 U14517 ( .A1(n14465), .A2(n11510), .ZN(n11511) );
  NOR2_X1 U14518 ( .A1(n15986), .A2(n11511), .ZN(n11512) );
  XNOR2_X1 U14519 ( .A(n16009), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14455) );
  NAND3_X1 U14520 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14527) );
  INV_X1 U14521 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11514) );
  INV_X1 U14522 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20932) );
  NAND2_X1 U14523 ( .A1(n11514), .A2(n20932), .ZN(n11515) );
  NAND2_X1 U14524 ( .A1(n11516), .A2(n14501), .ZN(n14595) );
  INV_X1 U14525 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14429) );
  NAND3_X1 U14526 ( .A1(n14530), .A2(n14429), .A3(n16053), .ZN(n14377) );
  NOR2_X1 U14527 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14557) );
  NAND3_X1 U14528 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14515) );
  AND2_X1 U14529 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14556) );
  AOI21_X1 U14530 ( .B1(n20162), .B2(n10437), .A(n14015), .ZN(n11519) );
  NAND2_X1 U14531 ( .A1(n20829), .A2(n11520), .ZN(n20847) );
  AND2_X1 U14532 ( .A1(n20847), .A2(n9880), .ZN(n11521) );
  NAND2_X1 U14533 ( .A1(n9880), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15813) );
  NAND2_X1 U14534 ( .A1(n20814), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11522) );
  NAND2_X1 U14535 ( .A1(n15813), .A2(n11522), .ZN(n20131) );
  NAND2_X1 U14536 ( .A1(n20135), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14523) );
  NAND2_X1 U14537 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11523) );
  OAI211_X1 U14538 ( .C1(n16029), .C2(n13744), .A(n14523), .B(n11523), .ZN(
        n11524) );
  MUX2_X1 U14539 ( .A(n19949), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12180) );
  NAND2_X1 U14540 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19958), .ZN(
        n12142) );
  INV_X1 U14541 ( .A(n12142), .ZN(n11525) );
  NAND2_X1 U14542 ( .A1(n12180), .A2(n11525), .ZN(n11527) );
  NAND2_X1 U14543 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19949), .ZN(
        n11526) );
  NAND2_X1 U14544 ( .A1(n11527), .A2(n11526), .ZN(n11606) );
  NAND2_X1 U14545 ( .A1(n16435), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U14546 ( .A1(n11606), .A2(n11605), .ZN(n11604) );
  NAND2_X1 U14547 ( .A1(n11604), .A2(n11529), .ZN(n11608) );
  AND2_X2 U14548 ( .A1(n11530), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11540) );
  AND2_X4 U14549 ( .A1(n11540), .A2(n16435), .ZN(n11723) );
  AOI22_X1 U14550 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11536) );
  AND2_X4 U14551 ( .A1(n12900), .A2(n11537), .ZN(n12730) );
  AND2_X2 U14552 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11544) );
  AND2_X4 U14553 ( .A1(n11544), .A2(n11532), .ZN(n11720) );
  INV_X1 U14554 ( .A(n11720), .ZN(n12897) );
  AND2_X2 U14555 ( .A1(n11531), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11899) );
  AOI22_X1 U14556 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11535) );
  AND2_X2 U14557 ( .A1(n11718), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12413) );
  AND2_X2 U14558 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14559 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11534) );
  AND2_X2 U14560 ( .A1(n12870), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11634) );
  AND2_X4 U14561 ( .A1(n11544), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11719) );
  AND2_X2 U14562 ( .A1(n13871), .A2(n11537), .ZN(n11898) );
  AOI22_X1 U14563 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11533) );
  NAND4_X1 U14564 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11550) );
  AND2_X2 U14565 ( .A1(n12902), .A2(n11537), .ZN(n11633) );
  AOI22_X1 U14566 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11548) );
  INV_X1 U14567 ( .A(n11722), .ZN(n12894) );
  AND2_X2 U14568 ( .A1(n11722), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12736) );
  AND2_X1 U14569 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14570 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11547) );
  AND2_X2 U14571 ( .A1(n11540), .A2(n12710), .ZN(n12737) );
  NOR2_X1 U14572 ( .A1(n14010), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11541) );
  AOI22_X1 U14573 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11904), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14574 ( .A1(n11586), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11545) );
  NAND4_X1 U14575 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11549) );
  AOI22_X1 U14576 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14577 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14578 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14579 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11552) );
  NAND4_X1 U14580 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11561) );
  AOI22_X1 U14581 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14582 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14583 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14584 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11556) );
  NAND4_X1 U14585 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n11560) );
  MUX2_X2 U14586 ( .A(n11561), .B(n11560), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12283) );
  AOI22_X1 U14587 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14588 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11564) );
  INV_X2 U14589 ( .A(n12829), .ZN(n12903) );
  AOI22_X1 U14590 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14591 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9750), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11562) );
  NAND4_X1 U14592 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11571) );
  AOI22_X1 U14593 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14594 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14595 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14596 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11566) );
  NAND4_X1 U14597 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11570) );
  MUX2_X2 U14598 ( .A(n11571), .B(n11570), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12973) );
  MUX2_X1 U14599 ( .A(n12140), .B(n12318), .S(n11774), .Z(n11580) );
  AOI22_X1 U14600 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12903), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14601 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14602 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14603 ( .A1(n11720), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14604 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11672), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14605 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14606 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14607 ( .A1(n12902), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11576) );
  MUX2_X1 U14608 ( .A(n11580), .B(P2_EBX_REG_4__SCAN_IN), .S(n19302), .Z(
        n11966) );
  AOI22_X1 U14609 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14610 ( .A1(n11899), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12735), .ZN(n11583) );
  AOI22_X1 U14611 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12736), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14612 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11634), .B1(
        n12413), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11581) );
  NAND4_X1 U14613 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11592) );
  AOI22_X1 U14614 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11904), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14615 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12737), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14616 ( .A1(n12383), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14617 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11587) );
  NAND4_X1 U14618 ( .A1(n11590), .A2(n11589), .A3(n11588), .A4(n11587), .ZN(
        n11591) );
  NOR2_X1 U14619 ( .A1(n11592), .A2(n11591), .ZN(n12298) );
  INV_X1 U14620 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13764) );
  INV_X1 U14621 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13085) );
  NAND2_X1 U14622 ( .A1(n13764), .A2(n13085), .ZN(n11593) );
  MUX2_X1 U14623 ( .A(n12298), .B(n11593), .S(n11765), .Z(n11957) );
  AOI22_X1 U14624 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n11896), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14625 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12730), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14626 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11633), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14627 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11594) );
  NAND4_X1 U14628 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11603) );
  AOI22_X1 U14629 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14630 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14631 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14632 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12737), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11598) );
  NAND4_X1 U14633 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11602) );
  OAI21_X1 U14634 ( .B1(n11606), .B2(n11605), .A(n11604), .ZN(n12186) );
  INV_X1 U14635 ( .A(n12186), .ZN(n12179) );
  AND2_X1 U14636 ( .A1(n12587), .A2(n12179), .ZN(n12189) );
  INV_X4 U14637 ( .A(n11765), .ZN(n12130) );
  NOR2_X1 U14638 ( .A1(n11608), .A2(n11607), .ZN(n11609) );
  INV_X1 U14639 ( .A(n12139), .ZN(n11621) );
  AOI22_X1 U14640 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14641 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14642 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14643 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11611) );
  NAND4_X1 U14644 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        n11620) );
  AOI22_X1 U14645 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14646 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14647 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14648 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11615) );
  NAND4_X1 U14649 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11619) );
  MUX2_X1 U14650 ( .A(n11621), .B(n11869), .S(n11774), .Z(n11622) );
  INV_X1 U14651 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13651) );
  MUX2_X1 U14652 ( .A(n11622), .B(n13651), .S(n19302), .Z(n11952) );
  NAND2_X1 U14653 ( .A1(n11953), .A2(n11952), .ZN(n11964) );
  INV_X1 U14654 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U14655 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14656 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14657 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14658 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14659 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11632) );
  AOI22_X1 U14660 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14661 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14662 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14663 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11627) );
  NAND4_X1 U14664 ( .A1(n11630), .A2(n11629), .A3(n11628), .A4(n11627), .ZN(
        n11631) );
  MUX2_X1 U14665 ( .A(n13213), .B(n11942), .S(n12130), .Z(n11946) );
  AOI22_X1 U14666 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12730), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14667 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14668 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14669 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11635) );
  NAND4_X1 U14670 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11644) );
  AOI22_X1 U14671 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14672 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12735), .ZN(n11641) );
  AOI22_X1 U14673 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12737), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14674 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11904), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11639) );
  NAND4_X1 U14675 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11643) );
  MUX2_X1 U14676 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12326), .S(n12130), .Z(
        n12003) );
  NAND2_X1 U14677 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11648) );
  NAND2_X1 U14678 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11647) );
  NAND2_X1 U14679 ( .A1(n12383), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11646) );
  NAND2_X1 U14680 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11645) );
  AOI22_X1 U14681 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12735), .ZN(n11651) );
  AOI22_X1 U14682 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12737), .B1(
        n11904), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14683 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11586), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14684 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11657) );
  NAND2_X1 U14685 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11655) );
  NAND2_X1 U14686 ( .A1(n11899), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11654) );
  NAND2_X1 U14687 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11653) );
  NAND2_X1 U14688 ( .A1(n11898), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11652) );
  INV_X1 U14689 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13514) );
  INV_X1 U14690 ( .A(n12331), .ZN(n12134) );
  INV_X1 U14691 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U14692 ( .A1(n19302), .A2(n13314), .ZN(n11660) );
  NAND2_X1 U14693 ( .A1(n12134), .A2(n11660), .ZN(n12013) );
  NAND2_X1 U14694 ( .A1(n19302), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12010) );
  NAND2_X1 U14695 ( .A1(n12114), .A2(n11661), .ZN(n12033) );
  NAND2_X1 U14696 ( .A1(n19302), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12039) );
  INV_X1 U14697 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12526) );
  NOR2_X1 U14698 ( .A1(n12130), .A2(n12526), .ZN(n12043) );
  INV_X1 U14699 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n20874) );
  NOR2_X1 U14700 ( .A1(n12130), .A2(n20874), .ZN(n12059) );
  NAND2_X1 U14701 ( .A1(n19302), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12056) );
  INV_X1 U14702 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11662) );
  NOR2_X1 U14703 ( .A1(n12130), .A2(n11662), .ZN(n12052) );
  OR2_X2 U14704 ( .A1(n12058), .A2(n12052), .ZN(n12051) );
  INV_X1 U14705 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12532) );
  NOR2_X1 U14706 ( .A1(n12130), .A2(n12532), .ZN(n12049) );
  NOR2_X1 U14707 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n11663) );
  NOR2_X1 U14708 ( .A1(n12130), .A2(n11663), .ZN(n11664) );
  INV_X1 U14709 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12544) );
  INV_X1 U14710 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12548) );
  NAND2_X1 U14711 ( .A1(n19302), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11665) );
  INV_X1 U14712 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11666) );
  NOR2_X1 U14713 ( .A1(n12130), .A2(n11666), .ZN(n12096) );
  XNOR2_X1 U14714 ( .A(n12097), .B(n12096), .ZN(n16253) );
  NOR2_X1 U14715 ( .A1(n16253), .A2(n10051), .ZN(n12095) );
  INV_X1 U14716 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14717 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14718 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14719 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n11722), .ZN(n11668) );
  AOI22_X1 U14720 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11667) );
  NAND4_X1 U14721 ( .A1(n11670), .A2(n11669), .A3(n11668), .A4(n11667), .ZN(
        n11671) );
  NAND2_X1 U14722 ( .A1(n11671), .A2(n11537), .ZN(n11679) );
  AOI22_X1 U14723 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14724 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14725 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14726 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11673) );
  NAND4_X1 U14727 ( .A1(n11676), .A2(n11675), .A3(n11674), .A4(n11673), .ZN(
        n11677) );
  AOI22_X1 U14728 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14729 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14730 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14731 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11680) );
  NAND2_X1 U14732 ( .A1(n11684), .A2(n11537), .ZN(n11690) );
  AOI22_X1 U14733 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14734 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14735 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14736 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11687) );
  NAND2_X1 U14737 ( .A1(n11690), .A2(n11689), .ZN(n11744) );
  AOI22_X1 U14738 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14739 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14740 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14741 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11691) );
  NAND4_X1 U14742 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11695) );
  NAND2_X1 U14743 ( .A1(n11695), .A2(n11537), .ZN(n11702) );
  AOI22_X1 U14744 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14745 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14746 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14747 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11696) );
  NAND4_X1 U14748 ( .A1(n11699), .A2(n11698), .A3(n11697), .A4(n11696), .ZN(
        n11700) );
  NAND2_X1 U14749 ( .A1(n11700), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11701) );
  NAND2_X1 U14750 ( .A1(n11702), .A2(n11701), .ZN(n11732) );
  AOI22_X1 U14751 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14752 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14753 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14754 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14755 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14756 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14757 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14758 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9750), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11708) );
  MUX2_X2 U14759 ( .A(n11713), .B(n11712), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19290) );
  AOI22_X1 U14760 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14761 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14762 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14763 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11714) );
  NAND4_X1 U14764 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11729) );
  AOI22_X1 U14765 ( .A1(n11551), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14766 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11719), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14767 ( .A1(n11721), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14768 ( .A1(n11723), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11722), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11724) );
  NAND4_X1 U14769 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n11728) );
  NAND2_X1 U14770 ( .A1(n11735), .A2(n11757), .ZN(n12159) );
  BUF_X4 U14771 ( .A(n12283), .Z(n15585) );
  NAND3_X1 U14772 ( .A1(n12159), .A2(n19290), .A3(n15585), .ZN(n11731) );
  NOR2_X1 U14773 ( .A1(n12169), .A2(n12928), .ZN(n11730) );
  NAND2_X1 U14774 ( .A1(n11731), .A2(n12175), .ZN(n12465) );
  MUX2_X1 U14775 ( .A(n12928), .B(n12929), .S(n12169), .Z(n11734) );
  NAND2_X1 U14776 ( .A1(n11742), .A2(n12255), .ZN(n11768) );
  AOI21_X1 U14777 ( .B1(n12928), .B2(n11743), .A(n12247), .ZN(n11733) );
  NAND3_X1 U14778 ( .A1(n11734), .A2(n11768), .A3(n11733), .ZN(n11737) );
  AND2_X1 U14779 ( .A1(n11751), .A2(n12247), .ZN(n11736) );
  NAND2_X1 U14780 ( .A1(n11735), .A2(n11736), .ZN(n12164) );
  NAND3_X1 U14781 ( .A1(n11737), .A2(n12164), .A3(n11750), .ZN(n12251) );
  NOR2_X1 U14782 ( .A1(n11743), .A2(n12929), .ZN(n11738) );
  NAND2_X1 U14783 ( .A1(n11739), .A2(n11738), .ZN(n11746) );
  AND3_X1 U14784 ( .A1(n11776), .A2(n11742), .A3(n11746), .ZN(n12243) );
  INV_X1 U14785 ( .A(n12243), .ZN(n11740) );
  NAND2_X1 U14786 ( .A1(n12166), .A2(n19297), .ZN(n12170) );
  NAND2_X1 U14787 ( .A1(n11745), .A2(n12170), .ZN(n12252) );
  NAND2_X1 U14788 ( .A1(n12252), .A2(n12255), .ZN(n11748) );
  NAND2_X1 U14789 ( .A1(n11748), .A2(n11747), .ZN(n11785) );
  OAI21_X2 U14790 ( .B1(n11784), .B2(n11749), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11801) );
  AND2_X2 U14791 ( .A1(n11751), .A2(n19290), .ZN(n11773) );
  NAND2_X1 U14792 ( .A1(n11754), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11760) );
  NOR2_X1 U14793 ( .A1(n12255), .A2(n21158), .ZN(n11755) );
  NAND4_X1 U14794 ( .A1(n11735), .A2(n11750), .A3(n11755), .A4(n12247), .ZN(
        n11759) );
  AND2_X1 U14795 ( .A1(n19297), .A2(n12973), .ZN(n11756) );
  NOR2_X1 U14796 ( .A1(n12928), .A2(n21158), .ZN(n12605) );
  NAND4_X1 U14797 ( .A1(n11754), .A2(n11757), .A3(n11756), .A4(n12605), .ZN(
        n11758) );
  NAND2_X1 U14798 ( .A1(n21158), .A2(n16467), .ZN(n14679) );
  NOR2_X1 U14799 ( .A1(n14679), .A2(n19949), .ZN(n11761) );
  NOR2_X1 U14800 ( .A1(n11771), .A2(n11761), .ZN(n11762) );
  OAI21_X2 U14801 ( .B1(n11801), .B2(n14010), .A(n11762), .ZN(n11798) );
  NAND3_X1 U14802 ( .A1(n11765), .A2(n11776), .A3(n19307), .ZN(n11766) );
  NAND2_X1 U14803 ( .A1(n11766), .A2(n11751), .ZN(n11767) );
  NAND2_X1 U14804 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  INV_X1 U14805 ( .A(n11746), .ZN(n11775) );
  NAND2_X1 U14806 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U14807 ( .A1(n12973), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12196) );
  NOR2_X1 U14808 ( .A1(n12196), .A2(n11776), .ZN(n11777) );
  NAND2_X1 U14809 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11780) );
  AND2_X1 U14810 ( .A1(n14679), .A2(n11780), .ZN(n11782) );
  AOI21_X1 U14811 ( .B1(n11803), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11783), .ZN(n11788) );
  AND2_X1 U14812 ( .A1(n11785), .A2(n11740), .ZN(n11786) );
  OAI21_X1 U14813 ( .B1(n11784), .B2(n11786), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11787) );
  NAND2_X1 U14814 ( .A1(n11788), .A2(n11787), .ZN(n11822) );
  NAND2_X1 U14815 ( .A1(n11825), .A2(n11821), .ZN(n11800) );
  INV_X1 U14816 ( .A(n11796), .ZN(n11797) );
  NAND2_X1 U14817 ( .A1(n11800), .A2(n11799), .ZN(n11816) );
  AOI21_X1 U14818 ( .B1(n21158), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U14819 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11806) );
  OAI211_X1 U14820 ( .C1(n11804), .C2(n10206), .A(n11806), .B(n11805), .ZN(
        n11807) );
  INV_X1 U14821 ( .A(n11817), .ZN(n11808) );
  NAND2_X1 U14822 ( .A1(n11818), .A2(n11808), .ZN(n11809) );
  NAND2_X1 U14823 ( .A1(n11816), .A2(n11809), .ZN(n11812) );
  INV_X1 U14824 ( .A(n11818), .ZN(n11810) );
  NAND2_X2 U14825 ( .A1(n11812), .A2(n11811), .ZN(n12497) );
  OAI22_X1 U14826 ( .A1(n11801), .A2(n11537), .B1(n14679), .B2(n19933), .ZN(
        n12500) );
  NAND2_X1 U14827 ( .A1(n12574), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11814) );
  NAND2_X1 U14828 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11813) );
  OAI211_X1 U14829 ( .C1(n11804), .C2(n13651), .A(n11814), .B(n11813), .ZN(
        n11815) );
  XNOR2_X1 U14830 ( .A(n11818), .B(n11817), .ZN(n11819) );
  INV_X1 U14831 ( .A(n11845), .ZN(n11820) );
  INV_X1 U14832 ( .A(n13607), .ZN(n19118) );
  AND2_X1 U14833 ( .A1(n19118), .A2(n11830), .ZN(n11855) );
  INV_X1 U14834 ( .A(n11855), .ZN(n11827) );
  INV_X1 U14835 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11828) );
  OAI22_X1 U14836 ( .A1(n11829), .A2(n19502), .B1(n19384), .B2(n11828), .ZN(
        n11834) );
  INV_X1 U14837 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11832) );
  OR2_X1 U14838 ( .A1(n11830), .A2(n13607), .ZN(n11853) );
  XNOR2_X2 U14839 ( .A(n11830), .B(n11821), .ZN(n14005) );
  OR2_X1 U14840 ( .A1(n14005), .A2(n19118), .ZN(n11841) );
  INV_X1 U14841 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11831) );
  OAI22_X1 U14842 ( .A1(n11832), .A2(n19325), .B1(n19416), .B2(n11831), .ZN(
        n11833) );
  NOR2_X1 U14843 ( .A1(n11834), .A2(n11833), .ZN(n11868) );
  INV_X1 U14844 ( .A(n14005), .ZN(n13098) );
  INV_X1 U14845 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11835) );
  NOR2_X1 U14846 ( .A1(n19733), .A2(n11835), .ZN(n11840) );
  INV_X1 U14847 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11838) );
  NAND2_X1 U14848 ( .A1(n14005), .A2(n13607), .ZN(n11842) );
  INV_X1 U14849 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11837) );
  OAI22_X1 U14850 ( .A1(n11838), .A2(n19444), .B1(n19475), .B2(n11837), .ZN(
        n11839) );
  NOR2_X1 U14851 ( .A1(n11840), .A2(n11839), .ZN(n11867) );
  INV_X1 U14852 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11844) );
  INV_X1 U14853 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12796) );
  OAI22_X1 U14854 ( .A1(n11844), .A2(n19275), .B1(n19350), .B2(n12796), .ZN(
        n11851) );
  INV_X1 U14855 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11849) );
  INV_X1 U14856 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12804) );
  OAI22_X1 U14857 ( .A1(n11849), .A2(n11934), .B1(n19602), .B2(n12804), .ZN(
        n11850) );
  NOR2_X1 U14858 ( .A1(n11851), .A2(n11850), .ZN(n11866) );
  INV_X1 U14859 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11852) );
  NOR2_X1 U14860 ( .A1(n11917), .A2(n11852), .ZN(n11864) );
  INV_X1 U14861 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11857) );
  INV_X1 U14862 ( .A(n11853), .ZN(n11854) );
  OR2_X2 U14863 ( .A1(n11859), .A2(n13176), .ZN(n19633) );
  INV_X1 U14864 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11856) );
  OAI22_X1 U14865 ( .A1(n11857), .A2(n11921), .B1(n19633), .B2(n11856), .ZN(
        n11863) );
  INV_X1 U14866 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11861) );
  OR2_X2 U14867 ( .A1(n11858), .A2(n11820), .ZN(n19689) );
  OR2_X2 U14868 ( .A1(n11859), .A2(n11820), .ZN(n19770) );
  INV_X1 U14869 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11860) );
  OAI22_X1 U14870 ( .A1(n11861), .A2(n19689), .B1(n19770), .B2(n11860), .ZN(
        n11862) );
  NOR3_X1 U14871 ( .A1(n11864), .A2(n11863), .A3(n11862), .ZN(n11865) );
  INV_X1 U14872 ( .A(n11869), .ZN(n12315) );
  NAND2_X1 U14873 ( .A1(n12315), .A2(n11776), .ZN(n11870) );
  INV_X1 U14874 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11872) );
  INV_X1 U14875 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11871) );
  OAI22_X1 U14876 ( .A1(n11872), .A2(n19325), .B1(n19384), .B2(n11871), .ZN(
        n11876) );
  INV_X1 U14877 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11874) );
  INV_X1 U14878 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11873) );
  OAI22_X1 U14879 ( .A1(n11874), .A2(n19416), .B1(n19475), .B2(n11873), .ZN(
        n11875) );
  NOR2_X1 U14880 ( .A1(n11876), .A2(n11875), .ZN(n11895) );
  INV_X1 U14881 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11879) );
  INV_X1 U14882 ( .A(n11921), .ZN(n11877) );
  OAI211_X1 U14883 ( .C1(n19444), .C2(n11879), .A(n11878), .B(n15585), .ZN(
        n11886) );
  INV_X1 U14884 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11881) );
  INV_X1 U14885 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11880) );
  OAI22_X1 U14886 ( .A1(n11881), .A2(n19689), .B1(n19633), .B2(n11880), .ZN(
        n11885) );
  INV_X1 U14887 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11883) );
  INV_X1 U14888 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11882) );
  OAI22_X1 U14889 ( .A1(n19770), .A2(n11883), .B1(n11934), .B2(n11882), .ZN(
        n11884) );
  INV_X1 U14890 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n21007) );
  INV_X1 U14891 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12748) );
  OAI22_X1 U14892 ( .A1(n21007), .A2(n19502), .B1(n19350), .B2(n12748), .ZN(
        n11888) );
  INV_X1 U14893 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12612) );
  INV_X1 U14894 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12755) );
  OAI22_X1 U14895 ( .A1(n12612), .A2(n19275), .B1(n19602), .B2(n12755), .ZN(
        n11887) );
  NOR2_X1 U14896 ( .A1(n11888), .A2(n11887), .ZN(n11893) );
  INV_X1 U14897 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11890) );
  INV_X1 U14898 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11889) );
  INV_X1 U14899 ( .A(n11891), .ZN(n11892) );
  AOI22_X1 U14900 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11897), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11903) );
  INV_X1 U14901 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n21152) );
  AOI22_X1 U14902 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14903 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14904 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11900) );
  NAND4_X1 U14905 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n11910) );
  AOI22_X1 U14906 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14907 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U14908 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14909 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11905) );
  NAND4_X1 U14910 ( .A1(n11908), .A2(n11907), .A3(n11906), .A4(n11905), .ZN(
        n11909) );
  OR2_X2 U14911 ( .A1(n11910), .A2(n11909), .ZN(n12291) );
  NAND2_X1 U14912 ( .A1(n11776), .A2(n12291), .ZN(n13100) );
  OR2_X1 U14913 ( .A1(n12298), .A2(n13100), .ZN(n12214) );
  INV_X1 U14914 ( .A(n12216), .ZN(n12303) );
  NAND2_X1 U14915 ( .A1(n12214), .A2(n12303), .ZN(n11911) );
  INV_X1 U14916 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11914) );
  INV_X1 U14917 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11913) );
  OAI22_X1 U14918 ( .A1(n11914), .A2(n19444), .B1(n19384), .B2(n11913), .ZN(
        n11916) );
  INV_X1 U14919 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13269) );
  INV_X1 U14920 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12846) );
  OAI22_X1 U14921 ( .A1(n13269), .A2(n19275), .B1(n19350), .B2(n12846), .ZN(
        n11915) );
  NOR2_X1 U14922 ( .A1(n11916), .A2(n11915), .ZN(n11941) );
  INV_X1 U14923 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11918) );
  NOR2_X1 U14924 ( .A1(n11917), .A2(n11918), .ZN(n11926) );
  INV_X1 U14925 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11920) );
  INV_X1 U14926 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11919) );
  OAI22_X1 U14927 ( .A1(n11920), .A2(n19689), .B1(n19770), .B2(n11919), .ZN(
        n11925) );
  INV_X1 U14928 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11923) );
  INV_X1 U14929 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11922) );
  OAI22_X1 U14930 ( .A1(n11923), .A2(n11921), .B1(n19633), .B2(n11922), .ZN(
        n11924) );
  NOR3_X1 U14931 ( .A1(n11926), .A2(n11925), .A3(n11924), .ZN(n11940) );
  INV_X1 U14932 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11927) );
  NOR2_X1 U14933 ( .A1(n19733), .A2(n11927), .ZN(n11931) );
  INV_X1 U14934 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11929) );
  INV_X1 U14935 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11928) );
  OAI22_X1 U14936 ( .A1(n11929), .A2(n19325), .B1(n19475), .B2(n11928), .ZN(
        n11930) );
  NOR2_X1 U14937 ( .A1(n11931), .A2(n11930), .ZN(n11939) );
  INV_X1 U14938 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11933) );
  INV_X1 U14939 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11932) );
  OAI22_X1 U14940 ( .A1(n11933), .A2(n19502), .B1(n19416), .B2(n11932), .ZN(
        n11937) );
  INV_X1 U14941 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11935) );
  INV_X1 U14942 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12853) );
  OAI22_X1 U14943 ( .A1(n11935), .A2(n11934), .B1(n19602), .B2(n12853), .ZN(
        n11936) );
  NOR2_X1 U14944 ( .A1(n11937), .A2(n11936), .ZN(n11938) );
  NAND4_X1 U14945 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11944) );
  INV_X1 U14946 ( .A(n11942), .ZN(n12322) );
  NAND2_X1 U14947 ( .A1(n12322), .A2(n11776), .ZN(n11943) );
  NAND2_X1 U14948 ( .A1(n12208), .A2(n10051), .ZN(n11948) );
  OAI21_X1 U14949 ( .B1(n11947), .B2(n11946), .A(n12004), .ZN(n13639) );
  INV_X1 U14950 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16404) );
  NAND2_X1 U14951 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  OAI21_X1 U14952 ( .B1(n11953), .B2(n11952), .A(n11964), .ZN(n13647) );
  XNOR2_X1 U14953 ( .A(n11957), .B(n11954), .ZN(n13813) );
  XNOR2_X1 U14954 ( .A(n13813), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13056) );
  AND2_X1 U14955 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11955) );
  NAND2_X1 U14956 ( .A1(n19302), .A2(n11955), .ZN(n11956) );
  NAND2_X1 U14957 ( .A1(n11957), .A2(n11956), .ZN(n13760) );
  INV_X1 U14958 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13868) );
  OAI21_X1 U14959 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19958), .A(
        n12142), .ZN(n12181) );
  INV_X1 U14960 ( .A(n12291), .ZN(n11958) );
  MUX2_X1 U14961 ( .A(n12181), .B(n11958), .S(n11774), .Z(n12154) );
  INV_X1 U14962 ( .A(n12154), .ZN(n11959) );
  MUX2_X1 U14963 ( .A(n11959), .B(P2_EBX_REG_0__SCAN_IN), .S(n19302), .Z(
        n19124) );
  NAND2_X1 U14964 ( .A1(n19124), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13101) );
  OAI21_X1 U14965 ( .B1(n13760), .B2(n13868), .A(n13101), .ZN(n11961) );
  NAND2_X1 U14966 ( .A1(n13760), .A2(n13868), .ZN(n11960) );
  AND2_X1 U14967 ( .A1(n11961), .A2(n11960), .ZN(n13057) );
  NAND2_X1 U14968 ( .A1(n13056), .A2(n13057), .ZN(n13132) );
  INV_X1 U14969 ( .A(n13813), .ZN(n11962) );
  NAND2_X1 U14970 ( .A1(n11962), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11963) );
  AND2_X1 U14971 ( .A1(n13132), .A2(n11963), .ZN(n13670) );
  INV_X1 U14972 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12264) );
  INV_X1 U14973 ( .A(n11964), .ZN(n11965) );
  XNOR2_X1 U14974 ( .A(n11966), .B(n11965), .ZN(n19098) );
  XNOR2_X1 U14975 ( .A(n19098), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13843) );
  INV_X1 U14976 ( .A(n19098), .ZN(n11967) );
  INV_X1 U14977 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16405) );
  NAND2_X1 U14978 ( .A1(n16333), .A2(n16334), .ZN(n11970) );
  NAND2_X1 U14979 ( .A1(n11968), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11969) );
  NAND2_X1 U14980 ( .A1(n11970), .A2(n11969), .ZN(n13917) );
  INV_X1 U14981 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11972) );
  INV_X1 U14982 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11971) );
  OAI22_X1 U14983 ( .A1(n11972), .A2(n19325), .B1(n19384), .B2(n11971), .ZN(
        n11975) );
  INV_X1 U14984 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11973) );
  INV_X1 U14985 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12631) );
  OAI22_X1 U14986 ( .A1(n11973), .A2(n19444), .B1(n19275), .B2(n12631), .ZN(
        n11974) );
  NOR2_X1 U14987 ( .A1(n11975), .A2(n11974), .ZN(n11996) );
  INV_X1 U14988 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11976) );
  NOR2_X1 U14989 ( .A1(n19733), .A2(n11976), .ZN(n11983) );
  INV_X1 U14990 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11978) );
  INV_X1 U14991 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11977) );
  OAI22_X1 U14992 ( .A1(n11978), .A2(n11921), .B1(n19689), .B2(n11977), .ZN(
        n11982) );
  INV_X1 U14993 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11980) );
  INV_X1 U14994 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11979) );
  OAI22_X1 U14995 ( .A1(n11980), .A2(n19770), .B1(n19633), .B2(n11979), .ZN(
        n11981) );
  NOR3_X1 U14996 ( .A1(n11983), .A2(n11982), .A3(n11981), .ZN(n11995) );
  INV_X1 U14997 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11984) );
  NOR2_X1 U14998 ( .A1(n11917), .A2(n11984), .ZN(n11988) );
  INV_X1 U14999 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11986) );
  INV_X1 U15000 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11985) );
  OAI22_X1 U15001 ( .A1(n11986), .A2(n19416), .B1(n19475), .B2(n11985), .ZN(
        n11987) );
  NOR2_X1 U15002 ( .A1(n11988), .A2(n11987), .ZN(n11994) );
  INV_X1 U15003 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11989) );
  INV_X1 U15004 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12864) );
  OAI22_X1 U15005 ( .A1(n11989), .A2(n19502), .B1(n19350), .B2(n12864), .ZN(
        n11992) );
  INV_X1 U15006 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11990) );
  INV_X1 U15007 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12873) );
  OAI22_X1 U15008 ( .A1(n11990), .A2(n11934), .B1(n19602), .B2(n12873), .ZN(
        n11991) );
  NOR2_X1 U15009 ( .A1(n11992), .A2(n11991), .ZN(n11993) );
  NAND4_X1 U15010 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n11998) );
  NAND2_X1 U15011 ( .A1(n12326), .A2(n11776), .ZN(n11997) );
  NAND2_X1 U15012 ( .A1(n11998), .A2(n11997), .ZN(n12226) );
  OAI21_X1 U15013 ( .B1(n12001), .B2(n11999), .A(n12226), .ZN(n12002) );
  NOR2_X1 U15014 ( .A1(n11999), .A2(n12226), .ZN(n12000) );
  AND2_X1 U15015 ( .A1(n12004), .A2(n12003), .ZN(n12005) );
  OR2_X1 U15016 ( .A1(n12005), .A2(n12015), .ZN(n19089) );
  INV_X1 U15017 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12006) );
  XNOR2_X1 U15018 ( .A(n12007), .B(n12006), .ZN(n13918) );
  NAND2_X1 U15019 ( .A1(n13917), .A2(n13918), .ZN(n12009) );
  NAND2_X1 U15020 ( .A1(n12007), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12008) );
  NOR2_X1 U15021 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  OR2_X1 U15022 ( .A1(n12022), .A2(n12012), .ZN(n19073) );
  NOR2_X1 U15023 ( .A1(n19073), .A2(n10051), .ZN(n12016) );
  AND2_X1 U15024 ( .A1(n12016), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15077) );
  INV_X1 U15025 ( .A(n12013), .ZN(n12014) );
  XNOR2_X1 U15026 ( .A(n12015), .B(n12014), .ZN(n13727) );
  AND2_X1 U15027 ( .A1(n13727), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15324) );
  INV_X1 U15028 ( .A(n12016), .ZN(n12017) );
  INV_X1 U15029 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20961) );
  NAND2_X1 U15030 ( .A1(n12017), .A2(n20961), .ZN(n15078) );
  INV_X1 U15031 ( .A(n13727), .ZN(n12019) );
  INV_X1 U15032 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12018) );
  NAND2_X1 U15033 ( .A1(n12019), .A2(n12018), .ZN(n15323) );
  AND2_X1 U15034 ( .A1(n15078), .A2(n15323), .ZN(n12020) );
  NOR2_X1 U15035 ( .A1(n12022), .A2(n12512), .ZN(n12021) );
  MUX2_X1 U15036 ( .A(n12022), .B(n12021), .S(n19302), .Z(n12024) );
  INV_X1 U15037 ( .A(n12025), .ZN(n12023) );
  NOR2_X1 U15038 ( .A1(n12024), .A2(n12023), .ZN(n13655) );
  NAND2_X1 U15039 ( .A1(n13655), .A2(n12131), .ZN(n12034) );
  INV_X1 U15040 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16369) );
  AND2_X1 U15041 ( .A1(n12034), .A2(n16369), .ZN(n15310) );
  OR2_X1 U15042 ( .A1(n12025), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12029) );
  NAND2_X1 U15043 ( .A1(n12025), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12026) );
  OAI21_X1 U15044 ( .B1(n12026), .B2(n12130), .A(n12114), .ZN(n12027) );
  INV_X1 U15045 ( .A(n12027), .ZN(n12028) );
  NAND2_X1 U15046 ( .A1(n12029), .A2(n12028), .ZN(n19060) );
  INV_X1 U15047 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12030) );
  OAI21_X1 U15048 ( .B1(n19060), .B2(n10051), .A(n12030), .ZN(n15069) );
  NAND2_X1 U15049 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12029), .ZN(n12031) );
  NOR2_X1 U15050 ( .A1(n12130), .A2(n12031), .ZN(n12032) );
  NOR2_X1 U15051 ( .A1(n12033), .A2(n12032), .ZN(n13717) );
  AOI21_X1 U15052 ( .B1(n13717), .B2(n12131), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16300) );
  OR2_X1 U15053 ( .A1(n12034), .A2(n16369), .ZN(n15066) );
  INV_X1 U15054 ( .A(n19060), .ZN(n12036) );
  AND2_X1 U15055 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12035) );
  NAND2_X1 U15056 ( .A1(n12036), .A2(n12035), .ZN(n15068) );
  AND2_X1 U15057 ( .A1(n15066), .A2(n15068), .ZN(n16298) );
  AND2_X1 U15058 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12037) );
  OR2_X1 U15059 ( .A1(n12039), .A2(n12038), .ZN(n12040) );
  NAND2_X1 U15060 ( .A1(n12044), .A2(n12040), .ZN(n19050) );
  INV_X1 U15061 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12041) );
  OR3_X1 U15062 ( .A1(n19050), .A2(n10051), .A3(n12041), .ZN(n15057) );
  INV_X1 U15063 ( .A(n15057), .ZN(n12042) );
  OAI21_X1 U15064 ( .B1(n19050), .B2(n10051), .A(n12041), .ZN(n15058) );
  NAND2_X1 U15065 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  NAND2_X1 U15066 ( .A1(n12060), .A2(n12045), .ZN(n13895) );
  NOR2_X1 U15067 ( .A1(n13895), .A2(n10051), .ZN(n12080) );
  NOR2_X1 U15068 ( .A1(n12080), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16282) );
  NAND2_X1 U15069 ( .A1(n19302), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12046) );
  NOR2_X1 U15070 ( .A1(n12063), .A2(n12046), .ZN(n12047) );
  NOR2_X1 U15071 ( .A1(n12048), .A2(n12047), .ZN(n12076) );
  AOI21_X1 U15072 ( .B1(n12076), .B2(n12131), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14979) );
  INV_X1 U15073 ( .A(n12049), .ZN(n12050) );
  XNOR2_X1 U15074 ( .A(n12051), .B(n12050), .ZN(n14703) );
  AOI21_X1 U15075 ( .B1(n14703), .B2(n12131), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15024) );
  INV_X1 U15076 ( .A(n12052), .ZN(n12053) );
  MUX2_X1 U15077 ( .A(P2_EBX_REG_16__SCAN_IN), .B(n12053), .S(n12058), .Z(
        n12054) );
  NAND2_X1 U15078 ( .A1(n12054), .A2(n12114), .ZN(n19011) );
  OR2_X1 U15079 ( .A1(n19011), .A2(n10051), .ZN(n12055) );
  INV_X1 U15080 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15033) );
  XNOR2_X1 U15081 ( .A(n12055), .B(n15033), .ZN(n14971) );
  OR2_X1 U15082 ( .A1(n9811), .A2(n12056), .ZN(n12057) );
  NAND2_X1 U15083 ( .A1(n12058), .A2(n12057), .ZN(n19030) );
  INV_X1 U15084 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15291) );
  OAI21_X1 U15085 ( .B1(n19030), .B2(n10051), .A(n15291), .ZN(n15281) );
  XNOR2_X1 U15086 ( .A(n12060), .B(n12059), .ZN(n12081) );
  INV_X1 U15087 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16344) );
  OAI21_X1 U15088 ( .B1(n12081), .B2(n10051), .A(n16344), .ZN(n15279) );
  NAND2_X1 U15089 ( .A1(n15281), .A2(n15279), .ZN(n14969) );
  NOR4_X1 U15090 ( .A1(n14979), .A2(n15024), .A3(n14971), .A4(n14969), .ZN(
        n12074) );
  NOR2_X1 U15091 ( .A1(n12066), .A2(n12544), .ZN(n12061) );
  MUX2_X1 U15092 ( .A(n12066), .B(n12061), .S(n19302), .Z(n12062) );
  INV_X1 U15093 ( .A(n12062), .ZN(n12065) );
  INV_X1 U15094 ( .A(n12063), .ZN(n12064) );
  NAND2_X1 U15095 ( .A1(n12065), .A2(n12064), .ZN(n18978) );
  INV_X1 U15096 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15219) );
  OAI21_X1 U15097 ( .B1(n18978), .B2(n10051), .A(n15219), .ZN(n14976) );
  INV_X1 U15098 ( .A(n12066), .ZN(n12068) );
  INV_X1 U15099 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12536) );
  NAND2_X1 U15100 ( .A1(n10216), .A2(n12536), .ZN(n12071) );
  NAND3_X1 U15101 ( .A1(n12071), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n19302), 
        .ZN(n12067) );
  NAND2_X1 U15102 ( .A1(n12068), .A2(n12067), .ZN(n18987) );
  OR2_X1 U15103 ( .A1(n18987), .A2(n10051), .ZN(n12078) );
  INV_X1 U15104 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15230) );
  NAND2_X1 U15105 ( .A1(n12078), .A2(n15230), .ZN(n14997) );
  NAND2_X1 U15106 ( .A1(n12069), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12070) );
  MUX2_X1 U15107 ( .A(n12070), .B(n12069), .S(n12130), .Z(n12072) );
  NAND2_X1 U15108 ( .A1(n12072), .A2(n12071), .ZN(n12086) );
  INV_X1 U15109 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15240) );
  AND2_X1 U15110 ( .A1(n14997), .A2(n15016), .ZN(n14974) );
  INV_X1 U15111 ( .A(n12076), .ZN(n14701) );
  NAND2_X1 U15112 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12077) );
  NOR2_X1 U15113 ( .A1(n14701), .A2(n12077), .ZN(n14978) );
  INV_X1 U15114 ( .A(n12078), .ZN(n12079) );
  NAND2_X1 U15115 ( .A1(n12079), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14998) );
  NAND2_X1 U15116 ( .A1(n12080), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16280) );
  INV_X1 U15117 ( .A(n12081), .ZN(n19036) );
  AND2_X1 U15118 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12082) );
  NAND2_X1 U15119 ( .A1(n19036), .A2(n12082), .ZN(n15046) );
  AND2_X1 U15120 ( .A1(n16280), .A2(n15046), .ZN(n15045) );
  NAND2_X1 U15121 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12083) );
  OR2_X1 U15122 ( .A1(n19030), .A2(n12083), .ZN(n15282) );
  AND2_X1 U15123 ( .A1(n15045), .A2(n15282), .ZN(n14970) );
  AND2_X1 U15124 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12084) );
  NAND2_X1 U15125 ( .A1(n14703), .A2(n12084), .ZN(n15025) );
  OR3_X1 U15126 ( .A1(n19011), .A2(n10051), .A3(n15033), .ZN(n14972) );
  NAND4_X1 U15127 ( .A1(n14998), .A2(n14970), .A3(n15025), .A4(n14972), .ZN(
        n12085) );
  NOR2_X1 U15128 ( .A1(n14978), .A2(n12085), .ZN(n12089) );
  INV_X1 U15129 ( .A(n12086), .ZN(n19002) );
  AND2_X1 U15130 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12087) );
  NAND2_X1 U15131 ( .A1(n19002), .A2(n12087), .ZN(n15013) );
  NAND2_X1 U15132 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12088) );
  INV_X1 U15133 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n14778) );
  NOR2_X1 U15134 ( .A1(n12130), .A2(n14778), .ZN(n12091) );
  NAND2_X1 U15135 ( .A1(n12092), .A2(n12091), .ZN(n12093) );
  AND2_X1 U15136 ( .A1(n12097), .A2(n12093), .ZN(n15778) );
  NAND2_X1 U15137 ( .A1(n15778), .A2(n12131), .ZN(n12094) );
  INV_X1 U15138 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U15139 ( .A1(n12094), .A2(n15194), .ZN(n14959) );
  NOR2_X1 U15140 ( .A1(n12094), .A2(n15194), .ZN(n14961) );
  XNOR2_X1 U15141 ( .A(n12095), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13974) );
  NAND3_X1 U15142 ( .A1(n12098), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n19302), 
        .ZN(n12099) );
  NAND2_X1 U15143 ( .A1(n12099), .A2(n12114), .ZN(n12100) );
  OR2_X1 U15144 ( .A1(n9785), .A2(n12100), .ZN(n16245) );
  INV_X1 U15145 ( .A(n16245), .ZN(n12101) );
  NAND2_X1 U15146 ( .A1(n12101), .A2(n12131), .ZN(n12103) );
  INV_X1 U15147 ( .A(n12103), .ZN(n12102) );
  NAND2_X1 U15148 ( .A1(n12102), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14948) );
  INV_X1 U15149 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15168) );
  AND2_X1 U15150 ( .A1(n12103), .A2(n15168), .ZN(n14949) );
  INV_X1 U15151 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12564) );
  NAND3_X1 U15152 ( .A1(n19302), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n12104), 
        .ZN(n12105) );
  AND2_X1 U15153 ( .A1(n12131), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12106) );
  NAND2_X1 U15154 ( .A1(n16217), .A2(n12106), .ZN(n12124) );
  INV_X1 U15155 ( .A(n16217), .ZN(n12107) );
  INV_X1 U15156 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15144) );
  OAI21_X1 U15157 ( .B1(n12107), .B2(n10051), .A(n15144), .ZN(n12108) );
  NAND2_X1 U15158 ( .A1(n19302), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12110) );
  INV_X1 U15159 ( .A(n12110), .ZN(n12111) );
  NAND2_X1 U15160 ( .A1(n12111), .A2(n9781), .ZN(n12112) );
  NAND2_X1 U15161 ( .A1(n12119), .A2(n12112), .ZN(n16209) );
  INV_X1 U15162 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15134) );
  NAND2_X1 U15163 ( .A1(n19302), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12113) );
  MUX2_X1 U15164 ( .A(n12113), .B(P2_EBX_REG_25__SCAN_IN), .S(n9785), .Z(
        n12115) );
  NAND2_X1 U15165 ( .A1(n12115), .A2(n12114), .ZN(n16228) );
  INV_X1 U15166 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15158) );
  NOR2_X1 U15167 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12121) );
  INV_X1 U15168 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12117) );
  NOR2_X1 U15169 ( .A1(n12130), .A2(n12117), .ZN(n12118) );
  NAND2_X1 U15170 ( .A1(n12119), .A2(n12118), .ZN(n12120) );
  NAND2_X1 U15171 ( .A1(n12129), .A2(n12120), .ZN(n16198) );
  NAND2_X1 U15172 ( .A1(n12125), .A2(n10267), .ZN(n12126) );
  INV_X1 U15173 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12581) );
  NOR2_X1 U15174 ( .A1(n12130), .A2(n12581), .ZN(n12128) );
  XNOR2_X1 U15175 ( .A(n10218), .B(n12128), .ZN(n12133) );
  AOI21_X1 U15176 ( .B1(n12133), .B2(n12131), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14896) );
  INV_X1 U15177 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12585) );
  INV_X1 U15178 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15092) );
  OAI21_X1 U15179 ( .B1(n16187), .B2(n10051), .A(n15092), .ZN(n14888) );
  AND3_X1 U15180 ( .A1(n12132), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12131), .ZN(n14887) );
  INV_X1 U15181 ( .A(n12133), .ZN(n12990) );
  INV_X1 U15182 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14901) );
  NOR3_X1 U15183 ( .A1(n12990), .A2(n10051), .A3(n14901), .ZN(n14897) );
  NOR2_X1 U15184 ( .A1(n12135), .A2(n12134), .ZN(n12136) );
  NOR2_X1 U15185 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15858), .ZN(
        n12137) );
  INV_X1 U15186 ( .A(n12197), .ZN(n12144) );
  INV_X1 U15187 ( .A(n12192), .ZN(n12141) );
  NOR2_X1 U15188 ( .A1(n12141), .A2(n12186), .ZN(n12145) );
  XNOR2_X1 U15189 ( .A(n12180), .B(n12142), .ZN(n12182) );
  NAND2_X1 U15190 ( .A1(n12145), .A2(n12182), .ZN(n12143) );
  INV_X1 U15191 ( .A(n12181), .ZN(n12183) );
  AOI21_X1 U15192 ( .B1(n12183), .B2(n12145), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n12146) );
  INV_X1 U15193 ( .A(n12146), .ZN(n12147) );
  OR2_X1 U15194 ( .A1(n16445), .A2(n12147), .ZN(n12151) );
  NAND2_X1 U15195 ( .A1(n11538), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12148) );
  NAND2_X1 U15196 ( .A1(n12148), .A2(n15589), .ZN(n16452) );
  INV_X1 U15197 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12149) );
  OAI21_X1 U15198 ( .B1(n12383), .B2(n16452), .A(n12149), .ZN(n12150) );
  NAND2_X1 U15199 ( .A1(n12150), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19950) );
  NAND2_X1 U15200 ( .A1(n12151), .A2(n19950), .ZN(n16466) );
  NAND2_X1 U15201 ( .A1(n16466), .A2(n15585), .ZN(n12158) );
  INV_X1 U15202 ( .A(n12180), .ZN(n12153) );
  OAI21_X1 U15203 ( .B1(n12154), .B2(n12153), .A(n12152), .ZN(n12155) );
  AND2_X1 U15204 ( .A1(n12192), .A2(n12155), .ZN(n12156) );
  OR2_X1 U15205 ( .A1(n12197), .A2(n12156), .ZN(n19961) );
  AND2_X1 U15206 ( .A1(n11776), .A2(n12973), .ZN(n12253) );
  NAND2_X1 U15207 ( .A1(n12158), .A2(n12157), .ZN(n12161) );
  INV_X1 U15208 ( .A(n16456), .ZN(n12160) );
  NAND2_X1 U15209 ( .A1(n12161), .A2(n12160), .ZN(n13045) );
  NAND2_X1 U15210 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n15853) );
  INV_X1 U15211 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18948) );
  NOR2_X1 U15212 ( .A1(n18948), .A2(n19866), .ZN(n19858) );
  NOR2_X1 U15213 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19859) );
  NOR3_X1 U15214 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19858), .A3(n19859), 
        .ZN(n19850) );
  NAND2_X1 U15215 ( .A1(n15853), .A2(n19850), .ZN(n13203) );
  INV_X1 U15216 ( .A(n13203), .ZN(n13043) );
  NAND2_X1 U15217 ( .A1(n12162), .A2(n13043), .ZN(n12163) );
  OR2_X1 U15218 ( .A1(n16445), .A2(n12163), .ZN(n12174) );
  INV_X1 U15219 ( .A(n12164), .ZN(n12165) );
  NAND2_X1 U15220 ( .A1(n12165), .A2(n11750), .ZN(n16451) );
  NAND2_X1 U15221 ( .A1(n12166), .A2(n12253), .ZN(n12168) );
  NAND3_X1 U15222 ( .A1(n12168), .A2(n19290), .A3(n12167), .ZN(n12173) );
  NAND2_X1 U15223 ( .A1(n12169), .A2(n11776), .ZN(n12240) );
  INV_X1 U15224 ( .A(n12929), .ZN(n19316) );
  AOI21_X1 U15225 ( .B1(n12240), .B2(n11750), .A(n19316), .ZN(n12171) );
  INV_X1 U15226 ( .A(n11773), .ZN(n12245) );
  OAI211_X1 U15227 ( .C1(n12171), .C2(n12247), .A(n12170), .B(n12245), .ZN(
        n12172) );
  AOI21_X1 U15228 ( .B1(n16451), .B2(n12173), .A(n12172), .ZN(n12242) );
  NAND2_X1 U15229 ( .A1(n12174), .A2(n12242), .ZN(n13197) );
  MUX2_X1 U15230 ( .A(n12175), .B(n19290), .S(n11776), .Z(n12176) );
  OR2_X1 U15231 ( .A1(n12176), .A2(n19857), .ZN(n12177) );
  NOR2_X1 U15232 ( .A1(n16445), .A2(n12177), .ZN(n12178) );
  NOR2_X1 U15233 ( .A1(n13197), .A2(n12178), .ZN(n12205) );
  AOI21_X1 U15234 ( .B1(n12196), .B2(n15585), .A(n12179), .ZN(n12188) );
  OAI21_X1 U15235 ( .B1(n12181), .B2(n12153), .A(n11774), .ZN(n12185) );
  OAI211_X1 U15236 ( .C1(n15585), .C2(n12183), .A(n11750), .B(n12182), .ZN(
        n12184) );
  OAI211_X1 U15237 ( .C1(n11763), .C2(n12186), .A(n12185), .B(n12184), .ZN(
        n12187) );
  OAI21_X1 U15238 ( .B1(n12189), .B2(n12188), .A(n12187), .ZN(n12190) );
  NAND2_X1 U15239 ( .A1(n12192), .A2(n12190), .ZN(n12191) );
  OAI21_X1 U15240 ( .B1(n12192), .B2(n11774), .A(n12191), .ZN(n12193) );
  INV_X1 U15241 ( .A(n12193), .ZN(n12194) );
  MUX2_X1 U15242 ( .A(n12195), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n21158), .Z(n12200) );
  NAND2_X1 U15243 ( .A1(n12197), .A2(n19187), .ZN(n12198) );
  AND2_X1 U15244 ( .A1(n16449), .A2(n15585), .ZN(n19183) );
  NOR2_X1 U15245 ( .A1(n19290), .A2(n13203), .ZN(n12199) );
  NAND2_X1 U15246 ( .A1(n19183), .A2(n12199), .ZN(n12204) );
  INV_X1 U15247 ( .A(n19183), .ZN(n12202) );
  AOI21_X1 U15248 ( .B1(n12200), .B2(n11750), .A(n19297), .ZN(n12201) );
  NAND2_X1 U15249 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  NAND4_X1 U15250 ( .A1(n13045), .A2(n12205), .A3(n12204), .A4(n12203), .ZN(
        n12207) );
  NAND2_X1 U15251 ( .A1(n16467), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12983) );
  INV_X1 U15252 ( .A(n12983), .ZN(n12206) );
  NOR2_X1 U15253 ( .A1(n16456), .A2(n12587), .ZN(n19963) );
  NAND2_X1 U15254 ( .A1(n12209), .A2(n16404), .ZN(n16328) );
  NAND2_X1 U15255 ( .A1(n13835), .A2(n16405), .ZN(n12221) );
  NAND2_X1 U15256 ( .A1(n13100), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13099) );
  INV_X1 U15257 ( .A(n13099), .ZN(n12211) );
  XNOR2_X1 U15258 ( .A(n12298), .B(n12291), .ZN(n12212) );
  NAND2_X1 U15259 ( .A1(n12211), .A2(n12212), .ZN(n12213) );
  XNOR2_X1 U15260 ( .A(n13099), .B(n12212), .ZN(n13032) );
  NAND2_X1 U15261 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13032), .ZN(
        n13031) );
  NAND2_X1 U15262 ( .A1(n12213), .A2(n13031), .ZN(n12217) );
  XOR2_X1 U15263 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12217), .Z(
        n13062) );
  INV_X1 U15264 ( .A(n12214), .ZN(n12215) );
  XNOR2_X1 U15265 ( .A(n12216), .B(n12215), .ZN(n13061) );
  NAND2_X1 U15266 ( .A1(n13062), .A2(n13061), .ZN(n13060) );
  NAND2_X1 U15267 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12217), .ZN(
        n12218) );
  NAND2_X1 U15268 ( .A1(n13060), .A2(n12218), .ZN(n12219) );
  XNOR2_X1 U15269 ( .A(n12219), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13671) );
  NAND2_X1 U15270 ( .A1(n12219), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12220) );
  INV_X1 U15271 ( .A(n13835), .ZN(n12222) );
  NAND2_X1 U15272 ( .A1(n12222), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12223) );
  NAND2_X1 U15273 ( .A1(n12224), .A2(n12223), .ZN(n16330) );
  NAND2_X2 U15274 ( .A1(n16328), .A2(n16330), .ZN(n12230) );
  INV_X1 U15275 ( .A(n12225), .ZN(n12231) );
  INV_X1 U15276 ( .A(n12226), .ZN(n12227) );
  OR2_X1 U15277 ( .A1(n16329), .A2(n12227), .ZN(n12229) );
  OAI211_X2 U15278 ( .C1(n12230), .C2(n12231), .A(n12229), .B(n12228), .ZN(
        n13920) );
  NAND2_X1 U15279 ( .A1(n13920), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13919) );
  NAND2_X1 U15280 ( .A1(n12230), .A2(n16329), .ZN(n12232) );
  NAND2_X1 U15281 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  NAND2_X1 U15282 ( .A1(n12234), .A2(n10051), .ZN(n12235) );
  NAND2_X1 U15283 ( .A1(n12236), .A2(n12235), .ZN(n15327) );
  XNOR2_X1 U15284 ( .A(n12236), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15083) );
  NAND2_X1 U15285 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16340) );
  NOR2_X1 U15286 ( .A1(n16340), .A2(n16344), .ZN(n12239) );
  NAND2_X1 U15287 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16370) );
  INV_X1 U15288 ( .A(n16370), .ZN(n12238) );
  AND2_X1 U15289 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n12238), .ZN(
        n15296) );
  AND2_X1 U15290 ( .A1(n12239), .A2(n15296), .ZN(n12266) );
  AND2_X1 U15291 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15253) );
  AND2_X1 U15292 ( .A1(n15253), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15239) );
  NAND2_X1 U15293 ( .A1(n15239), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15215) );
  NAND2_X1 U15294 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15207) );
  INV_X1 U15295 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13976) );
  AND2_X1 U15296 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15140) );
  INV_X1 U15297 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15117) );
  NOR2_X1 U15298 ( .A1(n16456), .A2(n16469), .ZN(n19962) );
  INV_X1 U15299 ( .A(n12240), .ZN(n12241) );
  NAND2_X1 U15300 ( .A1(n12598), .A2(n16441), .ZN(n15259) );
  NOR2_X1 U15301 ( .A1(n12243), .A2(n12245), .ZN(n12244) );
  NAND2_X1 U15302 ( .A1(n11785), .A2(n12244), .ZN(n12259) );
  NAND2_X1 U15303 ( .A1(n12245), .A2(n19297), .ZN(n12248) );
  INV_X1 U15304 ( .A(n12246), .ZN(n13042) );
  AOI22_X1 U15305 ( .A1(n12248), .A2(n13042), .B1(n12973), .B2(n12247), .ZN(
        n12250) );
  INV_X1 U15306 ( .A(n12249), .ZN(n12593) );
  NAND2_X1 U15307 ( .A1(n11740), .A2(n12593), .ZN(n12912) );
  AND3_X1 U15308 ( .A1(n12251), .A2(n12250), .A3(n12912), .ZN(n12258) );
  NAND2_X1 U15309 ( .A1(n12252), .A2(n15585), .ZN(n13608) );
  OAI21_X1 U15310 ( .B1(n12166), .B2(n19316), .A(n12253), .ZN(n12254) );
  NAND2_X1 U15311 ( .A1(n13608), .A2(n12254), .ZN(n12256) );
  NAND2_X1 U15312 ( .A1(n12256), .A2(n12255), .ZN(n12257) );
  INV_X1 U15313 ( .A(n12260), .ZN(n13184) );
  NAND2_X1 U15314 ( .A1(n13606), .A2(n13184), .ZN(n12261) );
  NAND2_X1 U15315 ( .A1(n12598), .A2(n12261), .ZN(n15264) );
  NAND2_X1 U15316 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13069) );
  INV_X1 U15317 ( .A(n13069), .ZN(n13051) );
  INV_X1 U15318 ( .A(n12598), .ZN(n12262) );
  INV_X2 U15319 ( .A(n19255), .ZN(n19058) );
  NAND2_X1 U15320 ( .A1(n12262), .A2(n19058), .ZN(n13112) );
  OAI21_X1 U15321 ( .B1(n15264), .B2(n13051), .A(n13112), .ZN(n13070) );
  NOR2_X1 U15322 ( .A1(n15264), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12263) );
  NOR2_X1 U15323 ( .A1(n13070), .A2(n12263), .ZN(n13837) );
  NAND2_X1 U15324 ( .A1(n13837), .A2(n15265), .ZN(n15297) );
  INV_X1 U15325 ( .A(n15297), .ZN(n16362) );
  INV_X1 U15326 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U15327 ( .A1(n12468), .A2(n13069), .ZN(n13838) );
  INV_X1 U15328 ( .A(n13838), .ZN(n12469) );
  NAND2_X1 U15329 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15339) );
  INV_X1 U15330 ( .A(n15339), .ZN(n16402) );
  NAND2_X1 U15331 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16402), .ZN(
        n15331) );
  NOR2_X1 U15332 ( .A1(n12018), .A2(n20961), .ZN(n16384) );
  INV_X1 U15333 ( .A(n16384), .ZN(n12470) );
  NOR3_X1 U15334 ( .A1(n12469), .A2(n15331), .A3(n12470), .ZN(n12265) );
  NAND2_X1 U15335 ( .A1(n15330), .A2(n12264), .ZN(n16411) );
  OAI211_X1 U15336 ( .C1(n15265), .C2(n12265), .A(n13837), .B(n16411), .ZN(
        n15314) );
  INV_X1 U15337 ( .A(n12266), .ZN(n12471) );
  OR2_X1 U15338 ( .A1(n15314), .A2(n12471), .ZN(n15262) );
  INV_X1 U15339 ( .A(n15215), .ZN(n12472) );
  INV_X1 U15340 ( .A(n15207), .ZN(n15218) );
  NAND3_X1 U15341 ( .A1(n12472), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15218), .ZN(n12267) );
  OAI21_X1 U15342 ( .B1(n15262), .B2(n12267), .A(n15297), .ZN(n15178) );
  NOR2_X1 U15343 ( .A1(n15194), .A2(n13976), .ZN(n15184) );
  OAI21_X1 U15344 ( .B1(n15265), .B2(n15184), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12268) );
  INV_X1 U15345 ( .A(n12268), .ZN(n12269) );
  NAND2_X1 U15346 ( .A1(n15178), .A2(n12269), .ZN(n15166) );
  NAND2_X1 U15347 ( .A1(n15166), .A2(n15297), .ZN(n15159) );
  OAI21_X1 U15348 ( .B1(n15140), .B2(n16362), .A(n15159), .ZN(n15103) );
  AND2_X1 U15349 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15104) );
  AOI21_X1 U15350 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15104), .A(
        n16362), .ZN(n12270) );
  NOR2_X1 U15351 ( .A1(n15103), .A2(n12270), .ZN(n15091) );
  OAI21_X1 U15352 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15265), .A(
        n15091), .ZN(n12599) );
  NOR2_X2 U15353 ( .A1(n12283), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15354 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15355 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15356 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15357 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12271) );
  NAND4_X1 U15358 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12280) );
  AOI22_X1 U15359 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15360 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15361 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15362 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12275) );
  NAND4_X1 U15363 ( .A1(n12278), .A2(n12277), .A3(n12276), .A4(n12275), .ZN(
        n12279) );
  INV_X1 U15364 ( .A(n13589), .ZN(n12285) );
  INV_X2 U15365 ( .A(n12296), .ZN(n12443) );
  AND2_X2 U15366 ( .A1(n15585), .A2(n19509), .ZN(n12293) );
  AOI22_X1 U15367 ( .A1(n12443), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12284) );
  OAI21_X1 U15368 ( .B1(n12285), .B2(n12281), .A(n12284), .ZN(n12286) );
  AOI21_X1 U15369 ( .B1(n12459), .B2(P2_REIP_REG_11__SCAN_IN), .A(n12286), 
        .ZN(n13373) );
  AOI222_X1 U15370 ( .A1(n12459), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12443), .C2(
        P2_EAX_REG_7__SCAN_IN), .ZN(n13729) );
  INV_X1 U15371 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n12290) );
  INV_X1 U15372 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19254) );
  NAND2_X1 U15373 ( .A1(n15585), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12287) );
  OAI211_X1 U15374 ( .C1(n12929), .C2(n19254), .A(n12287), .B(n19509), .ZN(
        n12288) );
  INV_X1 U15375 ( .A(n12288), .ZN(n12289) );
  OAI21_X1 U15376 ( .B1(n12450), .B2(n12290), .A(n12289), .ZN(n13109) );
  INV_X1 U15377 ( .A(n12281), .ZN(n12292) );
  INV_X1 U15378 ( .A(n11742), .ZN(n12916) );
  NAND2_X1 U15379 ( .A1(n12916), .A2(n12293), .ZN(n12304) );
  NAND2_X1 U15380 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12294) );
  NAND4_X1 U15381 ( .A1(n12295), .A2(n12296), .A3(n12304), .A4(n12294), .ZN(
        n13108) );
  NAND2_X1 U15382 ( .A1(n13109), .A2(n13108), .ZN(n13107) );
  AOI22_X1 U15383 ( .A1(n12282), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12293), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12297) );
  XNOR2_X1 U15384 ( .A(n13107), .B(n9787), .ZN(n13026) );
  OR2_X1 U15385 ( .A1(n12298), .A2(n12281), .ZN(n12301) );
  NAND2_X1 U15386 ( .A1(n11742), .A2(n12929), .ZN(n12299) );
  MUX2_X1 U15387 ( .A(n12299), .B(n19949), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12300) );
  NAND2_X1 U15388 ( .A1(n12301), .A2(n12300), .ZN(n13025) );
  OR2_X2 U15389 ( .A1(n13026), .A2(n13025), .ZN(n13028) );
  NAND2_X1 U15390 ( .A1(n9787), .A2(n13107), .ZN(n12302) );
  NAND2_X1 U15391 ( .A1(n13028), .A2(n12302), .ZN(n12309) );
  OR2_X1 U15392 ( .A1(n12281), .A2(n12303), .ZN(n12305) );
  OAI211_X1 U15393 ( .C1(n19940), .C2(n19509), .A(n12305), .B(n12304), .ZN(
        n12308) );
  XNOR2_X1 U15394 ( .A(n12309), .B(n12308), .ZN(n13054) );
  NAND2_X1 U15395 ( .A1(n12459), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15396 ( .A1(n12443), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12458), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12306) );
  AND2_X1 U15397 ( .A1(n12307), .A2(n12306), .ZN(n13053) );
  INV_X1 U15398 ( .A(n12308), .ZN(n12310) );
  NAND2_X1 U15399 ( .A1(n12310), .A2(n12309), .ZN(n12311) );
  INV_X1 U15400 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19872) );
  NAND2_X1 U15401 ( .A1(n12282), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12313) );
  NAND2_X1 U15402 ( .A1(n12293), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12312) );
  OAI211_X1 U15403 ( .C1(n19509), .C2(n19933), .A(n12313), .B(n12312), .ZN(
        n12314) );
  INV_X1 U15404 ( .A(n12314), .ZN(n12317) );
  OR2_X1 U15405 ( .A1(n12281), .A2(n12315), .ZN(n12316) );
  OAI211_X1 U15406 ( .C1(n12450), .C2(n19872), .A(n12317), .B(n12316), .ZN(
        n13531) );
  INV_X1 U15407 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15408 ( .A1(n12443), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12458), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12320) );
  OR2_X1 U15409 ( .A1(n12281), .A2(n12318), .ZN(n12319) );
  OAI211_X1 U15410 ( .C1(n12450), .C2(n12321), .A(n12320), .B(n12319), .ZN(
        n13535) );
  INV_X1 U15411 ( .A(n13536), .ZN(n13636) );
  INV_X1 U15412 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15413 ( .A1(n12443), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12458), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12324) );
  OR2_X1 U15414 ( .A1(n12281), .A2(n12322), .ZN(n12323) );
  OAI211_X1 U15415 ( .C1(n12450), .C2(n12325), .A(n12324), .B(n12323), .ZN(
        n13637) );
  NAND2_X1 U15416 ( .A1(n13636), .A2(n13637), .ZN(n13635) );
  OR2_X1 U15417 ( .A1(n12281), .A2(n12326), .ZN(n12327) );
  INV_X1 U15418 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15419 ( .A1(n12443), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12458), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12328) );
  OAI21_X1 U15420 ( .B1(n12450), .B2(n12329), .A(n12328), .ZN(n15342) );
  AND2_X2 U15421 ( .A1(n15343), .A2(n15342), .ZN(n15345) );
  AOI21_X1 U15422 ( .B1(n12331), .B2(n12330), .A(n15345), .ZN(n13730) );
  INV_X1 U15423 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15424 ( .A1(n12443), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12458), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15425 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15426 ( .A1(n12383), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15427 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15428 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12332) );
  NAND4_X1 U15429 ( .A1(n12335), .A2(n12334), .A3(n12333), .A4(n12332), .ZN(
        n12341) );
  AOI22_X1 U15430 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15431 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15432 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15433 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12336) );
  NAND4_X1 U15434 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12340) );
  INV_X1 U15435 ( .A(n13394), .ZN(n12342) );
  OR2_X1 U15436 ( .A1(n12281), .A2(n12342), .ZN(n12343) );
  OAI211_X1 U15437 ( .C1(n12450), .C2(n12345), .A(n12344), .B(n12343), .ZN(
        n13124) );
  NAND2_X1 U15438 ( .A1(n13123), .A2(n13124), .ZN(n13217) );
  AOI22_X1 U15439 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12383), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15440 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12730), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15441 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11898), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15442 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12346) );
  NAND4_X1 U15443 ( .A1(n12349), .A2(n12348), .A3(n12347), .A4(n12346), .ZN(
        n12355) );
  AOI22_X1 U15444 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15445 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15446 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15447 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12737), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12350) );
  NAND4_X1 U15448 ( .A1(n12353), .A2(n12352), .A3(n12351), .A4(n12350), .ZN(
        n12354) );
  NOR2_X1 U15449 ( .A1(n12355), .A2(n12354), .ZN(n13552) );
  AOI22_X1 U15450 ( .A1(n12443), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12458), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12356) );
  OAI21_X1 U15451 ( .B1(n13552), .B2(n12281), .A(n12356), .ZN(n12357) );
  AOI21_X1 U15452 ( .B1(n12459), .B2(P2_REIP_REG_9__SCAN_IN), .A(n12357), .ZN(
        n13218) );
  AOI22_X1 U15453 ( .A1(n12443), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15454 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12383), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15455 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12730), .B1(
        n12729), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15456 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12414), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15457 ( .A1(n11634), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12358) );
  NAND4_X1 U15458 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12367) );
  AOI22_X1 U15459 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15460 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15461 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15462 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11586), .B1(
        n11904), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12362) );
  NAND4_X1 U15463 ( .A1(n12365), .A2(n12364), .A3(n12363), .A4(n12362), .ZN(
        n12366) );
  NOR2_X1 U15464 ( .A1(n12367), .A2(n12366), .ZN(n13555) );
  OR2_X1 U15465 ( .A1(n12281), .A2(n13555), .ZN(n12368) );
  OAI211_X1 U15466 ( .C1(n12450), .C2(n19880), .A(n12369), .B(n12368), .ZN(
        n13262) );
  AOI22_X1 U15467 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U15468 ( .A1(n12383), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15469 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15470 ( .A1(n11899), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12370) );
  NAND4_X1 U15471 ( .A1(n12373), .A2(n12372), .A3(n12371), .A4(n12370), .ZN(
        n12379) );
  AOI22_X1 U15472 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15473 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15474 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15475 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12374) );
  NAND4_X1 U15476 ( .A1(n12377), .A2(n12376), .A3(n12375), .A4(n12374), .ZN(
        n12378) );
  OR2_X1 U15477 ( .A1(n12379), .A2(n12378), .ZN(n13588) );
  INV_X1 U15478 ( .A(n13588), .ZN(n12382) );
  NAND2_X1 U15479 ( .A1(n12459), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15480 ( .A1(n12443), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12380) );
  OAI211_X1 U15481 ( .C1(n12382), .C2(n12281), .A(n12381), .B(n12380), .ZN(
        n15300) );
  AOI22_X1 U15482 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15483 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15484 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15485 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12384) );
  NAND4_X1 U15486 ( .A1(n12387), .A2(n12386), .A3(n12385), .A4(n12384), .ZN(
        n12393) );
  AOI22_X1 U15487 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12391) );
  AOI22_X1 U15488 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12390) );
  AOI22_X1 U15489 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15490 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12388) );
  NAND4_X1 U15491 ( .A1(n12391), .A2(n12390), .A3(n12389), .A4(n12388), .ZN(
        n12392) );
  INV_X1 U15492 ( .A(n13524), .ZN(n12634) );
  AOI22_X1 U15493 ( .A1(n12443), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12394) );
  OAI21_X1 U15494 ( .B1(n12634), .B2(n12281), .A(n12394), .ZN(n12395) );
  AOI21_X1 U15495 ( .B1(n12459), .B2(P2_REIP_REG_13__SCAN_IN), .A(n12395), 
        .ZN(n13509) );
  INV_X1 U15496 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15497 ( .A1(n12443), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15498 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12383), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15499 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12730), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15500 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15501 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11899), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12396) );
  NAND4_X1 U15502 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12405) );
  AOI22_X1 U15503 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15504 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12735), .ZN(n12402) );
  AOI22_X1 U15505 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12737), .B1(
        n11904), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15506 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11586), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12400) );
  NAND4_X1 U15507 ( .A1(n12403), .A2(n12402), .A3(n12401), .A4(n12400), .ZN(
        n12404) );
  NOR2_X1 U15508 ( .A1(n12405), .A2(n12404), .ZN(n12632) );
  OR2_X1 U15509 ( .A1(n12281), .A2(n12632), .ZN(n12406) );
  OAI211_X1 U15510 ( .C1(n12450), .C2(n12408), .A(n12407), .B(n12406), .ZN(
        n13528) );
  AOI22_X1 U15511 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12383), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15512 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12730), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15513 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11898), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15514 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12409) );
  NAND4_X1 U15515 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12409), .ZN(
        n12425) );
  INV_X1 U15516 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12418) );
  INV_X1 U15517 ( .A(n12413), .ZN(n12417) );
  INV_X1 U15518 ( .A(n12414), .ZN(n12416) );
  INV_X1 U15519 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12415) );
  OAI22_X1 U15520 ( .A1(n12418), .A2(n12417), .B1(n12416), .B2(n12415), .ZN(
        n12419) );
  INV_X1 U15521 ( .A(n12419), .ZN(n12423) );
  AOI22_X1 U15522 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15523 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15524 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12737), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12420) );
  NAND4_X1 U15525 ( .A1(n12423), .A2(n12422), .A3(n12421), .A4(n12420), .ZN(
        n12424) );
  NOR2_X1 U15526 ( .A1(n12425), .A2(n12424), .ZN(n13791) );
  OR2_X1 U15527 ( .A1(n12281), .A2(n13791), .ZN(n12427) );
  AOI22_X1 U15528 ( .A1(n12443), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12426) );
  AND2_X1 U15529 ( .A1(n12427), .A2(n12426), .ZN(n12429) );
  NAND2_X1 U15530 ( .A1(n12459), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12428) );
  INV_X1 U15531 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U15532 ( .A1(n12443), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12430) );
  OAI21_X1 U15533 ( .B1(n12450), .B2(n19890), .A(n12430), .ZN(n13804) );
  INV_X1 U15534 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15535 ( .A1(n12443), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12431) );
  OAI21_X1 U15536 ( .B1(n12450), .B2(n12432), .A(n12431), .ZN(n13901) );
  AND2_X2 U15537 ( .A1(n13802), .A2(n13901), .ZN(n13934) );
  INV_X1 U15538 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19893) );
  AOI22_X1 U15539 ( .A1(n12443), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12433) );
  OAI21_X1 U15540 ( .B1(n12450), .B2(n19893), .A(n12433), .ZN(n13933) );
  NAND2_X1 U15541 ( .A1(n13934), .A2(n13933), .ZN(n13935) );
  INV_X1 U15542 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U15543 ( .A1(n12443), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12434) );
  OAI21_X1 U15544 ( .B1(n12450), .B2(n15005), .A(n12434), .ZN(n14877) );
  INV_X1 U15545 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19896) );
  AOI22_X1 U15546 ( .A1(n12443), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12435) );
  OAI21_X1 U15547 ( .B1(n12450), .B2(n19896), .A(n12435), .ZN(n12436) );
  INV_X1 U15548 ( .A(n12436), .ZN(n14868) );
  INV_X1 U15549 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15550 ( .A1(n12443), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12437) );
  OAI21_X1 U15551 ( .B1(n12450), .B2(n12438), .A(n12437), .ZN(n12439) );
  INV_X1 U15552 ( .A(n12439), .ZN(n14694) );
  INV_X1 U15553 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20948) );
  AOI22_X1 U15554 ( .A1(n12443), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12440) );
  OAI21_X1 U15555 ( .B1(n12450), .B2(n20948), .A(n12440), .ZN(n14852) );
  AND2_X2 U15556 ( .A1(n14853), .A2(n14852), .ZN(n15179) );
  INV_X1 U15557 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n13979) );
  AOI22_X1 U15558 ( .A1(n12443), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12441) );
  OAI21_X1 U15559 ( .B1(n12450), .B2(n13979), .A(n12441), .ZN(n15180) );
  AND2_X2 U15560 ( .A1(n15179), .A2(n15180), .ZN(n15182) );
  INV_X1 U15561 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U15562 ( .A1(n12443), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12442) );
  OAI21_X1 U15563 ( .B1(n12450), .B2(n19901), .A(n12442), .ZN(n14843) );
  NAND2_X1 U15564 ( .A1(n12459), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15565 ( .A1(n12443), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12444) );
  AND2_X1 U15566 ( .A1(n12445), .A2(n12444), .ZN(n14833) );
  NAND2_X1 U15567 ( .A1(n12459), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15568 ( .A1(n12443), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12446) );
  INV_X1 U15569 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15570 ( .A1(n12443), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12448) );
  OAI21_X1 U15571 ( .B1(n12450), .B2(n12449), .A(n12448), .ZN(n14819) );
  NAND2_X1 U15572 ( .A1(n12459), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15573 ( .A1(n12443), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12451) );
  AND2_X1 U15574 ( .A1(n12452), .A2(n12451), .ZN(n14811) );
  INV_X1 U15575 ( .A(n12453), .ZN(n14810) );
  NAND2_X1 U15576 ( .A1(n12459), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15577 ( .A1(n12443), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12454) );
  AND2_X1 U15578 ( .A1(n12455), .A2(n12454), .ZN(n12972) );
  OR2_X2 U15579 ( .A1(n14810), .A2(n12972), .ZN(n12970) );
  NAND2_X1 U15580 ( .A1(n12459), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15581 ( .A1(n12443), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12293), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12456) );
  AND2_X1 U15582 ( .A1(n12457), .A2(n12456), .ZN(n12926) );
  NOR2_X2 U15583 ( .A1(n12970), .A2(n12926), .ZN(n12462) );
  AOI222_X1 U15584 ( .A1(n12459), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12458), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12443), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n12460) );
  INV_X1 U15585 ( .A(n12460), .ZN(n12461) );
  NAND2_X1 U15586 ( .A1(n12162), .A2(n12973), .ZN(n12463) );
  AND2_X1 U15587 ( .A1(n12465), .A2(n12464), .ZN(n16442) );
  INV_X1 U15588 ( .A(n16442), .ZN(n12466) );
  OAI21_X1 U15589 ( .B1(n11776), .B2(n16443), .A(n12466), .ZN(n12467) );
  NAND2_X1 U15590 ( .A1(n19103), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n13988) );
  INV_X1 U15591 ( .A(n13988), .ZN(n12477) );
  INV_X1 U15592 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12473) );
  OAI22_X1 U15593 ( .A1(n15259), .A2(n12469), .B1(n13069), .B2(n12468), .ZN(
        n16415) );
  NAND3_X1 U15594 ( .A1(n15330), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n16415), .ZN(n16403) );
  NAND2_X1 U15595 ( .A1(n15286), .A2(n12472), .ZN(n15231) );
  NOR3_X1 U15596 ( .A1(n12473), .A2(n15207), .A3(n15231), .ZN(n15195) );
  NAND2_X1 U15597 ( .A1(n15184), .A2(n15195), .ZN(n15169) );
  INV_X1 U15598 ( .A(n15169), .ZN(n12474) );
  NAND2_X1 U15599 ( .A1(n15140), .A2(n15153), .ZN(n15130) );
  INV_X1 U15600 ( .A(n15104), .ZN(n12475) );
  NOR2_X1 U15601 ( .A1(n15130), .A2(n12475), .ZN(n15105) );
  INV_X1 U15602 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U15603 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12481) );
  AOI22_X1 U15604 ( .A1(n12574), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n12479) );
  INV_X1 U15605 ( .A(n12533), .ZN(n12588) );
  NAND2_X1 U15606 ( .A1(n12588), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12478) );
  AND2_X1 U15607 ( .A1(n12479), .A2(n12478), .ZN(n12480) );
  NAND2_X1 U15608 ( .A1(n12481), .A2(n12480), .ZN(n13794) );
  AOI22_X1 U15609 ( .A1(n12574), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12482) );
  OAI21_X1 U15610 ( .B1(n12533), .B2(n20874), .A(n12482), .ZN(n12483) );
  AOI21_X1 U15611 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21178), .A(
        n12483), .ZN(n13545) );
  NAND2_X1 U15612 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12488) );
  NAND2_X1 U15613 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12485) );
  NAND2_X1 U15614 ( .A1(n12574), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12484) );
  OAI211_X1 U15615 ( .C1(n12533), .C2(n13314), .A(n12485), .B(n12484), .ZN(
        n12486) );
  INV_X1 U15616 ( .A(n12486), .ZN(n12487) );
  NAND2_X1 U15617 ( .A1(n12488), .A2(n12487), .ZN(n13312) );
  INV_X1 U15618 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n20895) );
  NAND2_X1 U15619 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12490) );
  NAND2_X1 U15620 ( .A1(n12574), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12489) );
  OAI211_X1 U15621 ( .C1(n12533), .C2(n20895), .A(n12490), .B(n12489), .ZN(
        n12492) );
  AOI21_X1 U15622 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n12492), .ZN(n13266) );
  INV_X1 U15623 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12495) );
  NAND2_X1 U15624 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12494) );
  NAND2_X1 U15625 ( .A1(n12574), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12493) );
  OAI211_X1 U15626 ( .C1(n12533), .C2(n12495), .A(n12494), .B(n12493), .ZN(
        n12496) );
  AOI21_X1 U15627 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12496), .ZN(n13167) );
  INV_X1 U15628 ( .A(n12498), .ZN(n12499) );
  OR2_X1 U15629 ( .A1(n12500), .A2(n12499), .ZN(n12501) );
  NAND2_X1 U15630 ( .A1(n12502), .A2(n12501), .ZN(n13168) );
  NAND2_X1 U15631 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12504) );
  AOI22_X1 U15632 ( .A1(n12574), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12503) );
  OAI211_X1 U15633 ( .C1(n13213), .C2(n12533), .A(n12504), .B(n12503), .ZN(
        n13212) );
  INV_X1 U15634 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12507) );
  NAND2_X1 U15635 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12506) );
  NAND2_X1 U15636 ( .A1(n12574), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12505) );
  OAI211_X1 U15637 ( .C1(n12533), .C2(n12507), .A(n12506), .B(n12505), .ZN(
        n12508) );
  AOI21_X1 U15638 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12508), .ZN(n13390) );
  NAND2_X1 U15639 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12511) );
  NAND2_X1 U15640 ( .A1(n12574), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12510) );
  OAI211_X1 U15641 ( .C1(n12533), .C2(n12512), .A(n12511), .B(n12510), .ZN(
        n12513) );
  AOI21_X1 U15642 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12513), .ZN(n13398) );
  NOR2_X2 U15643 ( .A1(n13397), .A2(n13398), .ZN(n13558) );
  INV_X1 U15644 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12516) );
  NAND2_X1 U15645 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12515) );
  AOI22_X1 U15646 ( .A1(n12574), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12514) );
  OAI211_X1 U15647 ( .C1(n12516), .C2(n12533), .A(n12515), .B(n12514), .ZN(
        n13557) );
  NAND2_X1 U15648 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12518) );
  NAND2_X1 U15649 ( .A1(n12574), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12517) );
  OAI211_X1 U15650 ( .C1(n12533), .C2(n13514), .A(n12518), .B(n12517), .ZN(
        n12519) );
  AOI21_X1 U15651 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12519), .ZN(n13512) );
  INV_X1 U15652 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12522) );
  NAND2_X1 U15653 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U15654 ( .A1(n12574), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12520) );
  OAI211_X1 U15655 ( .C1(n12533), .C2(n12522), .A(n12521), .B(n12520), .ZN(
        n12523) );
  AOI21_X1 U15656 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12523), .ZN(n13584) );
  NAND2_X1 U15657 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12525) );
  AOI22_X1 U15658 ( .A1(n12574), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12524) );
  OAI211_X1 U15659 ( .C1(n12526), .C2(n12533), .A(n12525), .B(n12524), .ZN(
        n13525) );
  NOR2_X2 U15660 ( .A1(n13545), .A2(n13544), .ZN(n13793) );
  NAND2_X1 U15661 ( .A1(n13794), .A2(n13793), .ZN(n13849) );
  NAND2_X1 U15662 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U15663 ( .A1(n12574), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12527) );
  OAI211_X1 U15664 ( .C1(n12533), .C2(n11662), .A(n12528), .B(n12527), .ZN(
        n12529) );
  AOI21_X1 U15665 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12529), .ZN(n13848) );
  NAND2_X1 U15666 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12531) );
  AOI22_X1 U15667 ( .A1(n12574), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12530) );
  OAI211_X1 U15668 ( .C1(n12533), .C2(n12532), .A(n12531), .B(n12530), .ZN(
        n13827) );
  NAND2_X1 U15669 ( .A1(n13851), .A2(n13827), .ZN(n13929) );
  NAND2_X1 U15670 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U15671 ( .A1(n12574), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12534) );
  OAI211_X1 U15672 ( .C1(n12533), .C2(n12536), .A(n12535), .B(n12534), .ZN(
        n12537) );
  AOI21_X1 U15673 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12537), .ZN(n13928) );
  INV_X1 U15674 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12540) );
  NAND2_X1 U15675 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12539) );
  NAND2_X1 U15676 ( .A1(n12574), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12538) );
  OAI211_X1 U15677 ( .C1(n12533), .C2(n12540), .A(n12539), .B(n12538), .ZN(
        n12541) );
  AOI21_X1 U15678 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12541), .ZN(n14791) );
  NAND2_X1 U15679 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12543) );
  NAND2_X1 U15680 ( .A1(n12574), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12542) );
  OAI211_X1 U15681 ( .C1(n12533), .C2(n12544), .A(n12543), .B(n12542), .ZN(
        n12545) );
  AOI21_X1 U15682 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12545), .ZN(n14786) );
  NAND2_X1 U15683 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U15684 ( .A1(n12574), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12546) );
  OAI211_X1 U15685 ( .C1(n12533), .C2(n12548), .A(n12547), .B(n12546), .ZN(
        n12549) );
  AOI21_X1 U15686 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12549), .ZN(n14693) );
  NAND2_X1 U15687 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12553) );
  AOI22_X1 U15688 ( .A1(n12574), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12551) );
  NAND2_X1 U15689 ( .A1(n12588), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12550) );
  AND2_X1 U15690 ( .A1(n12551), .A2(n12550), .ZN(n12552) );
  NAND2_X1 U15691 ( .A1(n12553), .A2(n12552), .ZN(n14772) );
  AND2_X2 U15692 ( .A1(n14773), .A2(n14772), .ZN(n14775) );
  NAND2_X1 U15693 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12557) );
  AOI22_X1 U15694 ( .A1(n12574), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12555) );
  NAND2_X1 U15695 ( .A1(n12588), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12554) );
  AND2_X1 U15696 ( .A1(n12555), .A2(n12554), .ZN(n12556) );
  NAND2_X1 U15697 ( .A1(n12557), .A2(n12556), .ZN(n13977) );
  AND2_X2 U15698 ( .A1(n14775), .A2(n13977), .ZN(n14761) );
  NAND2_X1 U15699 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12561) );
  AOI22_X1 U15700 ( .A1(n12574), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12559) );
  NAND2_X1 U15701 ( .A1(n12588), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12558) );
  AND2_X1 U15702 ( .A1(n12559), .A2(n12558), .ZN(n12560) );
  NAND2_X1 U15703 ( .A1(n12561), .A2(n12560), .ZN(n14760) );
  NAND2_X1 U15704 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12563) );
  NAND2_X1 U15705 ( .A1(n12574), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12562) );
  OAI211_X1 U15706 ( .C1(n12533), .C2(n12564), .A(n12563), .B(n12562), .ZN(
        n12565) );
  AOI21_X1 U15707 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12565), .ZN(n14750) );
  OR2_X2 U15708 ( .A1(n14759), .A2(n14750), .ZN(n14752) );
  INV_X1 U15709 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12568) );
  NAND2_X1 U15710 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U15711 ( .A1(n12574), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12566) );
  OAI211_X1 U15712 ( .C1(n12533), .C2(n12568), .A(n12567), .B(n12566), .ZN(
        n12569) );
  AOI21_X1 U15713 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12569), .ZN(n14744) );
  NAND2_X1 U15714 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12573) );
  AOI22_X1 U15715 ( .A1(n12574), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12571) );
  NAND2_X1 U15716 ( .A1(n12588), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12570) );
  AND2_X1 U15717 ( .A1(n12571), .A2(n12570), .ZN(n12572) );
  NAND2_X1 U15718 ( .A1(n12573), .A2(n12572), .ZN(n14731) );
  NAND2_X1 U15719 ( .A1(n21178), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12578) );
  AOI22_X1 U15720 ( .A1(n12574), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12576) );
  NAND2_X1 U15721 ( .A1(n12588), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12575) );
  AND2_X1 U15722 ( .A1(n12576), .A2(n12575), .ZN(n12577) );
  NAND2_X1 U15723 ( .A1(n12578), .A2(n12577), .ZN(n14726) );
  NAND2_X1 U15724 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12580) );
  NAND2_X1 U15725 ( .A1(n12574), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12579) );
  OAI211_X1 U15726 ( .C1(n12533), .C2(n12581), .A(n12580), .B(n12579), .ZN(
        n12582) );
  AOI21_X1 U15727 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12582), .ZN(n12979) );
  NAND2_X1 U15728 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12584) );
  NAND2_X1 U15729 ( .A1(n12574), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12583) );
  OAI211_X1 U15730 ( .C1(n12533), .C2(n12585), .A(n12584), .B(n12583), .ZN(
        n12586) );
  AOI21_X1 U15731 ( .B1(n21178), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12586), .ZN(n14011) );
  NAND2_X1 U15732 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U15733 ( .A1(n12574), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12590) );
  NAND2_X1 U15734 ( .A1(n12588), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12589) );
  OAI211_X1 U15735 ( .C1(n11774), .C2(n12937), .A(n12590), .B(n12589), .ZN(
        n12591) );
  NAND2_X1 U15736 ( .A1(n12593), .A2(n11754), .ZN(n12594) );
  NAND2_X1 U15737 ( .A1(n16443), .A2(n12594), .ZN(n13876) );
  NAND2_X1 U15738 ( .A1(n13876), .A2(n11776), .ZN(n12596) );
  NAND2_X1 U15739 ( .A1(n12596), .A2(n12595), .ZN(n12597) );
  NAND2_X1 U15740 ( .A1(n11845), .A2(n12619), .ZN(n12604) );
  NAND2_X1 U15741 ( .A1(n12928), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12600) );
  NAND2_X1 U15742 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19629) );
  NAND2_X1 U15743 ( .A1(n19629), .A2(n19940), .ZN(n12602) );
  NAND2_X1 U15744 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19771) );
  INV_X1 U15745 ( .A(n19771), .ZN(n12601) );
  NAND2_X1 U15746 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12601), .ZN(
        n19274) );
  AND2_X1 U15747 ( .A1(n12602), .A2(n19274), .ZN(n19412) );
  AOI22_X1 U15748 ( .A1(n12622), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19928), .B2(n19412), .ZN(n12603) );
  INV_X1 U15749 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12606) );
  NAND2_X1 U15750 ( .A1(n12622), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12608) );
  NAND2_X1 U15751 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19949), .ZN(
        n19564) );
  NAND2_X1 U15752 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19958), .ZN(
        n19597) );
  AND2_X1 U15753 ( .A1(n19564), .A2(n19597), .ZN(n19411) );
  INV_X1 U15754 ( .A(n19411), .ZN(n12607) );
  NAND2_X1 U15755 ( .A1(n19928), .A2(n12607), .ZN(n19600) );
  NAND2_X1 U15756 ( .A1(n12608), .A2(n19600), .ZN(n12609) );
  INV_X1 U15757 ( .A(n12619), .ZN(n16471) );
  AOI22_X1 U15758 ( .A1(n12622), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19928), .B2(n19958), .ZN(n12610) );
  XNOR2_X1 U15759 ( .A(n13612), .B(n12613), .ZN(n13076) );
  NAND2_X1 U15760 ( .A1(n13075), .A2(n13076), .ZN(n13078) );
  NAND2_X1 U15761 ( .A1(n13084), .A2(n12613), .ZN(n12614) );
  INV_X1 U15762 ( .A(n12615), .ZN(n12616) );
  NAND2_X1 U15763 ( .A1(n12617), .A2(n12616), .ZN(n12618) );
  NAND2_X1 U15764 ( .A1(n13120), .A2(n12619), .ZN(n12624) );
  NAND2_X1 U15765 ( .A1(n19274), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12620) );
  NOR2_X1 U15766 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19771), .ZN(
        n19512) );
  NAND2_X1 U15767 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19512), .ZN(
        n19506) );
  NAND2_X1 U15768 ( .A1(n12620), .A2(n19506), .ZN(n12621) );
  AOI22_X1 U15769 ( .A1(n12622), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19928), .B2(n12621), .ZN(n12623) );
  NAND2_X1 U15770 ( .A1(n12628), .A2(n12625), .ZN(n13162) );
  NAND2_X1 U15771 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12928), .ZN(
        n12627) );
  AND2_X1 U15772 ( .A1(n12628), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12629) );
  NAND2_X2 U15773 ( .A1(n12630), .A2(n13163), .ZN(n13270) );
  INV_X1 U15774 ( .A(n13791), .ZN(n12636) );
  INV_X1 U15775 ( .A(n12632), .ZN(n13548) );
  OR2_X1 U15776 ( .A1(n13555), .A2(n13552), .ZN(n13511) );
  NAND2_X1 U15777 ( .A1(n13589), .A2(n13588), .ZN(n12633) );
  NOR2_X1 U15778 ( .A1(n12634), .A2(n13523), .ZN(n12635) );
  AND2_X1 U15779 ( .A1(n12635), .A2(n13394), .ZN(n13546) );
  AOI22_X1 U15780 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U15781 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U15782 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12639) );
  AOI22_X1 U15783 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12638) );
  NAND4_X1 U15784 ( .A1(n12641), .A2(n12640), .A3(n12639), .A4(n12638), .ZN(
        n12647) );
  AOI22_X1 U15785 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U15786 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12644) );
  AOI22_X1 U15787 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U15788 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12642) );
  NAND4_X1 U15789 ( .A1(n12645), .A2(n12644), .A3(n12643), .A4(n12642), .ZN(
        n12646) );
  NAND2_X1 U15790 ( .A1(n13801), .A2(n13800), .ZN(n13799) );
  AOI22_X1 U15791 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12383), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15792 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12730), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15793 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11633), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15794 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12648) );
  NAND4_X1 U15795 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        n12657) );
  AOI22_X1 U15796 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15797 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U15798 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15799 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12737), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12652) );
  NAND4_X1 U15800 ( .A1(n12655), .A2(n12654), .A3(n12653), .A4(n12652), .ZN(
        n12656) );
  NOR2_X1 U15801 ( .A1(n12657), .A2(n12656), .ZN(n13831) );
  NAND2_X1 U15802 ( .A1(n12659), .A2(n12658), .ZN(n13926) );
  AOI22_X1 U15803 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12383), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15804 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12730), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U15805 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11633), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15806 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12660) );
  NAND4_X1 U15807 ( .A1(n12663), .A2(n12662), .A3(n12661), .A4(n12660), .ZN(
        n12669) );
  AOI22_X1 U15808 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U15809 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U15810 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15811 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12737), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12664) );
  NAND4_X1 U15812 ( .A1(n12667), .A2(n12666), .A3(n12665), .A4(n12664), .ZN(
        n12668) );
  NOR2_X1 U15813 ( .A1(n12669), .A2(n12668), .ZN(n13927) );
  OR2_X2 U15814 ( .A1(n13926), .A2(n13927), .ZN(n14796) );
  AOI22_X1 U15815 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15816 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15817 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U15818 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12670) );
  NAND4_X1 U15819 ( .A1(n12673), .A2(n12672), .A3(n12671), .A4(n12670), .ZN(
        n12679) );
  AOI22_X1 U15820 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12677) );
  AOI22_X1 U15821 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U15822 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U15823 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12674) );
  NAND4_X1 U15824 ( .A1(n12677), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        n12678) );
  NOR2_X1 U15825 ( .A1(n12679), .A2(n12678), .ZN(n14797) );
  AOI22_X1 U15826 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U15827 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15828 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15829 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12680) );
  NAND4_X1 U15830 ( .A1(n12683), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12689) );
  AOI22_X1 U15831 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U15832 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15833 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U15834 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12684) );
  NAND4_X1 U15835 ( .A1(n12687), .A2(n12686), .A3(n12685), .A4(n12684), .ZN(
        n12688) );
  OR2_X1 U15836 ( .A1(n12689), .A2(n12688), .ZN(n14784) );
  AOI22_X1 U15837 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U15838 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U15839 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U15840 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12690) );
  NAND4_X1 U15841 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12699) );
  AOI22_X1 U15842 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U15843 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15844 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U15845 ( .A1(n12737), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12694) );
  NAND4_X1 U15846 ( .A1(n12697), .A2(n12696), .A3(n12695), .A4(n12694), .ZN(
        n12698) );
  OR2_X1 U15847 ( .A1(n12699), .A2(n12698), .ZN(n14780) );
  AOI22_X1 U15848 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12383), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15849 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12730), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15850 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11633), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15851 ( .A1(n12729), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12700) );
  NAND4_X1 U15852 ( .A1(n12703), .A2(n12702), .A3(n12701), .A4(n12700), .ZN(
        n12709) );
  AOI22_X1 U15853 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12414), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15854 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11586), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U15855 ( .A1(n11904), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12735), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15856 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12737), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12704) );
  NAND4_X1 U15857 ( .A1(n12707), .A2(n12706), .A3(n12705), .A4(n12704), .ZN(
        n12708) );
  NOR2_X1 U15858 ( .A1(n12709), .A2(n12708), .ZN(n14771) );
  AOI22_X1 U15859 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U15860 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12718) );
  INV_X2 U15861 ( .A(n13185), .ZN(n13871) );
  AOI22_X1 U15862 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12717) );
  INV_X1 U15863 ( .A(n12902), .ZN(n12891) );
  INV_X1 U15864 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U15865 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12713) );
  INV_X1 U15866 ( .A(n12710), .ZN(n12712) );
  NAND2_X1 U15867 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U15868 ( .A1(n12712), .A2(n12711), .ZN(n12892) );
  OAI211_X1 U15869 ( .C1(n12891), .C2(n12714), .A(n12713), .B(n12892), .ZN(
        n12715) );
  INV_X1 U15870 ( .A(n12715), .ZN(n12716) );
  NAND4_X1 U15871 ( .A1(n12719), .A2(n12718), .A3(n12717), .A4(n12716), .ZN(
        n12728) );
  AOI22_X1 U15872 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15873 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15874 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12724) );
  INV_X1 U15875 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12721) );
  NAND2_X1 U15876 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12720) );
  OAI211_X1 U15877 ( .C1(n12891), .C2(n12721), .A(n12720), .B(n12871), .ZN(
        n12722) );
  INV_X1 U15878 ( .A(n12722), .ZN(n12723) );
  NAND4_X1 U15879 ( .A1(n12726), .A2(n12725), .A3(n12724), .A4(n12723), .ZN(
        n12727) );
  NAND2_X1 U15880 ( .A1(n15585), .A2(n12763), .ZN(n12744) );
  AOI22_X1 U15881 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12383), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U15882 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12729), .B1(
        n11634), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15883 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U15884 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12414), .B1(
        n11898), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12731) );
  NAND4_X1 U15885 ( .A1(n12734), .A2(n12733), .A3(n12732), .A4(n12731), .ZN(
        n12743) );
  AOI22_X1 U15886 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11899), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15887 ( .A1(n12736), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12735), .ZN(n12740) );
  AOI22_X1 U15888 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12737), .B1(
        n11904), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U15889 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11586), .B1(
        n11585), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12738) );
  NAND4_X1 U15890 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12742) );
  OR2_X1 U15891 ( .A1(n12743), .A2(n12742), .ZN(n12764) );
  XNOR2_X1 U15892 ( .A(n12744), .B(n12764), .ZN(n12769) );
  XNOR2_X2 U15893 ( .A(n12745), .B(n12769), .ZN(n14765) );
  INV_X1 U15894 ( .A(n12763), .ZN(n12767) );
  NOR2_X1 U15895 ( .A1(n15585), .A2(n12767), .ZN(n14764) );
  AOI22_X1 U15896 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U15897 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U15898 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U15899 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12747) );
  OAI211_X1 U15900 ( .C1(n12891), .C2(n12748), .A(n12747), .B(n12892), .ZN(
        n12749) );
  INV_X1 U15901 ( .A(n12749), .ZN(n12750) );
  NAND4_X1 U15902 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12762) );
  AOI22_X1 U15903 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15904 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15905 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12758) );
  NAND2_X1 U15906 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12754) );
  OAI211_X1 U15907 ( .C1(n12891), .C2(n12755), .A(n12754), .B(n12871), .ZN(
        n12756) );
  INV_X1 U15908 ( .A(n12756), .ZN(n12757) );
  NAND4_X1 U15909 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  NAND2_X1 U15910 ( .A1(n12762), .A2(n12761), .ZN(n12771) );
  NAND2_X1 U15911 ( .A1(n12764), .A2(n12763), .ZN(n12772) );
  XOR2_X1 U15912 ( .A(n12771), .B(n12772), .Z(n12765) );
  NAND2_X1 U15913 ( .A1(n12765), .A2(n12839), .ZN(n14755) );
  INV_X1 U15914 ( .A(n12771), .ZN(n12766) );
  NAND2_X1 U15915 ( .A1(n11776), .A2(n12766), .ZN(n14758) );
  NOR2_X1 U15916 ( .A1(n14758), .A2(n12767), .ZN(n12768) );
  NOR2_X1 U15917 ( .A1(n12772), .A2(n12771), .ZN(n12789) );
  AOI22_X1 U15918 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U15919 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U15920 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12777) );
  INV_X1 U15921 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12774) );
  NAND2_X1 U15922 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12773) );
  OAI211_X1 U15923 ( .C1(n12891), .C2(n12774), .A(n12773), .B(n12892), .ZN(
        n12775) );
  INV_X1 U15924 ( .A(n12775), .ZN(n12776) );
  NAND4_X1 U15925 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n12788) );
  AOI22_X1 U15926 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U15927 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U15928 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12784) );
  INV_X1 U15929 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12781) );
  NAND2_X1 U15930 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12780) );
  OAI211_X1 U15931 ( .C1(n12891), .C2(n12781), .A(n12780), .B(n12871), .ZN(
        n12782) );
  INV_X1 U15932 ( .A(n12782), .ZN(n12783) );
  NAND4_X1 U15933 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n12787) );
  NAND2_X1 U15934 ( .A1(n12789), .A2(n12791), .ZN(n12813) );
  OAI211_X1 U15935 ( .C1(n12789), .C2(n12791), .A(n12813), .B(n12839), .ZN(
        n12793) );
  INV_X1 U15936 ( .A(n12793), .ZN(n12790) );
  INV_X1 U15937 ( .A(n12791), .ZN(n12792) );
  NOR2_X1 U15938 ( .A1(n15585), .A2(n12792), .ZN(n14748) );
  NAND2_X1 U15939 ( .A1(n14749), .A2(n14748), .ZN(n14747) );
  NAND2_X1 U15940 ( .A1(n14747), .A2(n10265), .ZN(n12817) );
  AOI22_X1 U15941 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U15942 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U15943 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U15944 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12795) );
  OAI211_X1 U15945 ( .C1(n12891), .C2(n12796), .A(n12795), .B(n12892), .ZN(
        n12797) );
  INV_X1 U15946 ( .A(n12797), .ZN(n12798) );
  NAND4_X1 U15947 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12811) );
  AOI22_X1 U15948 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U15949 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U15950 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U15951 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12803) );
  OAI211_X1 U15952 ( .C1(n12891), .C2(n12804), .A(n12803), .B(n12871), .ZN(
        n12805) );
  INV_X1 U15953 ( .A(n12805), .ZN(n12806) );
  NAND4_X1 U15954 ( .A1(n12809), .A2(n12808), .A3(n12807), .A4(n12806), .ZN(
        n12810) );
  NAND2_X1 U15955 ( .A1(n12811), .A2(n12810), .ZN(n12815) );
  AOI21_X1 U15956 ( .B1(n12813), .B2(n12815), .A(n12812), .ZN(n12814) );
  INV_X1 U15957 ( .A(n12815), .ZN(n12816) );
  NAND2_X1 U15958 ( .A1(n11776), .A2(n12816), .ZN(n14740) );
  INV_X1 U15959 ( .A(n12838), .ZN(n12840) );
  AOI22_X1 U15960 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U15961 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U15962 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12824) );
  INV_X1 U15963 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12821) );
  NAND2_X1 U15964 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12820) );
  OAI211_X1 U15965 ( .C1(n12819), .C2(n12821), .A(n12892), .B(n12820), .ZN(
        n12822) );
  INV_X1 U15966 ( .A(n12822), .ZN(n12823) );
  NAND4_X1 U15967 ( .A1(n12826), .A2(n12825), .A3(n12824), .A4(n12823), .ZN(
        n12836) );
  AOI22_X1 U15968 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U15969 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U15970 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9750), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12832) );
  INV_X1 U15971 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U15972 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12827) );
  OAI211_X1 U15973 ( .C1(n12829), .C2(n12828), .A(n12871), .B(n12827), .ZN(
        n12830) );
  INV_X1 U15974 ( .A(n12830), .ZN(n12831) );
  NAND4_X1 U15975 ( .A1(n12834), .A2(n12833), .A3(n12832), .A4(n12831), .ZN(
        n12835) );
  NAND2_X1 U15976 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  INV_X1 U15977 ( .A(n12837), .ZN(n12844) );
  OR2_X1 U15978 ( .A1(n12838), .A2(n12837), .ZN(n14722) );
  OAI211_X1 U15979 ( .C1(n12840), .C2(n12844), .A(n14722), .B(n12839), .ZN(
        n12841) );
  INV_X1 U15980 ( .A(n12861), .ZN(n14723) );
  NAND2_X1 U15981 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  NAND2_X1 U15982 ( .A1(n14723), .A2(n12843), .ZN(n14736) );
  NAND2_X1 U15983 ( .A1(n11776), .A2(n12844), .ZN(n14735) );
  NOR2_X2 U15984 ( .A1(n14736), .A2(n14735), .ZN(n14734) );
  AOI22_X1 U15985 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U15986 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U15987 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12849) );
  NAND2_X1 U15988 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12845) );
  OAI211_X1 U15989 ( .C1(n12891), .C2(n12846), .A(n12845), .B(n12892), .ZN(
        n12847) );
  INV_X1 U15990 ( .A(n12847), .ZN(n12848) );
  NAND4_X1 U15991 ( .A1(n12851), .A2(n12850), .A3(n12849), .A4(n12848), .ZN(
        n12860) );
  AOI22_X1 U15992 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U15993 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12857) );
  AOI22_X1 U15994 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12856) );
  NAND2_X1 U15995 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12852) );
  OAI211_X1 U15996 ( .C1(n12891), .C2(n12853), .A(n12852), .B(n12871), .ZN(
        n12854) );
  INV_X1 U15997 ( .A(n12854), .ZN(n12855) );
  NAND4_X1 U15998 ( .A1(n12858), .A2(n12857), .A3(n12856), .A4(n12855), .ZN(
        n12859) );
  AND2_X1 U15999 ( .A1(n12860), .A2(n12859), .ZN(n14724) );
  OAI21_X1 U16000 ( .B1(n14734), .B2(n12861), .A(n14724), .ZN(n14719) );
  NAND2_X1 U16001 ( .A1(n15585), .A2(n14724), .ZN(n12862) );
  NOR2_X1 U16002 ( .A1(n14722), .A2(n12862), .ZN(n12882) );
  AOI22_X1 U16003 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U16004 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11531), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U16005 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12867) );
  NAND2_X1 U16006 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12863) );
  OAI211_X1 U16007 ( .C1(n12891), .C2(n12864), .A(n12863), .B(n12892), .ZN(
        n12865) );
  INV_X1 U16008 ( .A(n12865), .ZN(n12866) );
  NAND4_X1 U16009 ( .A1(n12869), .A2(n12868), .A3(n12867), .A4(n12866), .ZN(
        n12880) );
  AOI22_X1 U16010 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U16011 ( .A1(n12870), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11531), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12877) );
  AOI22_X1 U16012 ( .A1(n12802), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12876) );
  NAND2_X1 U16013 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12872) );
  OAI211_X1 U16014 ( .C1(n12891), .C2(n12873), .A(n12872), .B(n12871), .ZN(
        n12874) );
  INV_X1 U16015 ( .A(n12874), .ZN(n12875) );
  NAND4_X1 U16016 ( .A1(n12878), .A2(n12877), .A3(n12876), .A4(n12875), .ZN(
        n12879) );
  AND2_X1 U16017 ( .A1(n12880), .A2(n12879), .ZN(n12881) );
  NAND2_X1 U16018 ( .A1(n12882), .A2(n12881), .ZN(n12883) );
  OAI21_X1 U16019 ( .B1(n12882), .B2(n12881), .A(n12883), .ZN(n14718) );
  NOR2_X1 U16020 ( .A1(n14719), .A2(n14718), .ZN(n14717) );
  INV_X1 U16021 ( .A(n12883), .ZN(n12884) );
  NOR2_X1 U16022 ( .A1(n14717), .A2(n12884), .ZN(n12911) );
  AOI22_X1 U16023 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U16024 ( .A1(n11531), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13871), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12885) );
  NAND2_X1 U16025 ( .A1(n12886), .A2(n12885), .ZN(n12909) );
  INV_X1 U16026 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16027 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12802), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12889) );
  AOI21_X1 U16028 ( .B1(n12887), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n12892), .ZN(n12888) );
  OAI211_X1 U16029 ( .C1(n12891), .C2(n12890), .A(n12889), .B(n12888), .ZN(
        n12908) );
  INV_X1 U16030 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12893) );
  OAI21_X1 U16031 ( .B1(n12894), .B2(n12893), .A(n12892), .ZN(n12899) );
  INV_X1 U16032 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12896) );
  INV_X1 U16033 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12895) );
  OAI22_X1 U16034 ( .A1(n12897), .A2(n12896), .B1(n13185), .B2(n12895), .ZN(
        n12898) );
  AOI211_X1 U16035 ( .C1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(n12802), .A(
        n12899), .B(n12898), .ZN(n12906) );
  AOI22_X1 U16036 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12900), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16037 ( .A1(n12903), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12902), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12904) );
  NAND3_X1 U16038 ( .A1(n12906), .A2(n12905), .A3(n12904), .ZN(n12907) );
  OAI21_X1 U16039 ( .B1(n12909), .B2(n12908), .A(n12907), .ZN(n12910) );
  XNOR2_X1 U16040 ( .A(n12911), .B(n12910), .ZN(n14014) );
  INV_X1 U16041 ( .A(n19838), .ZN(n16479) );
  AND2_X1 U16042 ( .A1(n12246), .A2(n15853), .ZN(n13196) );
  NAND2_X1 U16043 ( .A1(n18951), .A2(n13196), .ZN(n12915) );
  NAND2_X1 U16044 ( .A1(n16449), .A2(n16441), .ZN(n13198) );
  NAND2_X1 U16045 ( .A1(n13198), .A2(n12912), .ZN(n12913) );
  NOR4_X1 U16046 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12920) );
  NOR4_X1 U16047 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12919) );
  NOR4_X1 U16048 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12918) );
  NOR4_X1 U16049 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12917) );
  NAND4_X1 U16050 ( .A1(n12920), .A2(n12919), .A3(n12918), .A4(n12917), .ZN(
        n12925) );
  NOR4_X1 U16051 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12923) );
  NOR4_X1 U16052 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12922) );
  NOR4_X1 U16053 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n12921) );
  NAND4_X1 U16054 ( .A1(n12923), .A2(n12922), .A3(n12921), .A4(n19871), .ZN(
        n12924) );
  AOI22_X1 U16055 ( .A1(n19270), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19268), .ZN(n13530) );
  INV_X1 U16056 ( .A(n13530), .ZN(n13234) );
  INV_X1 U16057 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n19189) );
  OAI22_X1 U16058 ( .A1(n16267), .A2(n16189), .B1(n14836), .B2(n19189), .ZN(
        n12927) );
  AOI21_X1 U16059 ( .B1(n16265), .B2(n13234), .A(n12927), .ZN(n12932) );
  AND2_X1 U16060 ( .A1(n12929), .A2(n12928), .ZN(n12930) );
  AOI22_X1 U16061 ( .A1(n19134), .A2(BUF2_REG_30__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12931) );
  AND2_X1 U16062 ( .A1(n12932), .A2(n12931), .ZN(n12933) );
  OAI21_X1 U16063 ( .B1(n14014), .B2(n19168), .A(n12933), .ZN(P2_U2889) );
  NAND2_X1 U16064 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U16065 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n12945), .ZN(
        n12944) );
  NAND2_X1 U16066 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n12965), .ZN(
        n12966) );
  INV_X1 U16067 ( .A(n12966), .ZN(n12934) );
  AOI21_X1 U16068 ( .B1(n14902), .B2(n12967), .A(n12935), .ZN(n14904) );
  NAND2_X1 U16069 ( .A1(n12935), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12936) );
  INV_X1 U16070 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14684) );
  AOI21_X1 U16071 ( .B1(n12938), .B2(n13980), .A(n12963), .ZN(n13982) );
  INV_X1 U16072 ( .A(n13982), .ZN(n16259) );
  OAI21_X1 U16073 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12960), .A(
        n12938), .ZN(n15784) );
  AOI21_X1 U16074 ( .B1(n9773), .B2(n15006), .A(n12955), .ZN(n15008) );
  INV_X1 U16075 ( .A(n15008), .ZN(n18994) );
  AOI21_X1 U16076 ( .B1(n14705), .B2(n9823), .A(n12954), .ZN(n15028) );
  AOI21_X1 U16077 ( .B1(n19025), .B2(n12950), .A(n12952), .ZN(n19021) );
  AOI21_X1 U16078 ( .B1(n16291), .B2(n12948), .A(n12951), .ZN(n16279) );
  AOI21_X1 U16079 ( .B1(n16308), .B2(n12946), .A(n12949), .ZN(n16292) );
  AOI21_X1 U16080 ( .B1(n16315), .B2(n12944), .A(n12947), .ZN(n16309) );
  AOI21_X1 U16081 ( .B1(n16325), .B2(n12943), .A(n12945), .ZN(n16316) );
  AOI21_X1 U16082 ( .B1(n16339), .B2(n12941), .A(n9761), .ZN(n16326) );
  AOI21_X1 U16083 ( .B1(n13673), .B2(n12940), .A(n12942), .ZN(n13675) );
  OAI22_X1 U16084 ( .A1(n21158), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n13758) );
  INV_X1 U16085 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13761) );
  OAI22_X1 U16086 ( .A1(n21158), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13761), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13757) );
  AND2_X1 U16087 ( .A1(n13758), .A2(n13757), .ZN(n13756) );
  OAI21_X1 U16088 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12940), .ZN(n13819) );
  NAND2_X1 U16089 ( .A1(n13756), .A2(n13819), .ZN(n13644) );
  NOR2_X1 U16090 ( .A1(n13675), .A2(n13644), .ZN(n19107) );
  OAI21_X1 U16091 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12942), .A(
        n12941), .ZN(n19266) );
  NAND2_X1 U16092 ( .A1(n19107), .A2(n19266), .ZN(n13632) );
  NOR2_X1 U16093 ( .A1(n16326), .A2(n13632), .ZN(n19085) );
  OAI21_X1 U16094 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9761), .A(
        n12943), .ZN(n19086) );
  NAND2_X1 U16095 ( .A1(n19085), .A2(n19086), .ZN(n13725) );
  NOR2_X1 U16096 ( .A1(n16316), .A2(n13725), .ZN(n19075) );
  OAI21_X1 U16097 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12945), .A(
        n12944), .ZN(n19076) );
  NAND2_X1 U16098 ( .A1(n19075), .A2(n19076), .ZN(n13656) );
  NOR2_X1 U16099 ( .A1(n16309), .A2(n13656), .ZN(n19063) );
  OAI21_X1 U16100 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12947), .A(
        n12946), .ZN(n19064) );
  NAND2_X1 U16101 ( .A1(n19063), .A2(n19064), .ZN(n13715) );
  NOR2_X1 U16102 ( .A1(n16292), .A2(n13715), .ZN(n19046) );
  OAI21_X1 U16103 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12949), .A(
        n12948), .ZN(n19047) );
  NAND2_X1 U16104 ( .A1(n19046), .A2(n19047), .ZN(n13897) );
  NOR2_X1 U16105 ( .A1(n16279), .A2(n13897), .ZN(n13896) );
  OAI21_X1 U16106 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12951), .A(
        n12950), .ZN(n19039) );
  NAND2_X1 U16107 ( .A1(n13896), .A2(n19039), .ZN(n19020) );
  NOR2_X1 U16108 ( .A1(n19021), .A2(n19020), .ZN(n19009) );
  OAI21_X1 U16109 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12952), .A(
        n9823), .ZN(n19010) );
  AND2_X1 U16110 ( .A1(n19009), .A2(n19010), .ZN(n12953) );
  OAI21_X1 U16111 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12954), .A(
        n9773), .ZN(n19005) );
  NAND2_X1 U16112 ( .A1(n12939), .A2(n19003), .ZN(n18993) );
  NAND2_X1 U16113 ( .A1(n18994), .A2(n18993), .ZN(n18992) );
  INV_X1 U16114 ( .A(n12962), .ZN(n12959) );
  INV_X1 U16115 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12957) );
  INV_X1 U16116 ( .A(n12955), .ZN(n12956) );
  NAND2_X1 U16117 ( .A1(n12957), .A2(n12956), .ZN(n12958) );
  NAND2_X1 U16118 ( .A1(n12959), .A2(n12958), .ZN(n18982) );
  NAND2_X1 U16119 ( .A1(n12939), .A2(n18980), .ZN(n14692) );
  INV_X1 U16120 ( .A(n12960), .ZN(n12961) );
  OAI21_X1 U16121 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12962), .A(
        n12961), .ZN(n14983) );
  NAND2_X1 U16122 ( .A1(n15784), .A2(n15783), .ZN(n15782) );
  NAND2_X1 U16123 ( .A1(n12939), .A2(n15782), .ZN(n16258) );
  NAND2_X1 U16124 ( .A1(n16259), .A2(n16258), .ZN(n16257) );
  OAI21_X1 U16125 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12963), .A(
        n12964), .ZN(n16249) );
  AOI21_X1 U16126 ( .B1(n16227), .B2(n12964), .A(n12965), .ZN(n14940) );
  INV_X1 U16127 ( .A(n14940), .ZN(n16235) );
  OAI21_X1 U16128 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n12965), .A(
        n12966), .ZN(n16222) );
  INV_X1 U16129 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14923) );
  AOI21_X1 U16130 ( .B1(n12966), .B2(n14923), .A(n12968), .ZN(n16207) );
  OAI21_X1 U16131 ( .B1(n12968), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12967), .ZN(n16195) );
  NOR2_X1 U16132 ( .A1(n19108), .A2(n16205), .ZN(n12969) );
  NOR2_X1 U16133 ( .A1(n12969), .A2(n14904), .ZN(n16183) );
  NOR3_X1 U16134 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15855) );
  NAND2_X1 U16135 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15855), .ZN(n19841) );
  AOI211_X1 U16136 ( .C1(n14904), .C2(n12969), .A(n16183), .B(n19841), .ZN(
        n12991) );
  INV_X1 U16137 ( .A(n12970), .ZN(n12971) );
  AOI21_X1 U16138 ( .B1(n12972), .B2(n14810), .A(n12971), .ZN(n15109) );
  NAND2_X1 U16139 ( .A1(n12973), .A2(n19838), .ZN(n13044) );
  INV_X1 U16140 ( .A(n13044), .ZN(n12974) );
  NAND2_X1 U16141 ( .A1(n12162), .A2(n12974), .ZN(n12975) );
  NAND2_X1 U16142 ( .A1(n13043), .A2(n19661), .ZN(n16468) );
  INV_X1 U16143 ( .A(n16468), .ZN(n12976) );
  NAND2_X1 U16144 ( .A1(n18951), .A2(n11774), .ZN(n12981) );
  INV_X1 U16145 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12978) );
  AND2_X1 U16146 ( .A1(n15853), .A2(n19661), .ZN(n12977) );
  NAND2_X1 U16147 ( .A1(n14728), .A2(n12979), .ZN(n12980) );
  NAND2_X1 U16148 ( .A1(n9780), .A2(n12980), .ZN(n15112) );
  NOR2_X1 U16149 ( .A1(n19509), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19504) );
  INV_X1 U16150 ( .A(n19504), .ZN(n12982) );
  NOR2_X1 U16151 ( .A1(n12983), .A2(n12982), .ZN(n16464) );
  INV_X1 U16152 ( .A(n16464), .ZN(n12984) );
  NAND3_X1 U16153 ( .A1(n12984), .A2(n19841), .A3(n19058), .ZN(n12985) );
  INV_X2 U16154 ( .A(n19185), .ZN(n13258) );
  NAND2_X1 U16155 ( .A1(n13258), .A2(n16468), .ZN(n14685) );
  INV_X1 U16156 ( .A(n13179), .ZN(n13180) );
  AOI21_X1 U16157 ( .B1(n19661), .B2(n15853), .A(P2_EBX_REG_31__SCAN_IN), .ZN(
        n12986) );
  NAND2_X1 U16158 ( .A1(n13180), .A2(n12986), .ZN(n12987) );
  AOI22_X1 U16159 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19117), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19122), .ZN(n12988) );
  OAI21_X1 U16160 ( .B1(n14902), .B2(n19024), .A(n12988), .ZN(n12989) );
  NAND2_X1 U16161 ( .A1(n13324), .A2(n10451), .ZN(n13352) );
  NAND3_X1 U16162 ( .A1(n13412), .A2(n13303), .A3(n20848), .ZN(n12993) );
  NAND2_X1 U16163 ( .A1(n13352), .A2(n12993), .ZN(n12994) );
  NAND2_X1 U16164 ( .A1(n14032), .A2(n12994), .ZN(n12997) );
  NAND2_X1 U16165 ( .A1(n13136), .A2(n10451), .ZN(n12995) );
  NAND3_X1 U16166 ( .A1(n14023), .A2(n13464), .A3(n20848), .ZN(n12996) );
  NAND4_X1 U16167 ( .A1(n20224), .A2(n20199), .A3(n13420), .A4(n12998), .ZN(
        n12999) );
  NOR2_X1 U16168 ( .A1(n13348), .A2(n12999), .ZN(n13300) );
  NAND2_X1 U16169 ( .A1(n13300), .A2(n10451), .ZN(n13000) );
  AND2_X1 U16170 ( .A1(n15972), .A2(n20224), .ZN(n13002) );
  NAND2_X1 U16171 ( .A1(n13003), .A2(n13002), .ZN(n13020) );
  NOR4_X1 U16172 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13007) );
  NOR4_X1 U16173 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13006) );
  NOR4_X1 U16174 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13005) );
  NOR4_X1 U16175 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13004) );
  AND4_X1 U16176 ( .A1(n13007), .A2(n13006), .A3(n13005), .A4(n13004), .ZN(
        n13012) );
  NOR4_X1 U16177 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13010) );
  NOR4_X1 U16178 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13009) );
  NOR4_X1 U16179 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n13008) );
  INV_X1 U16180 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20766) );
  AND4_X1 U16181 ( .A1(n13010), .A2(n13009), .A3(n13008), .A4(n20766), .ZN(
        n13011) );
  NAND2_X1 U16182 ( .A1(n13012), .A2(n13011), .ZN(n13013) );
  INV_X1 U16183 ( .A(n13337), .ZN(n13409) );
  NOR3_X1 U16184 ( .A1(n14348), .A2(n20156), .A3(n13409), .ZN(n13014) );
  AOI22_X1 U16185 ( .A1(n14343), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14348), .ZN(n13015) );
  INV_X1 U16186 ( .A(n13015), .ZN(n13018) );
  INV_X1 U16187 ( .A(n20156), .ZN(n20157) );
  NOR2_X1 U16188 ( .A1(n13409), .A2(n20157), .ZN(n13016) );
  NAND2_X1 U16189 ( .A1(n15972), .A2(n13016), .ZN(n14306) );
  INV_X1 U16190 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20221) );
  NOR2_X1 U16191 ( .A1(n14306), .A2(n20221), .ZN(n13017) );
  NAND2_X1 U16192 ( .A1(n13020), .A2(n13019), .ZN(P1_U2873) );
  INV_X1 U16193 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20844) );
  NOR3_X1 U16194 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20844), .ZN(n13022) );
  NOR4_X1 U16195 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13021) );
  NAND4_X1 U16196 ( .A1(n20156), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13022), .A4(
        n13021), .ZN(U214) );
  NOR4_X1 U16197 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13023) );
  NAND3_X1 U16198 ( .A1(P2_W_R_N_REG_SCAN_IN), .A2(P2_M_IO_N_REG_SCAN_IN), 
        .A3(n13023), .ZN(n13024) );
  NAND3_X1 U16199 ( .A1(n16569), .A2(n19270), .A3(U214), .ZN(U212) );
  INV_X2 U16200 ( .A(n16642), .ZN(U215) );
  NAND2_X1 U16201 ( .A1(n13026), .A2(n13025), .ZN(n13027) );
  XNOR2_X1 U16202 ( .A(n13101), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13029) );
  XNOR2_X1 U16203 ( .A(n13029), .B(n13760), .ZN(n13090) );
  NAND2_X1 U16204 ( .A1(n16423), .A2(n13090), .ZN(n13030) );
  NAND2_X1 U16205 ( .A1(n19103), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13093) );
  OAI211_X1 U16206 ( .C1(n19165), .C2(n16413), .A(n13030), .B(n13093), .ZN(
        n13036) );
  INV_X1 U16207 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21038) );
  AOI211_X1 U16208 ( .C1(n21038), .C2(n13868), .A(n13051), .B(n15265), .ZN(
        n13035) );
  OAI21_X1 U16209 ( .B1(n13032), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13031), .ZN(n13094) );
  OAI22_X1 U16210 ( .A1(n16420), .A2(n13094), .B1(n13112), .B2(n13868), .ZN(
        n13034) );
  NOR2_X1 U16211 ( .A1(n16388), .A2(n13098), .ZN(n13033) );
  OR4_X1 U16212 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        P2_U3045) );
  NOR2_X1 U16213 ( .A1(n16445), .A2(n19181), .ZN(n13824) );
  INV_X1 U16214 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13038) );
  INV_X1 U16215 ( .A(n19928), .ZN(n19728) );
  NOR2_X1 U16216 ( .A1(n19728), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13039) );
  INV_X1 U16217 ( .A(n13039), .ZN(n13037) );
  OAI211_X1 U16218 ( .C1(n13824), .C2(n13038), .A(n13179), .B(n13037), .ZN(
        P2_U2814) );
  INV_X1 U16219 ( .A(n18951), .ZN(n13041) );
  OAI21_X1 U16220 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n13039), .A(n13041), 
        .ZN(n13040) );
  OAI21_X1 U16221 ( .B1(n13042), .B2(n13041), .A(n13040), .ZN(P2_U3612) );
  NOR3_X1 U16222 ( .A1(n13200), .A2(n13196), .A3(n13043), .ZN(n16450) );
  NOR2_X1 U16223 ( .A1(n16450), .A2(n16479), .ZN(n19967) );
  OAI21_X1 U16224 ( .B1(n19967), .B2(n12149), .A(n13092), .ZN(P2_U2819) );
  AND2_X1 U16225 ( .A1(n20813), .A2(n11284), .ZN(n13048) );
  AOI21_X1 U16226 ( .B1(n13046), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13048), 
        .ZN(n13047) );
  NAND2_X1 U16227 ( .A1(n13625), .A2(n13047), .ZN(P1_U2801) );
  NOR2_X1 U16228 ( .A1(n13048), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13050)
         );
  OAI21_X1 U16229 ( .B1(n10451), .B2(n14035), .A(n20846), .ZN(n13049) );
  OAI21_X1 U16230 ( .B1(n13050), .B2(n20846), .A(n13049), .ZN(P1_U3487) );
  NOR2_X1 U16231 ( .A1(n15259), .A2(n13838), .ZN(n13068) );
  NAND2_X1 U16232 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13051), .ZN(
        n13055) );
  OAI21_X1 U16233 ( .B1(n13054), .B2(n13053), .A(n13052), .ZN(n19938) );
  INV_X1 U16234 ( .A(n19938), .ZN(n13817) );
  OAI22_X1 U16235 ( .A1(n13055), .A2(n15259), .B1(n16413), .B2(n13817), .ZN(
        n13067) );
  INV_X1 U16236 ( .A(n13056), .ZN(n13059) );
  INV_X1 U16237 ( .A(n13057), .ZN(n13058) );
  NAND2_X1 U16238 ( .A1(n13059), .A2(n13058), .ZN(n13131) );
  NAND3_X1 U16239 ( .A1(n16423), .A2(n13132), .A3(n13131), .ZN(n13065) );
  OAI21_X1 U16240 ( .B1(n13062), .B2(n13061), .A(n13060), .ZN(n13063) );
  INV_X1 U16241 ( .A(n13063), .ZN(n13127) );
  NAND2_X1 U16242 ( .A1(n16400), .A2(n13127), .ZN(n13064) );
  NAND2_X1 U16243 ( .A1(n19103), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13128) );
  NAND3_X1 U16244 ( .A1(n13065), .A2(n13064), .A3(n13128), .ZN(n13066) );
  NOR3_X1 U16245 ( .A1(n13068), .A2(n13067), .A3(n13066), .ZN(n13074) );
  NOR2_X1 U16246 ( .A1(n15264), .A2(n13069), .ZN(n13071) );
  MUX2_X1 U16247 ( .A(n13071), .B(n13070), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13072) );
  INV_X1 U16248 ( .A(n13072), .ZN(n13073) );
  OAI211_X1 U16249 ( .C1(n16388), .C2(n11820), .A(n13074), .B(n13073), .ZN(
        P2_U3044) );
  OR2_X1 U16250 ( .A1(n13076), .A2(n13075), .ZN(n13077) );
  INV_X1 U16251 ( .A(n16449), .ZN(n13079) );
  NAND2_X1 U16252 ( .A1(n13079), .A2(n16442), .ZN(n13206) );
  NAND2_X1 U16253 ( .A1(n13206), .A2(n13184), .ZN(n13080) );
  MUX2_X1 U16254 ( .A(n13098), .B(n13764), .S(n14799), .Z(n13081) );
  OAI21_X1 U16255 ( .B1(n19943), .B2(n14785), .A(n13081), .ZN(P2_U2886) );
  NAND2_X1 U16256 ( .A1(n15585), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13082) );
  NAND4_X1 U16257 ( .A1(n19307), .A2(n13082), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19509), .ZN(n13083) );
  MUX2_X1 U16258 ( .A(n13607), .B(n13085), .S(n14799), .Z(n13086) );
  OAI21_X1 U16259 ( .B1(n19953), .B2(n14785), .A(n13086), .ZN(P2_U2887) );
  NAND2_X1 U16260 ( .A1(n16467), .A2(n19509), .ZN(n19924) );
  INV_X1 U16261 ( .A(n19924), .ZN(n13195) );
  OR2_X1 U16262 ( .A1(n19928), .A2(n13195), .ZN(n19941) );
  NAND2_X1 U16263 ( .A1(n19941), .A2(n21158), .ZN(n13087) );
  AND2_X1 U16264 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19942) );
  NAND2_X1 U16265 ( .A1(n19661), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13088) );
  NAND2_X1 U16266 ( .A1(n16471), .A2(n13088), .ZN(n13104) );
  INV_X1 U16267 ( .A(n13092), .ZN(n13089) );
  INV_X1 U16268 ( .A(n13090), .ZN(n13091) );
  OAI22_X1 U16269 ( .A1(n19259), .A2(n13091), .B1(n16338), .B2(n13761), .ZN(
        n13096) );
  OAI21_X1 U16270 ( .B1(n19257), .B2(n13094), .A(n13093), .ZN(n13095) );
  AOI211_X1 U16271 ( .C1(n16327), .C2(n13761), .A(n13096), .B(n13095), .ZN(
        n13097) );
  OAI21_X1 U16272 ( .B1(n13098), .B2(n16287), .A(n13097), .ZN(P2_U3013) );
  OAI21_X1 U16273 ( .B1(n13100), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13099), .ZN(n13110) );
  INV_X1 U16274 ( .A(n13110), .ZN(n13103) );
  AND2_X1 U16275 ( .A1(n19103), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13113) );
  OAI21_X1 U16276 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19124), .A(
        n13101), .ZN(n13111) );
  NOR2_X1 U16277 ( .A1(n19259), .A2(n13111), .ZN(n13102) );
  AOI211_X1 U16278 ( .C1(n9733), .C2(n13103), .A(n13113), .B(n13102), .ZN(
        n13106) );
  OAI21_X1 U16279 ( .B1(n19256), .B2(n13104), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13105) );
  OAI211_X1 U16280 ( .C1(n16287), .C2(n13607), .A(n13106), .B(n13105), .ZN(
        P2_U3014) );
  OAI21_X1 U16281 ( .B1(n13109), .B2(n13108), .A(n13107), .ZN(n19120) );
  OAI22_X1 U16282 ( .A1(n16420), .A2(n13110), .B1(n16413), .B2(n19120), .ZN(
        n13116) );
  NOR2_X1 U16283 ( .A1(n16388), .A2(n13607), .ZN(n13115) );
  OAI22_X1 U16284 ( .A1(n21038), .A2(n13112), .B1(n16393), .B2(n13111), .ZN(
        n13114) );
  NOR4_X1 U16285 ( .A1(n13116), .A2(n13115), .A3(n13114), .A4(n13113), .ZN(
        n13117) );
  OAI21_X1 U16286 ( .B1(n15265), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13117), .ZN(P2_U3046) );
  NAND2_X1 U16287 ( .A1(n14799), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13122) );
  NAND2_X1 U16288 ( .A1(n13120), .A2(n14790), .ZN(n13121) );
  OAI211_X1 U16289 ( .C1(n19565), .C2(n14785), .A(n13122), .B(n13121), .ZN(
        P2_U2884) );
  OR2_X1 U16290 ( .A1(n13124), .A2(n13123), .ZN(n13125) );
  NAND2_X1 U16291 ( .A1(n13125), .A2(n13217), .ZN(n19084) );
  INV_X1 U16292 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19234) );
  AOI22_X1 U16293 ( .A1(n19270), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19268), .ZN(n13238) );
  OAI222_X1 U16294 ( .A1(n19084), .A2(n19138), .B1(n14836), .B2(n19234), .C1(
        n19180), .C2(n13238), .ZN(P2_U2911) );
  INV_X1 U16295 ( .A(n13819), .ZN(n13821) );
  INV_X1 U16296 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U16297 ( .A1(n9733), .A2(n13127), .ZN(n13129) );
  OAI211_X1 U16298 ( .C1(n16338), .C2(n13130), .A(n13129), .B(n13128), .ZN(
        n13134) );
  AND3_X1 U16299 ( .A1(n16335), .A2(n13132), .A3(n13131), .ZN(n13133) );
  AOI211_X1 U16300 ( .C1(n16327), .C2(n13821), .A(n13134), .B(n13133), .ZN(
        n13135) );
  OAI21_X1 U16301 ( .B1(n11820), .B2(n16287), .A(n13135), .ZN(P2_U3012) );
  INV_X1 U16302 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13144) );
  NAND2_X1 U16303 ( .A1(n13136), .A2(n13296), .ZN(n13137) );
  NAND2_X1 U16304 ( .A1(n13412), .A2(n13138), .ZN(n15816) );
  INV_X1 U16305 ( .A(n15816), .ZN(n13140) );
  INV_X1 U16306 ( .A(n15842), .ZN(n13139) );
  OAI211_X1 U16307 ( .C1(n15789), .C2(n13140), .A(n13139), .B(n13420), .ZN(
        n13141) );
  INV_X1 U16308 ( .A(n13141), .ZN(n13142) );
  NAND2_X1 U16309 ( .A1(n20072), .A2(n13428), .ZN(n13388) );
  INV_X1 U16310 ( .A(n16179), .ZN(n16181) );
  NOR2_X1 U16311 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16181), .ZN(n20093) );
  NOR2_X4 U16312 ( .A1(n20072), .A2(n20849), .ZN(n15844) );
  AOI22_X1 U16313 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13143) );
  OAI21_X1 U16314 ( .B1(n13144), .B2(n13388), .A(n13143), .ZN(P1_U2912) );
  INV_X1 U16315 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13146) );
  AOI22_X1 U16316 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13145) );
  OAI21_X1 U16317 ( .B1(n13146), .B2(n13388), .A(n13145), .ZN(P1_U2913) );
  INV_X1 U16318 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13148) );
  AOI22_X1 U16319 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13147) );
  OAI21_X1 U16320 ( .B1(n13148), .B2(n13388), .A(n13147), .ZN(P1_U2914) );
  AOI22_X1 U16321 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13149) );
  OAI21_X1 U16322 ( .B1(n14291), .B2(n13388), .A(n13149), .ZN(P1_U2908) );
  INV_X1 U16323 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13151) );
  AOI22_X1 U16324 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13150) );
  OAI21_X1 U16325 ( .B1(n13151), .B2(n13388), .A(n13150), .ZN(P1_U2920) );
  INV_X1 U16326 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13153) );
  AOI22_X1 U16327 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13152) );
  OAI21_X1 U16328 ( .B1(n13153), .B2(n13388), .A(n13152), .ZN(P1_U2918) );
  INV_X1 U16329 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13155) );
  AOI22_X1 U16330 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13154) );
  OAI21_X1 U16331 ( .B1(n13155), .B2(n13388), .A(n13154), .ZN(P1_U2911) );
  INV_X1 U16332 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16333 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13156) );
  OAI21_X1 U16334 ( .B1(n13157), .B2(n13388), .A(n13156), .ZN(P1_U2909) );
  INV_X1 U16335 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13159) );
  AOI22_X1 U16336 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13158) );
  OAI21_X1 U16337 ( .B1(n13159), .B2(n13388), .A(n13158), .ZN(P1_U2917) );
  INV_X1 U16338 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13161) );
  AOI22_X1 U16339 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13160) );
  OAI21_X1 U16340 ( .B1(n13161), .B2(n13388), .A(n13160), .ZN(P1_U2919) );
  INV_X1 U16341 ( .A(n13162), .ZN(n13164) );
  OR3_X1 U16342 ( .A1(n13165), .A2(n13164), .A3(n13163), .ZN(n13166) );
  NAND2_X1 U16343 ( .A1(n13270), .A2(n13166), .ZN(n19148) );
  NAND2_X1 U16344 ( .A1(n13168), .A2(n13167), .ZN(n13170) );
  INV_X1 U16345 ( .A(n13211), .ZN(n13169) );
  AND2_X1 U16346 ( .A1(n13170), .A2(n13169), .ZN(n19262) );
  INV_X1 U16347 ( .A(n19262), .ZN(n19104) );
  MUX2_X1 U16348 ( .A(n12495), .B(n19104), .S(n14790), .Z(n13171) );
  OAI21_X1 U16349 ( .B1(n19148), .B2(n14785), .A(n13171), .ZN(P2_U2883) );
  INV_X1 U16350 ( .A(n19936), .ZN(n13825) );
  MUX2_X1 U16351 ( .A(n13176), .B(P2_EBX_REG_2__SCAN_IN), .S(n14799), .Z(
        n13177) );
  AOI21_X1 U16352 ( .B1(n13825), .B2(n14798), .A(n13177), .ZN(n13178) );
  INV_X1 U16353 ( .A(n13178), .ZN(P2_U2885) );
  NOR3_X4 U16354 ( .A1(n13179), .A2(n11776), .A3(n19857), .ZN(n13276) );
  INV_X1 U16355 ( .A(n13276), .ZN(n13182) );
  AOI22_X1 U16356 ( .A1(n19270), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19268), .ZN(n13572) );
  AOI22_X1 U16357 ( .A1(P2_LWORD_REG_15__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n13181) );
  OAI21_X1 U16358 ( .B1(n13182), .B2(n13572), .A(n13181), .ZN(P2_U2982) );
  INV_X1 U16359 ( .A(n19565), .ZN(n19930) );
  INV_X1 U16360 ( .A(n13606), .ZN(n14004) );
  NAND2_X1 U16361 ( .A1(n13120), .A2(n14004), .ZN(n13194) );
  NOR2_X1 U16362 ( .A1(n16441), .A2(n16442), .ZN(n13872) );
  INV_X1 U16363 ( .A(n13872), .ZN(n13183) );
  NOR2_X1 U16364 ( .A1(n14000), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13189) );
  NAND2_X1 U16365 ( .A1(n13183), .A2(n13189), .ZN(n13878) );
  NAND2_X1 U16366 ( .A1(n12595), .A2(n13184), .ZN(n13870) );
  NAND2_X1 U16367 ( .A1(n13870), .A2(n13185), .ZN(n13187) );
  INV_X1 U16368 ( .A(n11538), .ZN(n13875) );
  NAND2_X1 U16369 ( .A1(n13876), .A2(n13875), .ZN(n13186) );
  NAND2_X1 U16370 ( .A1(n13187), .A2(n13186), .ZN(n13874) );
  INV_X1 U16371 ( .A(n13874), .ZN(n13188) );
  NAND2_X1 U16372 ( .A1(n13878), .A2(n13188), .ZN(n13191) );
  INV_X1 U16373 ( .A(n13876), .ZN(n13999) );
  OAI22_X1 U16374 ( .A1(n13872), .A2(n13189), .B1(n13999), .B2(n13875), .ZN(
        n13190) );
  MUX2_X1 U16375 ( .A(n13191), .B(n13190), .S(n11537), .Z(n13192) );
  NOR2_X1 U16376 ( .A1(n13192), .A2(n11898), .ZN(n13193) );
  NAND2_X1 U16377 ( .A1(n13194), .A2(n13193), .ZN(n16432) );
  AOI22_X1 U16378 ( .A1(n19930), .A2(n16474), .B1(n13195), .B2(n16432), .ZN(
        n13210) );
  NOR2_X1 U16379 ( .A1(n21158), .A2(n15857), .ZN(n16481) );
  INV_X1 U16380 ( .A(n13196), .ZN(n13201) );
  INV_X1 U16381 ( .A(n13197), .ZN(n13199) );
  OAI211_X1 U16382 ( .C1(n13201), .C2(n13200), .A(n13199), .B(n13198), .ZN(
        n13202) );
  INV_X1 U16383 ( .A(n13202), .ZN(n13207) );
  NOR2_X1 U16384 ( .A1(n16451), .A2(n13203), .ZN(n13204) );
  NAND2_X1 U16385 ( .A1(n19183), .A2(n13204), .ZN(n13205) );
  OAI22_X1 U16386 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19509), .B1(n16458), 
        .B2(n16479), .ZN(n13208) );
  AOI21_X1 U16387 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16481), .A(n13208), .ZN(
        n13995) );
  NAND2_X1 U16388 ( .A1(n13995), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13209) );
  OAI21_X1 U16389 ( .B1(n13210), .B2(n13995), .A(n13209), .ZN(P2_U3596) );
  XOR2_X1 U16390 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13270), .Z(n13215)
         );
  OAI21_X1 U16391 ( .B1(n13212), .B2(n13211), .A(n13265), .ZN(n16332) );
  MUX2_X1 U16392 ( .A(n16332), .B(n13213), .S(n14799), .Z(n13214) );
  OAI21_X1 U16393 ( .B1(n13215), .B2(n14785), .A(n13214), .ZN(P2_U2882) );
  AOI21_X1 U16394 ( .B1(n13218), .B2(n13217), .A(n13216), .ZN(n15317) );
  INV_X1 U16395 ( .A(n15317), .ZN(n13661) );
  INV_X1 U16396 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19232) );
  INV_X1 U16397 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20955) );
  OR2_X1 U16398 ( .A1(n19268), .A2(n20955), .ZN(n13220) );
  NAND2_X1 U16399 ( .A1(n19268), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13219) );
  NAND2_X1 U16400 ( .A1(n13220), .A2(n13219), .ZN(n14838) );
  INV_X1 U16401 ( .A(n14838), .ZN(n13221) );
  OAI222_X1 U16402 ( .A1(n13661), .A2(n19138), .B1(n14836), .B2(n19232), .C1(
        n19180), .C2(n13221), .ZN(P2_U2910) );
  AOI22_X1 U16403 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U16404 ( .A1(n19270), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19268), .ZN(n19280) );
  INV_X1 U16405 ( .A(n19280), .ZN(n13806) );
  NAND2_X1 U16406 ( .A1(n13276), .A2(n13806), .ZN(n13236) );
  NAND2_X1 U16407 ( .A1(n13222), .A2(n13236), .ZN(P2_U2952) );
  AOI22_X1 U16408 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U16409 ( .A1(n19270), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19268), .ZN(n19308) );
  INV_X1 U16410 ( .A(n19308), .ZN(n14856) );
  NAND2_X1 U16411 ( .A1(n13276), .A2(n14856), .ZN(n13240) );
  NAND2_X1 U16412 ( .A1(n13223), .A2(n13240), .ZN(P2_U2958) );
  AOI22_X1 U16413 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13224) );
  OAI22_X1 U16414 ( .A1(n19268), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19270), .ZN(n19318) );
  INV_X1 U16415 ( .A(n19318), .ZN(n16264) );
  NAND2_X1 U16416 ( .A1(n13276), .A2(n16264), .ZN(n13246) );
  NAND2_X1 U16417 ( .A1(n13224), .A2(n13246), .ZN(P2_U2959) );
  AOI22_X1 U16418 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U16419 ( .A1(n19270), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19268), .ZN(n19303) );
  INV_X1 U16420 ( .A(n19303), .ZN(n14862) );
  NAND2_X1 U16421 ( .A1(n13276), .A2(n14862), .ZN(n13232) );
  NAND2_X1 U16422 ( .A1(n13225), .A2(n13232), .ZN(P2_U2957) );
  AOI22_X1 U16423 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U16424 ( .A1(n19270), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19268), .ZN(n19287) );
  INV_X1 U16425 ( .A(n19287), .ZN(n13903) );
  NAND2_X1 U16426 ( .A1(n13276), .A2(n13903), .ZN(n13228) );
  NAND2_X1 U16427 ( .A1(n13226), .A2(n13228), .ZN(P2_U2968) );
  AOI22_X1 U16428 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U16429 ( .A1(n19270), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19268), .ZN(n19291) );
  INV_X1 U16430 ( .A(n19291), .ZN(n13937) );
  NAND2_X1 U16431 ( .A1(n13276), .A2(n13937), .ZN(n13230) );
  NAND2_X1 U16432 ( .A1(n13227), .A2(n13230), .ZN(P2_U2969) );
  AOI22_X1 U16433 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13229) );
  NAND2_X1 U16434 ( .A1(n13229), .A2(n13228), .ZN(P2_U2953) );
  AOI22_X1 U16435 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13231) );
  NAND2_X1 U16436 ( .A1(n13231), .A2(n13230), .ZN(P2_U2954) );
  AOI22_X1 U16437 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13233) );
  NAND2_X1 U16438 ( .A1(n13233), .A2(n13232), .ZN(P2_U2972) );
  AOI22_X1 U16439 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n13235) );
  NAND2_X1 U16440 ( .A1(n13276), .A2(n13234), .ZN(n13256) );
  NAND2_X1 U16441 ( .A1(n13235), .A2(n13256), .ZN(P2_U2966) );
  AOI22_X1 U16442 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U16443 ( .A1(n13237), .A2(n13236), .ZN(P2_U2967) );
  AOI22_X1 U16444 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13239) );
  INV_X1 U16445 ( .A(n13238), .ZN(n14846) );
  NAND2_X1 U16446 ( .A1(n13276), .A2(n14846), .ZN(n13248) );
  NAND2_X1 U16447 ( .A1(n13239), .A2(n13248), .ZN(P2_U2975) );
  AOI22_X1 U16448 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13241) );
  NAND2_X1 U16449 ( .A1(n13241), .A2(n13240), .ZN(P2_U2973) );
  AOI22_X1 U16450 ( .A1(P2_LWORD_REG_10__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n13242) );
  MUX2_X1 U16451 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n19268), .Z(n14828) );
  NAND2_X1 U16452 ( .A1(n13276), .A2(n14828), .ZN(n13252) );
  NAND2_X1 U16453 ( .A1(n13242), .A2(n13252), .ZN(P2_U2977) );
  AOI22_X1 U16454 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13243) );
  INV_X1 U16455 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16605) );
  INV_X1 U16456 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18297) );
  OAI22_X1 U16457 ( .A1(n19268), .A2(n16605), .B1(n18297), .B2(n19270), .ZN(
        n19298) );
  NAND2_X1 U16458 ( .A1(n13276), .A2(n19298), .ZN(n13254) );
  NAND2_X1 U16459 ( .A1(n13243), .A2(n13254), .ZN(P2_U2956) );
  AOI22_X1 U16460 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16461 ( .A1(n19270), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19268), .ZN(n19141) );
  INV_X1 U16462 ( .A(n19141), .ZN(n14812) );
  NAND2_X1 U16463 ( .A1(n13276), .A2(n14812), .ZN(n13250) );
  NAND2_X1 U16464 ( .A1(n13244), .A2(n13250), .ZN(P2_U2979) );
  AOI22_X1 U16465 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U16466 ( .A1(n19270), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19268), .ZN(n19294) );
  INV_X1 U16467 ( .A(n19294), .ZN(n14880) );
  NAND2_X1 U16468 ( .A1(n13276), .A2(n14880), .ZN(n13260) );
  NAND2_X1 U16469 ( .A1(n13245), .A2(n13260), .ZN(P2_U2970) );
  AOI22_X1 U16470 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13247) );
  NAND2_X1 U16471 ( .A1(n13247), .A2(n13246), .ZN(P2_U2974) );
  AOI22_X1 U16472 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13249) );
  NAND2_X1 U16473 ( .A1(n13249), .A2(n13248), .ZN(P2_U2960) );
  AOI22_X1 U16474 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U16475 ( .A1(n13251), .A2(n13250), .ZN(P2_U2964) );
  AOI22_X1 U16476 ( .A1(P2_UWORD_REG_10__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U16477 ( .A1(n13253), .A2(n13252), .ZN(P2_U2962) );
  AOI22_X1 U16478 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13255) );
  NAND2_X1 U16479 ( .A1(n13255), .A2(n13254), .ZN(P2_U2971) );
  AOI22_X1 U16480 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(n13282), .B1(n13258), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n13257) );
  NAND2_X1 U16481 ( .A1(n13257), .A2(n13256), .ZN(P2_U2981) );
  AOI22_X1 U16482 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n13259), .B1(n13258), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13261) );
  NAND2_X1 U16483 ( .A1(n13261), .A2(n13260), .ZN(P2_U2955) );
  OR2_X1 U16484 ( .A1(n13262), .A2(n13216), .ZN(n13263) );
  NAND2_X1 U16485 ( .A1(n13263), .A2(n13372), .ZN(n19071) );
  INV_X1 U16486 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19230) );
  INV_X1 U16487 ( .A(n14828), .ZN(n13264) );
  OAI222_X1 U16488 ( .A1(n19071), .A2(n19138), .B1(n14836), .B2(n19230), .C1(
        n19180), .C2(n13264), .ZN(P2_U2909) );
  NAND2_X1 U16489 ( .A1(n13266), .A2(n13265), .ZN(n13268) );
  INV_X1 U16490 ( .A(n13311), .ZN(n13267) );
  NAND2_X1 U16491 ( .A1(n13268), .A2(n13267), .ZN(n19092) );
  NOR2_X1 U16492 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  OAI211_X1 U16493 ( .C1(n13271), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14798), .B(n13310), .ZN(n13273) );
  NAND2_X1 U16494 ( .A1(n14799), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13272) );
  OAI211_X1 U16495 ( .C1(n19092), .C2(n14799), .A(n13273), .B(n13272), .ZN(
        P2_U2881) );
  INV_X1 U16496 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19195) );
  MUX2_X1 U16497 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n19268), .Z(n14821) );
  NAND2_X1 U16498 ( .A1(n13276), .A2(n14821), .ZN(n13281) );
  NAND2_X1 U16499 ( .A1(n13282), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13274) );
  OAI211_X1 U16500 ( .C1(n19195), .C2(n19185), .A(n13281), .B(n13274), .ZN(
        P2_U2963) );
  INV_X1 U16501 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19199) );
  NAND2_X1 U16502 ( .A1(n13276), .A2(n14838), .ZN(n13279) );
  NAND2_X1 U16503 ( .A1(n13282), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13275) );
  OAI211_X1 U16504 ( .C1(n19199), .C2(n19185), .A(n13279), .B(n13275), .ZN(
        P2_U2961) );
  INV_X1 U16505 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19224) );
  MUX2_X1 U16506 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n19268), .Z(n14804) );
  NAND2_X1 U16507 ( .A1(n13276), .A2(n14804), .ZN(n13284) );
  NAND2_X1 U16508 ( .A1(n13282), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13277) );
  OAI211_X1 U16509 ( .C1(n19224), .C2(n19185), .A(n13284), .B(n13277), .ZN(
        P2_U2980) );
  NAND2_X1 U16510 ( .A1(n13282), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13278) );
  OAI211_X1 U16511 ( .C1(n19232), .C2(n19185), .A(n13279), .B(n13278), .ZN(
        P2_U2976) );
  INV_X1 U16512 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19228) );
  NAND2_X1 U16513 ( .A1(n13282), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13280) );
  OAI211_X1 U16514 ( .C1(n19228), .C2(n19185), .A(n13281), .B(n13280), .ZN(
        P2_U2978) );
  INV_X1 U16515 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19191) );
  NAND2_X1 U16516 ( .A1(n13282), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13283) );
  OAI211_X1 U16517 ( .C1(n19191), .C2(n19185), .A(n13284), .B(n13283), .ZN(
        P2_U2965) );
  INV_X1 U16518 ( .A(n13285), .ZN(n13288) );
  OAI21_X1 U16519 ( .B1(n13288), .B2(n13287), .A(n13286), .ZN(n20138) );
  NAND2_X1 U16520 ( .A1(n10437), .A2(n14027), .ZN(n13289) );
  NAND2_X1 U16521 ( .A1(n20157), .A2(DATAI_0_), .ZN(n13291) );
  NAND2_X1 U16522 ( .A1(n20156), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13290) );
  AND2_X1 U16523 ( .A1(n13291), .A2(n13290), .ZN(n20163) );
  INV_X1 U16524 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20096) );
  OAI222_X1 U16525 ( .A1(n20138), .A2(n14354), .B1(n14353), .B2(n20163), .C1(
        n15972), .C2(n20096), .ZN(P1_U2904) );
  OAI21_X1 U16526 ( .B1(n13293), .B2(n13292), .A(n13377), .ZN(n14191) );
  NAND2_X1 U16527 ( .A1(n20157), .A2(DATAI_1_), .ZN(n13295) );
  NAND2_X1 U16528 ( .A1(n20156), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13294) );
  AND2_X1 U16529 ( .A1(n13295), .A2(n13294), .ZN(n20179) );
  OAI222_X1 U16530 ( .A1(n14191), .A2(n14354), .B1(n14353), .B2(n20179), .C1(
        n15972), .C2(n10562), .ZN(P1_U2903) );
  INV_X1 U16531 ( .A(n14191), .ZN(n13320) );
  NOR2_X1 U16532 ( .A1(n13366), .A2(n20177), .ZN(n13416) );
  NAND2_X1 U16533 ( .A1(n13296), .A2(n10435), .ZN(n13297) );
  INV_X1 U16534 ( .A(n14022), .ZN(n13299) );
  NAND2_X1 U16535 ( .A1(n13300), .A2(n13303), .ZN(n13301) );
  OR2_X1 U16536 ( .A1(n13304), .A2(n13303), .ZN(n13305) );
  NAND2_X1 U16537 ( .A1(n13306), .A2(n13305), .ZN(n13440) );
  INV_X1 U16538 ( .A(n13440), .ZN(n14185) );
  OAI22_X1 U16539 ( .A1(n14280), .A2(n14185), .B1(n13307), .B2(n14278), .ZN(
        n13308) );
  AOI21_X1 U16540 ( .B1(n13320), .B2(n13782), .A(n13308), .ZN(n13309) );
  INV_X1 U16541 ( .A(n13309), .ZN(P1_U2871) );
  XOR2_X1 U16542 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13310), .Z(n13316)
         );
  OR2_X1 U16543 ( .A1(n13312), .A2(n13311), .ZN(n13313) );
  AND2_X1 U16544 ( .A1(n13391), .A2(n13313), .ZN(n16318) );
  INV_X1 U16545 ( .A(n16318), .ZN(n15334) );
  MUX2_X1 U16546 ( .A(n15334), .B(n13314), .S(n14799), .Z(n13315) );
  OAI21_X1 U16547 ( .B1(n13316), .B2(n14785), .A(n13315), .ZN(P2_U2880) );
  XNOR2_X1 U16548 ( .A(n13317), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13443) );
  INV_X1 U16549 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20836) );
  NOR2_X1 U16550 ( .A1(n20042), .A2(n20836), .ZN(n13439) );
  AOI21_X1 U16551 ( .B1(n20132), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13439), .ZN(n13318) );
  OAI21_X1 U16552 ( .B1(n16029), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13318), .ZN(n13319) );
  AOI21_X1 U16553 ( .B1(n13320), .B2(n20158), .A(n13319), .ZN(n13321) );
  OAI21_X1 U16554 ( .B1(n13443), .B2(n19981), .A(n13321), .ZN(P1_U2998) );
  INV_X1 U16555 ( .A(n13322), .ZN(n13335) );
  INV_X1 U16556 ( .A(n20848), .ZN(n16173) );
  NOR2_X1 U16557 ( .A1(n15842), .A2(n16173), .ZN(n13323) );
  AND2_X1 U16558 ( .A1(n14032), .A2(n13323), .ZN(n15811) );
  OAI21_X1 U16559 ( .B1(n13412), .B2(n15789), .A(n15811), .ZN(n13334) );
  INV_X1 U16560 ( .A(n13324), .ZN(n13325) );
  NAND2_X1 U16561 ( .A1(n13325), .A2(n11276), .ZN(n13329) );
  AOI21_X1 U16562 ( .B1(n13326), .B2(n13626), .A(n20162), .ZN(n13327) );
  NAND2_X1 U16563 ( .A1(n13328), .A2(n13327), .ZN(n13346) );
  NAND2_X1 U16564 ( .A1(n13329), .A2(n13346), .ZN(n13415) );
  NOR2_X1 U16565 ( .A1(n13741), .A2(n13338), .ZN(n13330) );
  NOR2_X1 U16566 ( .A1(n13415), .A2(n13330), .ZN(n13331) );
  AND2_X1 U16567 ( .A1(n13332), .A2(n13331), .ZN(n13333) );
  INV_X1 U16568 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19982) );
  NAND2_X1 U16569 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16179), .ZN(n13471) );
  OR2_X1 U16570 ( .A1(n19982), .A2(n13471), .ZN(n13336) );
  OAI21_X1 U16571 ( .B1(n15792), .B2(n19976), .A(n13336), .ZN(n16166) );
  NAND2_X1 U16572 ( .A1(n13337), .A2(n20162), .ZN(n13339) );
  AOI22_X1 U16573 ( .A1(n13450), .A2(n13626), .B1(n13339), .B2(n13338), .ZN(
        n13340) );
  OAI211_X1 U16574 ( .C1(n13342), .C2(n11383), .A(n13341), .B(n13340), .ZN(
        n13343) );
  INV_X1 U16575 ( .A(n13343), .ZN(n13347) );
  NAND2_X1 U16576 ( .A1(n13344), .A2(n10451), .ZN(n13345) );
  AND3_X1 U16577 ( .A1(n13347), .A2(n13346), .A3(n13345), .ZN(n13427) );
  NAND2_X1 U16578 ( .A1(n13429), .A2(n13348), .ZN(n13349) );
  OR2_X1 U16579 ( .A1(n13349), .A2(n13412), .ZN(n13350) );
  NOR2_X1 U16580 ( .A1(n13464), .A2(n13350), .ZN(n13351) );
  AND2_X1 U16581 ( .A1(n13427), .A2(n13351), .ZN(n14653) );
  INV_X1 U16582 ( .A(n14653), .ZN(n13456) );
  NAND2_X1 U16583 ( .A1(n20817), .A2(n13456), .ZN(n13363) );
  INV_X1 U16584 ( .A(n13352), .ZN(n13423) );
  OR2_X1 U16585 ( .A1(n13423), .A2(n14022), .ZN(n13451) );
  INV_X1 U16586 ( .A(n10286), .ZN(n14654) );
  NAND2_X1 U16587 ( .A1(n14654), .A2(n9966), .ZN(n13447) );
  NAND2_X1 U16588 ( .A1(n13451), .A2(n13447), .ZN(n13358) );
  NAND2_X1 U16589 ( .A1(n15789), .A2(n13353), .ZN(n14658) );
  INV_X1 U16590 ( .A(n14658), .ZN(n13356) );
  INV_X1 U16591 ( .A(n13451), .ZN(n13354) );
  NOR2_X1 U16592 ( .A1(n13354), .A2(n13447), .ZN(n13355) );
  AOI211_X1 U16593 ( .C1(n15789), .C2(n9966), .A(n13356), .B(n13355), .ZN(
        n13357) );
  MUX2_X1 U16594 ( .A(n13358), .B(n13357), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13362) );
  NAND3_X1 U16595 ( .A1(n15789), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n13359), .ZN(n13361) );
  NAND3_X1 U16596 ( .A1(n14653), .A2(n13450), .A3(n9841), .ZN(n13360) );
  NAND4_X1 U16597 ( .A1(n13363), .A2(n13362), .A3(n13361), .A4(n13360), .ZN(
        n13444) );
  INV_X1 U16598 ( .A(n14671), .ZN(n15822) );
  AOI22_X1 U16599 ( .A1(n13444), .A2(n19975), .B1(n9841), .B2(n15822), .ZN(
        n13365) );
  NAND2_X1 U16600 ( .A1(n16165), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13364) );
  OAI21_X1 U16601 ( .B1(n16165), .B2(n13365), .A(n13364), .ZN(P1_U3469) );
  AOI21_X1 U16602 ( .B1(n15789), .B2(n19975), .A(n16165), .ZN(n13371) );
  NOR2_X1 U16603 ( .A1(n13366), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13367) );
  AOI21_X1 U16604 ( .B1(n10570), .B2(n13456), .A(n13367), .ZN(n15791) );
  OAI21_X1 U16605 ( .B1(n15791), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n11284), 
        .ZN(n13368) );
  NOR2_X1 U16606 ( .A1(n11284), .A2(n9916), .ZN(n14663) );
  INV_X1 U16607 ( .A(n14663), .ZN(n14668) );
  AOI22_X1 U16608 ( .A1(n13368), .A2(n14668), .B1(n13370), .B2(n15822), .ZN(
        n13369) );
  OAI22_X1 U16609 ( .A1(n13371), .A2(n13370), .B1(n16165), .B2(n13369), .ZN(
        P1_U3474) );
  AOI21_X1 U16610 ( .B1(n13373), .B2(n13372), .A(n9816), .ZN(n16363) );
  INV_X1 U16611 ( .A(n16363), .ZN(n13375) );
  INV_X1 U16612 ( .A(n14821), .ZN(n13374) );
  OAI222_X1 U16613 ( .A1(n13375), .A2(n19138), .B1(n14836), .B2(n19228), .C1(
        n19180), .C2(n13374), .ZN(P2_U2908) );
  OAI21_X1 U16614 ( .B1(n13376), .B2(n10576), .A(n13378), .ZN(n13755) );
  NAND2_X1 U16615 ( .A1(n20157), .A2(DATAI_2_), .ZN(n13380) );
  NAND2_X1 U16616 ( .A1(n20156), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13379) );
  AND2_X1 U16617 ( .A1(n13380), .A2(n13379), .ZN(n20185) );
  OAI222_X1 U16618 ( .A1(n13755), .A2(n14354), .B1(n14353), .B2(n20185), .C1(
        n15972), .C2(n10554), .ZN(P1_U2902) );
  INV_X1 U16619 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13382) );
  AOI22_X1 U16620 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13381) );
  OAI21_X1 U16621 ( .B1(n13382), .B2(n13388), .A(n13381), .ZN(P1_U2915) );
  AOI22_X1 U16622 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13383) );
  OAI21_X1 U16623 ( .B1(n14304), .B2(n13388), .A(n13383), .ZN(P1_U2910) );
  INV_X1 U16624 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U16625 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13384) );
  OAI21_X1 U16626 ( .B1(n13385), .B2(n13388), .A(n13384), .ZN(P1_U2916) );
  AOI22_X1 U16627 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13386) );
  OAI21_X1 U16628 ( .B1(n11185), .B2(n13388), .A(n13386), .ZN(P1_U2907) );
  INV_X1 U16629 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13389) );
  AOI22_X1 U16630 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20849), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15844), .ZN(n13387) );
  OAI21_X1 U16631 ( .B1(n13389), .B2(n13388), .A(n13387), .ZN(P1_U2906) );
  NAND2_X1 U16632 ( .A1(n13391), .A2(n13390), .ZN(n13392) );
  NAND2_X1 U16633 ( .A1(n13397), .A2(n13392), .ZN(n19078) );
  NAND2_X1 U16634 ( .A1(n13393), .A2(n13394), .ZN(n13553) );
  OAI211_X1 U16635 ( .C1(n13393), .C2(n13394), .A(n13553), .B(n14798), .ZN(
        n13396) );
  NAND2_X1 U16636 ( .A1(n14799), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13395) );
  OAI211_X1 U16637 ( .C1(n19078), .C2(n14799), .A(n13396), .B(n13395), .ZN(
        P2_U2879) );
  XNOR2_X1 U16638 ( .A(n13553), .B(n13552), .ZN(n13400) );
  AOI21_X1 U16639 ( .B1(n13398), .B2(n13397), .A(n13558), .ZN(n16310) );
  INV_X1 U16640 ( .A(n16310), .ZN(n15319) );
  MUX2_X1 U16641 ( .A(n15319), .B(n12512), .S(n14799), .Z(n13399) );
  OAI21_X1 U16642 ( .B1(n13400), .B2(n14785), .A(n13399), .ZN(P2_U2878) );
  INV_X1 U16643 ( .A(n13755), .ZN(n13489) );
  NAND2_X1 U16644 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  AND2_X1 U16645 ( .A1(n13504), .A2(n13403), .ZN(n13743) );
  INV_X1 U16646 ( .A(n13743), .ZN(n13405) );
  OAI22_X1 U16647 ( .A1(n14280), .A2(n13405), .B1(n13404), .B2(n14278), .ZN(
        n13406) );
  AOI21_X1 U16648 ( .B1(n13489), .B2(n13782), .A(n13406), .ZN(n13407) );
  INV_X1 U16649 ( .A(n13407), .ZN(P1_U2870) );
  AOI21_X1 U16650 ( .B1(n13626), .B2(n15842), .A(n16173), .ZN(n13408) );
  NAND2_X1 U16651 ( .A1(n14023), .A2(n13408), .ZN(n13414) );
  NAND3_X1 U16652 ( .A1(n13412), .A2(n13626), .A3(n20848), .ZN(n13410) );
  NAND3_X1 U16653 ( .A1(n13410), .A2(n13428), .A3(n13409), .ZN(n13411) );
  AOI22_X1 U16654 ( .A1(n15811), .A2(n13412), .B1(n14032), .B2(n13411), .ZN(
        n13413) );
  INV_X1 U16655 ( .A(n14032), .ZN(n13417) );
  AOI21_X1 U16656 ( .B1(n13417), .B2(n13416), .A(n13415), .ZN(n13418) );
  NAND2_X1 U16657 ( .A1(n13419), .A2(n13418), .ZN(n13421) );
  NOR2_X1 U16658 ( .A1(n13423), .A2(n13422), .ZN(n14021) );
  OAI211_X1 U16659 ( .C1(n20199), .C2(n13436), .A(n14021), .B(n13424), .ZN(
        n13425) );
  OAI211_X1 U16660 ( .C1(n13429), .C2(n13428), .A(n13427), .B(n13426), .ZN(
        n13430) );
  NAND2_X1 U16661 ( .A1(n13438), .A2(n13430), .ZN(n14598) );
  NAND2_X1 U16662 ( .A1(n14598), .A2(n14642), .ZN(n20139) );
  NAND2_X1 U16663 ( .A1(n13438), .A2(n15789), .ZN(n16089) );
  NOR2_X1 U16664 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20143), .ZN(
        n13492) );
  NOR2_X1 U16665 ( .A1(n16064), .A2(n13492), .ZN(n13433) );
  AOI21_X1 U16666 ( .B1(n9916), .B2(n20139), .A(n20142), .ZN(n13431) );
  INV_X1 U16667 ( .A(n13431), .ZN(n13432) );
  MUX2_X1 U16668 ( .A(n13433), .B(n13432), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13434) );
  INV_X1 U16669 ( .A(n13434), .ZN(n13442) );
  OAI21_X1 U16670 ( .B1(n13436), .B2(n13435), .A(n15816), .ZN(n13437) );
  AOI21_X1 U16671 ( .B1(n20145), .B2(n13440), .A(n13439), .ZN(n13441) );
  OAI211_X1 U16672 ( .C1(n13443), .C2(n16160), .A(n13442), .B(n13441), .ZN(
        P1_U3030) );
  NOR2_X1 U16673 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n11284), .ZN(n13467) );
  MUX2_X1 U16674 ( .A(n13444), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15792), .Z(n15802) );
  AOI22_X1 U16675 ( .A1(n13467), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n11284), .B2(n15802), .ZN(n13461) );
  OR2_X1 U16676 ( .A1(n13446), .A2(n14653), .ZN(n13459) );
  NAND2_X1 U16677 ( .A1(n13448), .A2(n13447), .ZN(n14672) );
  INV_X1 U16678 ( .A(n14672), .ZN(n13449) );
  NAND2_X1 U16679 ( .A1(n13450), .A2(n13449), .ZN(n13455) );
  NAND2_X1 U16680 ( .A1(n13451), .A2(n14672), .ZN(n13454) );
  NAND2_X1 U16681 ( .A1(n15789), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13452) );
  MUX2_X1 U16682 ( .A(n13452), .B(n14658), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13453) );
  OAI211_X1 U16683 ( .C1(n13456), .C2(n13455), .A(n13454), .B(n13453), .ZN(
        n13457) );
  INV_X1 U16684 ( .A(n13457), .ZN(n13458) );
  NAND2_X1 U16685 ( .A1(n13459), .A2(n13458), .ZN(n14666) );
  MUX2_X1 U16686 ( .A(n14666), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15792), .Z(n15798) );
  AOI22_X1 U16687 ( .A1(n15798), .A2(n11284), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13467), .ZN(n13460) );
  OR2_X1 U16688 ( .A1(n13461), .A2(n13460), .ZN(n13468) );
  INV_X1 U16689 ( .A(n20322), .ZN(n20559) );
  NOR2_X1 U16690 ( .A1(n13462), .A2(n20559), .ZN(n13463) );
  XNOR2_X1 U16691 ( .A(n13463), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20057) );
  INV_X1 U16692 ( .A(n13464), .ZN(n13465) );
  NOR2_X1 U16693 ( .A1(n20057), .A2(n13465), .ZN(n16167) );
  MUX2_X1 U16694 ( .A(n16167), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n15792), .Z(n13466) );
  AOI22_X1 U16695 ( .A1(n13467), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n13466), .B2(n11284), .ZN(n13469) );
  NAND2_X1 U16696 ( .A1(n13468), .A2(n13469), .ZN(n15806) );
  NAND2_X1 U16697 ( .A1(n13469), .A2(n14661), .ZN(n13470) );
  NAND2_X1 U16698 ( .A1(n15806), .A2(n13470), .ZN(n15817) );
  NAND2_X1 U16699 ( .A1(n15817), .A2(n19982), .ZN(n13473) );
  INV_X1 U16700 ( .A(n13471), .ZN(n13472) );
  NAND2_X1 U16701 ( .A1(n13473), .A2(n13472), .ZN(n13474) );
  NAND2_X1 U16702 ( .A1(n13474), .A2(n20328), .ZN(n20835) );
  NOR2_X1 U16703 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n11284), .ZN(n20828) );
  NAND2_X1 U16704 ( .A1(n20682), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20605) );
  INV_X1 U16705 ( .A(n20605), .ZN(n13475) );
  NAND2_X1 U16706 ( .A1(n20606), .A2(n13475), .ZN(n20818) );
  OR2_X1 U16707 ( .A1(n20606), .A2(n20829), .ZN(n13476) );
  NAND2_X1 U16708 ( .A1(n20813), .A2(n20814), .ZN(n20557) );
  AND2_X1 U16709 ( .A1(n13476), .A2(n20557), .ZN(n20527) );
  MUX2_X1 U16710 ( .A(n20818), .B(n20527), .S(n20431), .Z(n13477) );
  OAI21_X1 U16711 ( .B1(n20828), .B2(n13446), .A(n13477), .ZN(n13478) );
  NAND2_X1 U16712 ( .A1(n20835), .A2(n13478), .ZN(n13479) );
  OAI21_X1 U16713 ( .B1(n20835), .B2(n20562), .A(n13479), .ZN(P1_U3476) );
  OAI21_X1 U16714 ( .B1(n13482), .B2(n13481), .A(n13596), .ZN(n14181) );
  NAND2_X1 U16715 ( .A1(n20157), .A2(DATAI_3_), .ZN(n13484) );
  NAND2_X1 U16716 ( .A1(n20156), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13483) );
  AND2_X1 U16717 ( .A1(n13484), .A2(n13483), .ZN(n20193) );
  OAI222_X1 U16718 ( .A1(n14181), .A2(n14354), .B1(n14353), .B2(n20193), .C1(
        n15972), .C2(n10613), .ZN(P1_U2901) );
  INV_X1 U16719 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13486) );
  NOR2_X1 U16720 ( .A1(n20042), .A2(n13486), .ZN(n13494) );
  AOI21_X1 U16721 ( .B1(n20132), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13494), .ZN(n13487) );
  OAI21_X1 U16722 ( .B1(n16029), .B2(n13746), .A(n13487), .ZN(n13488) );
  AOI21_X1 U16723 ( .B1(n13489), .B2(n20158), .A(n13488), .ZN(n13490) );
  OAI21_X1 U16724 ( .B1(n19981), .B2(n13500), .A(n13490), .ZN(P1_U2997) );
  NAND2_X1 U16725 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13491) );
  NAND2_X1 U16726 ( .A1(n16089), .A2(n14598), .ZN(n16131) );
  INV_X1 U16727 ( .A(n14598), .ZN(n14626) );
  INV_X1 U16728 ( .A(n14513), .ZN(n14621) );
  AOI21_X1 U16729 ( .B1(n11288), .B2(n16131), .A(n14621), .ZN(n13576) );
  OAI21_X1 U16730 ( .B1(n14642), .B2(n13491), .A(n13576), .ZN(n13498) );
  NAND3_X1 U16731 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14643), .A3(
        n13493), .ZN(n13496) );
  INV_X1 U16732 ( .A(n14642), .ZN(n14623) );
  AOI21_X1 U16733 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14509) );
  NAND2_X1 U16734 ( .A1(n14623), .A2(n14509), .ZN(n13575) );
  AOI21_X1 U16735 ( .B1(n20145), .B2(n13743), .A(n13494), .ZN(n13495) );
  NAND3_X1 U16736 ( .A1(n13496), .A2(n13575), .A3(n13495), .ZN(n13497) );
  AOI21_X1 U16737 ( .B1(n13498), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13497), .ZN(n13499) );
  OAI21_X1 U16738 ( .B1(n16160), .B2(n13500), .A(n13499), .ZN(P1_U3029) );
  OR2_X1 U16739 ( .A1(n13501), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13503) );
  NAND2_X1 U16740 ( .A1(n13503), .A2(n13502), .ZN(n13774) );
  OAI222_X1 U16741 ( .A1(n13774), .A2(n14280), .B1(n14278), .B2(n11292), .C1(
        n20138), .C2(n14277), .ZN(P1_U2872) );
  AOI21_X1 U16742 ( .B1(n13505), .B2(n13504), .A(n13579), .ZN(n13621) );
  INV_X1 U16743 ( .A(n13621), .ZN(n14176) );
  INV_X1 U16744 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13506) );
  OAI222_X1 U16745 ( .A1(n14176), .A2(n14280), .B1(n13506), .B2(n14278), .C1(
        n14181), .C2(n14277), .ZN(P1_U2869) );
  AOI21_X1 U16746 ( .B1(n13509), .B2(n13508), .A(n13507), .ZN(n16352) );
  INV_X1 U16747 ( .A(n16352), .ZN(n13891) );
  INV_X1 U16748 ( .A(n14804), .ZN(n13510) );
  OAI222_X1 U16749 ( .A1(n13891), .A2(n19138), .B1(n14836), .B2(n19224), .C1(
        n19180), .C2(n13510), .ZN(P2_U2906) );
  NOR2_X1 U16750 ( .A1(n13553), .A2(n13511), .ZN(n13590) );
  XNOR2_X1 U16751 ( .A(n13590), .B(n13589), .ZN(n13516) );
  NAND2_X1 U16752 ( .A1(n13560), .A2(n13512), .ZN(n13513) );
  AND2_X1 U16753 ( .A1(n13585), .A2(n13513), .ZN(n16297) );
  INV_X1 U16754 ( .A(n16297), .ZN(n16364) );
  MUX2_X1 U16755 ( .A(n16364), .B(n13514), .S(n14799), .Z(n13515) );
  OAI21_X1 U16756 ( .B1(n13516), .B2(n14785), .A(n13515), .ZN(P2_U2876) );
  XNOR2_X1 U16757 ( .A(n13518), .B(n13517), .ZN(n13623) );
  INV_X1 U16758 ( .A(n14181), .ZN(n13521) );
  NAND2_X1 U16759 ( .A1(n20135), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13619) );
  NAND2_X1 U16760 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13519) );
  OAI211_X1 U16761 ( .C1(n16029), .C2(n14173), .A(n13619), .B(n13519), .ZN(
        n13520) );
  AOI21_X1 U16762 ( .B1(n13521), .B2(n20158), .A(n13520), .ZN(n13522) );
  OAI21_X1 U16763 ( .B1(n13623), .B2(n19981), .A(n13522), .ZN(P1_U2996) );
  NOR2_X1 U16764 ( .A1(n13553), .A2(n13523), .ZN(n13592) );
  XNOR2_X1 U16765 ( .A(n13592), .B(n13524), .ZN(n13527) );
  OAI21_X1 U16766 ( .B1(n13587), .B2(n13525), .A(n13544), .ZN(n16355) );
  MUX2_X1 U16767 ( .A(n12526), .B(n16355), .S(n14790), .Z(n13526) );
  OAI21_X1 U16768 ( .B1(n13527), .B2(n14785), .A(n13526), .ZN(P2_U2874) );
  OR2_X1 U16769 ( .A1(n13528), .A2(n13507), .ZN(n13529) );
  NAND2_X1 U16770 ( .A1(n13529), .A2(n13570), .ZN(n19045) );
  INV_X1 U16771 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19222) );
  OAI222_X1 U16772 ( .A1(n19045), .A2(n19138), .B1(n14836), .B2(n19222), .C1(
        n19180), .C2(n13530), .ZN(P2_U2905) );
  XNOR2_X1 U16773 ( .A(n19943), .B(n19165), .ZN(n19167) );
  NOR2_X1 U16774 ( .A1(n19953), .A2(n19120), .ZN(n19174) );
  NOR2_X1 U16775 ( .A1(n19167), .A2(n19174), .ZN(n19166) );
  AOI21_X1 U16776 ( .B1(n19165), .B2(n19943), .A(n19166), .ZN(n19160) );
  XNOR2_X1 U16777 ( .A(n19936), .B(n13817), .ZN(n19161) );
  NOR2_X1 U16778 ( .A1(n19160), .A2(n19161), .ZN(n19159) );
  AOI21_X1 U16779 ( .B1(n13817), .B2(n19936), .A(n19159), .ZN(n19154) );
  OR2_X1 U16780 ( .A1(n13531), .A2(n9838), .ZN(n13534) );
  INV_X1 U16781 ( .A(n13532), .ZN(n13533) );
  NAND2_X1 U16782 ( .A1(n13534), .A2(n13533), .ZN(n16412) );
  XNOR2_X1 U16783 ( .A(n19565), .B(n16412), .ZN(n19155) );
  NOR2_X1 U16784 ( .A1(n19154), .A2(n19155), .ZN(n19153) );
  INV_X1 U16785 ( .A(n16412), .ZN(n19929) );
  NOR2_X1 U16786 ( .A1(n19930), .A2(n19929), .ZN(n13538) );
  OR2_X1 U16787 ( .A1(n13535), .A2(n13532), .ZN(n13537) );
  NAND2_X1 U16788 ( .A1(n13537), .A2(n13536), .ZN(n19099) );
  OAI21_X1 U16789 ( .B1(n19153), .B2(n13538), .A(n19099), .ZN(n19150) );
  XOR2_X1 U16790 ( .A(n19148), .B(n19150), .Z(n13543) );
  INV_X1 U16791 ( .A(n19099), .ZN(n13539) );
  AOI22_X1 U16792 ( .A1(n19173), .A2(n13539), .B1(n19172), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13542) );
  INV_X1 U16793 ( .A(n19180), .ZN(n13540) );
  NAND2_X1 U16794 ( .A1(n13540), .A2(n19298), .ZN(n13541) );
  OAI211_X1 U16795 ( .C1(n13543), .C2(n19168), .A(n13542), .B(n13541), .ZN(
        P2_U2915) );
  AOI21_X1 U16796 ( .B1(n13545), .B2(n13544), .A(n13793), .ZN(n19041) );
  INV_X1 U16797 ( .A(n19041), .ZN(n15052) );
  AND2_X1 U16798 ( .A1(n13393), .A2(n13546), .ZN(n13549) );
  NAND2_X1 U16799 ( .A1(n13393), .A2(n13547), .ZN(n13792) );
  OAI211_X1 U16800 ( .C1(n13549), .C2(n13548), .A(n14798), .B(n13792), .ZN(
        n13551) );
  NAND2_X1 U16801 ( .A1(n14799), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13550) );
  OAI211_X1 U16802 ( .C1(n15052), .C2(n14799), .A(n13551), .B(n13550), .ZN(
        P2_U2873) );
  OR2_X1 U16803 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  AOI211_X1 U16804 ( .C1(n13555), .C2(n13554), .A(n14785), .B(n13590), .ZN(
        n13556) );
  INV_X1 U16805 ( .A(n13556), .ZN(n13562) );
  OR2_X1 U16806 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  NAND2_X1 U16807 ( .A1(n13560), .A2(n13559), .ZN(n19066) );
  OR2_X1 U16808 ( .A1(n14799), .A2(n19066), .ZN(n13561) );
  OAI211_X1 U16809 ( .C1(n14790), .C2(n12516), .A(n13562), .B(n13561), .ZN(
        P2_U2877) );
  AND2_X1 U16810 ( .A1(n13595), .A2(n13563), .ZN(n13564) );
  OR2_X1 U16811 ( .A1(n13712), .A2(n13564), .ZN(n16032) );
  NAND2_X1 U16812 ( .A1(n13577), .A2(n13565), .ZN(n13566) );
  AND2_X1 U16813 ( .A1(n13787), .A2(n13566), .ZN(n20037) );
  AOI22_X1 U16814 ( .A1(n14268), .A2(n20037), .B1(n14267), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13567) );
  OAI21_X1 U16815 ( .B1(n16032), .B2(n14277), .A(n13567), .ZN(P1_U2867) );
  NAND2_X1 U16816 ( .A1(n20157), .A2(DATAI_5_), .ZN(n13569) );
  NAND2_X1 U16817 ( .A1(n20156), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13568) );
  AND2_X1 U16818 ( .A1(n13569), .A2(n13568), .ZN(n20208) );
  INV_X1 U16819 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20087) );
  OAI222_X1 U16820 ( .A1(n16032), .A2(n14354), .B1(n14353), .B2(n20208), .C1(
        n15972), .C2(n20087), .ZN(P1_U2899) );
  XNOR2_X1 U16821 ( .A(n13571), .B(n13570), .ZN(n19035) );
  INV_X1 U16822 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19220) );
  OAI222_X1 U16823 ( .A1(n19035), .A2(n19138), .B1(n14836), .B2(n19220), .C1(
        n13572), .C2(n19180), .ZN(P2_U2904) );
  XNOR2_X1 U16824 ( .A(n13574), .B(n13573), .ZN(n13603) );
  OAI211_X1 U16825 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n16113), .A(
        n13576), .B(n13575), .ZN(n13617) );
  OAI21_X1 U16826 ( .B1(n13579), .B2(n13578), .A(n13577), .ZN(n20061) );
  NAND3_X1 U16827 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14643), .ZN(n16132) );
  NAND2_X1 U16828 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14510) );
  OAI211_X1 U16829 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n16156), .B(n14510), .ZN(n13581) );
  INV_X1 U16830 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20765) );
  NOR2_X1 U16831 ( .A1(n20042), .A2(n20765), .ZN(n13599) );
  INV_X1 U16832 ( .A(n13599), .ZN(n13580) );
  OAI211_X1 U16833 ( .C1(n16135), .C2(n20061), .A(n13581), .B(n13580), .ZN(
        n13582) );
  AOI21_X1 U16834 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13617), .A(
        n13582), .ZN(n13583) );
  OAI21_X1 U16835 ( .B1(n16160), .B2(n13603), .A(n13583), .ZN(P1_U3027) );
  AND2_X1 U16836 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  OR2_X1 U16837 ( .A1(n13587), .A2(n13586), .ZN(n19052) );
  AOI21_X1 U16838 ( .B1(n13590), .B2(n13589), .A(n13588), .ZN(n13591) );
  OR3_X1 U16839 ( .A1(n13592), .A2(n13591), .A3(n14785), .ZN(n13594) );
  NAND2_X1 U16840 ( .A1(n14799), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13593) );
  OAI211_X1 U16841 ( .C1(n19052), .C2(n14799), .A(n13594), .B(n13593), .ZN(
        P2_U2875) );
  AOI21_X1 U16842 ( .B1(n13597), .B2(n13596), .A(n9975), .ZN(n20068) );
  INV_X1 U16843 ( .A(n13598), .ZN(n20055) );
  AOI21_X1 U16844 ( .B1(n20132), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13599), .ZN(n13600) );
  OAI21_X1 U16845 ( .B1(n16029), .B2(n20055), .A(n13600), .ZN(n13601) );
  AOI21_X1 U16846 ( .B1(n20068), .B2(n20158), .A(n13601), .ZN(n13602) );
  OAI21_X1 U16847 ( .B1(n19981), .B2(n13603), .A(n13602), .ZN(P1_U2995) );
  INV_X1 U16848 ( .A(n20068), .ZN(n13737) );
  NAND2_X1 U16849 ( .A1(n20157), .A2(DATAI_4_), .ZN(n13605) );
  NAND2_X1 U16850 ( .A1(n20156), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13604) );
  AND2_X1 U16851 ( .A1(n13605), .A2(n13604), .ZN(n20200) );
  INV_X1 U16852 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20089) );
  OAI222_X1 U16853 ( .A1(n13737), .A2(n14354), .B1(n14353), .B2(n20200), .C1(
        n20089), .C2(n15972), .ZN(P1_U2900) );
  INV_X1 U16854 ( .A(n13758), .ZN(n19116) );
  AOI22_X1 U16855 ( .A1(n19108), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19116), .B2(n12939), .ZN(n13869) );
  OR2_X1 U16856 ( .A1(n13607), .A2(n13606), .ZN(n13611) );
  INV_X1 U16857 ( .A(n12464), .ZN(n13609) );
  AND2_X1 U16858 ( .A1(n13609), .A2(n13608), .ZN(n14001) );
  MUX2_X1 U16859 ( .A(n14001), .B(n13999), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13610) );
  AND2_X1 U16860 ( .A1(n13611), .A2(n13610), .ZN(n16427) );
  INV_X1 U16861 ( .A(n16474), .ZN(n14006) );
  OAI22_X1 U16862 ( .A1(n16427), .A2(n19924), .B1(n13612), .B2(n14006), .ZN(
        n13613) );
  AOI21_X1 U16863 ( .B1(n13869), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n13613), 
        .ZN(n13615) );
  NAND2_X1 U16864 ( .A1(n13995), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13614) );
  OAI21_X1 U16865 ( .B1(n13615), .B2(n13995), .A(n13614), .ZN(P2_U3601) );
  AOI22_X1 U16866 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13617), .B1(
        n16156), .B2(n13616), .ZN(n13618) );
  NAND2_X1 U16867 ( .A1(n13619), .A2(n13618), .ZN(n13620) );
  AOI21_X1 U16868 ( .B1(n20145), .B2(n13621), .A(n13620), .ZN(n13622) );
  OAI21_X1 U16869 ( .B1(n13623), .B2(n16160), .A(n13622), .ZN(P1_U3028) );
  INV_X1 U16870 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13631) );
  INV_X1 U16871 ( .A(n20110), .ZN(n13630) );
  INV_X1 U16872 ( .A(DATAI_15_), .ZN(n13628) );
  INV_X1 U16873 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13627) );
  MUX2_X1 U16874 ( .A(n13628), .B(n13627), .S(n20156), .Z(n14346) );
  INV_X1 U16875 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13629) );
  OAI222_X1 U16876 ( .A1(n13680), .A2(n13631), .B1(n13630), .B2(n14346), .C1(
        n13629), .C2(n13681), .ZN(P1_U2967) );
  NAND2_X1 U16877 ( .A1(n12939), .A2(n13632), .ZN(n13633) );
  XNOR2_X1 U16878 ( .A(n16326), .B(n13633), .ZN(n13634) );
  NAND2_X1 U16879 ( .A1(n13634), .A2(n19080), .ZN(n13643) );
  OAI21_X1 U16880 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n16395) );
  AOI22_X1 U16881 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19130), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19117), .ZN(n13638) );
  OAI211_X1 U16882 ( .C1(n19100), .C2(n16395), .A(n13638), .B(n19058), .ZN(
        n13641) );
  OAI22_X1 U16883 ( .A1(n13639), .A2(n19090), .B1(n19105), .B2(n16332), .ZN(
        n13640) );
  AOI211_X1 U16884 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19122), .A(n13641), .B(
        n13640), .ZN(n13642) );
  NAND2_X1 U16885 ( .A1(n13643), .A2(n13642), .ZN(P2_U2850) );
  INV_X1 U16886 ( .A(n13824), .ZN(n19123) );
  NAND2_X1 U16887 ( .A1(n12939), .A2(n13644), .ZN(n13645) );
  XNOR2_X1 U16888 ( .A(n13675), .B(n13645), .ZN(n13646) );
  NAND2_X1 U16889 ( .A1(n13646), .A2(n19080), .ZN(n13654) );
  OAI22_X1 U16890 ( .A1(n13673), .A2(n19024), .B1(n19872), .B2(n19059), .ZN(
        n13649) );
  NOR2_X1 U16891 ( .A1(n19090), .A2(n13647), .ZN(n13648) );
  AOI211_X1 U16892 ( .C1(n19929), .C2(n19121), .A(n13649), .B(n13648), .ZN(
        n13650) );
  OAI21_X1 U16893 ( .B1(n19101), .B2(n13651), .A(n13650), .ZN(n13652) );
  AOI21_X1 U16894 ( .B1(n13120), .B2(n19119), .A(n13652), .ZN(n13653) );
  OAI211_X1 U16895 ( .C1(n19565), .C2(n19123), .A(n13654), .B(n13653), .ZN(
        P2_U2852) );
  INV_X1 U16896 ( .A(n13655), .ZN(n13666) );
  NAND2_X1 U16897 ( .A1(n12939), .A2(n13656), .ZN(n13657) );
  XNOR2_X1 U16898 ( .A(n16309), .B(n13657), .ZN(n13658) );
  NAND2_X1 U16899 ( .A1(n13658), .A2(n19080), .ZN(n13665) );
  INV_X1 U16900 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U16901 ( .B1(n19878), .B2(n19059), .A(n19058), .ZN(n13659) );
  AOI21_X1 U16902 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19130), .A(
        n13659), .ZN(n13660) );
  OAI21_X1 U16903 ( .B1(n19100), .B2(n13661), .A(n13660), .ZN(n13663) );
  NOR2_X1 U16904 ( .A1(n19101), .A2(n12512), .ZN(n13662) );
  AOI211_X1 U16905 ( .C1(n16310), .C2(n19119), .A(n13663), .B(n13662), .ZN(
        n13664) );
  OAI211_X1 U16906 ( .C1(n19090), .C2(n13666), .A(n13665), .B(n13664), .ZN(
        P2_U2846) );
  NAND2_X1 U16907 ( .A1(n13668), .A2(n13667), .ZN(n13669) );
  XOR2_X1 U16908 ( .A(n13670), .B(n13669), .Z(n16424) );
  XNOR2_X1 U16909 ( .A(n13672), .B(n13671), .ZN(n16421) );
  OAI22_X1 U16910 ( .A1(n16338), .A2(n13673), .B1(n19872), .B2(n19058), .ZN(
        n13674) );
  AOI21_X1 U16911 ( .B1(n16327), .B2(n13675), .A(n13674), .ZN(n13677) );
  NAND2_X1 U16912 ( .A1(n13120), .A2(n19263), .ZN(n13676) );
  OAI211_X1 U16913 ( .C1(n16421), .C2(n19257), .A(n13677), .B(n13676), .ZN(
        n13678) );
  AOI21_X1 U16914 ( .B1(n16424), .B2(n16335), .A(n13678), .ZN(n13679) );
  INV_X1 U16915 ( .A(n13679), .ZN(P2_U3011) );
  AOI22_X1 U16916 ( .A1(n20119), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20118), .ZN(n13684) );
  NAND2_X1 U16917 ( .A1(n20157), .A2(DATAI_6_), .ZN(n13683) );
  NAND2_X1 U16918 ( .A1(n20156), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13682) );
  AND2_X1 U16919 ( .A1(n13683), .A2(n13682), .ZN(n20215) );
  INV_X1 U16920 ( .A(n20215), .ZN(n14320) );
  NAND2_X1 U16921 ( .A1(n20110), .A2(n14320), .ZN(n13704) );
  NAND2_X1 U16922 ( .A1(n13684), .A2(n13704), .ZN(P1_U2958) );
  AOI22_X1 U16923 ( .A1(n20119), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20118), .ZN(n13685) );
  INV_X1 U16924 ( .A(n20193), .ZN(n14330) );
  NAND2_X1 U16925 ( .A1(n20110), .A2(n14330), .ZN(n13698) );
  NAND2_X1 U16926 ( .A1(n13685), .A2(n13698), .ZN(P1_U2955) );
  AOI22_X1 U16927 ( .A1(n20119), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20118), .ZN(n13686) );
  INV_X1 U16928 ( .A(n20185), .ZN(n14333) );
  NAND2_X1 U16929 ( .A1(n20110), .A2(n14333), .ZN(n13696) );
  NAND2_X1 U16930 ( .A1(n13686), .A2(n13696), .ZN(P1_U2939) );
  AOI22_X1 U16931 ( .A1(n20119), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20118), .ZN(n13687) );
  INV_X1 U16932 ( .A(n20208), .ZN(n14324) );
  NAND2_X1 U16933 ( .A1(n20110), .A2(n14324), .ZN(n13702) );
  NAND2_X1 U16934 ( .A1(n13687), .A2(n13702), .ZN(P1_U2957) );
  AOI22_X1 U16935 ( .A1(n20119), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20118), .ZN(n13688) );
  INV_X1 U16936 ( .A(n20200), .ZN(n14327) );
  NAND2_X1 U16937 ( .A1(n20110), .A2(n14327), .ZN(n13700) );
  NAND2_X1 U16938 ( .A1(n13688), .A2(n13700), .ZN(P1_U2941) );
  AOI22_X1 U16939 ( .A1(n20119), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20118), .ZN(n13691) );
  NAND2_X1 U16940 ( .A1(n20157), .A2(DATAI_7_), .ZN(n13690) );
  NAND2_X1 U16941 ( .A1(n20156), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13689) );
  INV_X1 U16942 ( .A(n20227), .ZN(n14316) );
  NAND2_X1 U16943 ( .A1(n20110), .A2(n14316), .ZN(n13706) );
  NAND2_X1 U16944 ( .A1(n13691), .A2(n13706), .ZN(P1_U2959) );
  AOI22_X1 U16945 ( .A1(n20119), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20118), .ZN(n13692) );
  INV_X1 U16946 ( .A(n20163), .ZN(n14341) );
  NAND2_X1 U16947 ( .A1(n20110), .A2(n14341), .ZN(n13693) );
  NAND2_X1 U16948 ( .A1(n13692), .A2(n13693), .ZN(P1_U2952) );
  AOI22_X1 U16949 ( .A1(n20119), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20118), .ZN(n13694) );
  NAND2_X1 U16950 ( .A1(n13694), .A2(n13693), .ZN(P1_U2937) );
  AOI22_X1 U16951 ( .A1(n20119), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20118), .ZN(n13695) );
  INV_X1 U16952 ( .A(n20179), .ZN(n14337) );
  NAND2_X1 U16953 ( .A1(n20110), .A2(n14337), .ZN(n13708) );
  NAND2_X1 U16954 ( .A1(n13695), .A2(n13708), .ZN(P1_U2938) );
  AOI22_X1 U16955 ( .A1(n20119), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20118), .ZN(n13697) );
  NAND2_X1 U16956 ( .A1(n13697), .A2(n13696), .ZN(P1_U2954) );
  AOI22_X1 U16957 ( .A1(n20119), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20118), .ZN(n13699) );
  NAND2_X1 U16958 ( .A1(n13699), .A2(n13698), .ZN(P1_U2940) );
  AOI22_X1 U16959 ( .A1(n20119), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20118), .ZN(n13701) );
  NAND2_X1 U16960 ( .A1(n13701), .A2(n13700), .ZN(P1_U2956) );
  AOI22_X1 U16961 ( .A1(n20119), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20118), .ZN(n13703) );
  NAND2_X1 U16962 ( .A1(n13703), .A2(n13702), .ZN(P1_U2942) );
  AOI22_X1 U16963 ( .A1(n20119), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20118), .ZN(n13705) );
  NAND2_X1 U16964 ( .A1(n13705), .A2(n13704), .ZN(P1_U2943) );
  AOI22_X1 U16965 ( .A1(n20119), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20118), .ZN(n13707) );
  NAND2_X1 U16966 ( .A1(n13707), .A2(n13706), .ZN(P1_U2944) );
  AOI22_X1 U16967 ( .A1(n20119), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20118), .ZN(n13709) );
  NAND2_X1 U16968 ( .A1(n13709), .A2(n13708), .ZN(P1_U2953) );
  OR2_X1 U16969 ( .A1(n13712), .A2(n13711), .ZN(n13713) );
  AND2_X1 U16970 ( .A1(n13710), .A2(n13713), .ZN(n20032) );
  INV_X1 U16971 ( .A(n20032), .ZN(n13738) );
  XNOR2_X1 U16972 ( .A(n13787), .B(n13783), .ZN(n20026) );
  AOI22_X1 U16973 ( .A1(n20026), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n13714) );
  OAI21_X1 U16974 ( .B1(n13738), .B2(n14270), .A(n13714), .ZN(P1_U2866) );
  NAND2_X1 U16975 ( .A1(n12939), .A2(n13715), .ZN(n13716) );
  XNOR2_X1 U16976 ( .A(n16292), .B(n13716), .ZN(n13723) );
  INV_X1 U16977 ( .A(n19090), .ZN(n19125) );
  AOI22_X1 U16978 ( .A1(n13717), .A2(n19125), .B1(P2_EBX_REG_11__SCAN_IN), 
        .B2(n19117), .ZN(n13718) );
  OAI21_X1 U16979 ( .B1(n16308), .B2(n19024), .A(n13718), .ZN(n13722) );
  AOI21_X1 U16980 ( .B1(n19121), .B2(n16363), .A(n19103), .ZN(n13720) );
  NAND2_X1 U16981 ( .A1(n19122), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n13719) );
  OAI211_X1 U16982 ( .C1(n16364), .C2(n19105), .A(n13720), .B(n13719), .ZN(
        n13721) );
  AOI211_X1 U16983 ( .C1(n13723), .C2(n19080), .A(n13722), .B(n13721), .ZN(
        n13724) );
  INV_X1 U16984 ( .A(n13724), .ZN(P2_U2844) );
  NAND2_X1 U16985 ( .A1(n12939), .A2(n13725), .ZN(n13726) );
  XNOR2_X1 U16986 ( .A(n16316), .B(n13726), .ZN(n13735) );
  AOI22_X1 U16987 ( .A1(n19125), .A2(n13727), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19117), .ZN(n13728) );
  OAI21_X1 U16988 ( .B1(n16325), .B2(n19024), .A(n13728), .ZN(n13734) );
  AOI21_X1 U16989 ( .B1(n13730), .B2(n13729), .A(n13123), .ZN(n19142) );
  INV_X1 U16990 ( .A(n19142), .ZN(n15333) );
  OAI21_X1 U16991 ( .B1(n19100), .B2(n15333), .A(n19058), .ZN(n13731) );
  AOI21_X1 U16992 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n19122), .A(n13731), .ZN(
        n13732) );
  OAI21_X1 U16993 ( .B1(n19105), .B2(n15334), .A(n13732), .ZN(n13733) );
  AOI211_X1 U16994 ( .C1(n13735), .C2(n19080), .A(n13734), .B(n13733), .ZN(
        n13736) );
  INV_X1 U16995 ( .A(n13736), .ZN(P2_U2848) );
  OAI222_X1 U16996 ( .A1(n20061), .A2(n14280), .B1(n14278), .B2(n11301), .C1(
        n14277), .C2(n13737), .ZN(P1_U2868) );
  OAI222_X1 U16997 ( .A1(n13738), .A2(n14354), .B1(n14353), .B2(n20215), .C1(
        n15972), .C2(n10690), .ZN(P1_U2898) );
  INV_X1 U16998 ( .A(n10451), .ZN(n13739) );
  NOR2_X1 U16999 ( .A1(n13742), .A2(n13739), .ZN(n13740) );
  OR2_X1 U17000 ( .A1(n20031), .A2(n13740), .ZN(n20067) );
  OAI21_X1 U17001 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20021), .A(n14158), .ZN(
        n14169) );
  OR2_X1 U17002 ( .A1(n13742), .A2(n13741), .ZN(n20056) );
  NOR2_X1 U17003 ( .A1(n13446), .A2(n20056), .ZN(n13753) );
  NAND2_X1 U17004 ( .A1(n20027), .A2(n13743), .ZN(n13751) );
  NAND2_X1 U17005 ( .A1(n20046), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13750) );
  NAND2_X1 U17006 ( .A1(n20019), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20063) );
  NOR2_X1 U17007 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20063), .ZN(n14170) );
  AOI21_X1 U17008 ( .B1(n20059), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14170), .ZN(n13749) );
  AND2_X1 U17009 ( .A1(n13744), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13745) );
  INV_X1 U17010 ( .A(n13746), .ZN(n13747) );
  NAND2_X1 U17011 ( .A1(n20040), .A2(n13747), .ZN(n13748) );
  NAND4_X1 U17012 ( .A1(n13751), .A2(n13750), .A3(n13749), .A4(n13748), .ZN(
        n13752) );
  AOI211_X1 U17013 ( .C1(n14169), .C2(P1_REIP_REG_2__SCAN_IN), .A(n13753), .B(
        n13752), .ZN(n13754) );
  OAI21_X1 U17014 ( .B1(n14190), .B2(n13755), .A(n13754), .ZN(P1_U2838) );
  NOR2_X1 U17015 ( .A1(n19108), .A2(n13756), .ZN(n13820) );
  OAI21_X1 U17016 ( .B1(n13758), .B2(n13757), .A(n13820), .ZN(n13867) );
  OAI21_X1 U17017 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12939), .A(
        n13867), .ZN(n13759) );
  NAND2_X1 U17018 ( .A1(n13759), .A2(n19080), .ZN(n13768) );
  INV_X1 U17019 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19867) );
  OAI22_X1 U17020 ( .A1(n19165), .A2(n19100), .B1(n19867), .B2(n19059), .ZN(
        n13766) );
  INV_X1 U17021 ( .A(n13760), .ZN(n13762) );
  AOI22_X1 U17022 ( .A1(n19125), .A2(n13762), .B1(n19130), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13763) );
  OAI21_X1 U17023 ( .B1(n19101), .B2(n13764), .A(n13763), .ZN(n13765) );
  AOI211_X1 U17024 ( .C1(n19119), .C2(n14005), .A(n13766), .B(n13765), .ZN(
        n13767) );
  OAI211_X1 U17025 ( .C1(n19943), .C2(n19123), .A(n13768), .B(n13767), .ZN(
        P2_U2854) );
  NAND2_X1 U17026 ( .A1(n13710), .A2(n13770), .ZN(n13771) );
  AND2_X1 U17027 ( .A1(n13769), .A2(n13771), .ZN(n20022) );
  INV_X1 U17028 ( .A(n20022), .ZN(n13773) );
  OAI222_X1 U17029 ( .A1(n13773), .A2(n14354), .B1(n14353), .B2(n20227), .C1(
        n13772), .C2(n15972), .ZN(P1_U2897) );
  INV_X1 U17030 ( .A(n13774), .ZN(n20144) );
  INV_X1 U17031 ( .A(n10570), .ZN(n20827) );
  NAND2_X1 U17032 ( .A1(n20046), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13776) );
  OAI21_X1 U17033 ( .B1(n20059), .B2(n20040), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13775) );
  OAI211_X1 U17034 ( .C1(n20056), .C2(n20827), .A(n13776), .B(n13775), .ZN(
        n13780) );
  INV_X1 U17035 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13777) );
  NOR2_X1 U17036 ( .A1(n13778), .A2(n13777), .ZN(n13779) );
  AOI211_X1 U17037 ( .C1(n20144), .C2(n20027), .A(n13780), .B(n13779), .ZN(
        n13781) );
  OAI21_X1 U17038 ( .B1(n14190), .B2(n20138), .A(n13781), .ZN(P1_U2840) );
  NAND2_X1 U17039 ( .A1(n20022), .A2(n13782), .ZN(n13790) );
  INV_X1 U17040 ( .A(n13783), .ZN(n13786) );
  INV_X1 U17041 ( .A(n13784), .ZN(n13785) );
  OAI21_X1 U17042 ( .B1(n13787), .B2(n13786), .A(n13785), .ZN(n13788) );
  AND2_X1 U17043 ( .A1(n13788), .A2(n13858), .ZN(n20016) );
  NAND2_X1 U17044 ( .A1(n20016), .A2(n14268), .ZN(n13789) );
  OAI211_X1 U17045 ( .C1(n20011), .C2(n14278), .A(n13790), .B(n13789), .ZN(
        P1_U2865) );
  XNOR2_X1 U17046 ( .A(n13792), .B(n13791), .ZN(n13798) );
  OR2_X1 U17047 ( .A1(n13794), .A2(n13793), .ZN(n13795) );
  AND2_X1 U17048 ( .A1(n13849), .A2(n13795), .ZN(n16275) );
  INV_X1 U17049 ( .A(n16275), .ZN(n19023) );
  INV_X1 U17050 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13796) );
  MUX2_X1 U17051 ( .A(n19023), .B(n13796), .S(n14799), .Z(n13797) );
  OAI21_X1 U17052 ( .B1(n13798), .B2(n14785), .A(n13797), .ZN(P2_U2872) );
  OAI21_X1 U17053 ( .B1(n13801), .B2(n13800), .A(n13830), .ZN(n13853) );
  NOR2_X1 U17054 ( .A1(n13804), .A2(n13803), .ZN(n13805) );
  OR2_X1 U17055 ( .A1(n13802), .A2(n13805), .ZN(n19015) );
  AOI22_X1 U17056 ( .A1(n19134), .A2(BUF2_REG_16__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U17057 ( .A1(n16265), .A2(n13806), .B1(n19172), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n13807) );
  OAI211_X1 U17058 ( .C1(n16267), .C2(n19015), .A(n13808), .B(n13807), .ZN(
        n13809) );
  INV_X1 U17059 ( .A(n13809), .ZN(n13810) );
  OAI21_X1 U17060 ( .B1(n13853), .B2(n19168), .A(n13810), .ZN(P2_U2903) );
  AOI22_X1 U17061 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19130), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19122), .ZN(n13812) );
  NAND2_X1 U17062 ( .A1(n19117), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n13811) );
  OAI211_X1 U17063 ( .C1(n19090), .C2(n13813), .A(n13812), .B(n13811), .ZN(
        n13814) );
  INV_X1 U17064 ( .A(n13814), .ZN(n13816) );
  NAND2_X1 U17065 ( .A1(n13176), .A2(n19119), .ZN(n13815) );
  OAI211_X1 U17066 ( .C1(n13817), .C2(n19100), .A(n13816), .B(n13815), .ZN(
        n13823) );
  INV_X1 U17067 ( .A(n13820), .ZN(n13818) );
  AOI221_X1 U17068 ( .B1(n13821), .B2(n13820), .C1(n13819), .C2(n13818), .A(
        n19841), .ZN(n13822) );
  AOI211_X1 U17069 ( .C1(n13825), .C2(n13824), .A(n13823), .B(n13822), .ZN(
        n13826) );
  INV_X1 U17070 ( .A(n13826), .ZN(P2_U2853) );
  OR2_X1 U17071 ( .A1(n13851), .A2(n13827), .ZN(n13828) );
  AND2_X1 U17072 ( .A1(n13929), .A2(n13828), .ZN(n15032) );
  INV_X1 U17073 ( .A(n15032), .ZN(n15252) );
  INV_X1 U17074 ( .A(n13926), .ZN(n13829) );
  AOI21_X1 U17075 ( .B1(n13831), .B2(n13830), .A(n13829), .ZN(n13907) );
  NAND2_X1 U17076 ( .A1(n13907), .A2(n14798), .ZN(n13833) );
  NAND2_X1 U17077 ( .A1(n14799), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13832) );
  OAI211_X1 U17078 ( .C1(n15252), .C2(n14799), .A(n13833), .B(n13832), .ZN(
        P2_U2870) );
  XNOR2_X1 U17079 ( .A(n13834), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13836) );
  XNOR2_X1 U17080 ( .A(n13836), .B(n13835), .ZN(n19258) );
  OAI21_X1 U17081 ( .B1(n15259), .B2(n13838), .A(n13837), .ZN(n13839) );
  INV_X1 U17082 ( .A(n13839), .ZN(n16426) );
  NAND2_X1 U17083 ( .A1(n16426), .A2(n16411), .ZN(n16397) );
  INV_X1 U17084 ( .A(n16403), .ZN(n13841) );
  OAI22_X1 U17085 ( .A1(n16413), .A2(n19099), .B1(n12321), .B2(n19058), .ZN(
        n13840) );
  AOI21_X1 U17086 ( .B1(n13841), .B2(n16405), .A(n13840), .ZN(n13842) );
  OAI21_X1 U17087 ( .B1(n16388), .B2(n19104), .A(n13842), .ZN(n13846) );
  XNOR2_X1 U17088 ( .A(n13844), .B(n13843), .ZN(n19260) );
  NOR2_X1 U17089 ( .A1(n19260), .A2(n16393), .ZN(n13845) );
  AOI211_X1 U17090 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n16397), .A(
        n13846), .B(n13845), .ZN(n13847) );
  OAI21_X1 U17091 ( .B1(n16420), .B2(n19258), .A(n13847), .ZN(P2_U3042) );
  AND2_X1 U17092 ( .A1(n13849), .A2(n13848), .ZN(n13850) );
  OR2_X1 U17093 ( .A1(n13851), .A2(n13850), .ZN(n19014) );
  MUX2_X1 U17094 ( .A(n19014), .B(n11662), .S(n14799), .Z(n13852) );
  OAI21_X1 U17095 ( .B1(n13853), .B2(n14785), .A(n13852), .ZN(P2_U2871) );
  INV_X1 U17096 ( .A(n13854), .ZN(n13855) );
  AOI21_X1 U17097 ( .B1(n13856), .B2(n13769), .A(n13855), .ZN(n13915) );
  INV_X1 U17098 ( .A(n13915), .ZN(n13889) );
  OAI21_X1 U17099 ( .B1(n20021), .B2(n20000), .A(n14158), .ZN(n20005) );
  AND2_X1 U17100 ( .A1(n13858), .A2(n13857), .ZN(n13859) );
  OR2_X1 U17101 ( .A1(n13859), .A2(n13946), .ZN(n16136) );
  NOR2_X1 U17102 ( .A1(n20021), .A2(n20018), .ZN(n20038) );
  NOR2_X1 U17103 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13860), .ZN(n13861) );
  AOI22_X1 U17104 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20059), .B1(
        n20038), .B2(n13861), .ZN(n13862) );
  OAI211_X1 U17105 ( .C1(n20062), .C2(n16136), .A(n13862), .B(n20042), .ZN(
        n13863) );
  AOI21_X1 U17106 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20005), .A(n13863), .ZN(
        n13866) );
  INV_X1 U17107 ( .A(n13913), .ZN(n13864) );
  AOI22_X1 U17108 ( .A1(n20046), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n13864), .B2(
        n20040), .ZN(n13865) );
  OAI211_X1 U17109 ( .C1(n13889), .C2(n15890), .A(n13866), .B(n13865), .ZN(
        P1_U2832) );
  OAI21_X1 U17110 ( .B1(n12939), .B2(n13868), .A(n13867), .ZN(n13998) );
  NOR2_X1 U17111 ( .A1(n13869), .A2(n16467), .ZN(n13996) );
  NAND2_X1 U17112 ( .A1(n13870), .A2(n14000), .ZN(n13873) );
  MUX2_X1 U17113 ( .A(n13873), .B(n13872), .S(n13871), .Z(n13880) );
  NAND2_X1 U17114 ( .A1(n13874), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13879) );
  NAND3_X1 U17115 ( .A1(n13876), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n13875), .ZN(n13877) );
  NAND4_X1 U17116 ( .A1(n13880), .A2(n13879), .A3(n13878), .A4(n13877), .ZN(
        n13881) );
  AOI21_X1 U17117 ( .B1(n13176), .B2(n14004), .A(n13881), .ZN(n16434) );
  OAI22_X1 U17118 ( .A1(n19936), .A2(n14006), .B1(n19924), .B2(n16434), .ZN(
        n13882) );
  AOI21_X1 U17119 ( .B1(n13998), .B2(n13996), .A(n13882), .ZN(n13883) );
  MUX2_X1 U17120 ( .A(n13883), .B(n16435), .S(n13995), .Z(n13884) );
  INV_X1 U17121 ( .A(n13884), .ZN(P2_U3599) );
  INV_X1 U17122 ( .A(DATAI_8_), .ZN(n13886) );
  NAND2_X1 U17123 ( .A1(n20156), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13885) );
  OAI21_X1 U17124 ( .B1(n20156), .B2(n13886), .A(n13885), .ZN(n20097) );
  INV_X1 U17125 ( .A(n20097), .ZN(n13888) );
  OAI222_X1 U17126 ( .A1(n13889), .A2(n14354), .B1(n14353), .B2(n13888), .C1(
        n13887), .C2(n15972), .ZN(P1_U2896) );
  OAI222_X1 U17127 ( .A1(n16136), .A2(n14280), .B1(n14278), .B2(n11319), .C1(
        n14277), .C2(n13889), .ZN(P1_U2864) );
  NOR2_X1 U17128 ( .A1(n19841), .A2(n12939), .ZN(n19022) );
  AOI22_X1 U17129 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19130), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19122), .ZN(n13890) );
  OAI211_X1 U17130 ( .C1(n19100), .C2(n13891), .A(n13890), .B(n19058), .ZN(
        n13893) );
  NOR2_X1 U17131 ( .A1(n16355), .A2(n19105), .ZN(n13892) );
  AOI211_X1 U17132 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n19117), .A(n13893), .B(
        n13892), .ZN(n13894) );
  OAI21_X1 U17133 ( .B1(n13895), .B2(n19090), .A(n13894), .ZN(n13899) );
  OR2_X1 U17134 ( .A1(n19108), .A2(n13896), .ZN(n19040) );
  AOI211_X1 U17135 ( .C1(n16279), .C2(n13897), .A(n19841), .B(n19040), .ZN(
        n13898) );
  AOI211_X1 U17136 ( .C1(n19022), .C2(n16279), .A(n13899), .B(n13898), .ZN(
        n13900) );
  INV_X1 U17137 ( .A(n13900), .ZN(P2_U2842) );
  NOR2_X1 U17138 ( .A1(n13802), .A2(n13901), .ZN(n13902) );
  NOR2_X1 U17139 ( .A1(n13934), .A2(n13902), .ZN(n15258) );
  INV_X1 U17140 ( .A(n15258), .ZN(n14706) );
  AOI22_X1 U17141 ( .A1(n19134), .A2(BUF2_REG_17__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13905) );
  AOI22_X1 U17142 ( .A1(n16265), .A2(n13903), .B1(n19172), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13904) );
  OAI211_X1 U17143 ( .C1(n16267), .C2(n14706), .A(n13905), .B(n13904), .ZN(
        n13906) );
  AOI21_X1 U17144 ( .B1(n13907), .B2(n19175), .A(n13906), .ZN(n13908) );
  INV_X1 U17145 ( .A(n13908), .ZN(P2_U2902) );
  XOR2_X1 U17146 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13909), .Z(
        n13910) );
  XNOR2_X1 U17147 ( .A(n13911), .B(n13910), .ZN(n16134) );
  AOI22_X1 U17148 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13912) );
  OAI21_X1 U17149 ( .B1(n16029), .B2(n13913), .A(n13912), .ZN(n13914) );
  AOI21_X1 U17150 ( .B1(n13915), .B2(n20158), .A(n13914), .ZN(n13916) );
  OAI21_X1 U17151 ( .B1(n16134), .B2(n19981), .A(n13916), .ZN(P1_U2991) );
  XNOR2_X1 U17152 ( .A(n13917), .B(n13918), .ZN(n15351) );
  OAI21_X1 U17153 ( .B1(n13920), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13919), .ZN(n15338) );
  INV_X1 U17154 ( .A(n15338), .ZN(n13924) );
  OAI22_X1 U17155 ( .A1(n12329), .A2(n19058), .B1(n19267), .B2(n19086), .ZN(
        n13923) );
  INV_X1 U17156 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13921) );
  OAI22_X1 U17157 ( .A1(n16287), .A2(n19092), .B1(n16338), .B2(n13921), .ZN(
        n13922) );
  AOI211_X1 U17158 ( .C1(n13924), .C2(n9733), .A(n13923), .B(n13922), .ZN(
        n13925) );
  OAI21_X1 U17159 ( .B1(n19259), .B2(n15351), .A(n13925), .ZN(P2_U3008) );
  AOI21_X1 U17160 ( .B1(n13927), .B2(n13926), .A(n10178), .ZN(n13941) );
  INV_X1 U17161 ( .A(n13941), .ZN(n13932) );
  NAND2_X1 U17162 ( .A1(n13929), .A2(n13928), .ZN(n13930) );
  NAND2_X1 U17163 ( .A1(n14792), .A2(n13930), .ZN(n18998) );
  MUX2_X1 U17164 ( .A(n18998), .B(n12536), .S(n14799), .Z(n13931) );
  OAI21_X1 U17165 ( .B1(n13932), .B2(n14785), .A(n13931), .ZN(P2_U2869) );
  OR2_X1 U17166 ( .A1(n13934), .A2(n13933), .ZN(n13936) );
  NAND2_X1 U17167 ( .A1(n13936), .A2(n13935), .ZN(n19008) );
  AOI22_X1 U17168 ( .A1(n19134), .A2(BUF2_REG_18__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17169 ( .A1(n16265), .A2(n13937), .B1(n19172), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n13938) );
  OAI211_X1 U17170 ( .C1(n16267), .C2(n19008), .A(n13939), .B(n13938), .ZN(
        n13940) );
  AOI21_X1 U17171 ( .B1(n13941), .B2(n19175), .A(n13940), .ZN(n13942) );
  INV_X1 U17172 ( .A(n13942), .ZN(P2_U2901) );
  AOI21_X1 U17173 ( .B1(n13944), .B2(n13854), .A(n13943), .ZN(n20006) );
  INV_X1 U17174 ( .A(n20006), .ZN(n13969) );
  INV_X1 U17175 ( .A(n13945), .ZN(n13948) );
  INV_X1 U17176 ( .A(n13946), .ZN(n13947) );
  AOI21_X1 U17177 ( .B1(n13948), .B2(n13947), .A(n13957), .ZN(n19999) );
  AOI22_X1 U17178 ( .A1(n19999), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n13949) );
  OAI21_X1 U17179 ( .B1(n13969), .B2(n14277), .A(n13949), .ZN(P1_U2863) );
  INV_X1 U17180 ( .A(DATAI_9_), .ZN(n13951) );
  NAND2_X1 U17181 ( .A1(n20156), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13950) );
  OAI21_X1 U17182 ( .B1(n20156), .B2(n13951), .A(n13950), .ZN(n20099) );
  AOI22_X1 U17183 ( .A1(n15969), .A2(n20099), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14348), .ZN(n13952) );
  OAI21_X1 U17184 ( .B1(n13969), .B2(n14354), .A(n13952), .ZN(P1_U2895) );
  NOR2_X1 U17185 ( .A1(n13943), .A2(n13954), .ZN(n13955) );
  OR2_X1 U17186 ( .A1(n13953), .A2(n13955), .ZN(n15960) );
  OR2_X1 U17187 ( .A1(n13957), .A2(n13956), .ZN(n13958) );
  NAND2_X1 U17188 ( .A1(n14272), .A2(n13958), .ZN(n16116) );
  OAI22_X1 U17189 ( .A1(n16116), .A2(n14280), .B1(n13959), .B2(n14278), .ZN(
        n13960) );
  INV_X1 U17190 ( .A(n13960), .ZN(n13961) );
  OAI21_X1 U17191 ( .B1(n15960), .B2(n14277), .A(n13961), .ZN(P1_U2862) );
  INV_X1 U17192 ( .A(n20158), .ZN(n20137) );
  XNOR2_X1 U17193 ( .A(n16009), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13962) );
  XNOR2_X1 U17194 ( .A(n13963), .B(n13962), .ZN(n16122) );
  NAND2_X1 U17195 ( .A1(n16122), .A2(n20134), .ZN(n13968) );
  INV_X1 U17196 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13964) );
  NOR2_X1 U17197 ( .A1(n20042), .A2(n13964), .ZN(n16121) );
  NOR2_X1 U17198 ( .A1(n16029), .A2(n13965), .ZN(n13966) );
  AOI211_X1 U17199 ( .C1(n20132), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16121), .B(n13966), .ZN(n13967) );
  OAI211_X1 U17200 ( .C1(n20137), .C2(n13969), .A(n13968), .B(n13967), .ZN(
        P1_U2990) );
  INV_X1 U17201 ( .A(DATAI_10_), .ZN(n13971) );
  NAND2_X1 U17202 ( .A1(n20156), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13970) );
  OAI21_X1 U17203 ( .B1(n20156), .B2(n13971), .A(n13970), .ZN(n20101) );
  INV_X1 U17204 ( .A(n20101), .ZN(n13973) );
  OAI222_X1 U17205 ( .A1(n15960), .A2(n14354), .B1(n14353), .B2(n13973), .C1(
        n13972), .C2(n15972), .ZN(P1_U2894) );
  NAND2_X1 U17206 ( .A1(n13975), .A2(n13974), .ZN(n15177) );
  NAND2_X1 U17207 ( .A1(n15177), .A2(n16335), .ZN(n13986) );
  AOI21_X1 U17208 ( .B1(n13976), .B2(n14963), .A(n14945), .ZN(n15175) );
  NOR2_X1 U17209 ( .A1(n14775), .A2(n13977), .ZN(n13978) );
  OR2_X1 U17210 ( .A1(n14761), .A2(n13978), .ZN(n16255) );
  OAI22_X1 U17211 ( .A1(n16338), .A2(n13980), .B1(n13979), .B2(n19058), .ZN(
        n13981) );
  AOI21_X1 U17212 ( .B1(n16327), .B2(n13982), .A(n13981), .ZN(n13983) );
  OAI21_X1 U17213 ( .B1(n16255), .B2(n16287), .A(n13983), .ZN(n13984) );
  AOI21_X1 U17214 ( .B1(n15175), .B2(n9733), .A(n13984), .ZN(n13985) );
  OAI21_X1 U17215 ( .B1(n15176), .B2(n13986), .A(n13985), .ZN(P2_U2991) );
  NOR2_X1 U17216 ( .A1(n14714), .A2(n16287), .ZN(n13991) );
  NAND2_X1 U17217 ( .A1(n19256), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13987) );
  OAI211_X1 U17218 ( .C1(n19267), .C2(n13989), .A(n13988), .B(n13987), .ZN(
        n13990) );
  OAI21_X1 U17219 ( .B1(n13994), .B2(n19259), .A(n13993), .ZN(P2_U2983) );
  INV_X1 U17220 ( .A(n13995), .ZN(n15590) );
  INV_X1 U17221 ( .A(n13996), .ZN(n13997) );
  NOR2_X1 U17222 ( .A1(n13998), .A2(n13997), .ZN(n14008) );
  NOR2_X1 U17223 ( .A1(n13999), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14003) );
  NOR3_X1 U17224 ( .A1(n14001), .A2(n11543), .A3(n14000), .ZN(n14002) );
  AOI211_X1 U17225 ( .C1(n14005), .C2(n14004), .A(n14003), .B(n14002), .ZN(
        n16428) );
  OAI22_X1 U17226 ( .A1(n19943), .A2(n14006), .B1(n19924), .B2(n16428), .ZN(
        n14007) );
  OAI21_X1 U17227 ( .B1(n14008), .B2(n14007), .A(n15590), .ZN(n14009) );
  OAI21_X1 U17228 ( .B1(n15590), .B2(n14010), .A(n14009), .ZN(P2_U3600) );
  XNOR2_X1 U17229 ( .A(n9780), .B(n14011), .ZN(n16190) );
  NOR2_X1 U17230 ( .A1(n16190), .A2(n14799), .ZN(n14012) );
  AOI21_X1 U17231 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14799), .A(n14012), .ZN(
        n14013) );
  OAI21_X1 U17232 ( .B1(n14014), .B2(n14785), .A(n14013), .ZN(P2_U2857) );
  INV_X1 U17233 ( .A(n14015), .ZN(n14019) );
  INV_X1 U17234 ( .A(n14016), .ZN(n14018) );
  NAND3_X1 U17235 ( .A1(n14019), .A2(n14018), .A3(n14017), .ZN(n14020) );
  AND2_X1 U17236 ( .A1(n14021), .A2(n14020), .ZN(n14026) );
  NAND2_X1 U17237 ( .A1(n14032), .A2(n14022), .ZN(n14025) );
  OR2_X1 U17238 ( .A1(n14023), .A2(n11276), .ZN(n14024) );
  OAI211_X1 U17239 ( .C1(n14032), .C2(n14026), .A(n14025), .B(n14024), .ZN(
        n14028) );
  AND2_X1 U17240 ( .A1(n14028), .A2(n14027), .ZN(n15804) );
  INV_X1 U17241 ( .A(n14029), .ZN(n14031) );
  OAI22_X1 U17242 ( .A1(n14032), .A2(n10451), .B1(n14031), .B2(n14030), .ZN(
        n19977) );
  INV_X1 U17243 ( .A(n14033), .ZN(n14034) );
  AOI21_X1 U17244 ( .B1(n14034), .B2(n15842), .A(n16173), .ZN(n20850) );
  NOR2_X1 U17245 ( .A1(n19977), .A2(n20850), .ZN(n15807) );
  NOR2_X1 U17246 ( .A1(n15807), .A2(n19976), .ZN(n19983) );
  MUX2_X1 U17247 ( .A(P1_MORE_REG_SCAN_IN), .B(n15804), .S(n19983), .Z(
        P1_U3484) );
  NAND2_X1 U17248 ( .A1(n14055), .A2(n14035), .ZN(n14039) );
  INV_X1 U17249 ( .A(n14036), .ZN(n14037) );
  NAND2_X1 U17250 ( .A1(n14068), .A2(n14037), .ZN(n14038) );
  NAND2_X1 U17251 ( .A1(n14039), .A2(n14038), .ZN(n14042) );
  INV_X1 U17252 ( .A(n14040), .ZN(n14041) );
  XNOR2_X1 U17253 ( .A(n14042), .B(n14041), .ZN(n14537) );
  AOI21_X1 U17254 ( .B1(n14044), .B2(n14057), .A(n14043), .ZN(n14365) );
  NAND2_X1 U17255 ( .A1(n14365), .A2(n20031), .ZN(n14052) );
  OAI22_X1 U17256 ( .A1(n14045), .A2(n20044), .B1(n20054), .B2(n14363), .ZN(
        n14050) );
  AOI21_X1 U17257 ( .B1(n14063), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14048) );
  INV_X1 U17258 ( .A(n14046), .ZN(n14047) );
  NOR2_X1 U17259 ( .A1(n14048), .A2(n14047), .ZN(n14049) );
  AOI211_X1 U17260 ( .C1(n20046), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14050), .B(
        n14049), .ZN(n14051) );
  OAI211_X1 U17261 ( .C1(n20062), .C2(n14537), .A(n14052), .B(n14051), .ZN(
        P1_U2810) );
  OR2_X1 U17262 ( .A1(n14068), .A2(n14053), .ZN(n14054) );
  NAND2_X1 U17263 ( .A1(n14055), .A2(n14054), .ZN(n14552) );
  OAI21_X1 U17264 ( .B1(n14056), .B2(n14058), .A(n14057), .ZN(n14376) );
  INV_X1 U17265 ( .A(n14376), .ZN(n14059) );
  NAND2_X1 U17266 ( .A1(n14059), .A2(n20031), .ZN(n14065) );
  INV_X1 U17267 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14367) );
  AOI22_X1 U17268 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20059), .B1(
        n20040), .B2(n14369), .ZN(n14061) );
  NAND2_X1 U17269 ( .A1(n20046), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14060) );
  OAI211_X1 U17270 ( .C1(n14075), .C2(n14367), .A(n14061), .B(n14060), .ZN(
        n14062) );
  AOI21_X1 U17271 ( .B1(n14063), .B2(n14367), .A(n14062), .ZN(n14064) );
  OAI211_X1 U17272 ( .C1(n20062), .C2(n14552), .A(n14065), .B(n14064), .ZN(
        P1_U2811) );
  NOR2_X1 U17273 ( .A1(n9782), .A2(n14066), .ZN(n14067) );
  NAND2_X1 U17274 ( .A1(n14387), .A2(n20031), .ZN(n14079) );
  INV_X1 U17275 ( .A(n14385), .ZN(n14071) );
  AOI22_X1 U17276 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20059), .B1(
        n20040), .B2(n14071), .ZN(n14073) );
  NAND2_X1 U17277 ( .A1(n20046), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14072) );
  OAI211_X1 U17278 ( .C1(n14074), .C2(P1_REIP_REG_28__SCAN_IN), .A(n14073), 
        .B(n14072), .ZN(n14077) );
  NOR2_X1 U17279 ( .A1(n14075), .A2(n14383), .ZN(n14076) );
  NOR2_X1 U17280 ( .A1(n14077), .A2(n14076), .ZN(n14078) );
  OAI211_X1 U17281 ( .C1(n14561), .C2(n20062), .A(n14079), .B(n14078), .ZN(
        P1_U2812) );
  INV_X1 U17282 ( .A(n14080), .ZN(n14081) );
  INV_X1 U17283 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U17284 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20059), .B1(
        n20040), .B2(n14394), .ZN(n14083) );
  OAI21_X1 U17285 ( .B1(n20060), .B2(n14084), .A(n14083), .ZN(n14086) );
  NOR3_X1 U17286 ( .A1(n14096), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n16045), 
        .ZN(n14085) );
  AOI211_X1 U17287 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14094), .A(n14086), 
        .B(n14085), .ZN(n14089) );
  AOI21_X1 U17288 ( .B1(n14087), .B2(n14099), .A(n9782), .ZN(n14565) );
  NAND2_X1 U17289 ( .A1(n14565), .A2(n20027), .ZN(n14088) );
  OAI211_X1 U17290 ( .C1(n14303), .C2(n15890), .A(n14089), .B(n14088), .ZN(
        P1_U2813) );
  INV_X1 U17291 ( .A(n14090), .ZN(n14091) );
  AOI21_X1 U17292 ( .B1(n14092), .B2(n14104), .A(n14091), .ZN(n14405) );
  INV_X1 U17293 ( .A(n14405), .ZN(n14310) );
  OAI22_X1 U17294 ( .A1(n14093), .A2(n20044), .B1(n20054), .B2(n14403), .ZN(
        n14098) );
  INV_X1 U17295 ( .A(n14094), .ZN(n14095) );
  AOI21_X1 U17296 ( .B1(n16045), .B2(n14096), .A(n14095), .ZN(n14097) );
  AOI211_X1 U17297 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20046), .A(n14098), .B(
        n14097), .ZN(n14103) );
  INV_X1 U17298 ( .A(n14099), .ZN(n14100) );
  AOI21_X1 U17299 ( .B1(n14101), .B2(n14110), .A(n14100), .ZN(n16038) );
  NAND2_X1 U17300 ( .A1(n16038), .A2(n20027), .ZN(n14102) );
  OAI211_X1 U17301 ( .C1(n14310), .C2(n15890), .A(n14103), .B(n14102), .ZN(
        P1_U2814) );
  OAI21_X1 U17302 ( .B1(n14116), .B2(n14105), .A(n14104), .ZN(n14410) );
  INV_X1 U17303 ( .A(n14137), .ZN(n14128) );
  INV_X1 U17304 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14198) );
  OAI211_X1 U17305 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n14119), .B(n14106), .ZN(n14109) );
  INV_X1 U17306 ( .A(n14412), .ZN(n14107) );
  AOI22_X1 U17307 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20059), .B1(
        n20040), .B2(n14107), .ZN(n14108) );
  OAI211_X1 U17308 ( .C1(n14198), .C2(n20060), .A(n14109), .B(n14108), .ZN(
        n14113) );
  OAI21_X1 U17309 ( .B1(n14125), .B2(n14111), .A(n14110), .ZN(n16048) );
  NOR2_X1 U17310 ( .A1(n16048), .A2(n20062), .ZN(n14112) );
  AOI211_X1 U17311 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14128), .A(n14113), 
        .B(n14112), .ZN(n14114) );
  OAI21_X1 U17312 ( .B1(n14410), .B2(n15890), .A(n14114), .ZN(P1_U2815) );
  INV_X1 U17313 ( .A(n14134), .ZN(n14117) );
  AOI21_X1 U17314 ( .B1(n10253), .B2(n14117), .A(n14116), .ZN(n14422) );
  INV_X1 U17315 ( .A(n14422), .ZN(n14315) );
  INV_X1 U17316 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U17317 ( .A1(n14119), .A2(n14118), .ZN(n14122) );
  INV_X1 U17318 ( .A(n14420), .ZN(n14120) );
  AOI22_X1 U17319 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20059), .B1(
        n20040), .B2(n14120), .ZN(n14121) );
  OAI211_X1 U17320 ( .C1(n14199), .C2(n20060), .A(n14122), .B(n14121), .ZN(
        n14127) );
  NOR2_X1 U17321 ( .A1(n14130), .A2(n14123), .ZN(n14124) );
  OR2_X1 U17322 ( .A1(n14125), .A2(n14124), .ZN(n14578) );
  NOR2_X1 U17323 ( .A1(n14578), .A2(n20062), .ZN(n14126) );
  AOI211_X1 U17324 ( .C1(n14128), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14127), 
        .B(n14126), .ZN(n14129) );
  OAI21_X1 U17325 ( .B1(n14315), .B2(n15890), .A(n14129), .ZN(P1_U2816) );
  INV_X1 U17326 ( .A(n14130), .ZN(n14131) );
  OAI21_X1 U17327 ( .B1(n14132), .B2(n14205), .A(n14131), .ZN(n14585) );
  AOI21_X1 U17328 ( .B1(n14135), .B2(n14133), .A(n14134), .ZN(n14431) );
  NAND2_X1 U17329 ( .A1(n14431), .A2(n20031), .ZN(n14142) );
  INV_X1 U17330 ( .A(n14434), .ZN(n14136) );
  OAI22_X1 U17331 ( .A1(n20941), .A2(n20044), .B1(n20054), .B2(n14136), .ZN(
        n14140) );
  AOI21_X1 U17332 ( .B1(n14432), .B2(n14138), .A(n14137), .ZN(n14139) );
  AOI211_X1 U17333 ( .C1(n20046), .C2(P1_EBX_REG_23__SCAN_IN), .A(n14140), .B(
        n14139), .ZN(n14141) );
  OAI211_X1 U17334 ( .C1(n14585), .C2(n20062), .A(n14142), .B(n14141), .ZN(
        P1_U2817) );
  INV_X1 U17335 ( .A(n14144), .ZN(n14145) );
  OAI21_X1 U17336 ( .B1(n14146), .B2(n14143), .A(n14145), .ZN(n14437) );
  XNOR2_X1 U17337 ( .A(n9774), .B(n14210), .ZN(n15848) );
  AOI22_X1 U17338 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20059), .B1(
        n20046), .B2(P1_EBX_REG_20__SCAN_IN), .ZN(n14147) );
  OAI21_X1 U17339 ( .B1(n14442), .B2(n20054), .A(n14147), .ZN(n14150) );
  INV_X1 U17340 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15868) );
  NAND2_X1 U17341 ( .A1(n20019), .A2(n14148), .ZN(n15867) );
  NAND2_X1 U17342 ( .A1(n14148), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15876) );
  INV_X1 U17343 ( .A(n14158), .ZN(n20017) );
  AOI21_X1 U17344 ( .B1(n20019), .B2(n15876), .A(n20017), .ZN(n15883) );
  AOI21_X1 U17345 ( .B1(n15868), .B2(n15867), .A(n15883), .ZN(n14149) );
  AOI211_X1 U17346 ( .C1(n20027), .C2(n15848), .A(n14150), .B(n14149), .ZN(
        n14151) );
  OAI21_X1 U17347 ( .B1(n14437), .B2(n15890), .A(n14151), .ZN(P1_U2820) );
  OR2_X1 U17348 ( .A1(n13953), .A2(n14153), .ZN(n14154) );
  NAND2_X1 U17349 ( .A1(n14152), .A2(n14154), .ZN(n14276) );
  INV_X1 U17350 ( .A(n14275), .ZN(n14155) );
  OAI21_X1 U17351 ( .B1(n14276), .B2(n14155), .A(n14152), .ZN(n14260) );
  AND2_X1 U17352 ( .A1(n14260), .A2(n14261), .ZN(n14262) );
  OAI21_X1 U17353 ( .B1(n14262), .B2(n14157), .A(n14156), .ZN(n14495) );
  NAND2_X1 U17354 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15906) );
  NAND2_X1 U17355 ( .A1(n14158), .A2(n14160), .ZN(n15950) );
  OAI21_X1 U17356 ( .B1(n15906), .B2(n15950), .A(n15951), .ZN(n14159) );
  INV_X1 U17357 ( .A(n14159), .ZN(n15946) );
  AOI21_X1 U17358 ( .B1(n9844), .B2(n10072), .A(n14256), .ZN(n16092) );
  INV_X1 U17359 ( .A(n14160), .ZN(n14161) );
  NOR2_X1 U17360 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15906), .ZN(n14162) );
  AOI22_X1 U17361 ( .A1(n20027), .A2(n16092), .B1(n15952), .B2(n14162), .ZN(
        n14163) );
  OAI21_X1 U17362 ( .B1(n14164), .B2(n20044), .A(n14163), .ZN(n14165) );
  AOI211_X1 U17363 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n15946), .A(n20135), 
        .B(n14165), .ZN(n14168) );
  INV_X1 U17364 ( .A(n14491), .ZN(n14166) );
  AOI22_X1 U17365 ( .A1(n20046), .A2(P1_EBX_REG_13__SCAN_IN), .B1(n20040), 
        .B2(n14166), .ZN(n14167) );
  OAI211_X1 U17366 ( .C1(n14495), .C2(n15890), .A(n14168), .B(n14167), .ZN(
        P1_U2827) );
  INV_X1 U17367 ( .A(n20056), .ZN(n14188) );
  OAI21_X1 U17368 ( .B1(n14170), .B2(n14169), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n14172) );
  NAND2_X1 U17369 ( .A1(n20059), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14171) );
  OAI211_X1 U17370 ( .C1(n20054), .C2(n14173), .A(n14172), .B(n14171), .ZN(
        n14174) );
  AOI21_X1 U17371 ( .B1(n20046), .B2(P1_EBX_REG_3__SCAN_IN), .A(n14174), .ZN(
        n14175) );
  OAI21_X1 U17372 ( .B1(n20062), .B2(n14176), .A(n14175), .ZN(n14179) );
  INV_X1 U17373 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20767) );
  NAND2_X1 U17374 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20767), .ZN(n14177) );
  NOR2_X1 U17375 ( .A1(n20063), .A2(n14177), .ZN(n14178) );
  AOI211_X1 U17376 ( .C1(n14188), .C2(n20817), .A(n14179), .B(n14178), .ZN(
        n14180) );
  OAI21_X1 U17377 ( .B1(n14190), .B2(n14181), .A(n14180), .ZN(P1_U2837) );
  NAND2_X1 U17378 ( .A1(n20046), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n14184) );
  AOI22_X1 U17379 ( .A1(n20059), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20017), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14183) );
  OAI211_X1 U17380 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20054), .A(
        n14184), .B(n14183), .ZN(n14187) );
  OAI22_X1 U17381 ( .A1(n20062), .A2(n14185), .B1(n20021), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14186) );
  AOI211_X1 U17382 ( .C1(n20647), .C2(n14188), .A(n14187), .B(n14186), .ZN(
        n14189) );
  OAI21_X1 U17383 ( .B1(n14191), .B2(n14190), .A(n14189), .ZN(P1_U2839) );
  INV_X1 U17384 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14192) );
  OAI22_X1 U17385 ( .A1(n14525), .A2(n14280), .B1(n14192), .B2(n14278), .ZN(
        P1_U2841) );
  INV_X1 U17386 ( .A(n14365), .ZN(n14286) );
  INV_X1 U17387 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14193) );
  OAI222_X1 U17388 ( .A1(n14270), .A2(n14286), .B1(n14278), .B2(n14193), .C1(
        n14537), .C2(n14280), .ZN(P1_U2842) );
  OAI222_X1 U17389 ( .A1(n14194), .A2(n14278), .B1(n14280), .B2(n14552), .C1(
        n14376), .C2(n14277), .ZN(P1_U2843) );
  INV_X1 U17390 ( .A(n14387), .ZN(n14298) );
  OAI222_X1 U17391 ( .A1(n14195), .A2(n14278), .B1(n14280), .B2(n14561), .C1(
        n14298), .C2(n14277), .ZN(P1_U2844) );
  AOI22_X1 U17392 ( .A1(n14565), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n14196) );
  OAI21_X1 U17393 ( .B1(n14303), .B2(n14270), .A(n14196), .ZN(P1_U2845) );
  AOI22_X1 U17394 ( .A1(n16038), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n14197) );
  OAI21_X1 U17395 ( .B1(n14310), .B2(n14270), .A(n14197), .ZN(P1_U2846) );
  OAI222_X1 U17396 ( .A1(n14198), .A2(n14278), .B1(n14280), .B2(n16048), .C1(
        n14410), .C2(n14277), .ZN(P1_U2847) );
  OAI222_X1 U17397 ( .A1(n14199), .A2(n14278), .B1(n14280), .B2(n14578), .C1(
        n14315), .C2(n14277), .ZN(P1_U2848) );
  INV_X1 U17398 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14200) );
  INV_X1 U17399 ( .A(n14431), .ZN(n14319) );
  OAI222_X1 U17400 ( .A1(n14585), .A2(n14280), .B1(n14278), .B2(n14200), .C1(
        n14277), .C2(n14319), .ZN(P1_U2849) );
  INV_X1 U17401 ( .A(n14133), .ZN(n14202) );
  AOI21_X1 U17402 ( .B1(n14203), .B2(n14201), .A(n14202), .ZN(n15974) );
  INV_X1 U17403 ( .A(n15974), .ZN(n14323) );
  AND2_X1 U17404 ( .A1(n14214), .A2(n14204), .ZN(n14206) );
  OR2_X1 U17405 ( .A1(n14206), .A2(n14205), .ZN(n15875) );
  OAI22_X1 U17406 ( .A1(n15875), .A2(n14280), .B1(n15869), .B2(n14278), .ZN(
        n14207) );
  INV_X1 U17407 ( .A(n14207), .ZN(n14208) );
  OAI21_X1 U17408 ( .B1(n14323), .B2(n14270), .A(n14208), .ZN(P1_U2850) );
  OAI21_X1 U17409 ( .B1(n14144), .B2(n14209), .A(n14201), .ZN(n15978) );
  INV_X1 U17410 ( .A(n14210), .ZN(n14213) );
  INV_X1 U17411 ( .A(n14211), .ZN(n14212) );
  OAI21_X1 U17412 ( .B1(n9774), .B2(n14213), .A(n14212), .ZN(n14215) );
  NAND2_X1 U17413 ( .A1(n14215), .A2(n14214), .ZN(n15877) );
  OAI22_X1 U17414 ( .A1(n15877), .A2(n14280), .B1(n14216), .B2(n14278), .ZN(
        n14217) );
  INV_X1 U17415 ( .A(n14217), .ZN(n14218) );
  OAI21_X1 U17416 ( .B1(n15978), .B2(n14270), .A(n14218), .ZN(P1_U2851) );
  AOI22_X1 U17417 ( .A1(n15848), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n14219) );
  OAI21_X1 U17418 ( .B1(n14437), .B2(n14270), .A(n14219), .ZN(P1_U2852) );
  AOI21_X1 U17419 ( .B1(n14220), .B2(n14228), .A(n14143), .ZN(n14452) );
  INV_X1 U17420 ( .A(n14452), .ZN(n15891) );
  NAND2_X1 U17421 ( .A1(n9822), .A2(n14221), .ZN(n14222) );
  NAND2_X1 U17422 ( .A1(n9774), .A2(n14222), .ZN(n15889) );
  INV_X1 U17423 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15888) );
  OAI22_X1 U17424 ( .A1(n15889), .A2(n14280), .B1(n15888), .B2(n14278), .ZN(
        n14223) );
  INV_X1 U17425 ( .A(n14223), .ZN(n14224) );
  OAI21_X1 U17426 ( .B1(n15891), .B2(n14270), .A(n14224), .ZN(P1_U2853) );
  NAND2_X1 U17427 ( .A1(n14225), .A2(n14226), .ZN(n14227) );
  AND2_X1 U17428 ( .A1(n14228), .A2(n14227), .ZN(n15903) );
  INV_X1 U17429 ( .A(n15903), .ZN(n14336) );
  OR2_X1 U17430 ( .A1(n14235), .A2(n14229), .ZN(n14230) );
  NAND2_X1 U17431 ( .A1(n9822), .A2(n14230), .ZN(n16055) );
  OAI22_X1 U17432 ( .A1(n16055), .A2(n14280), .B1(n15898), .B2(n14278), .ZN(
        n14231) );
  INV_X1 U17433 ( .A(n14231), .ZN(n14232) );
  OAI21_X1 U17434 ( .B1(n14336), .B2(n14270), .A(n14232), .ZN(P1_U2854) );
  NOR2_X1 U17435 ( .A1(n14241), .A2(n14233), .ZN(n14234) );
  OR2_X1 U17436 ( .A1(n14235), .A2(n14234), .ZN(n15916) );
  INV_X1 U17437 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14237) );
  OAI21_X1 U17438 ( .B1(n14239), .B2(n14236), .A(n14225), .ZN(n15905) );
  OAI222_X1 U17439 ( .A1(n15916), .A2(n14280), .B1(n14278), .B2(n14237), .C1(
        n14277), .C2(n15905), .ZN(P1_U2855) );
  AND2_X1 U17440 ( .A1(n14249), .A2(n14238), .ZN(n14240) );
  OR2_X1 U17441 ( .A1(n14240), .A2(n14239), .ZN(n15918) );
  AOI21_X1 U17442 ( .B1(n14242), .B2(n14247), .A(n14241), .ZN(n16066) );
  AOI22_X1 U17443 ( .A1(n16066), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14243) );
  OAI21_X1 U17444 ( .B1(n15918), .B2(n14270), .A(n14243), .ZN(P1_U2856) );
  NAND2_X1 U17445 ( .A1(n14245), .A2(n14244), .ZN(n14246) );
  NAND2_X1 U17446 ( .A1(n14247), .A2(n14246), .ZN(n16074) );
  INV_X1 U17447 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n20909) );
  INV_X1 U17448 ( .A(n14249), .ZN(n14250) );
  AOI21_X1 U17449 ( .B1(n14251), .B2(n14252), .A(n14250), .ZN(n15933) );
  INV_X1 U17450 ( .A(n15933), .ZN(n14482) );
  OAI222_X1 U17451 ( .A1(n16074), .A2(n14280), .B1(n14278), .B2(n20909), .C1(
        n14277), .C2(n14482), .ZN(P1_U2857) );
  INV_X1 U17452 ( .A(n14252), .ZN(n14253) );
  AOI21_X1 U17453 ( .B1(n9984), .B2(n14156), .A(n14253), .ZN(n16001) );
  INV_X1 U17454 ( .A(n16001), .ZN(n14258) );
  INV_X1 U17455 ( .A(n14254), .ZN(n14255) );
  XNOR2_X1 U17456 ( .A(n14256), .B(n14255), .ZN(n16083) );
  AOI22_X1 U17457 ( .A1(n16083), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14257) );
  OAI21_X1 U17458 ( .B1(n14258), .B2(n14270), .A(n14257), .ZN(P1_U2858) );
  AOI22_X1 U17459 ( .A1(n16092), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14259) );
  OAI21_X1 U17460 ( .B1(n14495), .B2(n14270), .A(n14259), .ZN(P1_U2859) );
  INV_X1 U17461 ( .A(n14260), .ZN(n14264) );
  INV_X1 U17462 ( .A(n14261), .ZN(n14263) );
  AOI21_X1 U17463 ( .B1(n14264), .B2(n14263), .A(n14262), .ZN(n16004) );
  INV_X1 U17464 ( .A(n16004), .ZN(n14350) );
  AOI21_X1 U17465 ( .B1(n14266), .B2(n14274), .A(n14265), .ZN(n15943) );
  AOI22_X1 U17466 ( .A1(n15943), .A2(n14268), .B1(n14267), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14269) );
  OAI21_X1 U17467 ( .B1(n14350), .B2(n14270), .A(n14269), .ZN(P1_U2860) );
  NAND2_X1 U17468 ( .A1(n14272), .A2(n14271), .ZN(n14273) );
  NAND2_X1 U17469 ( .A1(n14274), .A2(n14273), .ZN(n16104) );
  INV_X1 U17470 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14279) );
  XNOR2_X1 U17471 ( .A(n14276), .B(n14275), .ZN(n16014) );
  INV_X1 U17472 ( .A(n16014), .ZN(n14355) );
  OAI222_X1 U17473 ( .A1(n16104), .A2(n14280), .B1(n14279), .B2(n14278), .C1(
        n14277), .C2(n14355), .ZN(P1_U2861) );
  AOI22_X1 U17474 ( .A1(n14340), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14348), .ZN(n14285) );
  NOR3_X4 U17475 ( .A1(n14348), .A2(n20224), .A3(n14281), .ZN(n14342) );
  INV_X1 U17476 ( .A(DATAI_14_), .ZN(n14283) );
  NAND2_X1 U17477 ( .A1(n20156), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14282) );
  OAI21_X1 U17478 ( .B1(n20156), .B2(n14283), .A(n14282), .ZN(n20109) );
  AOI22_X1 U17479 ( .A1(n14343), .A2(DATAI_30_), .B1(n14342), .B2(n20109), 
        .ZN(n14284) );
  OAI211_X1 U17480 ( .C1(n14286), .C2(n14354), .A(n14285), .B(n14284), .ZN(
        P1_U2874) );
  AOI22_X1 U17481 ( .A1(n14340), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14348), .ZN(n14290) );
  INV_X1 U17482 ( .A(DATAI_13_), .ZN(n14288) );
  NAND2_X1 U17483 ( .A1(n20156), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14287) );
  OAI21_X1 U17484 ( .B1(n20156), .B2(n14288), .A(n14287), .ZN(n20107) );
  AOI22_X1 U17485 ( .A1(n14343), .A2(DATAI_29_), .B1(n14342), .B2(n20107), 
        .ZN(n14289) );
  OAI211_X1 U17486 ( .C1(n14376), .C2(n14354), .A(n14290), .B(n14289), .ZN(
        P1_U2875) );
  INV_X1 U17487 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n14292) );
  OAI22_X1 U17488 ( .A1(n14306), .A2(n14292), .B1(n14291), .B2(n15972), .ZN(
        n14293) );
  INV_X1 U17489 ( .A(n14293), .ZN(n14297) );
  INV_X1 U17490 ( .A(DATAI_12_), .ZN(n14295) );
  NAND2_X1 U17491 ( .A1(n20156), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14294) );
  OAI21_X1 U17492 ( .B1(n20156), .B2(n14295), .A(n14294), .ZN(n20105) );
  AOI22_X1 U17493 ( .A1(n14343), .A2(DATAI_28_), .B1(n14342), .B2(n20105), 
        .ZN(n14296) );
  OAI211_X1 U17494 ( .C1(n14298), .C2(n14354), .A(n14297), .B(n14296), .ZN(
        P1_U2876) );
  AOI22_X1 U17495 ( .A1(n14340), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14348), .ZN(n14302) );
  INV_X1 U17496 ( .A(DATAI_11_), .ZN(n14300) );
  NAND2_X1 U17497 ( .A1(n20156), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14299) );
  OAI21_X1 U17498 ( .B1(n20156), .B2(n14300), .A(n14299), .ZN(n20103) );
  AOI22_X1 U17499 ( .A1(n14343), .A2(DATAI_27_), .B1(n14342), .B2(n20103), 
        .ZN(n14301) );
  OAI211_X1 U17500 ( .C1(n14303), .C2(n14354), .A(n14302), .B(n14301), .ZN(
        P1_U2877) );
  INV_X1 U17501 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n14305) );
  OAI22_X1 U17502 ( .A1(n14306), .A2(n14305), .B1(n14304), .B2(n15972), .ZN(
        n14307) );
  INV_X1 U17503 ( .A(n14307), .ZN(n14309) );
  AOI22_X1 U17504 ( .A1(n14343), .A2(DATAI_26_), .B1(n14342), .B2(n20101), 
        .ZN(n14308) );
  OAI211_X1 U17505 ( .C1(n14310), .C2(n14354), .A(n14309), .B(n14308), .ZN(
        P1_U2878) );
  AOI22_X1 U17506 ( .A1(n14340), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14348), .ZN(n14312) );
  AOI22_X1 U17507 ( .A1(n14343), .A2(DATAI_25_), .B1(n14342), .B2(n20099), 
        .ZN(n14311) );
  OAI211_X1 U17508 ( .C1(n14410), .C2(n14354), .A(n14312), .B(n14311), .ZN(
        P1_U2879) );
  AOI22_X1 U17509 ( .A1(n14340), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14348), .ZN(n14314) );
  AOI22_X1 U17510 ( .A1(n14343), .A2(DATAI_24_), .B1(n14342), .B2(n20097), 
        .ZN(n14313) );
  OAI211_X1 U17511 ( .C1(n14315), .C2(n14354), .A(n14314), .B(n14313), .ZN(
        P1_U2880) );
  AOI22_X1 U17512 ( .A1(n14340), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14348), .ZN(n14318) );
  AOI22_X1 U17513 ( .A1(n14343), .A2(DATAI_23_), .B1(n14342), .B2(n14316), 
        .ZN(n14317) );
  OAI211_X1 U17514 ( .C1(n14319), .C2(n14354), .A(n14318), .B(n14317), .ZN(
        P1_U2881) );
  AOI22_X1 U17515 ( .A1(n14340), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14348), .ZN(n14322) );
  AOI22_X1 U17516 ( .A1(n14343), .A2(DATAI_22_), .B1(n14342), .B2(n14320), 
        .ZN(n14321) );
  OAI211_X1 U17517 ( .C1(n14323), .C2(n14354), .A(n14322), .B(n14321), .ZN(
        P1_U2882) );
  AOI22_X1 U17518 ( .A1(n14340), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14348), .ZN(n14326) );
  AOI22_X1 U17519 ( .A1(n14343), .A2(DATAI_21_), .B1(n14342), .B2(n14324), 
        .ZN(n14325) );
  OAI211_X1 U17520 ( .C1(n15978), .C2(n14354), .A(n14326), .B(n14325), .ZN(
        P1_U2883) );
  AOI22_X1 U17521 ( .A1(n14340), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14348), .ZN(n14329) );
  AOI22_X1 U17522 ( .A1(n14343), .A2(DATAI_20_), .B1(n14342), .B2(n14327), 
        .ZN(n14328) );
  OAI211_X1 U17523 ( .C1(n14437), .C2(n14354), .A(n14329), .B(n14328), .ZN(
        P1_U2884) );
  AOI22_X1 U17524 ( .A1(n14340), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14348), .ZN(n14332) );
  AOI22_X1 U17525 ( .A1(n14343), .A2(DATAI_19_), .B1(n14342), .B2(n14330), 
        .ZN(n14331) );
  OAI211_X1 U17526 ( .C1(n15891), .C2(n14354), .A(n14332), .B(n14331), .ZN(
        P1_U2885) );
  AOI22_X1 U17527 ( .A1(n14340), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14348), .ZN(n14335) );
  AOI22_X1 U17528 ( .A1(n14343), .A2(DATAI_18_), .B1(n14342), .B2(n14333), 
        .ZN(n14334) );
  OAI211_X1 U17529 ( .C1(n14336), .C2(n14354), .A(n14335), .B(n14334), .ZN(
        P1_U2886) );
  AOI22_X1 U17530 ( .A1(n14340), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14348), .ZN(n14339) );
  AOI22_X1 U17531 ( .A1(n14343), .A2(DATAI_17_), .B1(n14342), .B2(n14337), 
        .ZN(n14338) );
  OAI211_X1 U17532 ( .C1(n15905), .C2(n14354), .A(n14339), .B(n14338), .ZN(
        P1_U2887) );
  AOI22_X1 U17533 ( .A1(n14340), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14348), .ZN(n14345) );
  AOI22_X1 U17534 ( .A1(n14343), .A2(DATAI_16_), .B1(n14342), .B2(n14341), 
        .ZN(n14344) );
  OAI211_X1 U17535 ( .C1(n15918), .C2(n14354), .A(n14345), .B(n14344), .ZN(
        P1_U2888) );
  OAI222_X1 U17536 ( .A1(n14482), .A2(n14354), .B1(n14353), .B2(n14346), .C1(
        n15972), .C2(n13631), .ZN(P1_U2889) );
  AOI22_X1 U17537 ( .A1(n15969), .A2(n20107), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14348), .ZN(n14347) );
  OAI21_X1 U17538 ( .B1(n14495), .B2(n14354), .A(n14347), .ZN(P1_U2891) );
  AOI22_X1 U17539 ( .A1(n15969), .A2(n20105), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14348), .ZN(n14349) );
  OAI21_X1 U17540 ( .B1(n14350), .B2(n14354), .A(n14349), .ZN(P1_U2892) );
  INV_X1 U17541 ( .A(n20103), .ZN(n14352) );
  OAI222_X1 U17542 ( .A1(n14355), .A2(n14354), .B1(n14353), .B2(n14352), .C1(
        n14351), .C2(n15972), .ZN(P1_U2893) );
  OR2_X1 U17543 ( .A1(n14356), .A2(n14371), .ZN(n14359) );
  INV_X1 U17544 ( .A(n14370), .ZN(n14357) );
  NAND3_X1 U17545 ( .A1(n14390), .A2(n14556), .A3(n14357), .ZN(n14358) );
  NAND2_X1 U17546 ( .A1(n14359), .A2(n14358), .ZN(n14360) );
  XNOR2_X1 U17547 ( .A(n14360), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14546) );
  INV_X1 U17548 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14361) );
  NOR2_X1 U17549 ( .A1(n20042), .A2(n14361), .ZN(n14538) );
  AOI21_X1 U17550 ( .B1(n20132), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14538), .ZN(n14362) );
  OAI21_X1 U17551 ( .B1(n16029), .B2(n14363), .A(n14362), .ZN(n14364) );
  AOI21_X1 U17552 ( .B1(n14365), .B2(n20158), .A(n14364), .ZN(n14366) );
  OAI21_X1 U17553 ( .B1(n14546), .B2(n19981), .A(n14366), .ZN(P1_U2969) );
  NOR2_X1 U17554 ( .A1(n20042), .A2(n14367), .ZN(n14548) );
  NOR2_X1 U17555 ( .A1(n16037), .A2(n20944), .ZN(n14368) );
  AOI211_X1 U17556 ( .C1(n16033), .C2(n14369), .A(n14548), .B(n14368), .ZN(
        n14375) );
  NAND2_X1 U17557 ( .A1(n14371), .A2(n14370), .ZN(n14372) );
  XNOR2_X1 U17558 ( .A(n14373), .B(n14372), .ZN(n14554) );
  NAND2_X1 U17559 ( .A1(n14554), .A2(n20134), .ZN(n14374) );
  OAI211_X1 U17560 ( .C1(n14376), .C2(n20137), .A(n14375), .B(n14374), .ZN(
        P1_U2970) );
  OR4_X1 U17561 ( .A1(n14465), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(n14377), .ZN(n14380) );
  NAND3_X1 U17562 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14379) );
  INV_X1 U17563 ( .A(n14425), .ZN(n14408) );
  AOI21_X1 U17564 ( .B1(n14515), .B2(n16009), .A(n14408), .ZN(n14378) );
  MUX2_X1 U17565 ( .A(n14380), .B(n14379), .S(n14378), .Z(n14382) );
  NOR2_X1 U17566 ( .A1(n20042), .A2(n14383), .ZN(n14558) );
  AOI21_X1 U17567 ( .B1(n20132), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14558), .ZN(n14384) );
  OAI21_X1 U17568 ( .B1(n16029), .B2(n14385), .A(n14384), .ZN(n14386) );
  AOI21_X1 U17569 ( .B1(n14387), .B2(n20158), .A(n14386), .ZN(n14388) );
  OAI21_X1 U17570 ( .B1(n14562), .B2(n19981), .A(n14388), .ZN(P1_U2971) );
  NAND2_X1 U17571 ( .A1(n9808), .A2(n14389), .ZN(n14392) );
  INV_X1 U17572 ( .A(n14390), .ZN(n14391) );
  MUX2_X1 U17573 ( .A(n14392), .B(n14391), .S(n14465), .Z(n14393) );
  XOR2_X1 U17574 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14393), .Z(
        n14573) );
  NAND2_X1 U17575 ( .A1(n16033), .A2(n14394), .ZN(n14395) );
  NAND2_X1 U17576 ( .A1(n20135), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14566) );
  OAI211_X1 U17577 ( .C1(n16037), .C2(n14396), .A(n14395), .B(n14566), .ZN(
        n14397) );
  AOI21_X1 U17578 ( .B1(n14398), .B2(n20158), .A(n14397), .ZN(n14399) );
  OAI21_X1 U17579 ( .B1(n19981), .B2(n14573), .A(n14399), .ZN(P1_U2972) );
  NOR2_X1 U17580 ( .A1(n14408), .A2(n14515), .ZN(n14400) );
  MUX2_X1 U17581 ( .A(n9808), .B(n14400), .S(n14465), .Z(n14401) );
  XNOR2_X1 U17582 ( .A(n14401), .B(n16042), .ZN(n16041) );
  INV_X1 U17583 ( .A(n16041), .ZN(n14407) );
  AOI22_X1 U17584 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n14402) );
  OAI21_X1 U17585 ( .B1(n16029), .B2(n14403), .A(n14402), .ZN(n14404) );
  AOI21_X1 U17586 ( .B1(n14405), .B2(n20158), .A(n14404), .ZN(n14406) );
  OAI21_X1 U17587 ( .B1(n19981), .B2(n14407), .A(n14406), .ZN(P1_U2973) );
  INV_X1 U17588 ( .A(n14410), .ZN(n14414) );
  AOI22_X1 U17589 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n14411) );
  OAI21_X1 U17590 ( .B1(n16029), .B2(n14412), .A(n14411), .ZN(n14413) );
  AOI21_X1 U17591 ( .B1(n14414), .B2(n20158), .A(n14413), .ZN(n14415) );
  OAI21_X1 U17592 ( .B1(n16047), .B2(n19981), .A(n14415), .ZN(P1_U2974) );
  MUX2_X1 U17593 ( .A(n14424), .B(n14417), .S(n14416), .Z(n14418) );
  XNOR2_X1 U17594 ( .A(n14418), .B(n14530), .ZN(n14584) );
  NAND2_X1 U17595 ( .A1(n20135), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14577) );
  NAND2_X1 U17596 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14419) );
  OAI211_X1 U17597 ( .C1(n16029), .C2(n14420), .A(n14577), .B(n14419), .ZN(
        n14421) );
  AOI21_X1 U17598 ( .B1(n14422), .B2(n20158), .A(n14421), .ZN(n14423) );
  OAI21_X1 U17599 ( .B1(n14584), .B2(n19981), .A(n14423), .ZN(P1_U2975) );
  INV_X1 U17600 ( .A(n14424), .ZN(n14430) );
  NOR2_X1 U17601 ( .A1(n14501), .A2(n14429), .ZN(n14427) );
  MUX2_X1 U17602 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n14429), .S(
        n14465), .Z(n14426) );
  MUX2_X1 U17603 ( .A(n14427), .B(n14426), .S(n14425), .Z(n14428) );
  AOI21_X1 U17604 ( .B1(n14430), .B2(n14429), .A(n14428), .ZN(n14593) );
  NAND2_X1 U17605 ( .A1(n14431), .A2(n20158), .ZN(n14436) );
  NOR2_X1 U17606 ( .A1(n20042), .A2(n14432), .ZN(n14586) );
  NOR2_X1 U17607 ( .A1(n16037), .A2(n20941), .ZN(n14433) );
  AOI211_X1 U17608 ( .C1(n16033), .C2(n14434), .A(n14586), .B(n14433), .ZN(
        n14435) );
  OAI211_X1 U17609 ( .C1(n14593), .C2(n19981), .A(n14436), .B(n14435), .ZN(
        P1_U2976) );
  INV_X1 U17610 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14446) );
  INV_X1 U17611 ( .A(n14437), .ZN(n14438) );
  NAND2_X1 U17612 ( .A1(n14438), .A2(n20158), .ZN(n14445) );
  NOR2_X1 U17613 ( .A1(n20042), .A2(n15868), .ZN(n15845) );
  INV_X1 U17614 ( .A(n14439), .ZN(n14440) );
  INV_X1 U17615 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14609) );
  AOI21_X1 U17616 ( .B1(n14440), .B2(n14501), .A(n15826), .ZN(n14441) );
  AOI21_X1 U17617 ( .B1(n14441), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15827), .ZN(n15852) );
  OAI22_X1 U17618 ( .A1(n15852), .A2(n19981), .B1(n16029), .B2(n14442), .ZN(
        n14443) );
  NOR2_X1 U17619 ( .A1(n15845), .A2(n14443), .ZN(n14444) );
  OAI211_X1 U17620 ( .C1(n16037), .C2(n14446), .A(n14445), .B(n14444), .ZN(
        P1_U2979) );
  NOR2_X1 U17621 ( .A1(n14465), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14447) );
  MUX2_X1 U17622 ( .A(n14465), .B(n14447), .S(n14454), .Z(n14448) );
  XNOR2_X1 U17623 ( .A(n14448), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14619) );
  NAND2_X1 U17624 ( .A1(n16033), .A2(n15894), .ZN(n14449) );
  NAND2_X1 U17625 ( .A1(n20135), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14614) );
  OAI211_X1 U17626 ( .C1(n16037), .C2(n14450), .A(n14449), .B(n14614), .ZN(
        n14451) );
  AOI21_X1 U17627 ( .B1(n14452), .B2(n20158), .A(n14451), .ZN(n14453) );
  OAI21_X1 U17628 ( .B1(n14619), .B2(n19981), .A(n14453), .ZN(P1_U2980) );
  OAI21_X1 U17629 ( .B1(n14456), .B2(n14455), .A(n14454), .ZN(n16056) );
  AOI22_X1 U17630 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14457) );
  OAI21_X1 U17631 ( .B1(n16029), .B2(n15897), .A(n14457), .ZN(n14458) );
  AOI21_X1 U17632 ( .B1(n15903), .B2(n20158), .A(n14458), .ZN(n14459) );
  OAI21_X1 U17633 ( .B1(n19981), .B2(n16056), .A(n14459), .ZN(P1_U2981) );
  NOR2_X1 U17634 ( .A1(n16009), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14466) );
  INV_X1 U17635 ( .A(n14496), .ZN(n16010) );
  NOR2_X1 U17636 ( .A1(n14465), .A2(n14460), .ZN(n14483) );
  NOR2_X1 U17637 ( .A1(n14465), .A2(n14644), .ZN(n14486) );
  NOR3_X1 U17638 ( .A1(n16010), .A2(n14483), .A3(n14486), .ZN(n15997) );
  INV_X1 U17639 ( .A(n14461), .ZN(n14462) );
  AOI21_X1 U17640 ( .B1(n15997), .B2(n14463), .A(n14462), .ZN(n14464) );
  MUX2_X1 U17641 ( .A(n14466), .B(n14465), .S(n14464), .Z(n14467) );
  XNOR2_X1 U17642 ( .A(n14467), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14634) );
  NAND2_X1 U17643 ( .A1(n20135), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n14630) );
  OAI21_X1 U17644 ( .B1(n16037), .B2(n15908), .A(n14630), .ZN(n14469) );
  NOR2_X1 U17645 ( .A1(n15905), .A2(n20137), .ZN(n14468) );
  AOI211_X1 U17646 ( .C1(n16033), .C2(n15910), .A(n14469), .B(n14468), .ZN(
        n14470) );
  OAI21_X1 U17647 ( .B1(n14634), .B2(n19981), .A(n14470), .ZN(P1_U2982) );
  INV_X1 U17648 ( .A(n15928), .ZN(n14480) );
  AND2_X1 U17649 ( .A1(n14471), .A2(n15985), .ZN(n14476) );
  INV_X1 U17650 ( .A(n14472), .ZN(n14474) );
  NOR2_X1 U17651 ( .A1(n14496), .A2(n14473), .ZN(n15987) );
  NOR2_X1 U17652 ( .A1(n14474), .A2(n15987), .ZN(n14475) );
  XNOR2_X1 U17653 ( .A(n14476), .B(n14475), .ZN(n16076) );
  AOI22_X1 U17654 ( .A1(n20134), .A2(n16076), .B1(n20135), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n14477) );
  OAI21_X1 U17655 ( .B1(n16037), .B2(n14478), .A(n14477), .ZN(n14479) );
  AOI21_X1 U17656 ( .B1(n16033), .B2(n14480), .A(n14479), .ZN(n14481) );
  OAI21_X1 U17657 ( .B1(n14482), .B2(n20137), .A(n14481), .ZN(P1_U2984) );
  AOI21_X1 U17658 ( .B1(n16010), .B2(n14484), .A(n14483), .ZN(n14637) );
  INV_X1 U17659 ( .A(n14487), .ZN(n14485) );
  NOR2_X1 U17660 ( .A1(n14486), .A2(n14485), .ZN(n14636) );
  NAND2_X1 U17661 ( .A1(n14637), .A2(n14636), .ZN(n14635) );
  NAND2_X1 U17662 ( .A1(n14635), .A2(n14487), .ZN(n14488) );
  XOR2_X1 U17663 ( .A(n14489), .B(n14488), .Z(n16097) );
  NAND2_X1 U17664 ( .A1(n16097), .A2(n20134), .ZN(n14494) );
  INV_X1 U17665 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14490) );
  NOR2_X1 U17666 ( .A1(n20042), .A2(n14490), .ZN(n16091) );
  NOR2_X1 U17667 ( .A1(n16029), .A2(n14491), .ZN(n14492) );
  AOI211_X1 U17668 ( .C1(n20132), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16091), .B(n14492), .ZN(n14493) );
  OAI211_X1 U17669 ( .C1(n20137), .C2(n14495), .A(n14494), .B(n14493), .ZN(
        P1_U2986) );
  NAND2_X1 U17670 ( .A1(n14499), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14498) );
  XNOR2_X1 U17671 ( .A(n14496), .B(n14500), .ZN(n14497) );
  MUX2_X1 U17672 ( .A(n14498), .B(n14497), .S(n11423), .Z(n14503) );
  INV_X1 U17673 ( .A(n14499), .ZN(n14502) );
  NAND3_X1 U17674 ( .A1(n14502), .A2(n14501), .A3(n14500), .ZN(n16011) );
  NAND2_X1 U17675 ( .A1(n14503), .A2(n16011), .ZN(n16118) );
  NAND2_X1 U17676 ( .A1(n16118), .A2(n20134), .ZN(n14507) );
  OAI22_X1 U17677 ( .A1(n16037), .A2(n14504), .B1(n20042), .B2(n20775), .ZN(
        n14505) );
  AOI21_X1 U17678 ( .B1(n15959), .B2(n16033), .A(n14505), .ZN(n14506) );
  OAI211_X1 U17679 ( .C1(n20137), .C2(n15960), .A(n14507), .B(n14506), .ZN(
        P1_U2989) );
  NOR2_X1 U17680 ( .A1(n20932), .A2(n11365), .ZN(n14603) );
  NAND2_X1 U17681 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14514) );
  NAND3_X1 U17682 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14628) );
  NOR2_X1 U17683 ( .A1(n14627), .A2(n14628), .ZN(n16060) );
  NAND2_X1 U17684 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16060), .ZN(
        n14526) );
  OR2_X1 U17685 ( .A1(n16094), .A2(n14526), .ZN(n14612) );
  INV_X1 U17686 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14508) );
  INV_X1 U17687 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16138) );
  NAND2_X1 U17688 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16139) );
  NOR2_X1 U17689 ( .A1(n16138), .A2(n16139), .ZN(n16111) );
  NAND3_X1 U17690 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16111), .ZN(n14640) );
  NOR2_X1 U17691 ( .A1(n14508), .A2(n14640), .ZN(n14647) );
  NAND2_X1 U17692 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14647), .ZN(
        n14511) );
  INV_X1 U17693 ( .A(n14511), .ZN(n14620) );
  INV_X1 U17694 ( .A(n14510), .ZN(n16128) );
  NAND3_X1 U17695 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n16128), .ZN(n16130) );
  NOR2_X1 U17696 ( .A1(n11474), .A2(n16130), .ZN(n16112) );
  NAND2_X1 U17697 ( .A1(n14620), .A2(n16112), .ZN(n16101) );
  NOR2_X1 U17698 ( .A1(n14612), .A2(n16101), .ZN(n14601) );
  OR3_X1 U17699 ( .A1(n11474), .A2(n14510), .A3(n14509), .ZN(n14622) );
  OR2_X1 U17700 ( .A1(n14622), .A2(n14511), .ZN(n14528) );
  OAI21_X1 U17701 ( .B1(n14528), .B2(n14612), .A(n14623), .ZN(n14512) );
  OAI22_X1 U17702 ( .A1(n14514), .A2(n15846), .B1(n16133), .B2(n14621), .ZN(
        n15828) );
  OAI21_X1 U17703 ( .B1(n16064), .B2(n14603), .A(n15828), .ZN(n14591) );
  AOI21_X1 U17704 ( .B1(n14623), .B2(n14429), .A(n14591), .ZN(n14575) );
  INV_X1 U17705 ( .A(n14515), .ZN(n14516) );
  NAND2_X1 U17706 ( .A1(n14516), .A2(n14575), .ZN(n14517) );
  AND2_X1 U17707 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14531) );
  NAND2_X1 U17708 ( .A1(n14518), .A2(n14522), .ZN(n14568) );
  INV_X1 U17709 ( .A(n14556), .ZN(n14519) );
  NAND2_X1 U17710 ( .A1(n14522), .A2(n14519), .ZN(n14520) );
  NAND2_X1 U17711 ( .A1(n14568), .A2(n14520), .ZN(n14549) );
  INV_X1 U17712 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14547) );
  AND2_X1 U17713 ( .A1(n16133), .A2(n14547), .ZN(n14521) );
  NAND3_X1 U17714 ( .A1(n14542), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14522), .ZN(n14524) );
  OAI211_X1 U17715 ( .C1(n14525), .C2(n16135), .A(n14524), .B(n14523), .ZN(
        n14534) );
  INV_X1 U17716 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14530) );
  NOR3_X1 U17717 ( .A1(n11365), .A2(n14527), .A3(n14526), .ZN(n14574) );
  NOR2_X1 U17718 ( .A1(n14642), .A2(n14528), .ZN(n14599) );
  INV_X1 U17719 ( .A(n14599), .ZN(n14613) );
  INV_X1 U17720 ( .A(n16112), .ZN(n14639) );
  NAND2_X1 U17721 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14620), .ZN(
        n14529) );
  NOR2_X1 U17722 ( .A1(n14639), .A2(n14529), .ZN(n16090) );
  NAND2_X1 U17723 ( .A1(n14643), .A2(n16090), .ZN(n14576) );
  NAND2_X1 U17724 ( .A1(n14574), .A2(n16082), .ZN(n14579) );
  NOR3_X1 U17725 ( .A1(n14530), .A2(n14429), .A3(n14579), .ZN(n16046) );
  AND2_X1 U17726 ( .A1(n16046), .A2(n14531), .ZN(n14571) );
  AND2_X1 U17727 ( .A1(n14556), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14532) );
  NAND2_X1 U17728 ( .A1(n14571), .A2(n14532), .ZN(n14541) );
  NOR3_X1 U17729 ( .A1(n14541), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14540), .ZN(n14533) );
  NOR2_X1 U17730 ( .A1(n14534), .A2(n14533), .ZN(n14535) );
  INV_X1 U17731 ( .A(n14537), .ZN(n14539) );
  AOI21_X1 U17732 ( .B1(n14539), .B2(n20145), .A(n14538), .ZN(n14545) );
  NAND2_X1 U17733 ( .A1(n14541), .A2(n14540), .ZN(n14543) );
  NAND2_X1 U17734 ( .A1(n14543), .A2(n14542), .ZN(n14544) );
  OAI211_X1 U17735 ( .C1(n14546), .C2(n16160), .A(n14545), .B(n14544), .ZN(
        P1_U3001) );
  NAND3_X1 U17736 ( .A1(n14571), .A2(n14556), .A3(n14547), .ZN(n14551) );
  AOI21_X1 U17737 ( .B1(n14549), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14548), .ZN(n14550) );
  OAI211_X1 U17738 ( .C1(n14552), .C2(n16135), .A(n14551), .B(n14550), .ZN(
        n14553) );
  AOI21_X1 U17739 ( .B1(n14554), .B2(n20140), .A(n14553), .ZN(n14555) );
  INV_X1 U17740 ( .A(n14555), .ZN(P1_U3002) );
  NOR2_X1 U17741 ( .A1(n14557), .A2(n14556), .ZN(n14564) );
  INV_X1 U17742 ( .A(n14568), .ZN(n14559) );
  AOI21_X1 U17743 ( .B1(n14559), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14558), .ZN(n14560) );
  OAI21_X1 U17744 ( .B1(n14561), .B2(n16135), .A(n14560), .ZN(n14563) );
  INV_X1 U17745 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14570) );
  NAND2_X1 U17746 ( .A1(n14565), .A2(n20145), .ZN(n14567) );
  OAI211_X1 U17747 ( .C1(n14568), .C2(n14570), .A(n14567), .B(n14566), .ZN(
        n14569) );
  AOI21_X1 U17748 ( .B1(n14571), .B2(n14570), .A(n14569), .ZN(n14572) );
  OAI21_X1 U17749 ( .B1(n14573), .B2(n16160), .A(n14572), .ZN(P1_U3004) );
  NAND2_X1 U17750 ( .A1(n14574), .A2(n14429), .ZN(n14589) );
  OAI21_X1 U17751 ( .B1(n14576), .B2(n14589), .A(n14575), .ZN(n14582) );
  OAI21_X1 U17752 ( .B1(n14578), .B2(n16135), .A(n14577), .ZN(n14581) );
  NOR3_X1 U17753 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14429), .A3(
        n14579), .ZN(n14580) );
  AOI211_X1 U17754 ( .C1(n14582), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14581), .B(n14580), .ZN(n14583) );
  OAI21_X1 U17755 ( .B1(n14584), .B2(n16160), .A(n14583), .ZN(P1_U3007) );
  INV_X1 U17756 ( .A(n16082), .ZN(n14629) );
  INV_X1 U17757 ( .A(n14585), .ZN(n14587) );
  AOI21_X1 U17758 ( .B1(n14587), .B2(n20145), .A(n14586), .ZN(n14588) );
  OAI21_X1 U17759 ( .B1(n14629), .B2(n14589), .A(n14588), .ZN(n14590) );
  AOI21_X1 U17760 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14591), .A(
        n14590), .ZN(n14592) );
  OAI21_X1 U17761 ( .B1(n14593), .B2(n16160), .A(n14592), .ZN(P1_U3008) );
  NAND2_X1 U17762 ( .A1(n14595), .A2(n14594), .ZN(n14596) );
  XOR2_X1 U17763 ( .A(n11365), .B(n14596), .Z(n15973) );
  INV_X1 U17764 ( .A(n15973), .ZN(n14608) );
  INV_X1 U17765 ( .A(n15875), .ZN(n14606) );
  INV_X1 U17766 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14597) );
  OAI22_X1 U17767 ( .A1(n11365), .A2(n15828), .B1(n20042), .B2(n14597), .ZN(
        n14605) );
  NOR3_X1 U17768 ( .A1(n16101), .A2(n14598), .A3(n9916), .ZN(n14600) );
  NOR2_X1 U17769 ( .A1(n14600), .A2(n14599), .ZN(n16095) );
  NOR2_X1 U17770 ( .A1(n16095), .A2(n14612), .ZN(n14610) );
  AOI21_X1 U17771 ( .B1(n20143), .B2(n14601), .A(n14610), .ZN(n14602) );
  NOR2_X1 U17772 ( .A1(n14602), .A2(n14609), .ZN(n15849) );
  NAND2_X1 U17773 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15849), .ZN(
        n15829) );
  AOI211_X1 U17774 ( .C1(n20932), .C2(n11365), .A(n14603), .B(n15829), .ZN(
        n14604) );
  AOI211_X1 U17775 ( .C1(n20145), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n14607) );
  OAI21_X1 U17776 ( .B1(n14608), .B2(n16160), .A(n14607), .ZN(P1_U3009) );
  OAI21_X1 U17777 ( .B1(n20143), .B2(n14610), .A(n14609), .ZN(n14611) );
  INV_X1 U17778 ( .A(n14611), .ZN(n15847) );
  AOI21_X1 U17779 ( .B1(n16101), .B2(n14613), .A(n14612), .ZN(n14617) );
  NAND2_X1 U17780 ( .A1(n15846), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14615) );
  OAI211_X1 U17781 ( .C1(n16135), .C2(n15889), .A(n14615), .B(n14614), .ZN(
        n14616) );
  AOI21_X1 U17782 ( .B1(n15847), .B2(n14617), .A(n14616), .ZN(n14618) );
  OAI21_X1 U17783 ( .B1(n14619), .B2(n16160), .A(n14618), .ZN(P1_U3012) );
  OAI22_X1 U17784 ( .A1(n14620), .A2(n14642), .B1(n16090), .B2(n16089), .ZN(
        n14625) );
  AOI21_X1 U17785 ( .B1(n14623), .B2(n14622), .A(n14621), .ZN(n16114) );
  OAI21_X1 U17786 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16095), .A(
        n16114), .ZN(n14624) );
  AOI211_X1 U17787 ( .C1(n14626), .C2(n16101), .A(n14625), .B(n14624), .ZN(
        n16093) );
  OAI21_X1 U17788 ( .B1(n16064), .B2(n16060), .A(n16093), .ZN(n16058) );
  OAI21_X1 U17789 ( .B1(n14629), .B2(n14628), .A(n14627), .ZN(n14632) );
  OAI21_X1 U17790 ( .B1(n15916), .B2(n16135), .A(n14630), .ZN(n14631) );
  AOI21_X1 U17791 ( .B1(n16058), .B2(n14632), .A(n14631), .ZN(n14633) );
  OAI21_X1 U17792 ( .B1(n14634), .B2(n16160), .A(n14633), .ZN(P1_U3014) );
  NAND3_X1 U17793 ( .A1(n16128), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n16156), .ZN(n16153) );
  NOR2_X1 U17794 ( .A1(n16153), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14648) );
  OAI21_X1 U17795 ( .B1(n14637), .B2(n14636), .A(n14635), .ZN(n14638) );
  INV_X1 U17796 ( .A(n14638), .ZN(n16008) );
  NOR2_X1 U17797 ( .A1(n14640), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16102) );
  OAI21_X1 U17798 ( .B1(n14640), .B2(n14639), .A(n16131), .ZN(n14641) );
  OAI211_X1 U17799 ( .C1(n14647), .C2(n14642), .A(n16114), .B(n14641), .ZN(
        n16107) );
  AOI21_X1 U17800 ( .B1(n14643), .B2(n16102), .A(n16107), .ZN(n14645) );
  OAI22_X1 U17801 ( .A1(n16008), .A2(n16160), .B1(n14645), .B2(n14644), .ZN(
        n14646) );
  AOI21_X1 U17802 ( .B1(n14648), .B2(n14647), .A(n14646), .ZN(n14650) );
  AOI22_X1 U17803 ( .A1(n15943), .A2(n20145), .B1(n20135), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14649) );
  NAND2_X1 U17804 ( .A1(n14650), .A2(n14649), .ZN(P1_U3019) );
  MUX2_X1 U17805 ( .A(n20605), .B(n20557), .S(n20606), .Z(n14651) );
  OAI21_X1 U17806 ( .B1(n20828), .B2(n14182), .A(n14651), .ZN(n14652) );
  MUX2_X1 U17807 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14652), .S(
        n20835), .Z(P1_U3477) );
  OR2_X1 U17808 ( .A1(n14182), .A2(n14653), .ZN(n14660) );
  INV_X1 U17809 ( .A(n14661), .ZN(n14655) );
  NAND3_X1 U17810 ( .A1(n14656), .A2(n14655), .A3(n14654), .ZN(n14657) );
  AND2_X1 U17811 ( .A1(n14658), .A2(n14657), .ZN(n14659) );
  AND2_X1 U17812 ( .A1(n14660), .A2(n14659), .ZN(n15793) );
  INV_X1 U17813 ( .A(n19975), .ZN(n14670) );
  INV_X1 U17814 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20899) );
  AOI22_X1 U17815 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n11288), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20899), .ZN(n14667) );
  NOR3_X1 U17816 ( .A1(n14661), .A2(n10286), .A3(n14671), .ZN(n14662) );
  AOI21_X1 U17817 ( .B1(n14667), .B2(n14663), .A(n14662), .ZN(n14664) );
  OAI21_X1 U17818 ( .B1(n15793), .B2(n14670), .A(n14664), .ZN(n14665) );
  MUX2_X1 U17819 ( .A(n14665), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n16165), .Z(P1_U3473) );
  INV_X1 U17820 ( .A(n14666), .ZN(n14669) );
  OAI222_X1 U17821 ( .A1(n14672), .A2(n14671), .B1(n14670), .B2(n14669), .C1(
        n14668), .C2(n14667), .ZN(n14673) );
  MUX2_X1 U17822 ( .A(n14673), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16165), .Z(P1_U3472) );
  INV_X1 U17823 ( .A(n19850), .ZN(n14674) );
  OAI21_X1 U17824 ( .B1(n14674), .B2(n19661), .A(n19187), .ZN(n14676) );
  NAND3_X1 U17825 ( .A1(n11750), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14674), 
        .ZN(n14675) );
  MUX2_X1 U17826 ( .A(n14676), .B(n14675), .S(n15585), .Z(n14678) );
  OAI21_X1 U17827 ( .B1(n19857), .B2(n19951), .A(n16473), .ZN(n14677) );
  NAND2_X1 U17828 ( .A1(n14678), .A2(n14677), .ZN(n14682) );
  CLKBUF_X2 U17829 ( .A(n19244), .Z(n19251) );
  AOI21_X1 U17830 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n14679), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14680) );
  AOI211_X1 U17831 ( .C1(n15853), .C2(n19251), .A(n14680), .B(n18951), .ZN(
        n14681) );
  MUX2_X1 U17832 ( .A(n14682), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14681), 
        .Z(P2_U3610) );
  XNOR2_X1 U17833 ( .A(n12935), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16184) );
  NAND4_X1 U17834 ( .A1(n16183), .A2(n19080), .A3(n12939), .A4(n16184), .ZN(
        n14690) );
  NOR3_X1 U17835 ( .A1(n14683), .A2(P2_EBX_REG_30__SCAN_IN), .A3(n19090), .ZN(
        n14688) );
  INV_X1 U17836 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19914) );
  OAI22_X1 U17837 ( .A1(n14684), .A2(n19024), .B1(n19914), .B2(n19059), .ZN(
        n14687) );
  OAI22_X1 U17838 ( .A1(n19133), .A2(n19100), .B1(n12978), .B2(n14685), .ZN(
        n14686) );
  NOR3_X1 U17839 ( .A1(n14688), .A2(n14687), .A3(n14686), .ZN(n14689) );
  OAI211_X1 U17840 ( .C1(n14714), .C2(n19105), .A(n14690), .B(n14689), .ZN(
        P2_U2824) );
  OAI211_X1 U17841 ( .C1(n14692), .C2(n14983), .A(n19080), .B(n14691), .ZN(
        n14700) );
  AOI21_X1 U17842 ( .B1(n14693), .B2(n9783), .A(n14773), .ZN(n15203) );
  AND2_X1 U17843 ( .A1(n14870), .A2(n14694), .ZN(n14695) );
  OR2_X1 U17844 ( .A1(n14853), .A2(n14695), .ZN(n15206) );
  INV_X1 U17845 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14696) );
  OAI22_X1 U17846 ( .A1(n19100), .A2(n15206), .B1(n19024), .B2(n14696), .ZN(
        n14698) );
  OAI22_X1 U17847 ( .A1(n19101), .A2(n12548), .B1(n12438), .B2(n19059), .ZN(
        n14697) );
  AOI211_X1 U17848 ( .C1(n19119), .C2(n15203), .A(n14698), .B(n14697), .ZN(
        n14699) );
  OAI211_X1 U17849 ( .C1(n19090), .C2(n14701), .A(n14700), .B(n14699), .ZN(
        P2_U2834) );
  AOI21_X1 U17850 ( .B1(n15028), .B2(n14702), .A(n19841), .ZN(n14712) );
  AOI22_X1 U17851 ( .A1(n14703), .A2(n19125), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n19117), .ZN(n14704) );
  OAI21_X1 U17852 ( .B1(n14705), .B2(n19024), .A(n14704), .ZN(n14710) );
  OAI21_X1 U17853 ( .B1(n19100), .B2(n14706), .A(n19058), .ZN(n14707) );
  AOI21_X1 U17854 ( .B1(P2_REIP_REG_17__SCAN_IN), .B2(n19122), .A(n14707), 
        .ZN(n14708) );
  OAI21_X1 U17855 ( .B1(n15252), .B2(n19105), .A(n14708), .ZN(n14709) );
  AOI211_X1 U17856 ( .C1(n14712), .C2(n14711), .A(n14710), .B(n14709), .ZN(
        n14713) );
  INV_X1 U17857 ( .A(n14713), .ZN(P2_U2838) );
  INV_X1 U17858 ( .A(n14714), .ZN(n14715) );
  NAND2_X1 U17859 ( .A1(n14715), .A2(n14790), .ZN(n14716) );
  OAI21_X1 U17860 ( .B1(n14790), .B2(n12978), .A(n14716), .ZN(P2_U2856) );
  INV_X1 U17861 ( .A(n14717), .ZN(n14803) );
  NAND2_X1 U17862 ( .A1(n14719), .A2(n14718), .ZN(n14802) );
  NAND3_X1 U17863 ( .A1(n14803), .A2(n14798), .A3(n14802), .ZN(n14721) );
  NAND2_X1 U17864 ( .A1(n14799), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14720) );
  OAI211_X1 U17865 ( .C1(n14799), .C2(n15112), .A(n14721), .B(n14720), .ZN(
        P2_U2858) );
  NAND2_X1 U17866 ( .A1(n14723), .A2(n14722), .ZN(n14725) );
  XNOR2_X1 U17867 ( .A(n14725), .B(n14724), .ZN(n14817) );
  OR2_X1 U17868 ( .A1(n14733), .A2(n14726), .ZN(n14727) );
  NAND2_X1 U17869 ( .A1(n14728), .A2(n14727), .ZN(n15120) );
  NOR2_X1 U17870 ( .A1(n15120), .A2(n14799), .ZN(n14729) );
  AOI21_X1 U17871 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14799), .A(n14729), .ZN(
        n14730) );
  OAI21_X1 U17872 ( .B1(n14817), .B2(n14785), .A(n14730), .ZN(P2_U2859) );
  NOR2_X1 U17873 ( .A1(n14743), .A2(n14731), .ZN(n14732) );
  AOI21_X1 U17874 ( .B1(n14736), .B2(n14735), .A(n14734), .ZN(n14818) );
  NAND2_X1 U17875 ( .A1(n14818), .A2(n14798), .ZN(n14738) );
  NAND2_X1 U17876 ( .A1(n14799), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14737) );
  OAI211_X1 U17877 ( .C1(n14799), .C2(n15128), .A(n14738), .B(n14737), .ZN(
        P2_U2860) );
  AOI21_X1 U17878 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n14742) );
  INV_X1 U17879 ( .A(n14742), .ZN(n14831) );
  NAND2_X1 U17880 ( .A1(n14799), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14746) );
  AOI21_X1 U17881 ( .B1(n14744), .B2(n14752), .A(n14743), .ZN(n16219) );
  NAND2_X1 U17882 ( .A1(n16219), .A2(n14790), .ZN(n14745) );
  OAI211_X1 U17883 ( .C1(n14831), .C2(n14785), .A(n14746), .B(n14745), .ZN(
        P2_U2861) );
  OAI21_X1 U17884 ( .B1(n14749), .B2(n14748), .A(n14747), .ZN(n14832) );
  NAND2_X1 U17885 ( .A1(n14799), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U17886 ( .A1(n14759), .A2(n14750), .ZN(n14751) );
  NAND2_X1 U17887 ( .A1(n16232), .A2(n14790), .ZN(n14753) );
  OAI211_X1 U17888 ( .C1(n14832), .C2(n14785), .A(n14754), .B(n14753), .ZN(
        P2_U2862) );
  AOI21_X1 U17889 ( .B1(n14756), .B2(n14755), .A(n9803), .ZN(n14757) );
  XOR2_X1 U17890 ( .A(n14758), .B(n14757), .Z(n14851) );
  OAI21_X1 U17891 ( .B1(n14761), .B2(n14760), .A(n14759), .ZN(n14953) );
  NOR2_X1 U17892 ( .A1(n14953), .A2(n14799), .ZN(n14762) );
  AOI21_X1 U17893 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14799), .A(n14762), .ZN(
        n14763) );
  OAI21_X1 U17894 ( .B1(n14851), .B2(n14785), .A(n14763), .ZN(P2_U2863) );
  NOR2_X1 U17895 ( .A1(n14765), .A2(n14764), .ZN(n14766) );
  OR2_X1 U17896 ( .A1(n9786), .A2(n14766), .ZN(n16268) );
  NOR2_X1 U17897 ( .A1(n16255), .A2(n14799), .ZN(n14767) );
  AOI21_X1 U17898 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n14799), .A(n14767), .ZN(
        n14768) );
  OAI21_X1 U17899 ( .B1(n16268), .B2(n14785), .A(n14768), .ZN(P2_U2864) );
  AOI21_X1 U17900 ( .B1(n14771), .B2(n14769), .A(n14770), .ZN(n14860) );
  NAND2_X1 U17901 ( .A1(n14860), .A2(n14798), .ZN(n14777) );
  NOR2_X1 U17902 ( .A1(n14773), .A2(n14772), .ZN(n14774) );
  OR2_X1 U17903 ( .A1(n14775), .A2(n14774), .ZN(n15198) );
  INV_X1 U17904 ( .A(n15198), .ZN(n15781) );
  NAND2_X1 U17905 ( .A1(n15781), .A2(n14790), .ZN(n14776) );
  OAI211_X1 U17906 ( .C1(n14790), .C2(n14778), .A(n14777), .B(n14776), .ZN(
        P2_U2865) );
  OAI21_X1 U17907 ( .B1(n14779), .B2(n14780), .A(n14769), .ZN(n14867) );
  NOR2_X1 U17908 ( .A1(n14790), .A2(n12548), .ZN(n14781) );
  AOI21_X1 U17909 ( .B1(n15203), .B2(n14790), .A(n14781), .ZN(n14782) );
  OAI21_X1 U17910 ( .B1(n14867), .B2(n14785), .A(n14782), .ZN(P2_U2866) );
  INV_X1 U17911 ( .A(n14779), .ZN(n14783) );
  OAI21_X1 U17912 ( .B1(n14795), .B2(n14784), .A(n14783), .ZN(n14875) );
  OR2_X1 U17913 ( .A1(n14875), .A2(n14785), .ZN(n14789) );
  NAND2_X1 U17914 ( .A1(n14794), .A2(n14786), .ZN(n14787) );
  NAND2_X1 U17915 ( .A1(n9783), .A2(n14787), .ZN(n14992) );
  NAND2_X1 U17916 ( .A1(n18976), .A2(n14790), .ZN(n14788) );
  OAI211_X1 U17917 ( .C1(n14790), .C2(n12544), .A(n14789), .B(n14788), .ZN(
        P2_U2867) );
  NAND2_X1 U17918 ( .A1(n14792), .A2(n14791), .ZN(n14793) );
  AND2_X1 U17919 ( .A1(n14794), .A2(n14793), .ZN(n18991) );
  INV_X1 U17920 ( .A(n18991), .ZN(n15232) );
  AOI21_X1 U17921 ( .B1(n14797), .B2(n14796), .A(n14795), .ZN(n14884) );
  NAND2_X1 U17922 ( .A1(n14884), .A2(n14798), .ZN(n14801) );
  NAND2_X1 U17923 ( .A1(n14799), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14800) );
  OAI211_X1 U17924 ( .C1(n15232), .C2(n14799), .A(n14801), .B(n14800), .ZN(
        P2_U2868) );
  NAND3_X1 U17925 ( .A1(n14803), .A2(n19175), .A3(n14802), .ZN(n14808) );
  AOI22_X1 U17926 ( .A1(n19173), .A2(n15109), .B1(n19172), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n14807) );
  AOI22_X1 U17927 ( .A1(n19134), .A2(BUF2_REG_29__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14806) );
  NAND2_X1 U17928 ( .A1(n16265), .A2(n14804), .ZN(n14805) );
  NAND4_X1 U17929 ( .A1(n14808), .A2(n14807), .A3(n14806), .A4(n14805), .ZN(
        P2_U2890) );
  AOI21_X1 U17930 ( .B1(n14811), .B2(n14809), .A(n12453), .ZN(n16200) );
  INV_X1 U17931 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19193) );
  NAND2_X1 U17932 ( .A1(n16265), .A2(n14812), .ZN(n14813) );
  OAI21_X1 U17933 ( .B1(n19193), .B2(n14836), .A(n14813), .ZN(n14814) );
  AOI21_X1 U17934 ( .B1(n19173), .B2(n16200), .A(n14814), .ZN(n14816) );
  AOI22_X1 U17935 ( .A1(n19134), .A2(BUF2_REG_28__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14815) );
  OAI211_X1 U17936 ( .C1(n14817), .C2(n19168), .A(n14816), .B(n14815), .ZN(
        P2_U2891) );
  INV_X1 U17937 ( .A(n14818), .ZN(n14824) );
  OAI21_X1 U17938 ( .B1(n14825), .B2(n14819), .A(n14809), .ZN(n16211) );
  OAI22_X1 U17939 ( .A1(n16267), .A2(n16211), .B1(n14836), .B2(n19195), .ZN(
        n14820) );
  AOI21_X1 U17940 ( .B1(n16265), .B2(n14821), .A(n14820), .ZN(n14823) );
  AOI22_X1 U17941 ( .A1(n19134), .A2(BUF2_REG_27__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14822) );
  OAI211_X1 U17942 ( .C1(n14824), .C2(n19168), .A(n14823), .B(n14822), .ZN(
        P2_U2892) );
  AOI21_X1 U17943 ( .B1(n14826), .B2(n14835), .A(n14825), .ZN(n16218) );
  INV_X1 U17944 ( .A(n16218), .ZN(n15143) );
  INV_X1 U17945 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19197) );
  OAI22_X1 U17946 ( .A1(n16267), .A2(n15143), .B1(n14836), .B2(n19197), .ZN(
        n14827) );
  AOI21_X1 U17947 ( .B1(n16265), .B2(n14828), .A(n14827), .ZN(n14830) );
  AOI22_X1 U17948 ( .A1(n19134), .A2(BUF2_REG_26__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14829) );
  OAI211_X1 U17949 ( .C1(n14831), .C2(n19168), .A(n14830), .B(n14829), .ZN(
        P2_U2893) );
  OR2_X1 U17950 ( .A1(n14832), .A2(n19168), .ZN(n14842) );
  NAND2_X1 U17951 ( .A1(n14845), .A2(n14833), .ZN(n14834) );
  NAND2_X1 U17952 ( .A1(n14835), .A2(n14834), .ZN(n16230) );
  OAI22_X1 U17953 ( .A1(n16267), .A2(n16230), .B1(n14836), .B2(n19199), .ZN(
        n14837) );
  INV_X1 U17954 ( .A(n14837), .ZN(n14841) );
  AOI22_X1 U17955 ( .A1(n19134), .A2(BUF2_REG_25__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14840) );
  NAND2_X1 U17956 ( .A1(n16265), .A2(n14838), .ZN(n14839) );
  NAND4_X1 U17957 ( .A1(n14842), .A2(n14841), .A3(n14840), .A4(n14839), .ZN(
        P2_U2894) );
  OR2_X1 U17958 ( .A1(n15182), .A2(n14843), .ZN(n14844) );
  NAND2_X1 U17959 ( .A1(n14845), .A2(n14844), .ZN(n16252) );
  AOI22_X1 U17960 ( .A1(n19134), .A2(BUF2_REG_24__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14848) );
  AOI22_X1 U17961 ( .A1(n16265), .A2(n14846), .B1(n19172), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n14847) );
  OAI211_X1 U17962 ( .C1(n16267), .C2(n16252), .A(n14848), .B(n14847), .ZN(
        n14849) );
  INV_X1 U17963 ( .A(n14849), .ZN(n14850) );
  OAI21_X1 U17964 ( .B1(n14851), .B2(n19168), .A(n14850), .ZN(P2_U2895) );
  OR2_X1 U17965 ( .A1(n14853), .A2(n14852), .ZN(n14855) );
  INV_X1 U17966 ( .A(n15179), .ZN(n14854) );
  NAND2_X1 U17967 ( .A1(n14855), .A2(n14854), .ZN(n15779) );
  AOI22_X1 U17968 ( .A1(n19134), .A2(BUF2_REG_22__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14858) );
  AOI22_X1 U17969 ( .A1(n16265), .A2(n14856), .B1(n19172), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n14857) );
  OAI211_X1 U17970 ( .C1(n16267), .C2(n15779), .A(n14858), .B(n14857), .ZN(
        n14859) );
  AOI21_X1 U17971 ( .B1(n14860), .B2(n19175), .A(n14859), .ZN(n14861) );
  INV_X1 U17972 ( .A(n14861), .ZN(P2_U2897) );
  AOI22_X1 U17973 ( .A1(n19134), .A2(BUF2_REG_21__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14864) );
  AOI22_X1 U17974 ( .A1(n16265), .A2(n14862), .B1(n19172), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n14863) );
  OAI211_X1 U17975 ( .C1(n16267), .C2(n15206), .A(n14864), .B(n14863), .ZN(
        n14865) );
  INV_X1 U17976 ( .A(n14865), .ZN(n14866) );
  OAI21_X1 U17977 ( .B1(n14867), .B2(n19168), .A(n14866), .ZN(P2_U2898) );
  NAND2_X1 U17978 ( .A1(n14879), .A2(n14868), .ZN(n14869) );
  NAND2_X1 U17979 ( .A1(n14870), .A2(n14869), .ZN(n18985) );
  AOI22_X1 U17980 ( .A1(n19134), .A2(BUF2_REG_20__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14872) );
  AOI22_X1 U17981 ( .A1(n16265), .A2(n19298), .B1(n19172), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n14871) );
  OAI211_X1 U17982 ( .C1(n16267), .C2(n18985), .A(n14872), .B(n14871), .ZN(
        n14873) );
  INV_X1 U17983 ( .A(n14873), .ZN(n14874) );
  OAI21_X1 U17984 ( .B1(n14875), .B2(n19168), .A(n14874), .ZN(P2_U2899) );
  OR2_X1 U17985 ( .A1(n14877), .A2(n14876), .ZN(n14878) );
  NAND2_X1 U17986 ( .A1(n14879), .A2(n14878), .ZN(n18989) );
  AOI22_X1 U17987 ( .A1(n19134), .A2(BUF2_REG_19__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14882) );
  AOI22_X1 U17988 ( .A1(n16265), .A2(n14880), .B1(n19172), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14881) );
  OAI211_X1 U17989 ( .C1(n16267), .C2(n18989), .A(n14882), .B(n14881), .ZN(
        n14883) );
  AOI21_X1 U17990 ( .B1(n14884), .B2(n19175), .A(n14883), .ZN(n14885) );
  INV_X1 U17991 ( .A(n14885), .ZN(P2_U2900) );
  INV_X1 U17992 ( .A(n14887), .ZN(n14889) );
  NAND2_X1 U17993 ( .A1(n14889), .A2(n14888), .ZN(n14890) );
  XNOR2_X1 U17994 ( .A(n14891), .B(n14890), .ZN(n15102) );
  XNOR2_X1 U17995 ( .A(n14900), .B(n15092), .ZN(n15100) );
  NOR2_X1 U17996 ( .A1(n16190), .A2(n16287), .ZN(n14894) );
  NAND2_X1 U17997 ( .A1(n19103), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15093) );
  NAND2_X1 U17998 ( .A1(n19256), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14892) );
  OAI211_X1 U17999 ( .C1(n19267), .C2(n16184), .A(n15093), .B(n14892), .ZN(
        n14893) );
  OAI21_X1 U18000 ( .B1(n15102), .B2(n19259), .A(n14895), .ZN(P2_U2984) );
  NOR2_X1 U18001 ( .A1(n14897), .A2(n14896), .ZN(n14899) );
  XOR2_X1 U18002 ( .A(n14899), .B(n14898), .Z(n15116) );
  AOI21_X1 U18003 ( .B1(n14901), .B2(n14916), .A(n14900), .ZN(n15114) );
  NAND2_X1 U18004 ( .A1(n19103), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15106) );
  OAI21_X1 U18005 ( .B1(n16338), .B2(n14902), .A(n15106), .ZN(n14903) );
  AOI21_X1 U18006 ( .B1(n16327), .B2(n14904), .A(n14903), .ZN(n14905) );
  OAI21_X1 U18007 ( .B1(n15112), .B2(n16287), .A(n14905), .ZN(n14906) );
  AOI21_X1 U18008 ( .B1(n15114), .B2(n9733), .A(n14906), .ZN(n14907) );
  OAI21_X1 U18009 ( .B1(n15116), .B2(n19259), .A(n14907), .ZN(P2_U2985) );
  INV_X1 U18010 ( .A(n14908), .ZN(n14910) );
  XNOR2_X1 U18011 ( .A(n14911), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14912) );
  XNOR2_X1 U18012 ( .A(n14913), .B(n14912), .ZN(n15127) );
  INV_X1 U18013 ( .A(n15120), .ZN(n16201) );
  INV_X1 U18014 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19907) );
  NOR2_X1 U18015 ( .A1(n19058), .A2(n19907), .ZN(n15118) );
  AOI21_X1 U18016 ( .B1(n19256), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15118), .ZN(n14914) );
  OAI21_X1 U18017 ( .B1(n19267), .B2(n16195), .A(n14914), .ZN(n14918) );
  NAND2_X1 U18018 ( .A1(n14921), .A2(n15117), .ZN(n14915) );
  NAND2_X1 U18019 ( .A1(n14916), .A2(n14915), .ZN(n15121) );
  NOR2_X1 U18020 ( .A1(n15121), .A2(n19257), .ZN(n14917) );
  AOI211_X1 U18021 ( .C1(n16201), .C2(n19263), .A(n14918), .B(n14917), .ZN(
        n14919) );
  OAI21_X1 U18022 ( .B1(n15127), .B2(n19259), .A(n14919), .ZN(P2_U2986) );
  XNOR2_X1 U18023 ( .A(n14920), .B(n15134), .ZN(n15139) );
  INV_X1 U18024 ( .A(n14921), .ZN(n14922) );
  AOI21_X1 U18025 ( .B1(n15134), .B2(n14933), .A(n14922), .ZN(n15137) );
  NAND2_X1 U18026 ( .A1(n19103), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15129) );
  OAI21_X1 U18027 ( .B1(n16338), .B2(n14923), .A(n15129), .ZN(n14924) );
  AOI21_X1 U18028 ( .B1(n16327), .B2(n16207), .A(n14924), .ZN(n14925) );
  OAI21_X1 U18029 ( .B1(n15128), .B2(n16287), .A(n14925), .ZN(n14926) );
  AOI21_X1 U18030 ( .B1(n15137), .B2(n9733), .A(n14926), .ZN(n14927) );
  OAI21_X1 U18031 ( .B1(n15139), .B2(n19259), .A(n14927), .ZN(P2_U2987) );
  OAI21_X1 U18032 ( .B1(n9862), .B2(n14937), .A(n14938), .ZN(n14930) );
  XNOR2_X1 U18033 ( .A(n14930), .B(n14929), .ZN(n15150) );
  NAND2_X1 U18034 ( .A1(n19103), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15142) );
  NAND2_X1 U18035 ( .A1(n19256), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14931) );
  OAI211_X1 U18036 ( .C1(n19267), .C2(n16222), .A(n15142), .B(n14931), .ZN(
        n14935) );
  INV_X1 U18037 ( .A(n14947), .ZN(n14932) );
  NOR2_X1 U18038 ( .A1(n14932), .A2(n15158), .ZN(n15152) );
  OAI21_X1 U18039 ( .B1(n15152), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14933), .ZN(n15147) );
  NOR2_X1 U18040 ( .A1(n15147), .A2(n19257), .ZN(n14934) );
  AOI211_X1 U18041 ( .C1(n16219), .C2(n19263), .A(n14935), .B(n14934), .ZN(
        n14936) );
  OAI21_X1 U18042 ( .B1(n15150), .B2(n19259), .A(n14936), .ZN(P2_U2988) );
  NAND2_X1 U18043 ( .A1(n10055), .A2(n14938), .ZN(n14939) );
  XNOR2_X1 U18044 ( .A(n9862), .B(n14939), .ZN(n15163) );
  NAND2_X1 U18045 ( .A1(n16327), .A2(n14940), .ZN(n14941) );
  NAND2_X1 U18046 ( .A1(n19103), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15155) );
  OAI211_X1 U18047 ( .C1(n16338), .C2(n16227), .A(n14941), .B(n15155), .ZN(
        n14943) );
  NOR2_X1 U18048 ( .A1(n14947), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15151) );
  NOR3_X1 U18049 ( .A1(n15152), .A2(n15151), .A3(n19257), .ZN(n14942) );
  AOI211_X1 U18050 ( .C1(n19263), .C2(n16232), .A(n14943), .B(n14942), .ZN(
        n14944) );
  OAI21_X1 U18051 ( .B1(n15163), .B2(n19259), .A(n14944), .ZN(P2_U2989) );
  NOR2_X1 U18052 ( .A1(n14945), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14946) );
  OR2_X1 U18053 ( .A1(n14947), .A2(n14946), .ZN(n15174) );
  INV_X1 U18054 ( .A(n14948), .ZN(n14950) );
  NOR2_X1 U18055 ( .A1(n14950), .A2(n14949), .ZN(n14951) );
  XNOR2_X1 U18056 ( .A(n14952), .B(n14951), .ZN(n15164) );
  NAND2_X1 U18057 ( .A1(n15164), .A2(n16335), .ZN(n14957) );
  INV_X1 U18058 ( .A(n14953), .ZN(n16243) );
  NAND2_X1 U18059 ( .A1(n19255), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U18060 ( .A1(n19256), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14954) );
  OAI211_X1 U18061 ( .C1(n19267), .C2(n16249), .A(n15165), .B(n14954), .ZN(
        n14955) );
  AOI21_X1 U18062 ( .B1(n16243), .B2(n19263), .A(n14955), .ZN(n14956) );
  OAI211_X1 U18063 ( .C1(n15174), .C2(n19257), .A(n14957), .B(n14956), .ZN(
        P2_U2990) );
  INV_X1 U18064 ( .A(n14959), .ZN(n14960) );
  NOR2_X1 U18065 ( .A1(n14961), .A2(n14960), .ZN(n14962) );
  XNOR2_X1 U18066 ( .A(n14958), .B(n14962), .ZN(n15202) );
  INV_X1 U18067 ( .A(n14963), .ZN(n14964) );
  AOI21_X1 U18068 ( .B1(n15194), .B2(n14984), .A(n14964), .ZN(n15200) );
  OAI22_X1 U18069 ( .A1(n20948), .A2(n19058), .B1(n19267), .B2(n15784), .ZN(
        n14967) );
  INV_X1 U18070 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14965) );
  OAI22_X1 U18071 ( .A1(n15198), .A2(n16287), .B1(n14965), .B2(n16338), .ZN(
        n14966) );
  AOI211_X1 U18072 ( .C1(n15200), .C2(n9733), .A(n14967), .B(n14966), .ZN(
        n14968) );
  OAI21_X1 U18073 ( .B1(n15202), .B2(n19259), .A(n14968), .ZN(P2_U2992) );
  INV_X1 U18074 ( .A(n14971), .ZN(n15038) );
  NAND2_X1 U18075 ( .A1(n15039), .A2(n15038), .ZN(n15037) );
  INV_X1 U18076 ( .A(n15013), .ZN(n14973) );
  INV_X1 U18077 ( .A(n14974), .ZN(n14975) );
  AND2_X1 U18078 ( .A1(n14976), .A2(n14977), .ZN(n14989) );
  NAND2_X1 U18079 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  NAND2_X1 U18080 ( .A1(n14988), .A2(n14977), .ZN(n14981) );
  NOR2_X1 U18081 ( .A1(n14979), .A2(n14978), .ZN(n14980) );
  XNOR2_X1 U18082 ( .A(n14981), .B(n14980), .ZN(n15214) );
  NAND2_X1 U18083 ( .A1(n19255), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15204) );
  NAND2_X1 U18084 ( .A1(n19256), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14982) );
  OAI211_X1 U18085 ( .C1(n19267), .C2(n14983), .A(n15204), .B(n14982), .ZN(
        n14986) );
  OAI21_X1 U18086 ( .B1(n14991), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14984), .ZN(n15211) );
  NOR2_X1 U18087 ( .A1(n15211), .A2(n19257), .ZN(n14985) );
  AOI211_X1 U18088 ( .C1(n19263), .C2(n15203), .A(n14986), .B(n14985), .ZN(
        n14987) );
  OAI21_X1 U18089 ( .B1(n15214), .B2(n19259), .A(n14987), .ZN(P2_U2993) );
  OAI21_X1 U18090 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n15226) );
  INV_X1 U18091 ( .A(n15002), .ZN(n15020) );
  NAND2_X1 U18092 ( .A1(n15020), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15004) );
  AOI21_X1 U18093 ( .B1(n15219), .B2(n15004), .A(n14991), .ZN(n15223) );
  NOR2_X1 U18094 ( .A1(n16287), .A2(n14992), .ZN(n14995) );
  NAND2_X1 U18095 ( .A1(n19103), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15216) );
  NAND2_X1 U18096 ( .A1(n19256), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14993) );
  OAI211_X1 U18097 ( .C1(n19267), .C2(n18982), .A(n15216), .B(n14993), .ZN(
        n14994) );
  AOI211_X1 U18098 ( .C1(n15223), .C2(n9733), .A(n14995), .B(n14994), .ZN(
        n14996) );
  OAI21_X1 U18099 ( .B1(n15226), .B2(n19259), .A(n14996), .ZN(P2_U2994) );
  NAND2_X1 U18100 ( .A1(n14998), .A2(n14997), .ZN(n15001) );
  INV_X1 U18101 ( .A(n15016), .ZN(n14999) );
  XOR2_X1 U18102 ( .A(n15001), .B(n15000), .Z(n15227) );
  NAND2_X1 U18103 ( .A1(n15002), .A2(n15230), .ZN(n15003) );
  NAND2_X1 U18104 ( .A1(n15004), .A2(n15003), .ZN(n15237) );
  OAI22_X1 U18105 ( .A1(n16338), .A2(n15006), .B1(n15005), .B2(n19058), .ZN(
        n15007) );
  AOI21_X1 U18106 ( .B1(n16327), .B2(n15008), .A(n15007), .ZN(n15010) );
  NAND2_X1 U18107 ( .A1(n19263), .A2(n18991), .ZN(n15009) );
  OAI211_X1 U18108 ( .C1(n15237), .C2(n19257), .A(n15010), .B(n15009), .ZN(
        n15011) );
  INV_X1 U18109 ( .A(n15011), .ZN(n15012) );
  OAI21_X1 U18110 ( .B1(n15227), .B2(n19259), .A(n15012), .ZN(P2_U2995) );
  NAND2_X1 U18111 ( .A1(n15016), .A2(n15013), .ZN(n15014) );
  AOI22_X1 U18112 ( .A1(n15017), .A2(n15016), .B1(n15015), .B2(n15014), .ZN(
        n15250) );
  NAND2_X1 U18113 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15019) );
  OR2_X1 U18114 ( .A1(n15042), .A2(n15019), .ZN(n15034) );
  AOI21_X1 U18115 ( .B1(n15240), .B2(n15034), .A(n15020), .ZN(n15248) );
  OAI22_X1 U18116 ( .A1(n19893), .A2(n19058), .B1(n19267), .B2(n19005), .ZN(
        n15022) );
  OAI22_X1 U18117 ( .A1(n16287), .A2(n18998), .B1(n10115), .B2(n16338), .ZN(
        n15021) );
  AOI211_X1 U18118 ( .C1(n15248), .C2(n9733), .A(n15022), .B(n15021), .ZN(
        n15023) );
  OAI21_X1 U18119 ( .B1(n15250), .B2(n19259), .A(n15023), .ZN(P2_U2996) );
  NAND2_X1 U18120 ( .A1(n10007), .A2(n15025), .ZN(n15026) );
  XNOR2_X1 U18121 ( .A(n15027), .B(n15026), .ZN(n15269) );
  INV_X1 U18122 ( .A(n15028), .ZN(n15030) );
  NAND2_X1 U18123 ( .A1(n19103), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15251) );
  NAND2_X1 U18124 ( .A1(n19256), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15029) );
  OAI211_X1 U18125 ( .C1(n19267), .C2(n15030), .A(n15251), .B(n15029), .ZN(
        n15031) );
  AOI21_X1 U18126 ( .B1(n19263), .B2(n15032), .A(n15031), .ZN(n15036) );
  NOR2_X1 U18127 ( .A1(n15042), .A2(n15033), .ZN(n15254) );
  OAI211_X1 U18128 ( .C1(n15254), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n9733), .B(n15034), .ZN(n15035) );
  OAI211_X1 U18129 ( .C1(n15269), .C2(n19259), .A(n15036), .B(n15035), .ZN(
        P2_U2997) );
  OAI21_X1 U18130 ( .B1(n15039), .B2(n15038), .A(n15037), .ZN(n15278) );
  INV_X1 U18131 ( .A(n19014), .ZN(n15272) );
  NAND2_X1 U18132 ( .A1(n19103), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15270) );
  OAI21_X1 U18133 ( .B1(n16338), .B2(n10118), .A(n15270), .ZN(n15041) );
  NOR2_X1 U18134 ( .A1(n19267), .A2(n19010), .ZN(n15040) );
  AOI211_X1 U18135 ( .C1(n15272), .C2(n19263), .A(n15041), .B(n15040), .ZN(
        n15044) );
  INV_X1 U18136 ( .A(n15042), .ZN(n15285) );
  INV_X1 U18137 ( .A(n15254), .ZN(n15260) );
  OAI211_X1 U18138 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15285), .A(
        n15260), .B(n9733), .ZN(n15043) );
  OAI211_X1 U18139 ( .C1(n15278), .C2(n19259), .A(n15044), .B(n15043), .ZN(
        P2_U2998) );
  NAND3_X1 U18140 ( .A1(n9778), .A2(n15045), .A3(n15279), .ZN(n15280) );
  INV_X1 U18141 ( .A(n15280), .ZN(n15048) );
  AOI22_X1 U18142 ( .A1(n9778), .A2(n16280), .B1(n15279), .B2(n15046), .ZN(
        n15047) );
  NOR2_X1 U18143 ( .A1(n15048), .A2(n15047), .ZN(n16349) );
  NAND2_X1 U18144 ( .A1(n15049), .A2(n15296), .ZN(n16295) );
  OR2_X1 U18145 ( .A1(n16295), .A2(n16340), .ZN(n16285) );
  INV_X1 U18146 ( .A(n15018), .ZN(n15050) );
  AOI21_X1 U18147 ( .B1(n16344), .B2(n16285), .A(n15050), .ZN(n16346) );
  OAI22_X1 U18148 ( .A1(n12408), .A2(n19058), .B1(n19267), .B2(n19039), .ZN(
        n15054) );
  INV_X1 U18149 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15051) );
  OAI22_X1 U18150 ( .A1(n16287), .A2(n15052), .B1(n16338), .B2(n15051), .ZN(
        n15053) );
  AOI211_X1 U18151 ( .C1(n16346), .C2(n9733), .A(n15054), .B(n15053), .ZN(
        n15056) );
  OAI21_X1 U18152 ( .B1(n16349), .B2(n19259), .A(n15056), .ZN(P2_U3000) );
  NAND2_X1 U18153 ( .A1(n15058), .A2(n15057), .ZN(n15060) );
  XOR2_X1 U18154 ( .A(n15060), .B(n15059), .Z(n15306) );
  NOR2_X1 U18155 ( .A1(n16287), .A2(n19052), .ZN(n15062) );
  INV_X1 U18156 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19884) );
  OAI22_X1 U18157 ( .A1(n19884), .A2(n19058), .B1(n19267), .B2(n19047), .ZN(
        n15061) );
  AOI211_X1 U18158 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19256), .A(
        n15062), .B(n15061), .ZN(n15065) );
  NAND2_X1 U18159 ( .A1(n16295), .A2(n12041), .ZN(n15304) );
  NOR2_X1 U18160 ( .A1(n12041), .A2(n16295), .ZN(n16286) );
  INV_X1 U18161 ( .A(n16286), .ZN(n15063) );
  NAND3_X1 U18162 ( .A1(n15304), .A2(n9733), .A3(n15063), .ZN(n15064) );
  OAI211_X1 U18163 ( .C1(n15306), .C2(n19259), .A(n15065), .B(n15064), .ZN(
        P2_U3002) );
  INV_X1 U18164 ( .A(n15066), .ZN(n15311) );
  NOR2_X1 U18165 ( .A1(n15067), .A2(n15311), .ZN(n15071) );
  NAND2_X1 U18166 ( .A1(n15069), .A2(n15068), .ZN(n15070) );
  XNOR2_X1 U18167 ( .A(n15071), .B(n15070), .ZN(n16382) );
  NAND2_X1 U18168 ( .A1(n15049), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15307) );
  OR2_X1 U18169 ( .A1(n15307), .A2(n12030), .ZN(n16294) );
  NAND2_X1 U18170 ( .A1(n15307), .A2(n12030), .ZN(n15072) );
  AND2_X1 U18171 ( .A1(n16294), .A2(n15072), .ZN(n16379) );
  INV_X1 U18172 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19880) );
  OAI22_X1 U18173 ( .A1(n19880), .A2(n19058), .B1(n19267), .B2(n19064), .ZN(
        n15074) );
  OAI22_X1 U18174 ( .A1(n16287), .A2(n19066), .B1(n16338), .B2(n10123), .ZN(
        n15073) );
  AOI211_X1 U18175 ( .C1(n16379), .C2(n9733), .A(n15074), .B(n15073), .ZN(
        n15075) );
  OAI21_X1 U18176 ( .B1(n16382), .B2(n19259), .A(n15075), .ZN(P2_U3004) );
  AOI21_X1 U18177 ( .B1(n15076), .B2(n15323), .A(n15324), .ZN(n15081) );
  INV_X1 U18178 ( .A(n15077), .ZN(n15079) );
  NAND2_X1 U18179 ( .A1(n15079), .A2(n15078), .ZN(n15080) );
  XNOR2_X1 U18180 ( .A(n15081), .B(n15080), .ZN(n16394) );
  OAI21_X1 U18181 ( .B1(n15084), .B2(n15083), .A(n15082), .ZN(n16389) );
  INV_X1 U18182 ( .A(n16389), .ZN(n15088) );
  OAI22_X1 U18183 ( .A1(n12345), .A2(n19058), .B1(n19267), .B2(n19076), .ZN(
        n15087) );
  INV_X1 U18184 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15085) );
  OAI22_X1 U18185 ( .A1(n16287), .A2(n19078), .B1(n16338), .B2(n15085), .ZN(
        n15086) );
  AOI211_X1 U18186 ( .C1(n15088), .C2(n9733), .A(n15087), .B(n15086), .ZN(
        n15089) );
  OAI21_X1 U18187 ( .B1(n16394), .B2(n19259), .A(n15089), .ZN(P2_U3006) );
  INV_X1 U18188 ( .A(n16190), .ZN(n15090) );
  NAND3_X1 U18189 ( .A1(n15105), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15092), .ZN(n15094) );
  OAI211_X1 U18190 ( .C1(n16189), .C2(n16413), .A(n15094), .B(n15093), .ZN(
        n15095) );
  NAND3_X1 U18191 ( .A1(n15098), .A2(n15097), .A3(n15096), .ZN(n15099) );
  AOI21_X1 U18192 ( .B1(n15100), .B2(n16400), .A(n15099), .ZN(n15101) );
  OAI21_X1 U18193 ( .B1(n15102), .B2(n16393), .A(n15101), .ZN(P2_U3016) );
  INV_X1 U18194 ( .A(n15103), .ZN(n15135) );
  OAI21_X1 U18195 ( .B1(n15104), .B2(n15130), .A(n15135), .ZN(n15125) );
  NAND2_X1 U18196 ( .A1(n15125), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15111) );
  INV_X1 U18197 ( .A(n15105), .ZN(n15107) );
  OAI21_X1 U18198 ( .B1(n15107), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15106), .ZN(n15108) );
  AOI21_X1 U18199 ( .B1(n16396), .B2(n15109), .A(n15108), .ZN(n15110) );
  OAI211_X1 U18200 ( .C1(n16388), .C2(n15112), .A(n15111), .B(n15110), .ZN(
        n15113) );
  AOI21_X1 U18201 ( .B1(n15114), .B2(n16400), .A(n15113), .ZN(n15115) );
  OAI21_X1 U18202 ( .B1(n15116), .B2(n16393), .A(n15115), .ZN(P2_U3017) );
  OAI21_X1 U18203 ( .B1(n15130), .B2(n15134), .A(n15117), .ZN(n15124) );
  AOI21_X1 U18204 ( .B1(n16396), .B2(n16200), .A(n15118), .ZN(n15119) );
  OAI21_X1 U18205 ( .B1(n15120), .B2(n16388), .A(n15119), .ZN(n15123) );
  NOR2_X1 U18206 ( .A1(n15121), .A2(n16420), .ZN(n15122) );
  AOI211_X1 U18207 ( .C1(n15125), .C2(n15124), .A(n15123), .B(n15122), .ZN(
        n15126) );
  OAI21_X1 U18208 ( .B1(n15127), .B2(n16393), .A(n15126), .ZN(P2_U3018) );
  INV_X1 U18209 ( .A(n15128), .ZN(n16213) );
  NOR2_X1 U18210 ( .A1(n16413), .A2(n16211), .ZN(n15132) );
  OAI21_X1 U18211 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15130), .A(
        n15129), .ZN(n15131) );
  AOI211_X1 U18212 ( .C1(n16213), .C2(n16417), .A(n15132), .B(n15131), .ZN(
        n15133) );
  OAI21_X1 U18213 ( .B1(n15135), .B2(n15134), .A(n15133), .ZN(n15136) );
  AOI21_X1 U18214 ( .B1(n15137), .B2(n16400), .A(n15136), .ZN(n15138) );
  OAI21_X1 U18215 ( .B1(n15139), .B2(n16393), .A(n15138), .ZN(P2_U3019) );
  OAI211_X1 U18216 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n10199), .B(n15153), .ZN(
        n15141) );
  OAI211_X1 U18217 ( .C1(n16413), .C2(n15143), .A(n15142), .B(n15141), .ZN(
        n15146) );
  NOR2_X1 U18218 ( .A1(n15159), .A2(n15144), .ZN(n15145) );
  AOI211_X1 U18219 ( .C1(n16219), .C2(n16417), .A(n15146), .B(n15145), .ZN(
        n15149) );
  OR2_X1 U18220 ( .A1(n15147), .A2(n16420), .ZN(n15148) );
  OAI211_X1 U18221 ( .C1(n15150), .C2(n16393), .A(n15149), .B(n15148), .ZN(
        P2_U3020) );
  NOR3_X1 U18222 ( .A1(n15152), .A2(n15151), .A3(n16420), .ZN(n15161) );
  NAND2_X1 U18223 ( .A1(n15153), .A2(n15158), .ZN(n15154) );
  OAI211_X1 U18224 ( .C1(n16413), .C2(n16230), .A(n15155), .B(n15154), .ZN(
        n15156) );
  AOI21_X1 U18225 ( .B1(n16232), .B2(n16417), .A(n15156), .ZN(n15157) );
  OAI21_X1 U18226 ( .B1(n15159), .B2(n15158), .A(n15157), .ZN(n15160) );
  NOR2_X1 U18227 ( .A1(n15161), .A2(n15160), .ZN(n15162) );
  OAI21_X1 U18228 ( .B1(n15163), .B2(n16393), .A(n15162), .ZN(P2_U3021) );
  NAND2_X1 U18229 ( .A1(n15164), .A2(n16423), .ZN(n15173) );
  OAI21_X1 U18230 ( .B1(n16413), .B2(n16252), .A(n15165), .ZN(n15171) );
  INV_X1 U18231 ( .A(n15166), .ZN(n15167) );
  AOI21_X1 U18232 ( .B1(n15169), .B2(n15168), .A(n15167), .ZN(n15170) );
  AOI211_X1 U18233 ( .C1(n16417), .C2(n16243), .A(n15171), .B(n15170), .ZN(
        n15172) );
  OAI211_X1 U18234 ( .C1(n16420), .C2(n15174), .A(n15173), .B(n15172), .ZN(
        P2_U3022) );
  INV_X1 U18235 ( .A(n15175), .ZN(n15191) );
  NAND3_X1 U18236 ( .A1(n10229), .A2(n16423), .A3(n15177), .ZN(n15190) );
  INV_X1 U18237 ( .A(n15178), .ZN(n15210) );
  NOR2_X1 U18238 ( .A1(n15180), .A2(n15179), .ZN(n15181) );
  OR2_X1 U18239 ( .A1(n15182), .A2(n15181), .ZN(n16266) );
  INV_X1 U18240 ( .A(n16266), .ZN(n15186) );
  OAI21_X1 U18241 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n15195), .ZN(n15183) );
  OAI22_X1 U18242 ( .A1(n19058), .A2(n13979), .B1(n15184), .B2(n15183), .ZN(
        n15185) );
  AOI21_X1 U18243 ( .B1(n16396), .B2(n15186), .A(n15185), .ZN(n15187) );
  OAI21_X1 U18244 ( .B1(n16255), .B2(n16388), .A(n15187), .ZN(n15188) );
  AOI21_X1 U18245 ( .B1(n15210), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15188), .ZN(n15189) );
  OAI211_X1 U18246 ( .C1(n15191), .C2(n16420), .A(n15190), .B(n15189), .ZN(
        P2_U3023) );
  NAND2_X1 U18247 ( .A1(n15210), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15197) );
  NOR2_X1 U18248 ( .A1(n20948), .A2(n19058), .ZN(n15193) );
  NOR2_X1 U18249 ( .A1(n16413), .A2(n15779), .ZN(n15192) );
  AOI211_X1 U18250 ( .C1(n15195), .C2(n15194), .A(n15193), .B(n15192), .ZN(
        n15196) );
  OAI211_X1 U18251 ( .C1(n15198), .C2(n16388), .A(n15197), .B(n15196), .ZN(
        n15199) );
  AOI21_X1 U18252 ( .B1(n15200), .B2(n16400), .A(n15199), .ZN(n15201) );
  OAI21_X1 U18253 ( .B1(n15202), .B2(n16393), .A(n15201), .ZN(P2_U3024) );
  NAND2_X1 U18254 ( .A1(n15203), .A2(n16417), .ZN(n15205) );
  OAI211_X1 U18255 ( .C1(n16413), .C2(n15206), .A(n15205), .B(n15204), .ZN(
        n15209) );
  NOR3_X1 U18256 ( .A1(n15231), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15207), .ZN(n15208) );
  AOI211_X1 U18257 ( .C1(n15210), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15209), .B(n15208), .ZN(n15213) );
  OR2_X1 U18258 ( .A1(n15211), .A2(n16420), .ZN(n15212) );
  OAI211_X1 U18259 ( .C1(n15214), .C2(n16393), .A(n15213), .B(n15212), .ZN(
        P2_U3025) );
  OAI21_X1 U18260 ( .B1(n15262), .B2(n15215), .A(n15297), .ZN(n15229) );
  INV_X1 U18261 ( .A(n15229), .ZN(n15222) );
  NAND2_X1 U18262 ( .A1(n16417), .A2(n18976), .ZN(n15217) );
  OAI211_X1 U18263 ( .C1(n16413), .C2(n18985), .A(n15217), .B(n15216), .ZN(
        n15221) );
  AOI211_X1 U18264 ( .C1(n15219), .C2(n15230), .A(n15218), .B(n15231), .ZN(
        n15220) );
  AOI211_X1 U18265 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15222), .A(
        n15221), .B(n15220), .ZN(n15225) );
  NAND2_X1 U18266 ( .A1(n15223), .A2(n16400), .ZN(n15224) );
  OAI211_X1 U18267 ( .C1(n15226), .C2(n16393), .A(n15225), .B(n15224), .ZN(
        P2_U3026) );
  OR2_X1 U18268 ( .A1(n15227), .A2(n16393), .ZN(n15236) );
  NAND2_X1 U18269 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19103), .ZN(n15228) );
  OAI221_X1 U18270 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15231), 
        .C1(n15230), .C2(n15229), .A(n15228), .ZN(n15234) );
  OAI22_X1 U18271 ( .A1(n16388), .A2(n15232), .B1(n16413), .B2(n18989), .ZN(
        n15233) );
  NOR2_X1 U18272 ( .A1(n15234), .A2(n15233), .ZN(n15235) );
  OAI211_X1 U18273 ( .C1(n15237), .C2(n16420), .A(n15236), .B(n15235), .ZN(
        P2_U3027) );
  NOR2_X1 U18274 ( .A1(n16413), .A2(n19008), .ZN(n15247) );
  INV_X1 U18275 ( .A(n15262), .ZN(n15238) );
  AOI211_X1 U18276 ( .C1(n15239), .C2(n15238), .A(n16362), .B(n15240), .ZN(
        n15244) );
  INV_X1 U18277 ( .A(n15239), .ZN(n15242) );
  NAND2_X1 U18278 ( .A1(n15286), .A2(n15240), .ZN(n15241) );
  NOR2_X1 U18279 ( .A1(n15242), .A2(n15241), .ZN(n15243) );
  AOI211_X1 U18280 ( .C1(n19103), .C2(P2_REIP_REG_18__SCAN_IN), .A(n15244), 
        .B(n15243), .ZN(n15245) );
  OAI21_X1 U18281 ( .B1(n16388), .B2(n18998), .A(n15245), .ZN(n15246) );
  AOI211_X1 U18282 ( .C1(n15248), .C2(n16400), .A(n15247), .B(n15246), .ZN(
        n15249) );
  OAI21_X1 U18283 ( .B1(n15250), .B2(n16393), .A(n15249), .ZN(P2_U3028) );
  OAI21_X1 U18284 ( .B1(n16388), .B2(n15252), .A(n15251), .ZN(n15257) );
  AOI22_X1 U18285 ( .A1(n15254), .A2(n16400), .B1(n15253), .B2(n15286), .ZN(
        n15255) );
  NOR2_X1 U18286 ( .A1(n15255), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15256) );
  AOI211_X1 U18287 ( .C1(n16396), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        n15268) );
  INV_X1 U18288 ( .A(n15259), .ZN(n15261) );
  OAI21_X1 U18289 ( .B1(n16400), .B2(n15261), .A(n15260), .ZN(n15263) );
  NAND2_X1 U18290 ( .A1(n15262), .A2(n15297), .ZN(n15292) );
  OAI211_X1 U18291 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15264), .A(
        n15263), .B(n15292), .ZN(n15276) );
  NOR2_X1 U18292 ( .A1(n15265), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15266) );
  OAI21_X1 U18293 ( .B1(n15276), .B2(n15266), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15267) );
  OAI211_X1 U18294 ( .C1(n15269), .C2(n16393), .A(n15268), .B(n15267), .ZN(
        P2_U3029) );
  AOI22_X1 U18295 ( .A1(n15285), .A2(n16400), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15286), .ZN(n15274) );
  OAI21_X1 U18296 ( .B1(n16413), .B2(n19015), .A(n15270), .ZN(n15271) );
  AOI21_X1 U18297 ( .B1(n16417), .B2(n15272), .A(n15271), .ZN(n15273) );
  OAI21_X1 U18298 ( .B1(n15274), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15273), .ZN(n15275) );
  AOI21_X1 U18299 ( .B1(n15276), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15275), .ZN(n15277) );
  OAI21_X1 U18300 ( .B1(n15278), .B2(n16393), .A(n15277), .ZN(P2_U3030) );
  NAND2_X1 U18301 ( .A1(n15280), .A2(n15279), .ZN(n15284) );
  NAND2_X1 U18302 ( .A1(n15282), .A2(n15281), .ZN(n15283) );
  XNOR2_X1 U18303 ( .A(n15284), .B(n15283), .ZN(n16273) );
  AOI21_X1 U18304 ( .B1(n15291), .B2(n15018), .A(n15285), .ZN(n16274) );
  NAND2_X1 U18305 ( .A1(n15286), .A2(n15291), .ZN(n15290) );
  INV_X1 U18306 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19888) );
  NOR2_X1 U18307 ( .A1(n19888), .A2(n19058), .ZN(n15288) );
  NOR2_X1 U18308 ( .A1(n16413), .A2(n19035), .ZN(n15287) );
  AOI211_X1 U18309 ( .C1(n16275), .C2(n16417), .A(n15288), .B(n15287), .ZN(
        n15289) );
  OAI211_X1 U18310 ( .C1(n15292), .C2(n15291), .A(n15290), .B(n15289), .ZN(
        n15293) );
  AOI21_X1 U18311 ( .B1(n16274), .B2(n16400), .A(n15293), .ZN(n15294) );
  OAI21_X1 U18312 ( .B1(n16273), .B2(n16393), .A(n15294), .ZN(P2_U3031) );
  NOR2_X1 U18313 ( .A1(n16420), .A2(n16286), .ZN(n15303) );
  NAND2_X1 U18314 ( .A1(n15296), .A2(n15295), .ZN(n16351) );
  INV_X1 U18315 ( .A(n15296), .ZN(n15298) );
  OAI21_X1 U18316 ( .B1(n15298), .B2(n15314), .A(n15297), .ZN(n16341) );
  NAND2_X1 U18317 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19103), .ZN(n15299) );
  OAI221_X1 U18318 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16351), 
        .C1(n12041), .C2(n16341), .A(n15299), .ZN(n15302) );
  XNOR2_X1 U18319 ( .A(n15300), .B(n9816), .ZN(n19053) );
  OAI22_X1 U18320 ( .A1(n19053), .A2(n16413), .B1(n16388), .B2(n19052), .ZN(
        n15301) );
  AOI211_X1 U18321 ( .C1(n15304), .C2(n15303), .A(n15302), .B(n15301), .ZN(
        n15305) );
  OAI21_X1 U18322 ( .B1(n15306), .B2(n16393), .A(n15305), .ZN(P2_U3034) );
  INV_X1 U18323 ( .A(n15049), .ZN(n15309) );
  INV_X1 U18324 ( .A(n15307), .ZN(n15308) );
  AOI21_X1 U18325 ( .B1(n15309), .B2(n16369), .A(n15308), .ZN(n16312) );
  INV_X1 U18326 ( .A(n16312), .ZN(n15322) );
  NOR2_X1 U18327 ( .A1(n15311), .A2(n15310), .ZN(n15312) );
  XNOR2_X1 U18328 ( .A(n15313), .B(n15312), .ZN(n16311) );
  NOR2_X1 U18329 ( .A1(n16369), .A2(n15314), .ZN(n16361) );
  AOI21_X1 U18330 ( .B1(n16369), .B2(n16368), .A(n16361), .ZN(n15316) );
  NOR2_X1 U18331 ( .A1(n19058), .A2(n19878), .ZN(n15315) );
  AOI211_X1 U18332 ( .C1(n16396), .C2(n15317), .A(n15316), .B(n15315), .ZN(
        n15318) );
  OAI21_X1 U18333 ( .B1(n16388), .B2(n15319), .A(n15318), .ZN(n15320) );
  AOI21_X1 U18334 ( .B1(n16311), .B2(n16423), .A(n15320), .ZN(n15321) );
  OAI21_X1 U18335 ( .B1(n15322), .B2(n16420), .A(n15321), .ZN(P2_U3037) );
  INV_X1 U18336 ( .A(n15323), .ZN(n15325) );
  NOR2_X1 U18337 ( .A1(n15325), .A2(n15324), .ZN(n15326) );
  XNOR2_X1 U18338 ( .A(n15076), .B(n15326), .ZN(n16321) );
  XNOR2_X1 U18339 ( .A(n15327), .B(n12018), .ZN(n15328) );
  XNOR2_X1 U18340 ( .A(n15329), .B(n15328), .ZN(n16317) );
  AOI21_X1 U18341 ( .B1(n15331), .B2(n15330), .A(n16397), .ZN(n16385) );
  NAND2_X1 U18342 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19255), .ZN(n15332) );
  OAI221_X1 U18343 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16383), .C1(
        n12018), .C2(n16385), .A(n15332), .ZN(n15336) );
  OAI22_X1 U18344 ( .A1(n16388), .A2(n15334), .B1(n16413), .B2(n15333), .ZN(
        n15335) );
  AOI211_X1 U18345 ( .C1(n16317), .C2(n16400), .A(n15336), .B(n15335), .ZN(
        n15337) );
  OAI21_X1 U18346 ( .B1(n16321), .B2(n16393), .A(n15337), .ZN(P2_U3039) );
  NOR2_X1 U18347 ( .A1(n15338), .A2(n16420), .ZN(n15349) );
  NOR2_X1 U18348 ( .A1(n15339), .A2(n16403), .ZN(n15341) );
  INV_X1 U18349 ( .A(n16385), .ZN(n15340) );
  MUX2_X1 U18350 ( .A(n15341), .B(n15340), .S(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n15348) );
  NOR2_X1 U18351 ( .A1(n16388), .A2(n19092), .ZN(n15347) );
  NOR2_X1 U18352 ( .A1(n15343), .A2(n15342), .ZN(n15344) );
  OR2_X1 U18353 ( .A1(n15345), .A2(n15344), .ZN(n19093) );
  OAI22_X1 U18354 ( .A1(n16413), .A2(n19093), .B1(n12329), .B2(n19058), .ZN(
        n15346) );
  NOR4_X1 U18355 ( .A1(n15349), .A2(n15348), .A3(n15347), .A4(n15346), .ZN(
        n15350) );
  OAI21_X1 U18356 ( .B1(n16393), .B2(n15351), .A(n15350), .ZN(P2_U3040) );
  INV_X2 U18357 ( .A(n9777), .ZN(n17286) );
  AOI22_X1 U18358 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9737), .ZN(n15353) );
  OAI21_X1 U18359 ( .B1(n10262), .B2(n18285), .A(n15353), .ZN(n15363) );
  NOR2_X2 U18360 ( .A1(n15354), .A2(n18741), .ZN(n15460) );
  AOI22_X1 U18361 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15361) );
  INV_X2 U18362 ( .A(n15493), .ZN(n17214) );
  AOI22_X1 U18363 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15360) );
  CLKBUF_X3 U18364 ( .A(n15419), .Z(n17289) );
  INV_X4 U18365 ( .A(n9775), .ZN(n17275) );
  AOI22_X1 U18366 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15359) );
  AOI22_X1 U18367 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15358) );
  NAND4_X1 U18368 ( .A1(n15361), .A2(n15360), .A3(n15359), .A4(n15358), .ZN(
        n15362) );
  AOI211_X2 U18369 ( .C1(n17284), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n15363), .B(n15362), .ZN(n15364) );
  AOI22_X1 U18370 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15374) );
  AOI22_X1 U18371 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9738), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U18372 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15367) );
  OAI21_X1 U18373 ( .B1(n10262), .B2(n18282), .A(n15367), .ZN(n15372) );
  AOI22_X1 U18374 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15371) );
  INV_X2 U18375 ( .A(n9777), .ZN(n17227) );
  AOI22_X1 U18376 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15370) );
  AOI22_X1 U18377 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U18378 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U18379 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15378) );
  AOI22_X1 U18380 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17272), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15377) );
  AOI22_X1 U18381 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15376) );
  AOI22_X1 U18382 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15375) );
  NAND4_X1 U18383 ( .A1(n15378), .A2(n15377), .A3(n15376), .A4(n15375), .ZN(
        n15384) );
  AOI22_X1 U18384 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15382) );
  INV_X2 U18385 ( .A(n10262), .ZN(n17238) );
  AOI22_X1 U18386 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15381) );
  AOI22_X1 U18387 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15380) );
  AOI22_X1 U18388 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15379) );
  NAND4_X1 U18389 ( .A1(n15382), .A2(n15381), .A3(n15380), .A4(n15379), .ZN(
        n15383) );
  AOI22_X1 U18390 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15388) );
  AOI22_X1 U18391 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15387) );
  AOI22_X1 U18392 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9739), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15386) );
  AOI22_X1 U18393 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15385) );
  NAND4_X1 U18394 ( .A1(n15388), .A2(n15387), .A3(n15386), .A4(n15385), .ZN(
        n15394) );
  AOI22_X1 U18395 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9741), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15392) );
  AOI22_X1 U18396 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15391) );
  AOI22_X1 U18397 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15390) );
  AOI22_X1 U18398 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15389) );
  NAND4_X1 U18399 ( .A1(n15392), .A2(n15391), .A3(n15390), .A4(n15389), .ZN(
        n15393) );
  AOI22_X1 U18400 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15398) );
  AOI22_X1 U18401 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15397) );
  AOI22_X1 U18402 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15396) );
  AOI22_X1 U18403 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15395) );
  NAND4_X1 U18404 ( .A1(n15398), .A2(n15397), .A3(n15396), .A4(n15395), .ZN(
        n15404) );
  AOI22_X1 U18405 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U18406 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15401) );
  AOI22_X1 U18407 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9738), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15400) );
  AOI22_X1 U18408 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15399) );
  NAND4_X1 U18409 ( .A1(n15402), .A2(n15401), .A3(n15400), .A4(n15399), .ZN(
        n15403) );
  AOI22_X1 U18410 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U18411 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15412) );
  INV_X1 U18412 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18302) );
  AOI22_X1 U18413 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15405) );
  OAI21_X1 U18414 ( .B1(n10262), .B2(n18302), .A(n15405), .ZN(n15411) );
  AOI22_X1 U18415 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15409) );
  AOI22_X1 U18416 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U18417 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U18418 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15406) );
  NAND4_X1 U18419 ( .A1(n15409), .A2(n15408), .A3(n15407), .A4(n15406), .ZN(
        n15410) );
  AOI22_X1 U18420 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U18421 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15416) );
  AOI22_X1 U18422 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15415) );
  AOI22_X1 U18423 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15414) );
  NAND4_X1 U18424 ( .A1(n15417), .A2(n15416), .A3(n15415), .A4(n15414), .ZN(
        n15425) );
  AOI22_X1 U18425 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15423) );
  AOI22_X1 U18426 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U18427 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15421) );
  AOI22_X1 U18428 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15420) );
  NAND4_X1 U18429 ( .A1(n15423), .A2(n15422), .A3(n15421), .A4(n15420), .ZN(
        n15424) );
  AOI22_X1 U18430 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15429) );
  AOI22_X1 U18431 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U18432 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15427) );
  AOI22_X1 U18433 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15426) );
  NAND4_X1 U18434 ( .A1(n15429), .A2(n15428), .A3(n15427), .A4(n15426), .ZN(
        n15436) );
  AOI22_X1 U18435 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15434) );
  AOI22_X1 U18436 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15433) );
  AOI22_X1 U18437 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9741), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U18438 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15431) );
  NAND4_X1 U18439 ( .A1(n15434), .A2(n15433), .A3(n15432), .A4(n15431), .ZN(
        n15435) );
  NOR2_X1 U18440 ( .A1(n18303), .A2(n15551), .ZN(n15718) );
  NAND3_X1 U18441 ( .A1(n15566), .A2(n15572), .A3(n15718), .ZN(n15727) );
  NAND2_X1 U18442 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15439), .ZN(
        n15441) );
  OAI22_X1 U18443 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15439), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21010), .ZN(n15443) );
  AOI21_X1 U18444 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15441), .A(
        n15443), .ZN(n15440) );
  NOR2_X1 U18445 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21010), .ZN(
        n15442) );
  AOI22_X1 U18446 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15443), .B1(
        n15442), .B2(n15441), .ZN(n15447) );
  OAI21_X1 U18447 ( .B1(n15446), .B2(n15445), .A(n15447), .ZN(n15444) );
  AOI21_X1 U18448 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18910), .A(
        n15574), .ZN(n15714) );
  NAND3_X1 U18449 ( .A1(n15575), .A2(n15447), .A3(n15714), .ZN(n15448) );
  NAND3_X1 U18450 ( .A1(n15576), .A2(n15577), .A3(n15448), .ZN(n18752) );
  NAND2_X1 U18451 ( .A1(n17333), .A2(n18303), .ZN(n15549) );
  INV_X1 U18452 ( .A(n15549), .ZN(n15552) );
  INV_X1 U18453 ( .A(n18294), .ZN(n15548) );
  AOI22_X1 U18454 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9739), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U18455 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15452) );
  INV_X2 U18456 ( .A(n10254), .ZN(n17053) );
  AOI22_X1 U18457 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U18458 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15450) );
  NAND4_X1 U18459 ( .A1(n15453), .A2(n15452), .A3(n15451), .A4(n15450), .ZN(
        n15459) );
  AOI22_X1 U18460 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U18461 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U18462 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U18463 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15454) );
  NAND4_X1 U18464 ( .A1(n15457), .A2(n15456), .A3(n15455), .A4(n15454), .ZN(
        n15458) );
  NOR2_X1 U18465 ( .A1(n15459), .A2(n15458), .ZN(n17078) );
  AOI22_X1 U18466 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15464) );
  AOI22_X1 U18467 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15463) );
  AOI22_X1 U18468 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15462) );
  AOI22_X1 U18469 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15461) );
  NAND4_X1 U18470 ( .A1(n15464), .A2(n15463), .A3(n15462), .A4(n15461), .ZN(
        n15470) );
  AOI22_X1 U18471 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15468) );
  AOI22_X1 U18472 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15467) );
  AOI22_X1 U18473 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U18474 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15465) );
  NAND4_X1 U18475 ( .A1(n15468), .A2(n15467), .A3(n15466), .A4(n15465), .ZN(
        n15469) );
  NOR2_X1 U18476 ( .A1(n15470), .A2(n15469), .ZN(n17088) );
  AOI22_X1 U18477 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17275), .ZN(n15474) );
  AOI22_X1 U18478 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15473) );
  AOI22_X1 U18479 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9741), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U18480 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17267), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17289), .ZN(n15471) );
  NAND4_X1 U18481 ( .A1(n15474), .A2(n15473), .A3(n15472), .A4(n15471), .ZN(
        n15480) );
  AOI22_X1 U18482 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9738), .ZN(n15478) );
  AOI22_X1 U18483 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9743), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U18484 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U18485 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n15669), .ZN(n15475) );
  NAND4_X1 U18486 ( .A1(n15478), .A2(n15477), .A3(n15476), .A4(n15475), .ZN(
        n15479) );
  NOR2_X1 U18487 ( .A1(n15480), .A2(n15479), .ZN(n17097) );
  AOI22_X1 U18488 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15491) );
  AOI22_X1 U18489 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U18490 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15482) );
  OAI21_X1 U18491 ( .B1(n10254), .B2(n18282), .A(n15482), .ZN(n15488) );
  AOI22_X1 U18492 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9741), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15486) );
  AOI22_X1 U18493 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15485) );
  AOI22_X1 U18494 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15484) );
  AOI22_X1 U18495 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15483) );
  NAND4_X1 U18496 ( .A1(n15486), .A2(n15485), .A3(n15484), .A4(n15483), .ZN(
        n15487) );
  AOI211_X1 U18497 ( .C1(n15595), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n15488), .B(n15487), .ZN(n15489) );
  NAND3_X1 U18498 ( .A1(n15491), .A2(n15490), .A3(n15489), .ZN(n17101) );
  AOI22_X1 U18499 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U18500 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15503) );
  INV_X1 U18501 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20889) );
  AOI22_X1 U18502 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15492) );
  OAI21_X1 U18503 ( .B1(n15493), .B2(n20889), .A(n15492), .ZN(n15501) );
  AOI22_X1 U18504 ( .A1(n15669), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15499) );
  AOI22_X1 U18505 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15498) );
  AOI22_X1 U18506 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U18507 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15496) );
  NAND4_X1 U18508 ( .A1(n15499), .A2(n15498), .A3(n15497), .A4(n15496), .ZN(
        n15500) );
  AOI211_X1 U18509 ( .C1(n15595), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n15501), .B(n15500), .ZN(n15502) );
  NAND3_X1 U18510 ( .A1(n15504), .A2(n15503), .A3(n15502), .ZN(n17102) );
  NAND2_X1 U18511 ( .A1(n17101), .A2(n17102), .ZN(n17100) );
  NOR2_X1 U18512 ( .A1(n17097), .A2(n17100), .ZN(n17094) );
  AOI22_X1 U18513 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15514) );
  AOI22_X1 U18514 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15513) );
  INV_X1 U18515 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n20995) );
  AOI22_X1 U18516 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15505) );
  OAI21_X1 U18517 ( .B1(n10262), .B2(n20995), .A(n15505), .ZN(n15511) );
  AOI22_X1 U18518 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U18519 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15508) );
  AOI22_X1 U18520 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15507) );
  AOI22_X1 U18521 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15506) );
  NAND4_X1 U18522 ( .A1(n15509), .A2(n15508), .A3(n15507), .A4(n15506), .ZN(
        n15510) );
  AOI211_X1 U18523 ( .C1(n17286), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n15511), .B(n15510), .ZN(n15512) );
  NAND3_X1 U18524 ( .A1(n15514), .A2(n15513), .A3(n15512), .ZN(n17093) );
  NAND2_X1 U18525 ( .A1(n17094), .A2(n17093), .ZN(n17092) );
  NOR2_X1 U18526 ( .A1(n17088), .A2(n17092), .ZN(n17353) );
  AOI22_X1 U18527 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15524) );
  AOI22_X1 U18528 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15523) );
  AOI22_X1 U18529 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15515) );
  OAI21_X1 U18530 ( .B1(n10254), .B2(n18302), .A(n15515), .ZN(n15521) );
  AOI22_X1 U18531 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U18532 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U18533 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15517) );
  AOI22_X1 U18534 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15516) );
  NAND4_X1 U18535 ( .A1(n15519), .A2(n15518), .A3(n15517), .A4(n15516), .ZN(
        n15520) );
  AOI211_X1 U18536 ( .C1(n17272), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n15521), .B(n15520), .ZN(n15522) );
  NAND3_X1 U18537 ( .A1(n15524), .A2(n15523), .A3(n15522), .ZN(n17352) );
  NAND2_X1 U18538 ( .A1(n17353), .A2(n17352), .ZN(n17351) );
  XNOR2_X1 U18539 ( .A(n17078), .B(n17351), .ZN(n17350) );
  AND2_X1 U18540 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17082) );
  NAND2_X1 U18541 ( .A1(n18316), .A2(n17324), .ZN(n17327) );
  INV_X1 U18542 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21154) );
  INV_X1 U18543 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17044) );
  INV_X1 U18544 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17106) );
  INV_X1 U18545 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16812) );
  INV_X1 U18546 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17168) );
  INV_X1 U18547 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17305) );
  INV_X1 U18548 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17311) );
  INV_X1 U18549 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17316) );
  INV_X1 U18550 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17325) );
  INV_X1 U18551 ( .A(n17144), .ZN(n17157) );
  NAND2_X1 U18552 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17104), .ZN(n17091) );
  NAND2_X1 U18553 ( .A1(n17331), .A2(n17087), .ZN(n17086) );
  OAI21_X1 U18554 ( .B1(n17082), .B2(n17327), .A(n17086), .ZN(n17083) );
  INV_X1 U18555 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21125) );
  NOR3_X1 U18556 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21125), .A3(n17087), .ZN(
        n15525) );
  AOI21_X1 U18557 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17083), .A(n15525), .ZN(
        n15526) );
  OAI21_X1 U18558 ( .B1(n17331), .B2(n17350), .A(n15526), .ZN(P3_U2675) );
  AOI22_X1 U18559 ( .A1(n15481), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15530) );
  AOI22_X1 U18560 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15529) );
  AOI22_X1 U18561 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9741), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U18562 ( .A1(n15653), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15527) );
  NAND4_X1 U18563 ( .A1(n15530), .A2(n15529), .A3(n15528), .A4(n15527), .ZN(
        n15536) );
  AOI22_X1 U18564 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15534) );
  AOI22_X1 U18565 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15533) );
  AOI22_X1 U18566 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15460), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U18567 ( .A1(n17274), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15531) );
  NAND4_X1 U18568 ( .A1(n15534), .A2(n15533), .A3(n15532), .A4(n15531), .ZN(
        n15535) );
  NOR2_X1 U18569 ( .A1(n15536), .A2(n15535), .ZN(n17423) );
  OAI21_X1 U18570 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n15537), .A(n17195), .ZN(
        n15538) );
  AOI22_X1 U18571 ( .A1(n17323), .A2(n17423), .B1(n15538), .B2(n17318), .ZN(
        P3_U2690) );
  OAI21_X1 U18572 ( .B1(n18930), .B2(n18889), .A(n18880), .ZN(n18267) );
  INV_X1 U18573 ( .A(n18267), .ZN(n18924) );
  NOR2_X1 U18574 ( .A1(n18889), .A2(n16675), .ZN(n17850) );
  INV_X1 U18575 ( .A(n17850), .ZN(n17781) );
  NAND2_X1 U18576 ( .A1(n18924), .A2(n17781), .ZN(n15544) );
  NAND2_X1 U18577 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18272) );
  NOR3_X1 U18578 ( .A1(n18933), .A2(n18930), .A3(n18889), .ZN(n15540) );
  INV_X1 U18579 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15584) );
  OAI21_X1 U18580 ( .B1(n15539), .B2(n18903), .A(n15584), .ZN(n15582) );
  OR2_X1 U18581 ( .A1(n15582), .A2(n9737), .ZN(n18264) );
  NOR2_X1 U18582 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18936) );
  AOI21_X1 U18583 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n18936), .ZN(n18788) );
  INV_X1 U18584 ( .A(n18367), .ZN(n18576) );
  INV_X1 U18585 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18265) );
  INV_X1 U18586 ( .A(n15540), .ZN(n18878) );
  NOR2_X1 U18587 ( .A1(n18265), .A2(n18878), .ZN(n15581) );
  AOI211_X1 U18588 ( .C1(n15540), .C2(n18264), .A(n18576), .B(n15581), .ZN(
        n15546) );
  AOI21_X1 U18589 ( .B1(n15544), .B2(n18272), .A(n15546), .ZN(n15547) );
  INV_X1 U18590 ( .A(n15547), .ZN(n15542) );
  NAND3_X1 U18591 ( .A1(n18930), .A2(n18880), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18620) );
  INV_X1 U18592 ( .A(n18620), .ZN(n18572) );
  NOR2_X1 U18593 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18880), .ZN(
        n18322) );
  OR2_X1 U18594 ( .A1(n18725), .A2(n18322), .ZN(n18366) );
  NOR3_X1 U18595 ( .A1(n18572), .A2(n15546), .A3(n18366), .ZN(n15541) );
  AOI21_X1 U18596 ( .B1(n18725), .B2(n15542), .A(n15541), .ZN(P3_U2864) );
  NAND2_X1 U18597 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18503) );
  INV_X1 U18598 ( .A(n18503), .ZN(n15543) );
  AOI21_X1 U18599 ( .B1(n18880), .B2(n15544), .A(n15543), .ZN(n15545) );
  NOR3_X1 U18600 ( .A1(n18322), .A2(n15546), .A3(n15545), .ZN(n18270) );
  INV_X1 U18601 ( .A(n15546), .ZN(n18271) );
  AOI22_X1 U18602 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15547), .B1(
        n18572), .B2(n18271), .ZN(n18269) );
  AOI22_X1 U18603 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18270), .B1(
        n18269), .B2(n18746), .ZN(P3_U2865) );
  INV_X1 U18604 ( .A(n18303), .ZN(n17336) );
  NAND2_X1 U18605 ( .A1(n18287), .A2(n15726), .ZN(n15564) );
  NOR2_X1 U18606 ( .A1(n17333), .A2(n18303), .ZN(n18720) );
  OAI211_X1 U18607 ( .C1(n18298), .C2(n18720), .A(n15566), .B(n15549), .ZN(
        n15550) );
  NOR3_X1 U18608 ( .A1(n15552), .A2(n15558), .A3(n17485), .ZN(n15555) );
  INV_X1 U18609 ( .A(n18720), .ZN(n15863) );
  NOR2_X1 U18610 ( .A1(n18298), .A2(n18316), .ZN(n15553) );
  AOI22_X1 U18611 ( .A1(n15863), .A2(n18298), .B1(n15711), .B2(n15553), .ZN(
        n15554) );
  AOI211_X1 U18612 ( .C1(n18294), .C2(n15556), .A(n15555), .B(n15554), .ZN(
        n15561) );
  NAND2_X1 U18613 ( .A1(n17485), .A2(n9961), .ZN(n15725) );
  INV_X1 U18614 ( .A(n15725), .ZN(n15557) );
  NAND2_X1 U18615 ( .A1(n17450), .A2(n15863), .ZN(n15864) );
  NAND2_X1 U18616 ( .A1(n15557), .A2(n15864), .ZN(n15560) );
  OAI211_X1 U18617 ( .C1(n15567), .C2(n15724), .A(n15561), .B(n15560), .ZN(
        n15719) );
  AOI221_X1 U18618 ( .B1(n15718), .B2(n15560), .C1(n15559), .C2(n15560), .A(
        n18294), .ZN(n15563) );
  INV_X1 U18619 ( .A(n15561), .ZN(n15562) );
  NAND2_X1 U18620 ( .A1(n15565), .A2(n15571), .ZN(n15728) );
  INV_X1 U18621 ( .A(n15566), .ZN(n15569) );
  NAND3_X1 U18622 ( .A1(n15569), .A2(n18929), .A3(n15568), .ZN(n15570) );
  NAND2_X1 U18623 ( .A1(n15571), .A2(n15570), .ZN(n15729) );
  NOR2_X1 U18624 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18793) );
  NAND2_X1 U18625 ( .A1(n9961), .A2(n17523), .ZN(n18772) );
  NAND2_X1 U18626 ( .A1(n15568), .A2(n18772), .ZN(n15573) );
  XNOR2_X1 U18627 ( .A(n15575), .B(n15574), .ZN(n15578) );
  AOI211_X1 U18628 ( .C1(n15859), .C2(n17483), .A(n18931), .B(n18749), .ZN(
        n15579) );
  INV_X1 U18629 ( .A(n18761), .ZN(n18744) );
  NOR2_X1 U18630 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18880), .ZN(n18276) );
  INV_X1 U18631 ( .A(n18911), .ZN(n18908) );
  AND2_X1 U18632 ( .A1(n15582), .A2(n18736), .ZN(n18760) );
  NAND3_X1 U18633 ( .A1(n18908), .A2(n18906), .A3(n18760), .ZN(n15583) );
  OAI21_X1 U18634 ( .B1(n18908), .B2(n15584), .A(n15583), .ZN(P3_U3284) );
  INV_X1 U18635 ( .A(n16452), .ZN(n15586) );
  NOR4_X1 U18636 ( .A1(n16451), .A2(n15586), .A3(n19924), .A4(n15585), .ZN(
        n15587) );
  NAND2_X1 U18637 ( .A1(n15590), .A2(n15587), .ZN(n15588) );
  OAI21_X1 U18638 ( .B1(n15590), .B2(n15589), .A(n15588), .ZN(P2_U3595) );
  AOI22_X1 U18639 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15594) );
  AOI22_X1 U18640 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15593) );
  AOI22_X1 U18641 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15592) );
  AOI22_X1 U18642 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15591) );
  NAND4_X1 U18643 ( .A1(n15594), .A2(n15593), .A3(n15592), .A4(n15591), .ZN(
        n15601) );
  AOI22_X1 U18644 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U18645 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U18646 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15597) );
  AOI22_X1 U18647 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15596) );
  NAND4_X1 U18648 ( .A1(n15599), .A2(n15598), .A3(n15597), .A4(n15596), .ZN(
        n15600) );
  AOI22_X1 U18649 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15606) );
  AOI22_X1 U18650 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9739), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15605) );
  AOI22_X1 U18651 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15604) );
  AOI22_X1 U18652 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15603) );
  NAND4_X1 U18653 ( .A1(n15606), .A2(n15605), .A3(n15604), .A4(n15603), .ZN(
        n15612) );
  AOI22_X1 U18654 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15610) );
  AOI22_X1 U18655 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15609) );
  AOI22_X1 U18656 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17272), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15608) );
  AOI22_X1 U18657 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15607) );
  NAND4_X1 U18658 ( .A1(n15610), .A2(n15609), .A3(n15608), .A4(n15607), .ZN(
        n15611) );
  AOI22_X1 U18659 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15616) );
  AOI22_X1 U18660 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15615) );
  AOI22_X1 U18661 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U18662 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15613) );
  NAND4_X1 U18663 ( .A1(n15616), .A2(n15615), .A3(n15614), .A4(n15613), .ZN(
        n15622) );
  AOI22_X1 U18664 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15620) );
  AOI22_X1 U18665 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9739), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15619) );
  AOI22_X1 U18666 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U18667 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15617) );
  NAND4_X1 U18668 ( .A1(n15620), .A2(n15619), .A3(n15618), .A4(n15617), .ZN(
        n15621) );
  AOI22_X1 U18669 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15634) );
  AOI22_X1 U18670 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15633) );
  AOI22_X1 U18671 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15623) );
  OAI21_X1 U18672 ( .B1(n9779), .B2(n20995), .A(n15623), .ZN(n15631) );
  AOI22_X1 U18673 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15629) );
  AOI22_X1 U18674 ( .A1(n17273), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15628) );
  AOI22_X1 U18675 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15494), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U18676 ( .A1(n17267), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15625), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15626) );
  NAND4_X1 U18677 ( .A1(n15629), .A2(n15628), .A3(n15627), .A4(n15626), .ZN(
        n15630) );
  NAND3_X1 U18678 ( .A1(n15634), .A2(n15633), .A3(n15632), .ZN(n15741) );
  AOI22_X1 U18679 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17273), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15642) );
  AOI22_X1 U18680 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15625), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17275), .ZN(n15641) );
  INV_X1 U18681 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20859) );
  INV_X2 U18682 ( .A(n17288), .ZN(n17239) );
  AOI22_X1 U18683 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15635) );
  OAI21_X1 U18684 ( .B1(n10254), .B2(n20859), .A(n15635), .ZN(n15640) );
  AOI22_X1 U18685 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17227), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n15669), .ZN(n15639) );
  AOI22_X1 U18686 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n9741), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n15653), .ZN(n15638) );
  AOI22_X1 U18687 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15637) );
  AOI22_X1 U18688 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17196), .ZN(n15636) );
  NAND2_X1 U18689 ( .A1(n15741), .A2(n15681), .ZN(n15668) );
  AOI22_X1 U18690 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U18691 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15651) );
  INV_X1 U18692 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21008) );
  AOI22_X1 U18693 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15643) );
  OAI21_X1 U18694 ( .B1(n9777), .B2(n21008), .A(n15643), .ZN(n15649) );
  AOI22_X1 U18695 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9739), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15647) );
  AOI22_X1 U18696 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15646) );
  AOI22_X1 U18697 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15645) );
  AOI22_X1 U18698 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15644) );
  NAND4_X1 U18699 ( .A1(n15647), .A2(n15646), .A3(n15645), .A4(n15644), .ZN(
        n15648) );
  AOI211_X1 U18700 ( .C1(n9743), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n15649), .B(n15648), .ZN(n15650) );
  NAND3_X1 U18701 ( .A1(n15652), .A2(n15651), .A3(n15650), .ZN(n15737) );
  NAND2_X1 U18702 ( .A1(n15667), .A2(n15737), .ZN(n15666) );
  AOI22_X1 U18703 ( .A1(n17273), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15663) );
  AOI22_X1 U18704 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15662) );
  AOI22_X1 U18705 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15653), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15654) );
  OAI21_X1 U18706 ( .B1(n9775), .B2(n18313), .A(n15654), .ZN(n15660) );
  AOI22_X1 U18707 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15658) );
  AOI22_X1 U18708 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U18709 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18710 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15655) );
  NAND4_X1 U18711 ( .A1(n15658), .A2(n15657), .A3(n15656), .A4(n15655), .ZN(
        n15659) );
  AOI211_X1 U18712 ( .C1(n17272), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n15660), .B(n15659), .ZN(n15661) );
  NAND3_X1 U18713 ( .A1(n15663), .A2(n15662), .A3(n15661), .ZN(n15736) );
  NAND2_X1 U18714 ( .A1(n15664), .A2(n15736), .ZN(n16553) );
  NAND2_X1 U18715 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17856), .ZN(
        n16548) );
  INV_X1 U18716 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17626) );
  INV_X1 U18717 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18074) );
  NAND2_X1 U18718 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18142) );
  NOR2_X1 U18719 ( .A1(n18142), .A2(n17819), .ZN(n18113) );
  NAND2_X1 U18720 ( .A1(n18113), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18099) );
  NOR2_X1 U18721 ( .A1(n18099), .A2(n18095), .ZN(n18101) );
  AND2_X1 U18722 ( .A1(n18101), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18083) );
  NAND2_X1 U18723 ( .A1(n18083), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15732) );
  AOI21_X1 U18724 ( .B1(n17451), .B2(n16553), .A(n17856), .ZN(n15696) );
  XOR2_X1 U18725 ( .A(n15736), .B(n15664), .Z(n15665) );
  NAND2_X1 U18726 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15665), .ZN(
        n15694) );
  XOR2_X1 U18727 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15665), .Z(
        n17875) );
  INV_X1 U18728 ( .A(n17458), .ZN(n15738) );
  XNOR2_X1 U18729 ( .A(n15738), .B(n15666), .ZN(n15690) );
  XOR2_X1 U18730 ( .A(n15737), .B(n15667), .Z(n15688) );
  XOR2_X1 U18731 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15688), .Z(
        n17898) );
  XOR2_X1 U18732 ( .A(n17466), .B(n15668), .Z(n15684) );
  INV_X1 U18733 ( .A(n15681), .ZN(n17482) );
  NAND2_X1 U18734 ( .A1(n17482), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15680) );
  AOI22_X1 U18735 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15673) );
  AOI22_X1 U18736 ( .A1(n17273), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15672) );
  AOI22_X1 U18737 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15671) );
  AOI22_X1 U18738 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15670) );
  NAND4_X1 U18739 ( .A1(n15673), .A2(n15672), .A3(n15671), .A4(n15670), .ZN(
        n15679) );
  AOI22_X1 U18740 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15677) );
  AOI22_X1 U18741 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U18742 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U18743 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15674) );
  NAND4_X1 U18744 ( .A1(n15677), .A2(n15676), .A3(n15675), .A4(n15674), .ZN(
        n15678) );
  INV_X1 U18745 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18907) );
  NOR2_X1 U18746 ( .A1(n17939), .A2(n18907), .ZN(n17938) );
  NAND2_X1 U18747 ( .A1(n17932), .A2(n17938), .ZN(n17931) );
  NAND2_X1 U18748 ( .A1(n15680), .A2(n17931), .ZN(n17921) );
  XNOR2_X1 U18749 ( .A(n15741), .B(n15681), .ZN(n15682) );
  INV_X1 U18750 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18236) );
  OR2_X1 U18751 ( .A1(n18236), .A2(n15682), .ZN(n15683) );
  NAND2_X1 U18752 ( .A1(n15684), .A2(n15686), .ZN(n15687) );
  NAND2_X1 U18753 ( .A1(n15687), .A2(n17911), .ZN(n17897) );
  NAND2_X1 U18754 ( .A1(n17898), .A2(n17897), .ZN(n17896) );
  NAND2_X1 U18755 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15688), .ZN(
        n15689) );
  NAND2_X1 U18756 ( .A1(n15690), .A2(n15692), .ZN(n15693) );
  NAND2_X1 U18757 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17885), .ZN(
        n17884) );
  NAND2_X1 U18758 ( .A1(n15693), .A2(n17884), .ZN(n17874) );
  NAND2_X1 U18759 ( .A1(n15696), .A2(n15695), .ZN(n15697) );
  INV_X1 U18760 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17841) );
  INV_X1 U18761 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18132) );
  OAI221_X1 U18762 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17792), 
        .C1(n18074), .C2(n15700), .A(n15699), .ZN(n17733) );
  INV_X1 U18763 ( .A(n15699), .ZN(n15701) );
  NAND2_X1 U18764 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18054) );
  INV_X1 U18765 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18024) );
  NAND2_X1 U18766 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18023) );
  NOR2_X1 U18767 ( .A1(n18024), .A2(n18023), .ZN(n18007) );
  NAND2_X1 U18768 ( .A1(n18007), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17594) );
  INV_X1 U18769 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21129) );
  INV_X1 U18770 ( .A(n18054), .ZN(n17728) );
  NAND2_X1 U18771 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17728), .ZN(
        n18020) );
  INV_X1 U18772 ( .A(n18020), .ZN(n17700) );
  NAND2_X1 U18773 ( .A1(n17700), .A2(n18007), .ZN(n18005) );
  NAND2_X1 U18774 ( .A1(n18010), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17992) );
  NOR2_X1 U18775 ( .A1(n17992), .A2(n17998), .ZN(n17644) );
  INV_X1 U18776 ( .A(n17644), .ZN(n17959) );
  NAND2_X1 U18777 ( .A1(n21129), .A2(n17792), .ZN(n17721) );
  NOR2_X1 U18778 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17721), .ZN(
        n15702) );
  INV_X1 U18779 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18006) );
  NAND2_X1 U18780 ( .A1(n15702), .A2(n18006), .ZN(n17681) );
  NOR2_X1 U18781 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17681), .ZN(
        n17666) );
  INV_X1 U18782 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17950) );
  NAND3_X1 U18783 ( .A1(n17666), .A2(n17950), .A3(n17998), .ZN(n15703) );
  NAND3_X1 U18784 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17655), .A3(
        n17650), .ZN(n15706) );
  INV_X1 U18785 ( .A(n15706), .ZN(n17639) );
  NAND2_X1 U18786 ( .A1(n17792), .A2(n17650), .ZN(n17638) );
  NAND2_X1 U18787 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17949) );
  OR2_X1 U18788 ( .A1(n15706), .A2(n17949), .ZN(n15707) );
  NAND2_X1 U18789 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15709), .ZN(
        n16552) );
  INV_X1 U18790 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17597) );
  NAND3_X1 U18791 ( .A1(n16563), .A2(n17597), .A3(n17792), .ZN(n15833) );
  OAI21_X1 U18792 ( .B1(n16548), .B2(n16552), .A(n15833), .ZN(n15710) );
  INV_X1 U18793 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16531) );
  INV_X1 U18794 ( .A(n15711), .ZN(n15713) );
  AOI21_X1 U18795 ( .B1(n18287), .B2(n15713), .A(n15712), .ZN(n15722) );
  AOI21_X1 U18796 ( .B1(n15715), .B2(n15714), .A(n18749), .ZN(n18756) );
  NAND2_X1 U18797 ( .A1(n18287), .A2(n18929), .ZN(n15716) );
  NOR2_X1 U18798 ( .A1(n18310), .A2(n15716), .ZN(n15723) );
  XNOR2_X1 U18799 ( .A(n18929), .B(n18287), .ZN(n15717) );
  OAI21_X1 U18800 ( .B1(n15717), .B2(n18928), .A(n18796), .ZN(n16654) );
  NOR3_X1 U18801 ( .A1(n15718), .A2(n18749), .A3(n16654), .ZN(n15720) );
  AOI211_X1 U18802 ( .C1(n18756), .C2(n15723), .A(n15720), .B(n15719), .ZN(
        n15721) );
  AOI221_X4 U18803 ( .B1(n15722), .B2(n15721), .C1(n18752), .C2(n15721), .A(
        n18925), .ZN(n18254) );
  NOR2_X1 U18804 ( .A1(n17451), .A2(n18757), .ZN(n16551) );
  INV_X1 U18805 ( .A(n18906), .ZN(n18881) );
  NOR2_X1 U18806 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18881), .ZN(n18944) );
  INV_X2 U18807 ( .A(n18148), .ZN(n18255) );
  NAND2_X1 U18808 ( .A1(n15726), .A2(n15725), .ZN(n18942) );
  INV_X1 U18809 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17953) );
  OR3_X1 U18810 ( .A1(n17998), .A2(n17986), .A3(n17949), .ZN(n17596) );
  NOR2_X1 U18811 ( .A1(n17992), .A2(n17596), .ZN(n16513) );
  NAND3_X1 U18812 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18081) );
  INV_X1 U18813 ( .A(n18081), .ZN(n15731) );
  NAND3_X1 U18814 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18180) );
  NAND2_X1 U18815 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18209) );
  NOR2_X1 U18816 ( .A1(n18180), .A2(n18209), .ZN(n18165) );
  NAND2_X1 U18817 ( .A1(n15731), .A2(n18165), .ZN(n18069) );
  NOR2_X1 U18818 ( .A1(n18907), .A2(n18069), .ZN(n18137) );
  NAND2_X1 U18819 ( .A1(n18048), .A2(n18137), .ZN(n18071) );
  NOR2_X1 U18820 ( .A1(n17615), .A2(n18071), .ZN(n15770) );
  NOR2_X1 U18821 ( .A1(n15732), .A2(n18069), .ZN(n18051) );
  NAND2_X1 U18822 ( .A1(n16513), .A2(n18051), .ZN(n15773) );
  AOI21_X1 U18823 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18207) );
  NOR2_X1 U18824 ( .A1(n18207), .A2(n18180), .ZN(n18166) );
  NAND2_X1 U18825 ( .A1(n18166), .A2(n15731), .ZN(n18070) );
  NOR2_X1 U18826 ( .A1(n15732), .A2(n18070), .ZN(n18053) );
  NAND2_X1 U18827 ( .A1(n17700), .A2(n18053), .ZN(n18004) );
  OR2_X1 U18828 ( .A1(n18004), .A2(n17594), .ZN(n17983) );
  NOR2_X1 U18829 ( .A1(n17596), .A2(n17983), .ZN(n15771) );
  NOR2_X1 U18830 ( .A1(n15771), .A2(n18739), .ZN(n17948) );
  AOI211_X1 U18831 ( .C1(n18716), .C2(n15773), .A(n17948), .B(n18217), .ZN(
        n15733) );
  OAI221_X1 U18832 ( .B1(n18732), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n18732), .C2(n15770), .A(n15733), .ZN(n15835) );
  AOI21_X1 U18833 ( .B1(n15734), .B2(n17953), .A(n15835), .ZN(n16555) );
  INV_X2 U18834 ( .A(n15734), .ZN(n18151) );
  NAND2_X1 U18835 ( .A1(n17597), .A2(n18168), .ZN(n15768) );
  NAND2_X1 U18836 ( .A1(n17451), .A2(n18260), .ZN(n18179) );
  INV_X1 U18837 ( .A(n18179), .ZN(n18107) );
  NAND2_X1 U18838 ( .A1(n18101), .A2(n17809), .ZN(n17773) );
  NOR2_X1 U18839 ( .A1(n17597), .A2(n17953), .ZN(n16517) );
  NAND2_X1 U18840 ( .A1(n16517), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15836) );
  INV_X1 U18841 ( .A(n15836), .ZN(n16497) );
  NAND2_X1 U18842 ( .A1(n17945), .A2(n16497), .ZN(n16504) );
  INV_X1 U18843 ( .A(n15736), .ZN(n17455) );
  INV_X1 U18844 ( .A(n15737), .ZN(n17462) );
  NOR2_X1 U18845 ( .A1(n17939), .A2(n17482), .ZN(n15742) );
  NOR2_X1 U18846 ( .A1(n15741), .A2(n15742), .ZN(n15740) );
  NAND2_X1 U18847 ( .A1(n15739), .A2(n15738), .ZN(n15756) );
  NAND2_X1 U18848 ( .A1(n15760), .A2(n16545), .ZN(n15761) );
  XOR2_X1 U18849 ( .A(n15739), .B(n15738), .Z(n15753) );
  XNOR2_X1 U18850 ( .A(n15740), .B(n17466), .ZN(n15747) );
  INV_X1 U18851 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18220) );
  NOR2_X1 U18852 ( .A1(n15747), .A2(n18220), .ZN(n15748) );
  INV_X1 U18853 ( .A(n15741), .ZN(n17472) );
  XNOR2_X1 U18854 ( .A(n17472), .B(n15742), .ZN(n15743) );
  NOR2_X1 U18855 ( .A1(n15743), .A2(n18236), .ZN(n15746) );
  XOR2_X1 U18856 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15743), .Z(
        n18234) );
  NOR2_X1 U18857 ( .A1(n17482), .A2(n18907), .ZN(n15745) );
  NAND3_X1 U18858 ( .A1(n17939), .A2(n17482), .A3(n18907), .ZN(n15744) );
  OAI221_X1 U18859 ( .B1(n15745), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n17939), .C2(n17482), .A(n15744), .ZN(n18233) );
  NOR2_X1 U18860 ( .A1(n18234), .A2(n18233), .ZN(n17923) );
  NOR2_X1 U18861 ( .A1(n15746), .A2(n17923), .ZN(n17910) );
  XOR2_X1 U18862 ( .A(n15747), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n17909) );
  NOR2_X1 U18863 ( .A1(n17910), .A2(n17909), .ZN(n17908) );
  NOR2_X1 U18864 ( .A1(n15748), .A2(n17908), .ZN(n15750) );
  XNOR2_X1 U18865 ( .A(n15749), .B(n17462), .ZN(n15751) );
  NOR2_X1 U18866 ( .A1(n15750), .A2(n15751), .ZN(n15752) );
  INV_X1 U18867 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18210) );
  XNOR2_X1 U18868 ( .A(n15751), .B(n15750), .ZN(n17902) );
  NOR2_X1 U18869 ( .A1(n18210), .A2(n17902), .ZN(n17901) );
  NOR2_X1 U18870 ( .A1(n15752), .A2(n17901), .ZN(n17888) );
  INV_X1 U18871 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15754) );
  XOR2_X1 U18872 ( .A(n15754), .B(n15753), .Z(n17887) );
  NOR2_X1 U18873 ( .A1(n17888), .A2(n17887), .ZN(n17886) );
  XNOR2_X1 U18874 ( .A(n15756), .B(n17455), .ZN(n15758) );
  NOR2_X1 U18875 ( .A1(n15757), .A2(n15758), .ZN(n15759) );
  XNOR2_X1 U18876 ( .A(n15758), .B(n15757), .ZN(n17879) );
  INV_X1 U18877 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18195) );
  NOR2_X1 U18878 ( .A1(n15759), .A2(n17878), .ZN(n15762) );
  XOR2_X1 U18879 ( .A(n15760), .B(n17451), .Z(n15763) );
  NAND2_X1 U18880 ( .A1(n15762), .A2(n15763), .ZN(n17860) );
  NAND2_X1 U18881 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17860), .ZN(
        n15765) );
  NOR2_X1 U18882 ( .A1(n15761), .A2(n15765), .ZN(n15767) );
  INV_X1 U18883 ( .A(n15761), .ZN(n15766) );
  OR2_X1 U18884 ( .A1(n15763), .A2(n15762), .ZN(n17861) );
  OAI21_X1 U18885 ( .B1(n15766), .B2(n15765), .A(n17861), .ZN(n15764) );
  AOI21_X1 U18886 ( .B1(n15766), .B2(n15765), .A(n15764), .ZN(n17855) );
  NAND2_X1 U18887 ( .A1(n17946), .A2(n16497), .ZN(n16505) );
  AOI22_X1 U18888 ( .A1(n18107), .A2(n16504), .B1(n18258), .B2(n16505), .ZN(
        n15837) );
  OAI221_X1 U18889 ( .B1(n18255), .B2(n16555), .C1(n18255), .C2(n15768), .A(
        n15837), .ZN(n15769) );
  AOI22_X1 U18890 ( .A1(n18255), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15769), .ZN(n15777) );
  AOI22_X1 U18891 ( .A1(n17946), .A2(n18258), .B1(n17945), .B2(n18107), .ZN(
        n15775) );
  INV_X1 U18892 ( .A(n18732), .ZN(n18721) );
  AOI22_X1 U18893 ( .A1(n18751), .A2(n15771), .B1(n15770), .B2(n18721), .ZN(
        n15772) );
  OAI21_X1 U18894 ( .B1(n15773), .B2(n18722), .A(n15772), .ZN(n15774) );
  NAND2_X1 U18895 ( .A1(n15774), .A2(n18254), .ZN(n16533) );
  NAND2_X1 U18896 ( .A1(n15775), .A2(n16533), .ZN(n15839) );
  NAND3_X1 U18897 ( .A1(n16517), .A2(n16531), .A3(n15839), .ZN(n15776) );
  OAI211_X1 U18898 ( .C1(n16529), .C2(n18162), .A(n15777), .B(n15776), .ZN(
        P3_U2833) );
  AOI22_X1 U18899 ( .A1(n15778), .A2(n19125), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19130), .ZN(n15788) );
  AOI22_X1 U18900 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19117), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19122), .ZN(n15787) );
  INV_X1 U18901 ( .A(n15779), .ZN(n15780) );
  AOI22_X1 U18902 ( .A1(n15781), .A2(n19119), .B1(n19121), .B2(n15780), .ZN(
        n15786) );
  OAI211_X1 U18903 ( .C1(n15784), .C2(n15783), .A(n19080), .B(n15782), .ZN(
        n15785) );
  NAND4_X1 U18904 ( .A1(n15788), .A2(n15787), .A3(n15786), .A4(n15785), .ZN(
        P2_U2833) );
  AOI21_X1 U18905 ( .B1(n15789), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20834), .ZN(n15790) );
  AND2_X1 U18906 ( .A1(n15791), .A2(n15790), .ZN(n15794) );
  OAI22_X1 U18907 ( .A1(n15793), .A2(n15792), .B1(n15794), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15797) );
  INV_X1 U18908 ( .A(n15794), .ZN(n15795) );
  OR2_X1 U18909 ( .A1(n15795), .A2(n20490), .ZN(n15796) );
  AND2_X1 U18910 ( .A1(n15797), .A2(n15796), .ZN(n15799) );
  INV_X1 U18911 ( .A(n15799), .ZN(n15801) );
  OAI21_X1 U18912 ( .B1(n15799), .B2(n20562), .A(n15798), .ZN(n15800) );
  OAI21_X1 U18913 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15801), .A(
        n15800), .ZN(n15803) );
  AOI222_X1 U18914 ( .A1(n15803), .A2(n20825), .B1(n15803), .B2(n15802), .C1(
        n20825), .C2(n15802), .ZN(n15810) );
  NOR3_X1 U18915 ( .A1(n15806), .A2(n15805), .A3(n15804), .ZN(n15809) );
  OAI21_X1 U18916 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15807), .ZN(n15808) );
  OAI211_X1 U18917 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15810), .A(
        n15809), .B(n15808), .ZN(n15818) );
  NAND2_X1 U18918 ( .A1(n15811), .A2(n20814), .ZN(n15815) );
  OAI21_X1 U18919 ( .B1(n20848), .B2(n15813), .A(n15812), .ZN(n15814) );
  OAI21_X1 U18920 ( .B1(n15816), .B2(n15815), .A(n15814), .ZN(n16178) );
  AOI221_X1 U18921 ( .B1(n9880), .B2(n11284), .C1(n15818), .C2(n11284), .A(
        n16178), .ZN(n16180) );
  AND2_X1 U18922 ( .A1(n15817), .A2(n16179), .ZN(n20832) );
  AOI21_X1 U18923 ( .B1(n15819), .B2(n15818), .A(n20832), .ZN(n15820) );
  OAI211_X1 U18924 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20848), .A(n15820), 
        .B(n16174), .ZN(n15821) );
  NOR2_X1 U18925 ( .A1(n16180), .A2(n15821), .ZN(n15825) );
  NAND2_X1 U18926 ( .A1(n20852), .A2(n15822), .ZN(n15823) );
  NAND2_X1 U18927 ( .A1(n9880), .A2(n15823), .ZN(n15824) );
  OAI22_X1 U18928 ( .A1(n15825), .A2(n9880), .B1(n16180), .B2(n15824), .ZN(
        P1_U3161) );
  INV_X1 U18929 ( .A(n15877), .ZN(n15831) );
  NAND2_X1 U18930 ( .A1(n20135), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15982) );
  OAI221_X1 U18931 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15829), 
        .C1(n20932), .C2(n15828), .A(n15982), .ZN(n15830) );
  AOI21_X1 U18932 ( .B1(n15831), .B2(n20145), .A(n15830), .ZN(n15832) );
  OAI21_X1 U18933 ( .B1(n15979), .B2(n16160), .A(n15832), .ZN(P1_U3010) );
  NOR2_X1 U18934 ( .A1(n16495), .A2(n16494), .ZN(n15834) );
  XOR2_X1 U18935 ( .A(n15834), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16516) );
  NOR2_X1 U18936 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15836), .ZN(
        n16512) );
  NAND2_X1 U18937 ( .A1(n18168), .A2(n18254), .ZN(n18242) );
  INV_X1 U18938 ( .A(n18242), .ZN(n16538) );
  AOI22_X1 U18939 ( .A1(n16538), .A2(n15836), .B1(n18148), .B2(n15835), .ZN(
        n16535) );
  INV_X1 U18940 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16506) );
  AOI21_X1 U18941 ( .B1(n16535), .B2(n15837), .A(n16506), .ZN(n15838) );
  AOI21_X1 U18942 ( .B1(n16512), .B2(n15839), .A(n15838), .ZN(n15840) );
  NAND2_X1 U18943 ( .A1(n18255), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16507) );
  OAI211_X1 U18944 ( .C1(n16516), .C2(n18162), .A(n15840), .B(n16507), .ZN(
        P3_U2832) );
  INV_X1 U18945 ( .A(HOLD), .ZN(n19855) );
  NAND2_X1 U18946 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20762), .ZN(n20753) );
  NAND2_X1 U18947 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20755) );
  INV_X1 U18948 ( .A(n20755), .ZN(n15841) );
  NOR2_X1 U18949 ( .A1(n19972), .A2(n20848), .ZN(n20756) );
  AOI221_X1 U18950 ( .B1(n19855), .B2(n15841), .C1(n20762), .C2(n15841), .A(
        n20756), .ZN(n15843) );
  OAI211_X1 U18951 ( .C1(n19855), .C2(n20753), .A(n15843), .B(n15842), .ZN(
        P1_U3195) );
  AND2_X1 U18952 ( .A1(n15844), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI221_X1 U18953 ( .B1(n15847), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), 
        .C1(n15846), .C2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15845), .ZN(
        n15851) );
  AOI22_X1 U18954 ( .A1(n15849), .A2(n11514), .B1(n20145), .B2(n15848), .ZN(
        n15850) );
  OAI211_X1 U18955 ( .C1(n15852), .C2(n16160), .A(n15851), .B(n15850), .ZN(
        P1_U3011) );
  NOR2_X1 U18956 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15854) );
  NOR2_X1 U18957 ( .A1(n21158), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19839) );
  INV_X1 U18958 ( .A(n19839), .ZN(n18950) );
  NOR2_X1 U18959 ( .A1(n15853), .A2(n18950), .ZN(n16465) );
  NOR4_X1 U18960 ( .A1(n15855), .A2(n15854), .A3(n16465), .A4(n16481), .ZN(
        P2_U3178) );
  INV_X1 U18961 ( .A(n16466), .ZN(n19964) );
  INV_X1 U18962 ( .A(n16473), .ZN(n15856) );
  AOI221_X1 U18963 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16481), .C1(n19964), .C2(
        n16481), .A(n19731), .ZN(n19956) );
  INV_X1 U18964 ( .A(n19956), .ZN(n19957) );
  NOR2_X1 U18965 ( .A1(n15858), .A2(n19957), .ZN(P2_U3047) );
  AOI22_X1 U18966 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17478), .B1(
        P3_EAX_REG_0__SCAN_IN), .B2(n17479), .ZN(n15866) );
  NAND3_X1 U18967 ( .A1(n17332), .A2(n18316), .A3(n17553), .ZN(n15865) );
  OAI211_X1 U18968 ( .C1(n17939), .C2(n17473), .A(n15866), .B(n15865), .ZN(
        P3_U2735) );
  INV_X1 U18969 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15882) );
  NOR4_X1 U18970 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15882), .A3(n15868), 
        .A4(n15867), .ZN(n15871) );
  OAI22_X1 U18971 ( .A1(n20060), .A2(n15869), .B1(n20054), .B2(n15977), .ZN(
        n15870) );
  AOI211_X1 U18972 ( .C1(n20059), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15871), .B(n15870), .ZN(n15874) );
  OAI21_X1 U18973 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n20021), .A(n15883), 
        .ZN(n15872) );
  AOI22_X1 U18974 ( .A1(n15974), .A2(n20031), .B1(P1_REIP_REG_22__SCAN_IN), 
        .B2(n15872), .ZN(n15873) );
  OAI211_X1 U18975 ( .C1(n20062), .C2(n15875), .A(n15874), .B(n15873), .ZN(
        P1_U2818) );
  AOI22_X1 U18976 ( .A1(n20046), .A2(P1_EBX_REG_21__SCAN_IN), .B1(n20059), 
        .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15881) );
  NOR3_X1 U18977 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20021), .A3(n15876), 
        .ZN(n15879) );
  OAI22_X1 U18978 ( .A1(n15978), .A2(n15890), .B1(n20062), .B2(n15877), .ZN(
        n15878) );
  AOI211_X1 U18979 ( .C1(n20040), .C2(n15981), .A(n15879), .B(n15878), .ZN(
        n15880) );
  OAI211_X1 U18980 ( .C1(n15883), .C2(n15882), .A(n15881), .B(n15880), .ZN(
        P1_U2819) );
  AOI21_X1 U18981 ( .B1(n20019), .B2(n15884), .A(n20017), .ZN(n15907) );
  NAND3_X1 U18982 ( .A1(n15885), .A2(n15952), .A3(n16063), .ZN(n15900) );
  NAND4_X1 U18983 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15885), .A3(n15952), 
        .A4(n15896), .ZN(n15887) );
  AOI21_X1 U18984 ( .B1(n20059), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20135), .ZN(n15886) );
  OAI211_X1 U18985 ( .C1(n15888), .C2(n20060), .A(n15887), .B(n15886), .ZN(
        n15893) );
  OAI22_X1 U18986 ( .A1(n15891), .A2(n15890), .B1(n20062), .B2(n15889), .ZN(
        n15892) );
  AOI211_X1 U18987 ( .C1(n15894), .C2(n20040), .A(n15893), .B(n15892), .ZN(
        n15895) );
  OAI221_X1 U18988 ( .B1(n15896), .B2(n15907), .C1(n15896), .C2(n15900), .A(
        n15895), .ZN(P1_U2821) );
  OAI22_X1 U18989 ( .A1(n20060), .A2(n15898), .B1(n20054), .B2(n15897), .ZN(
        n15899) );
  AOI211_X1 U18990 ( .C1(n20059), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20135), .B(n15899), .ZN(n15901) );
  OAI211_X1 U18991 ( .C1(n15907), .C2(n16063), .A(n15901), .B(n15900), .ZN(
        n15902) );
  AOI21_X1 U18992 ( .B1(n15903), .B2(n20031), .A(n15902), .ZN(n15904) );
  OAI21_X1 U18993 ( .B1(n20062), .B2(n16055), .A(n15904), .ZN(P1_U2822) );
  INV_X1 U18994 ( .A(n15905), .ZN(n15914) );
  INV_X1 U18995 ( .A(n15906), .ZN(n15936) );
  NAND4_X1 U18996 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n15936), .A4(n15952), .ZN(n15935) );
  AOI221_X1 U18997 ( .B1(n15917), .B2(n20785), .C1(n15935), .C2(n20785), .A(
        n15907), .ZN(n15913) );
  OAI21_X1 U18998 ( .B1(n20044), .B2(n15908), .A(n20042), .ZN(n15909) );
  AOI21_X1 U18999 ( .B1(n20040), .B2(n15910), .A(n15909), .ZN(n15911) );
  OAI21_X1 U19000 ( .B1(n14237), .B2(n20060), .A(n15911), .ZN(n15912) );
  AOI211_X1 U19001 ( .C1(n15914), .C2(n20031), .A(n15913), .B(n15912), .ZN(
        n15915) );
  OAI21_X1 U19002 ( .B1(n20062), .B2(n15916), .A(n15915), .ZN(P1_U2823) );
  OAI21_X1 U19003 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15917), .ZN(n15926) );
  INV_X1 U19004 ( .A(n15918), .ZN(n15990) );
  OAI21_X1 U19005 ( .B1(n15919), .B2(n15950), .A(n15951), .ZN(n15937) );
  INV_X1 U19006 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20963) );
  NAND2_X1 U19007 ( .A1(n20059), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15920) );
  OAI211_X1 U19008 ( .C1(n20054), .C2(n15993), .A(n20042), .B(n15920), .ZN(
        n15921) );
  AOI21_X1 U19009 ( .B1(n20046), .B2(P1_EBX_REG_16__SCAN_IN), .A(n15921), .ZN(
        n15923) );
  NAND2_X1 U19010 ( .A1(n16066), .A2(n20027), .ZN(n15922) );
  OAI211_X1 U19011 ( .C1(n15937), .C2(n20963), .A(n15923), .B(n15922), .ZN(
        n15924) );
  AOI21_X1 U19012 ( .B1(n15990), .B2(n20031), .A(n15924), .ZN(n15925) );
  OAI21_X1 U19013 ( .B1(n15935), .B2(n15926), .A(n15925), .ZN(P1_U2824) );
  INV_X1 U19014 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n16073) );
  AOI21_X1 U19015 ( .B1(n20059), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20135), .ZN(n15927) );
  OAI21_X1 U19016 ( .B1(n15928), .B2(n20054), .A(n15927), .ZN(n15930) );
  NOR2_X1 U19017 ( .A1(n16074), .A2(n20062), .ZN(n15929) );
  AOI211_X1 U19018 ( .C1(n20046), .C2(P1_EBX_REG_15__SCAN_IN), .A(n15930), .B(
        n15929), .ZN(n15931) );
  OAI21_X1 U19019 ( .B1(n15937), .B2(n16073), .A(n15931), .ZN(n15932) );
  AOI21_X1 U19020 ( .B1(n15933), .B2(n20031), .A(n15932), .ZN(n15934) );
  OAI21_X1 U19021 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15935), .A(n15934), 
        .ZN(P1_U2825) );
  AOI22_X1 U19022 ( .A1(n16000), .A2(n20040), .B1(n20027), .B2(n16083), .ZN(
        n15942) );
  AOI22_X1 U19023 ( .A1(n20046), .A2(P1_EBX_REG_14__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20059), .ZN(n15941) );
  INV_X1 U19024 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20781) );
  NAND3_X1 U19025 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15936), .A3(n15952), 
        .ZN(n15938) );
  AOI21_X1 U19026 ( .B1(n20781), .B2(n15938), .A(n15937), .ZN(n15939) );
  AOI21_X1 U19027 ( .B1(n16001), .B2(n20031), .A(n15939), .ZN(n15940) );
  NAND4_X1 U19028 ( .A1(n15942), .A2(n15941), .A3(n15940), .A4(n20042), .ZN(
        P1_U2826) );
  AOI22_X1 U19029 ( .A1(n16005), .A2(n20040), .B1(n20027), .B2(n15943), .ZN(
        n15949) );
  AOI22_X1 U19030 ( .A1(n20046), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20059), .ZN(n15948) );
  INV_X1 U19031 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20779) );
  OAI21_X1 U19032 ( .B1(n16103), .B2(n15944), .A(n20779), .ZN(n15945) );
  AOI22_X1 U19033 ( .A1(n20031), .A2(n16004), .B1(n15946), .B2(n15945), .ZN(
        n15947) );
  NAND4_X1 U19034 ( .A1(n15949), .A2(n15948), .A3(n15947), .A4(n20042), .ZN(
        P1_U2828) );
  NAND2_X1 U19035 ( .A1(n15951), .A2(n15950), .ZN(n15964) );
  OAI22_X1 U19036 ( .A1(n16017), .A2(n20054), .B1(n20062), .B2(n16104), .ZN(
        n15956) );
  INV_X1 U19037 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15954) );
  AOI22_X1 U19038 ( .A1(n15952), .A2(n16103), .B1(n20046), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15953) );
  OAI211_X1 U19039 ( .C1(n20044), .C2(n15954), .A(n15953), .B(n20042), .ZN(
        n15955) );
  AOI211_X1 U19040 ( .C1(n20031), .C2(n16014), .A(n15956), .B(n15955), .ZN(
        n15957) );
  OAI21_X1 U19041 ( .B1(n16103), .B2(n15964), .A(n15957), .ZN(P1_U2829) );
  OAI22_X1 U19042 ( .A1(n14504), .A2(n20044), .B1(n20062), .B2(n16116), .ZN(
        n15958) );
  AOI211_X1 U19043 ( .C1(n20040), .C2(n15959), .A(n20135), .B(n15958), .ZN(
        n15968) );
  INV_X1 U19044 ( .A(n15960), .ZN(n15966) );
  NOR3_X1 U19045 ( .A1(n20021), .A2(P1_REIP_REG_10__SCAN_IN), .A3(n15961), 
        .ZN(n15962) );
  AOI21_X1 U19046 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(n20046), .A(n15962), .ZN(
        n15963) );
  OAI21_X1 U19047 ( .B1(n15964), .B2(n20775), .A(n15963), .ZN(n15965) );
  AOI21_X1 U19048 ( .B1(n15966), .B2(n20031), .A(n15965), .ZN(n15967) );
  NAND2_X1 U19049 ( .A1(n15968), .A2(n15967), .ZN(P1_U2830) );
  INV_X1 U19050 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20908) );
  AOI22_X1 U19051 ( .A1(n16001), .A2(n15970), .B1(n15969), .B2(n20109), .ZN(
        n15971) );
  OAI21_X1 U19052 ( .B1(n15972), .B2(n20908), .A(n15971), .ZN(P1_U2890) );
  AOI22_X1 U19053 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15976) );
  AOI22_X1 U19054 ( .A1(n15974), .A2(n20158), .B1(n20134), .B2(n15973), .ZN(
        n15975) );
  OAI211_X1 U19055 ( .C1(n16029), .C2(n15977), .A(n15976), .B(n15975), .ZN(
        P1_U2977) );
  AOI21_X1 U19056 ( .B1(n16033), .B2(n15981), .A(n15980), .ZN(n15983) );
  OAI211_X1 U19057 ( .C1(n15984), .C2(n16037), .A(n15983), .B(n15982), .ZN(
        P1_U2978) );
  AOI22_X1 U19058 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15992) );
  OAI21_X1 U19059 ( .B1(n15987), .B2(n15986), .A(n15985), .ZN(n15989) );
  XNOR2_X1 U19060 ( .A(n15989), .B(n15988), .ZN(n16070) );
  AOI22_X1 U19061 ( .A1(n16070), .A2(n20134), .B1(n15990), .B2(n20158), .ZN(
        n15991) );
  OAI211_X1 U19062 ( .C1(n16029), .C2(n15993), .A(n15992), .B(n15991), .ZN(
        P1_U2983) );
  INV_X1 U19063 ( .A(n15994), .ZN(n15996) );
  OAI21_X1 U19064 ( .B1(n15997), .B2(n15996), .A(n15995), .ZN(n15999) );
  XNOR2_X1 U19065 ( .A(n16009), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15998) );
  XNOR2_X1 U19066 ( .A(n15999), .B(n15998), .ZN(n16088) );
  AOI22_X1 U19067 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16003) );
  AOI22_X1 U19068 ( .A1(n16001), .A2(n20158), .B1(n16000), .B2(n16033), .ZN(
        n16002) );
  OAI211_X1 U19069 ( .C1(n16088), .C2(n19981), .A(n16003), .B(n16002), .ZN(
        P1_U2985) );
  AOI22_X1 U19070 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16007) );
  AOI22_X1 U19071 ( .A1(n16033), .A2(n16005), .B1(n20158), .B2(n16004), .ZN(
        n16006) );
  OAI211_X1 U19072 ( .C1(n16008), .C2(n19981), .A(n16007), .B(n16006), .ZN(
        P1_U2987) );
  AOI22_X1 U19073 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16016) );
  NAND3_X1 U19074 ( .A1(n16010), .A2(n16009), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16012) );
  NAND2_X1 U19075 ( .A1(n16012), .A2(n16011), .ZN(n16013) );
  XOR2_X1 U19076 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16013), .Z(
        n16106) );
  AOI22_X1 U19077 ( .A1(n20134), .A2(n16106), .B1(n20158), .B2(n16014), .ZN(
        n16015) );
  OAI211_X1 U19078 ( .C1(n16029), .C2(n16017), .A(n16016), .B(n16015), .ZN(
        P1_U2988) );
  AOI22_X1 U19079 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16022) );
  XNOR2_X1 U19080 ( .A(n16018), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16019) );
  XNOR2_X1 U19081 ( .A(n16020), .B(n16019), .ZN(n16143) );
  AOI22_X1 U19082 ( .A1(n16143), .A2(n20134), .B1(n20158), .B2(n20022), .ZN(
        n16021) );
  OAI211_X1 U19083 ( .C1(n16029), .C2(n20010), .A(n16022), .B(n16021), .ZN(
        P1_U2992) );
  AOI22_X1 U19084 ( .A1(n20132), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20135), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16028) );
  NAND2_X1 U19085 ( .A1(n16024), .A2(n16023), .ZN(n16025) );
  XNOR2_X1 U19086 ( .A(n16026), .B(n16025), .ZN(n16149) );
  AOI22_X1 U19087 ( .A1(n16149), .A2(n20134), .B1(n20158), .B2(n20032), .ZN(
        n16027) );
  OAI211_X1 U19088 ( .C1(n16029), .C2(n20025), .A(n16028), .B(n16027), .ZN(
        P1_U2993) );
  XNOR2_X1 U19089 ( .A(n16031), .B(n16030), .ZN(n16161) );
  INV_X1 U19090 ( .A(n16161), .ZN(n16034) );
  INV_X1 U19091 ( .A(n16032), .ZN(n20051) );
  AOI222_X1 U19092 ( .A1(n16034), .A2(n20134), .B1(n20158), .B2(n20051), .C1(
        n20039), .C2(n16033), .ZN(n16036) );
  INV_X1 U19093 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20053) );
  NOR2_X1 U19094 ( .A1(n20042), .A2(n20053), .ZN(n16157) );
  INV_X1 U19095 ( .A(n16157), .ZN(n16035) );
  OAI211_X1 U19096 ( .C1(n20043), .C2(n16037), .A(n16036), .B(n16035), .ZN(
        P1_U2994) );
  INV_X1 U19097 ( .A(n16038), .ZN(n16039) );
  OAI22_X1 U19098 ( .A1(n16039), .A2(n16135), .B1(n16042), .B2(n16054), .ZN(
        n16040) );
  AOI21_X1 U19099 ( .B1(n20140), .B2(n16041), .A(n16040), .ZN(n16044) );
  NAND3_X1 U19100 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n16046), .A3(
        n16042), .ZN(n16043) );
  OAI211_X1 U19101 ( .C1(n16045), .C2(n20042), .A(n16044), .B(n16043), .ZN(
        P1_U3005) );
  AOI22_X1 U19102 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n20135), .B1(n16046), 
        .B2(n16053), .ZN(n16052) );
  INV_X1 U19103 ( .A(n16048), .ZN(n16049) );
  AOI22_X1 U19104 ( .A1(n16050), .A2(n20140), .B1(n20145), .B2(n16049), .ZN(
        n16051) );
  OAI211_X1 U19105 ( .C1(n16054), .C2(n16053), .A(n16052), .B(n16051), .ZN(
        P1_U3006) );
  OAI22_X1 U19106 ( .A1(n16056), .A2(n16160), .B1(n16135), .B2(n16055), .ZN(
        n16057) );
  AOI21_X1 U19107 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16058), .A(
        n16057), .ZN(n16062) );
  NAND3_X1 U19108 ( .A1(n16060), .A2(n16059), .A3(n16082), .ZN(n16061) );
  OAI211_X1 U19109 ( .C1(n16063), .C2(n20042), .A(n16062), .B(n16061), .ZN(
        P1_U3013) );
  OAI21_X1 U19110 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16064), .A(
        n16093), .ZN(n16065) );
  INV_X1 U19111 ( .A(n16065), .ZN(n16078) );
  NAND2_X1 U19112 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16082), .ZN(
        n16080) );
  AOI221_X1 U19113 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n16079), .C2(n16072), .A(
        n16080), .ZN(n16069) );
  INV_X1 U19114 ( .A(n16066), .ZN(n16067) );
  OAI22_X1 U19115 ( .A1(n16067), .A2(n16135), .B1(n20963), .B2(n20042), .ZN(
        n16068) );
  AOI211_X1 U19116 ( .C1(n20140), .C2(n16070), .A(n16069), .B(n16068), .ZN(
        n16071) );
  OAI21_X1 U19117 ( .B1(n16078), .B2(n16072), .A(n16071), .ZN(P1_U3015) );
  OAI22_X1 U19118 ( .A1(n16074), .A2(n16135), .B1(n16073), .B2(n20042), .ZN(
        n16075) );
  AOI21_X1 U19119 ( .B1(n20140), .B2(n16076), .A(n16075), .ZN(n16077) );
  OAI221_X1 U19120 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16080), 
        .C1(n16079), .C2(n16078), .A(n16077), .ZN(P1_U3016) );
  INV_X1 U19121 ( .A(n16093), .ZN(n16081) );
  MUX2_X1 U19122 ( .A(n16082), .B(n16081), .S(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16086) );
  NAND2_X1 U19123 ( .A1(n16083), .A2(n20145), .ZN(n16084) );
  OAI21_X1 U19124 ( .B1(n20781), .B2(n20042), .A(n16084), .ZN(n16085) );
  NOR2_X1 U19125 ( .A1(n16086), .A2(n16085), .ZN(n16087) );
  OAI21_X1 U19126 ( .B1(n16088), .B2(n16160), .A(n16087), .ZN(P1_U3017) );
  OR2_X1 U19127 ( .A1(n16090), .A2(n16089), .ZN(n16100) );
  AOI21_X1 U19128 ( .B1(n16092), .B2(n20145), .A(n16091), .ZN(n16099) );
  AOI21_X1 U19129 ( .B1(n16095), .B2(n16094), .A(n16093), .ZN(n16096) );
  AOI21_X1 U19130 ( .B1(n16097), .B2(n20140), .A(n16096), .ZN(n16098) );
  OAI211_X1 U19131 ( .C1(n16101), .C2(n16100), .A(n16099), .B(n16098), .ZN(
        P1_U3018) );
  INV_X1 U19132 ( .A(n16102), .ZN(n16110) );
  INV_X1 U19133 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16103) );
  OAI22_X1 U19134 ( .A1(n16104), .A2(n16135), .B1(n20042), .B2(n16103), .ZN(
        n16105) );
  INV_X1 U19135 ( .A(n16105), .ZN(n16109) );
  AOI22_X1 U19136 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16107), .B1(
        n20140), .B2(n16106), .ZN(n16108) );
  OAI211_X1 U19137 ( .C1(n16153), .C2(n16110), .A(n16109), .B(n16108), .ZN(
        P1_U3020) );
  OAI21_X1 U19138 ( .B1(n16113), .B2(n16112), .A(n16111), .ZN(n16115) );
  INV_X1 U19139 ( .A(n16114), .ZN(n16129) );
  AOI21_X1 U19140 ( .B1(n16133), .B2(n16115), .A(n16129), .ZN(n16127) );
  OAI22_X1 U19141 ( .A1(n16135), .A2(n16116), .B1(n20775), .B2(n20042), .ZN(
        n16117) );
  AOI21_X1 U19142 ( .B1(n20140), .B2(n16118), .A(n16117), .ZN(n16120) );
  NOR3_X1 U19143 ( .A1(n16138), .A2(n16139), .A3(n16153), .ZN(n16123) );
  OAI221_X1 U19144 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14500), .C2(n16126), .A(
        n16123), .ZN(n16119) );
  OAI211_X1 U19145 ( .C1(n16127), .C2(n14500), .A(n16120), .B(n16119), .ZN(
        P1_U3021) );
  AOI21_X1 U19146 ( .B1(n19999), .B2(n20145), .A(n16121), .ZN(n16125) );
  AOI22_X1 U19147 ( .A1(n16123), .A2(n16126), .B1(n16122), .B2(n20140), .ZN(
        n16124) );
  OAI211_X1 U19148 ( .C1(n16127), .C2(n16126), .A(n16125), .B(n16124), .ZN(
        P1_U3022) );
  NAND2_X1 U19149 ( .A1(n16128), .A2(n11474), .ZN(n16154) );
  AOI21_X1 U19150 ( .B1(n16131), .B2(n16130), .A(n16129), .ZN(n16164) );
  OAI21_X1 U19151 ( .B1(n16132), .B2(n16154), .A(n16164), .ZN(n16150) );
  AOI21_X1 U19152 ( .B1(n16138), .B2(n16133), .A(n16150), .ZN(n16148) );
  INV_X1 U19153 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16142) );
  OAI222_X1 U19154 ( .A1(n16136), .A2(n16135), .B1(n20042), .B2(n20773), .C1(
        n16160), .C2(n16134), .ZN(n16137) );
  INV_X1 U19155 ( .A(n16137), .ZN(n16141) );
  NOR2_X1 U19156 ( .A1(n16138), .A2(n16153), .ZN(n16144) );
  OAI211_X1 U19157 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16144), .B(n16139), .ZN(n16140) );
  OAI211_X1 U19158 ( .C1(n16148), .C2(n16142), .A(n16141), .B(n16140), .ZN(
        P1_U3023) );
  INV_X1 U19159 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16147) );
  AOI22_X1 U19160 ( .A1(n20145), .A2(n20016), .B1(n20135), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16146) );
  AOI22_X1 U19161 ( .A1(n16144), .A2(n16147), .B1(n20140), .B2(n16143), .ZN(
        n16145) );
  OAI211_X1 U19162 ( .C1(n16148), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        P1_U3024) );
  AOI22_X1 U19163 ( .A1(n20145), .A2(n20026), .B1(n20135), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16152) );
  AOI22_X1 U19164 ( .A1(n16150), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20140), .B2(n16149), .ZN(n16151) );
  OAI211_X1 U19165 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16153), .A(
        n16152), .B(n16151), .ZN(P1_U3025) );
  INV_X1 U19166 ( .A(n16154), .ZN(n16155) );
  NAND2_X1 U19167 ( .A1(n16156), .A2(n16155), .ZN(n16159) );
  AOI21_X1 U19168 ( .B1(n20145), .B2(n20037), .A(n16157), .ZN(n16158) );
  OAI211_X1 U19169 ( .C1(n16161), .C2(n16160), .A(n16159), .B(n16158), .ZN(
        n16162) );
  INV_X1 U19170 ( .A(n16162), .ZN(n16163) );
  OAI21_X1 U19171 ( .B1(n16164), .B2(n11474), .A(n16163), .ZN(P1_U3026) );
  INV_X1 U19172 ( .A(n16165), .ZN(n16170) );
  NAND3_X1 U19173 ( .A1(n16167), .A2(n19975), .A3(n16166), .ZN(n16168) );
  OAI21_X1 U19174 ( .B1(n16170), .B2(n16169), .A(n16168), .ZN(P1_U3468) );
  NAND4_X1 U19175 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20260), .A4(n20848), .ZN(n16171) );
  NAND2_X1 U19176 ( .A1(n16172), .A2(n16171), .ZN(n20744) );
  NAND2_X1 U19177 ( .A1(n16173), .A2(n20260), .ZN(n16176) );
  OAI21_X1 U19178 ( .B1(n16180), .B2(n9880), .A(n11284), .ZN(n16175) );
  OAI211_X1 U19179 ( .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n16176), .A(n16175), 
        .B(n16174), .ZN(n16177) );
  AOI221_X1 U19180 ( .B1(n16179), .B2(n16178), .C1(n20744), .C2(n16178), .A(
        n16177), .ZN(P1_U3162) );
  INV_X1 U19181 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20568) );
  NOR2_X1 U19182 ( .A1(n16180), .A2(n9880), .ZN(n16182) );
  OAI22_X1 U19183 ( .A1(n20568), .A2(n16182), .B1(n16181), .B2(n9880), .ZN(
        P1_U3466) );
  NOR2_X1 U19184 ( .A1(n19108), .A2(n16183), .ZN(n16185) );
  XOR2_X1 U19185 ( .A(n16185), .B(n16184), .Z(n16194) );
  AOI22_X1 U19186 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19130), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19122), .ZN(n16186) );
  OAI21_X1 U19187 ( .B1(n16187), .B2(n19090), .A(n16186), .ZN(n16188) );
  AOI21_X1 U19188 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19117), .A(n16188), .ZN(
        n16193) );
  OAI22_X1 U19189 ( .A1(n16190), .A2(n19105), .B1(n16189), .B2(n19100), .ZN(
        n16191) );
  INV_X1 U19190 ( .A(n16191), .ZN(n16192) );
  OAI211_X1 U19191 ( .C1(n19841), .C2(n16194), .A(n16193), .B(n16192), .ZN(
        P2_U2825) );
  OAI21_X1 U19192 ( .B1(n16196), .B2(n16195), .A(n19080), .ZN(n16204) );
  AOI22_X1 U19193 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19130), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19122), .ZN(n16197) );
  OAI21_X1 U19194 ( .B1(n16198), .B2(n19090), .A(n16197), .ZN(n16199) );
  AOI21_X1 U19195 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19117), .A(n16199), .ZN(
        n16203) );
  AOI22_X1 U19196 ( .A1(n16201), .A2(n19119), .B1(n16200), .B2(n19121), .ZN(
        n16202) );
  OAI211_X1 U19197 ( .C1(n16205), .C2(n16204), .A(n16203), .B(n16202), .ZN(
        P2_U2827) );
  NAND2_X1 U19198 ( .A1(n16220), .A2(n12939), .ZN(n16206) );
  XOR2_X1 U19199 ( .A(n16207), .B(n16206), .Z(n16216) );
  AOI22_X1 U19200 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19130), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19122), .ZN(n16208) );
  OAI21_X1 U19201 ( .B1(n16209), .B2(n19090), .A(n16208), .ZN(n16210) );
  AOI21_X1 U19202 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19117), .A(n16210), .ZN(
        n16215) );
  INV_X1 U19203 ( .A(n16211), .ZN(n16212) );
  AOI22_X1 U19204 ( .A1(n16213), .A2(n19119), .B1(n16212), .B2(n19121), .ZN(
        n16214) );
  OAI211_X1 U19205 ( .C1(n19841), .C2(n16216), .A(n16215), .B(n16214), .ZN(
        P2_U2828) );
  AOI22_X1 U19206 ( .A1(n16217), .A2(n19125), .B1(P2_REIP_REG_26__SCAN_IN), 
        .B2(n19122), .ZN(n16226) );
  AOI22_X1 U19207 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19130), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19117), .ZN(n16225) );
  AOI22_X1 U19208 ( .A1(n16219), .A2(n19119), .B1(n16218), .B2(n19121), .ZN(
        n16224) );
  OAI211_X1 U19209 ( .C1(n16222), .C2(n16221), .A(n19080), .B(n16220), .ZN(
        n16223) );
  NAND4_X1 U19210 ( .A1(n16226), .A2(n16225), .A3(n16224), .A4(n16223), .ZN(
        P2_U2829) );
  OAI22_X1 U19211 ( .A1(n16228), .A2(n19090), .B1(n19024), .B2(n16227), .ZN(
        n16229) );
  INV_X1 U19212 ( .A(n16229), .ZN(n16239) );
  AOI22_X1 U19213 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19117), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19122), .ZN(n16238) );
  INV_X1 U19214 ( .A(n16230), .ZN(n16231) );
  AOI22_X1 U19215 ( .A1(n16232), .A2(n19119), .B1(n16231), .B2(n19121), .ZN(
        n16237) );
  OAI211_X1 U19216 ( .C1(n16235), .C2(n16234), .A(n19080), .B(n16233), .ZN(
        n16236) );
  NAND4_X1 U19217 ( .A1(n16239), .A2(n16238), .A3(n16237), .A4(n16236), .ZN(
        P2_U2830) );
  INV_X1 U19218 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n20973) );
  OAI22_X1 U19219 ( .A1(n19101), .A2(n20973), .B1(n19901), .B2(n19059), .ZN(
        n16242) );
  INV_X1 U19220 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16240) );
  NOR2_X1 U19221 ( .A1(n19024), .A2(n16240), .ZN(n16241) );
  AOI211_X1 U19222 ( .C1(n16243), .C2(n19119), .A(n16242), .B(n16241), .ZN(
        n16244) );
  OAI21_X1 U19223 ( .B1(n16245), .B2(n19090), .A(n16244), .ZN(n16246) );
  INV_X1 U19224 ( .A(n16246), .ZN(n16251) );
  OAI211_X1 U19225 ( .C1(n16249), .C2(n16248), .A(n19080), .B(n16247), .ZN(
        n16250) );
  OAI211_X1 U19226 ( .C1(n19100), .C2(n16252), .A(n16251), .B(n16250), .ZN(
        P2_U2831) );
  INV_X1 U19227 ( .A(n16253), .ZN(n16254) );
  AOI22_X1 U19228 ( .A1(n16254), .A2(n19125), .B1(P2_REIP_REG_23__SCAN_IN), 
        .B2(n19122), .ZN(n16263) );
  AOI22_X1 U19229 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19117), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19130), .ZN(n16262) );
  OAI22_X1 U19230 ( .A1(n16255), .A2(n19105), .B1(n19100), .B2(n16266), .ZN(
        n16256) );
  INV_X1 U19231 ( .A(n16256), .ZN(n16261) );
  OAI211_X1 U19232 ( .C1(n16259), .C2(n16258), .A(n19080), .B(n16257), .ZN(
        n16260) );
  NAND4_X1 U19233 ( .A1(n16263), .A2(n16262), .A3(n16261), .A4(n16260), .ZN(
        P2_U2832) );
  AOI22_X1 U19234 ( .A1(n16265), .A2(n16264), .B1(n19172), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16272) );
  AOI22_X1 U19235 ( .A1(n19134), .A2(BUF2_REG_23__SCAN_IN), .B1(n19135), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16271) );
  OAI22_X1 U19236 ( .A1(n16268), .A2(n19168), .B1(n16267), .B2(n16266), .ZN(
        n16269) );
  INV_X1 U19237 ( .A(n16269), .ZN(n16270) );
  NAND3_X1 U19238 ( .A1(n16272), .A2(n16271), .A3(n16270), .ZN(P2_U2896) );
  AOI22_X1 U19239 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19103), .B1(n16327), 
        .B2(n19021), .ZN(n16278) );
  INV_X1 U19240 ( .A(n16273), .ZN(n16276) );
  AOI222_X1 U19241 ( .A1(n16276), .A2(n16335), .B1(n19263), .B2(n16275), .C1(
        n9733), .C2(n16274), .ZN(n16277) );
  OAI211_X1 U19242 ( .C1(n19025), .C2(n16338), .A(n16278), .B(n16277), .ZN(
        P2_U2999) );
  AOI22_X1 U19243 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19103), .B1(n16327), 
        .B2(n16279), .ZN(n16290) );
  INV_X1 U19244 ( .A(n16280), .ZN(n16281) );
  NOR2_X1 U19245 ( .A1(n16282), .A2(n16281), .ZN(n16283) );
  XNOR2_X1 U19246 ( .A(n16284), .B(n16283), .ZN(n16358) );
  OAI21_X1 U19247 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16286), .A(
        n16285), .ZN(n16356) );
  OAI22_X1 U19248 ( .A1(n16287), .A2(n16355), .B1(n19257), .B2(n16356), .ZN(
        n16288) );
  AOI21_X1 U19249 ( .B1(n16358), .B2(n16335), .A(n16288), .ZN(n16289) );
  OAI211_X1 U19250 ( .C1(n16291), .C2(n16338), .A(n16290), .B(n16289), .ZN(
        P2_U3001) );
  AOI22_X1 U19251 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19103), .B1(n16327), 
        .B2(n16292), .ZN(n16307) );
  INV_X1 U19252 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16293) );
  NAND2_X1 U19253 ( .A1(n16294), .A2(n16293), .ZN(n16296) );
  NAND2_X1 U19254 ( .A1(n16296), .A2(n16295), .ZN(n16365) );
  NAND2_X1 U19255 ( .A1(n19263), .A2(n16297), .ZN(n16304) );
  NAND2_X1 U19256 ( .A1(n16299), .A2(n16298), .ZN(n16302) );
  OR2_X1 U19257 ( .A1(n16300), .A2(n9833), .ZN(n16301) );
  XNOR2_X1 U19258 ( .A(n16302), .B(n16301), .ZN(n16367) );
  NAND2_X1 U19259 ( .A1(n16367), .A2(n16335), .ZN(n16303) );
  OAI211_X1 U19260 ( .C1(n16365), .C2(n19257), .A(n16304), .B(n16303), .ZN(
        n16305) );
  INV_X1 U19261 ( .A(n16305), .ZN(n16306) );
  OAI211_X1 U19262 ( .C1(n16308), .C2(n16338), .A(n16307), .B(n16306), .ZN(
        P2_U3003) );
  AOI22_X1 U19263 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19103), .B1(n16327), 
        .B2(n16309), .ZN(n16314) );
  AOI222_X1 U19264 ( .A1(n16312), .A2(n9733), .B1(n16335), .B2(n16311), .C1(
        n19263), .C2(n16310), .ZN(n16313) );
  OAI211_X1 U19265 ( .C1(n16315), .C2(n16338), .A(n16314), .B(n16313), .ZN(
        P2_U3005) );
  AOI22_X1 U19266 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19255), .B1(n16327), 
        .B2(n16316), .ZN(n16324) );
  NAND2_X1 U19267 ( .A1(n16317), .A2(n9733), .ZN(n16320) );
  NAND2_X1 U19268 ( .A1(n19263), .A2(n16318), .ZN(n16319) );
  OAI211_X1 U19269 ( .C1(n16321), .C2(n19259), .A(n16320), .B(n16319), .ZN(
        n16322) );
  INV_X1 U19270 ( .A(n16322), .ZN(n16323) );
  OAI211_X1 U19271 ( .C1(n16325), .C2(n16338), .A(n16324), .B(n16323), .ZN(
        P2_U3007) );
  AOI22_X1 U19272 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19255), .B1(n16327), 
        .B2(n16326), .ZN(n16337) );
  NAND2_X1 U19273 ( .A1(n16329), .A2(n16328), .ZN(n16331) );
  XNOR2_X1 U19274 ( .A(n16331), .B(n16330), .ZN(n16401) );
  INV_X1 U19275 ( .A(n16332), .ZN(n16399) );
  XOR2_X1 U19276 ( .A(n16333), .B(n16334), .Z(n16398) );
  AOI222_X1 U19277 ( .A1(n16401), .A2(n9733), .B1(n19263), .B2(n16399), .C1(
        n16335), .C2(n16398), .ZN(n16336) );
  OAI211_X1 U19278 ( .C1(n16339), .C2(n16338), .A(n16337), .B(n16336), .ZN(
        P2_U3009) );
  NOR2_X1 U19279 ( .A1(n16340), .A2(n16351), .ZN(n16345) );
  INV_X1 U19280 ( .A(n16340), .ZN(n16342) );
  OAI21_X1 U19281 ( .B1(n16351), .B2(n16342), .A(n16341), .ZN(n16354) );
  OAI22_X1 U19282 ( .A1(n16413), .A2(n19045), .B1(n12408), .B2(n19058), .ZN(
        n16343) );
  AOI221_X1 U19283 ( .B1(n16345), .B2(n16344), .C1(n16354), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n16343), .ZN(n16348) );
  AOI22_X1 U19284 ( .A1(n16346), .A2(n16400), .B1(n16417), .B2(n19041), .ZN(
        n16347) );
  OAI211_X1 U19285 ( .C1(n16349), .C2(n16393), .A(n16348), .B(n16347), .ZN(
        P2_U3032) );
  INV_X1 U19286 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19886) );
  INV_X1 U19287 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16350) );
  OAI21_X1 U19288 ( .B1(n12041), .B2(n16351), .A(n16350), .ZN(n16353) );
  AOI22_X1 U19289 ( .A1(n16354), .A2(n16353), .B1(n16396), .B2(n16352), .ZN(
        n16360) );
  OAI22_X1 U19290 ( .A1(n16420), .A2(n16356), .B1(n16355), .B2(n16388), .ZN(
        n16357) );
  AOI21_X1 U19291 ( .B1(n16423), .B2(n16358), .A(n16357), .ZN(n16359) );
  OAI211_X1 U19292 ( .C1(n19886), .C2(n19058), .A(n16360), .B(n16359), .ZN(
        P2_U3033) );
  NOR2_X1 U19293 ( .A1(n16362), .A2(n16361), .ZN(n16377) );
  AOI22_X1 U19294 ( .A1(n16377), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16396), .B2(n16363), .ZN(n16374) );
  OAI22_X1 U19295 ( .A1(n16365), .A2(n16420), .B1(n16388), .B2(n16364), .ZN(
        n16366) );
  AOI21_X1 U19296 ( .B1(n16423), .B2(n16367), .A(n16366), .ZN(n16373) );
  NAND2_X1 U19297 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19103), .ZN(n16372) );
  NOR2_X1 U19298 ( .A1(n16369), .A2(n16368), .ZN(n16376) );
  OAI211_X1 U19299 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16376), .B(n16370), .ZN(
        n16371) );
  NAND4_X1 U19300 ( .A1(n16374), .A2(n16373), .A3(n16372), .A4(n16371), .ZN(
        P2_U3035) );
  OAI22_X1 U19301 ( .A1(n16413), .A2(n19071), .B1(n19880), .B2(n19058), .ZN(
        n16375) );
  AOI221_X1 U19302 ( .B1(n16377), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n16376), .C2(n12030), .A(n16375), .ZN(n16381) );
  NOR2_X1 U19303 ( .A1(n16388), .A2(n19066), .ZN(n16378) );
  AOI21_X1 U19304 ( .B1(n16379), .B2(n16400), .A(n16378), .ZN(n16380) );
  OAI211_X1 U19305 ( .C1(n16382), .C2(n16393), .A(n16381), .B(n16380), .ZN(
        P2_U3036) );
  AOI211_X1 U19306 ( .C1(n12018), .C2(n20961), .A(n16384), .B(n16383), .ZN(
        n16387) );
  OAI22_X1 U19307 ( .A1(n16385), .A2(n20961), .B1(n16413), .B2(n19084), .ZN(
        n16386) );
  AOI211_X1 U19308 ( .C1(n19103), .C2(P2_REIP_REG_8__SCAN_IN), .A(n16387), .B(
        n16386), .ZN(n16392) );
  OAI22_X1 U19309 ( .A1(n16389), .A2(n16420), .B1(n16388), .B2(n19078), .ZN(
        n16390) );
  INV_X1 U19310 ( .A(n16390), .ZN(n16391) );
  OAI211_X1 U19311 ( .C1(n16394), .C2(n16393), .A(n16392), .B(n16391), .ZN(
        P2_U3038) );
  INV_X1 U19312 ( .A(n16395), .ZN(n19146) );
  AOI22_X1 U19313 ( .A1(n16397), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n16396), .B2(n19146), .ZN(n16410) );
  AOI222_X1 U19314 ( .A1(n16401), .A2(n16400), .B1(n16417), .B2(n16399), .C1(
        n16423), .C2(n16398), .ZN(n16409) );
  NAND2_X1 U19315 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19103), .ZN(n16408) );
  AOI211_X1 U19316 ( .C1(n16405), .C2(n16404), .A(n16403), .B(n16402), .ZN(
        n16406) );
  INV_X1 U19317 ( .A(n16406), .ZN(n16407) );
  NAND4_X1 U19318 ( .A1(n16410), .A2(n16409), .A3(n16408), .A4(n16407), .ZN(
        P2_U3041) );
  INV_X1 U19319 ( .A(n16411), .ZN(n16416) );
  OAI22_X1 U19320 ( .A1(n16413), .A2(n16412), .B1(n19872), .B2(n19058), .ZN(
        n16414) );
  AOI21_X1 U19321 ( .B1(n16416), .B2(n16415), .A(n16414), .ZN(n16419) );
  NAND2_X1 U19322 ( .A1(n16417), .A2(n13120), .ZN(n16418) );
  OAI211_X1 U19323 ( .C1(n16421), .C2(n16420), .A(n16419), .B(n16418), .ZN(
        n16422) );
  AOI21_X1 U19324 ( .B1(n16424), .B2(n16423), .A(n16422), .ZN(n16425) );
  OAI21_X1 U19325 ( .B1(n16426), .B2(n12264), .A(n16425), .ZN(P2_U3043) );
  INV_X1 U19326 ( .A(n16428), .ZN(n16430) );
  OAI211_X1 U19327 ( .C1(n16428), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16427), .ZN(n16429) );
  INV_X1 U19328 ( .A(n16458), .ZN(n16433) );
  OAI211_X1 U19329 ( .C1(n16430), .C2(n19949), .A(n16429), .B(n16433), .ZN(
        n16431) );
  AOI21_X1 U19330 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16434), .A(
        n16431), .ZN(n16438) );
  MUX2_X1 U19331 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16432), .S(
        n16433), .Z(n16440) );
  MUX2_X1 U19332 ( .A(n16435), .B(n16434), .S(n16433), .Z(n16460) );
  NOR2_X1 U19333 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16460), .ZN(
        n16436) );
  OR3_X1 U19334 ( .A1(n16438), .A2(n16440), .A3(n16436), .ZN(n16437) );
  AOI22_X1 U19335 ( .A1(n16438), .A2(n16440), .B1(n19933), .B2(n16437), .ZN(
        n16439) );
  NOR2_X1 U19336 ( .A1(n16439), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n16463) );
  INV_X1 U19337 ( .A(n16440), .ZN(n16461) );
  INV_X1 U19338 ( .A(n16441), .ZN(n16448) );
  NAND2_X1 U19339 ( .A1(n16449), .A2(n16442), .ZN(n16447) );
  INV_X1 U19340 ( .A(n16443), .ZN(n16444) );
  NAND2_X1 U19341 ( .A1(n16445), .A2(n16444), .ZN(n16446) );
  OAI211_X1 U19342 ( .C1(n16449), .C2(n16448), .A(n16447), .B(n16446), .ZN(
        n19960) );
  OAI21_X1 U19343 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16450), .ZN(n16455) );
  INV_X1 U19344 ( .A(n16451), .ZN(n16453) );
  NAND3_X1 U19345 ( .A1(n16453), .A2(n11776), .A3(n16452), .ZN(n16454) );
  OAI211_X1 U19346 ( .C1(n11750), .C2(n16456), .A(n16455), .B(n16454), .ZN(
        n16457) );
  AOI211_X1 U19347 ( .C1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n16458), .A(
        n19960), .B(n16457), .ZN(n16459) );
  OAI21_X1 U19348 ( .B1(n16461), .B2(n16460), .A(n16459), .ZN(n16462) );
  NOR2_X1 U19349 ( .A1(n16463), .A2(n16462), .ZN(n16480) );
  AOI211_X1 U19350 ( .C1(n16481), .C2(n16466), .A(n16465), .B(n16464), .ZN(
        n16478) );
  NAND3_X1 U19351 ( .A1(n16480), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n16467), 
        .ZN(n16472) );
  NOR3_X1 U19352 ( .A1(n12175), .A2(n16469), .A3(n16468), .ZN(n16470) );
  OAI21_X1 U19353 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16474), .A(n16473), 
        .ZN(n16476) );
  NAND2_X1 U19354 ( .A1(n19843), .A2(n19857), .ZN(n16475) );
  AOI22_X1 U19355 ( .A1(n19843), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16476), 
        .B2(n16475), .ZN(n16477) );
  OAI211_X1 U19356 ( .C1(n16480), .C2(n16479), .A(n16478), .B(n16477), .ZN(
        P2_U3176) );
  AOI221_X1 U19357 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n21158), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19843), .A(n16481), .ZN(n16482) );
  INV_X1 U19358 ( .A(n16482), .ZN(P2_U3593) );
  INV_X1 U19359 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18890) );
  NAND3_X1 U19360 ( .A1(n17946), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16497), .ZN(n16483) );
  XNOR2_X1 U19361 ( .A(n18890), .B(n16483), .ZN(n16544) );
  INV_X1 U19362 ( .A(n18756), .ZN(n16484) );
  INV_X1 U19363 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16689) );
  INV_X1 U19364 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20970) );
  INV_X1 U19365 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16485) );
  NAND2_X1 U19366 ( .A1(n17872), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17849) );
  NAND2_X1 U19367 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17834) );
  INV_X1 U19368 ( .A(n17834), .ZN(n17847) );
  NAND4_X1 U19369 ( .A1(n17847), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17767) );
  NAND2_X1 U19370 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16859) );
  NAND3_X1 U19371 ( .A1(n17782), .A2(n17780), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17744) );
  NAND2_X1 U19372 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17748) );
  NAND2_X1 U19373 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17735), .ZN(
        n17711) );
  NAND2_X1 U19374 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17713) );
  NAND2_X1 U19375 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17673) );
  NAND2_X1 U19376 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17634) );
  NAND3_X1 U19377 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n16680), .ZN(n16525) );
  NAND2_X1 U19378 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16524), .ZN(
        n16486) );
  INV_X1 U19379 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18867) );
  NOR2_X1 U19380 ( .A1(n18148), .A2(n18867), .ZN(n16537) );
  INV_X1 U19381 ( .A(n16487), .ZN(n17623) );
  NOR2_X1 U19382 ( .A1(n20970), .A2(n17623), .ZN(n17602) );
  NAND3_X1 U19383 ( .A1(n17602), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16521) );
  NOR2_X1 U19384 ( .A1(n16720), .A2(n16521), .ZN(n16489) );
  NAND2_X1 U19385 ( .A1(n18933), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18791) );
  AOI21_X1 U19386 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16488), .A(
        n18662), .ZN(n17712) );
  INV_X1 U19387 ( .A(n17712), .ZN(n17746) );
  NAND2_X1 U19388 ( .A1(n16489), .A2(n17746), .ZN(n16509) );
  XNOR2_X1 U19389 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16492) );
  NOR2_X1 U19390 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17694), .ZN(
        n16526) );
  INV_X1 U19391 ( .A(n16525), .ZN(n16677) );
  OAI21_X1 U19392 ( .B1(n18365), .B2(n16489), .A(n17940), .ZN(n16490) );
  INV_X1 U19393 ( .A(n16490), .ZN(n16491) );
  OAI21_X1 U19394 ( .B1(n16677), .B2(n18791), .A(n16491), .ZN(n16523) );
  NOR2_X1 U19395 ( .A1(n16526), .A2(n16523), .ZN(n16508) );
  OAI22_X1 U19396 ( .A1(n16509), .A2(n16492), .B1(n16508), .B2(n16689), .ZN(
        n16493) );
  AOI211_X1 U19397 ( .C1(n17801), .C2(n16953), .A(n16537), .B(n16493), .ZN(
        n16503) );
  AOI22_X1 U19398 ( .A1(n17856), .A2(n18890), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17792), .ZN(n16496) );
  NOR2_X1 U19399 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18890), .ZN(
        n16539) );
  INV_X1 U19400 ( .A(n17945), .ZN(n16518) );
  NAND3_X1 U19401 ( .A1(n16497), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n18890), .ZN(n16534) );
  OAI21_X1 U19402 ( .B1(n16506), .B2(n16504), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16498) );
  OAI21_X1 U19403 ( .B1(n16518), .B2(n16534), .A(n16498), .ZN(n16540) );
  INV_X1 U19404 ( .A(n16540), .ZN(n16500) );
  NOR2_X2 U19405 ( .A1(n16545), .A2(n17943), .ZN(n17777) );
  OAI211_X1 U19406 ( .C1(n16544), .C2(n17944), .A(n16503), .B(n16502), .ZN(
        P3_U2799) );
  INV_X1 U19407 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16702) );
  XNOR2_X1 U19408 ( .A(n16702), .B(n16524), .ZN(n16700) );
  NAND2_X1 U19409 ( .A1(n17777), .A2(n16504), .ZN(n16520) );
  NAND2_X1 U19410 ( .A1(n9734), .A2(n16505), .ZN(n16532) );
  AOI21_X1 U19411 ( .B1(n16520), .B2(n16532), .A(n16506), .ZN(n16511) );
  OAI221_X1 U19412 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16509), .C1(
        n16702), .C2(n16508), .A(n16507), .ZN(n16510) );
  AOI211_X1 U19413 ( .C1(n17801), .C2(n16700), .A(n16511), .B(n16510), .ZN(
        n16515) );
  INV_X1 U19414 ( .A(n17809), .ZN(n18133) );
  OAI22_X2 U19415 ( .A1(n18135), .A2(n17944), .B1(n16499), .B2(n18133), .ZN(
        n17840) );
  INV_X1 U19416 ( .A(n17755), .ZN(n17729) );
  NAND3_X1 U19417 ( .A1(n16513), .A2(n17729), .A3(n16512), .ZN(n16514) );
  OAI211_X1 U19418 ( .C1(n16516), .C2(n17844), .A(n16515), .B(n16514), .ZN(
        P3_U2800) );
  NAND2_X1 U19419 ( .A1(n17946), .A2(n16517), .ZN(n16558) );
  INV_X1 U19420 ( .A(n16517), .ZN(n16519) );
  NOR2_X1 U19421 ( .A1(n16519), .A2(n16518), .ZN(n16554) );
  INV_X1 U19422 ( .A(n16520), .ZN(n16530) );
  OAI21_X1 U19423 ( .B1(n18365), .B2(n16521), .A(n16720), .ZN(n16522) );
  AOI22_X1 U19424 ( .A1(n18255), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n16523), 
        .B2(n16522), .ZN(n16528) );
  AOI21_X1 U19425 ( .B1(n16720), .B2(n16525), .A(n16524), .ZN(n16714) );
  OAI21_X1 U19426 ( .B1(n16526), .B2(n17801), .A(n16714), .ZN(n16527) );
  OAI22_X1 U19427 ( .A1(n16535), .A2(n18890), .B1(n16534), .B2(n16533), .ZN(
        n16536) );
  AOI211_X1 U19428 ( .C1(n16539), .C2(n16538), .A(n16537), .B(n16536), .ZN(
        n16543) );
  AOI22_X1 U19429 ( .A1(n18175), .A2(n16541), .B1(n18107), .B2(n16540), .ZN(
        n16542) );
  NOR2_X1 U19430 ( .A1(n16545), .A2(n18757), .ZN(n18134) );
  INV_X1 U19431 ( .A(n18134), .ZN(n18115) );
  NOR2_X1 U19432 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18716), .ZN(
        n18243) );
  NAND2_X1 U19433 ( .A1(n18722), .A2(n18732), .ZN(n18226) );
  NOR2_X1 U19434 ( .A1(n18243), .A2(n18164), .ZN(n18228) );
  AOI22_X1 U19435 ( .A1(n18751), .A2(n18053), .B1(n18051), .B2(n18228), .ZN(
        n17967) );
  NAND2_X1 U19436 ( .A1(n18750), .A2(n18001), .ZN(n16546) );
  OAI211_X1 U19437 ( .C1(n18079), .C2(n18115), .A(n17967), .B(n16546), .ZN(
        n18009) );
  NAND2_X1 U19438 ( .A1(n18254), .A2(n18009), .ZN(n18018) );
  NOR2_X1 U19439 ( .A1(n17615), .A2(n18018), .ZN(n17955) );
  INV_X1 U19440 ( .A(n16563), .ZN(n16547) );
  NAND2_X1 U19441 ( .A1(n16547), .A2(n16552), .ZN(n17609) );
  NOR2_X1 U19442 ( .A1(n17792), .A2(n17609), .ZN(n17608) );
  NOR2_X1 U19443 ( .A1(n16563), .A2(n17608), .ZN(n17593) );
  OAI21_X1 U19444 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17856), .A(
        n16548), .ZN(n17592) );
  NOR2_X1 U19445 ( .A1(n17591), .A2(n18162), .ZN(n16562) );
  AOI22_X1 U19446 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17955), .B1(
        n16549), .B2(n16562), .ZN(n16566) );
  INV_X1 U19447 ( .A(n17591), .ZN(n16550) );
  OAI211_X1 U19448 ( .C1(n16553), .C2(n16552), .A(n16551), .B(n16550), .ZN(
        n16560) );
  OR2_X1 U19449 ( .A1(n16554), .A2(n18115), .ZN(n16556) );
  AOI21_X1 U19450 ( .B1(n16558), .B2(n18750), .A(n16557), .ZN(n16559) );
  AOI22_X1 U19451 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18255), .B1(n16563), 
        .B2(n16562), .ZN(n16564) );
  OAI221_X1 U19452 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n16566), 
        .C1(n17597), .C2(n16565), .A(n16564), .ZN(P3_U2834) );
  NOR3_X1 U19453 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16568) );
  NOR4_X1 U19454 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16567) );
  NAND4_X1 U19455 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16568), .A3(n16567), .A4(
        U215), .ZN(U213) );
  INV_X1 U19456 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16645) );
  NAND2_X1 U19457 ( .A1(n19270), .A2(n16569), .ZN(n16570) );
  NAND2_X2 U19458 ( .A1(U214), .A2(n16570), .ZN(n16614) );
  INV_X1 U19459 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16571) );
  OAI222_X1 U19460 ( .A1(U212), .A2(n16645), .B1(n16614), .B2(n20221), .C1(
        U214), .C2(n16571), .ZN(U216) );
  INV_X1 U19461 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16646) );
  INV_X1 U19462 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20213) );
  INV_X1 U19463 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n21011) );
  OAI222_X1 U19464 ( .A1(U212), .A2(n16646), .B1(n16614), .B2(n20213), .C1(
        U214), .C2(n21011), .ZN(U217) );
  INV_X1 U19465 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20206) );
  INV_X2 U19466 ( .A(U214), .ZN(n16612) );
  INV_X2 U19467 ( .A(U212), .ZN(n16611) );
  AOI22_X1 U19468 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16611), .ZN(n16572) );
  OAI21_X1 U19469 ( .B1(n20206), .B2(n16614), .A(n16572), .ZN(U218) );
  AOI22_X1 U19470 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16611), .ZN(n16573) );
  OAI21_X1 U19471 ( .B1(n14292), .B2(n16614), .A(n16573), .ZN(U219) );
  INV_X1 U19472 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20191) );
  AOI22_X1 U19473 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16611), .ZN(n16574) );
  OAI21_X1 U19474 ( .B1(n20191), .B2(n16614), .A(n16574), .ZN(U220) );
  AOI22_X1 U19475 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16611), .ZN(n16575) );
  OAI21_X1 U19476 ( .B1(n14305), .B2(n16614), .A(n16575), .ZN(U221) );
  INV_X1 U19477 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n21113) );
  INV_X1 U19478 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20176) );
  INV_X1 U19479 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n16576) );
  OAI222_X1 U19480 ( .A1(U212), .A2(n21113), .B1(n16614), .B2(n20176), .C1(
        U214), .C2(n16576), .ZN(U222) );
  INV_X1 U19481 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20160) );
  AOI22_X1 U19482 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16611), .ZN(n16577) );
  OAI21_X1 U19483 ( .B1(n20160), .B2(n16614), .A(n16577), .ZN(U223) );
  INV_X1 U19484 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U19485 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16611), .ZN(n16578) );
  OAI21_X1 U19486 ( .B1(n20218), .B2(n16614), .A(n16578), .ZN(U224) );
  INV_X1 U19487 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n21037) );
  AOI22_X1 U19488 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16611), .ZN(n16579) );
  OAI21_X1 U19489 ( .B1(n21037), .B2(n16614), .A(n16579), .ZN(U225) );
  INV_X1 U19490 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20203) );
  AOI22_X1 U19491 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16611), .ZN(n16580) );
  OAI21_X1 U19492 ( .B1(n20203), .B2(n16614), .A(n16580), .ZN(U226) );
  INV_X1 U19493 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20196) );
  AOI22_X1 U19494 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16611), .ZN(n16581) );
  OAI21_X1 U19495 ( .B1(n20196), .B2(n16614), .A(n16581), .ZN(U227) );
  INV_X1 U19496 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20189) );
  AOI22_X1 U19497 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16611), .ZN(n16582) );
  OAI21_X1 U19498 ( .B1(n20189), .B2(n16614), .A(n16582), .ZN(U228) );
  INV_X1 U19499 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20182) );
  AOI22_X1 U19500 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16611), .ZN(n16583) );
  OAI21_X1 U19501 ( .B1(n20182), .B2(n16614), .A(n16583), .ZN(U229) );
  INV_X1 U19502 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20174) );
  AOI22_X1 U19503 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16611), .ZN(n16584) );
  OAI21_X1 U19504 ( .B1(n20174), .B2(n16614), .A(n16584), .ZN(U230) );
  INV_X1 U19505 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n21025) );
  INV_X1 U19506 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20169) );
  INV_X1 U19507 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n16585) );
  OAI222_X1 U19508 ( .A1(U212), .A2(n21025), .B1(n16614), .B2(n20169), .C1(
        U214), .C2(n16585), .ZN(U231) );
  AOI22_X1 U19509 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16611), .ZN(n16586) );
  OAI21_X1 U19510 ( .B1(n13627), .B2(n16614), .A(n16586), .ZN(U232) );
  INV_X1 U19511 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16588) );
  AOI22_X1 U19512 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16611), .ZN(n16587) );
  OAI21_X1 U19513 ( .B1(n16588), .B2(n16614), .A(n16587), .ZN(U233) );
  INV_X1 U19514 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16629) );
  INV_X1 U19515 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16589) );
  INV_X1 U19516 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n21013) );
  OAI222_X1 U19517 ( .A1(U212), .A2(n16629), .B1(n16614), .B2(n16589), .C1(
        U214), .C2(n21013), .ZN(U234) );
  INV_X1 U19518 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16591) );
  AOI22_X1 U19519 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16611), .ZN(n16590) );
  OAI21_X1 U19520 ( .B1(n16591), .B2(n16614), .A(n16590), .ZN(U235) );
  INV_X1 U19521 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16593) );
  AOI22_X1 U19522 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16611), .ZN(n16592) );
  OAI21_X1 U19523 ( .B1(n16593), .B2(n16614), .A(n16592), .ZN(U236) );
  INV_X1 U19524 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16595) );
  AOI22_X1 U19525 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16611), .ZN(n16594) );
  OAI21_X1 U19526 ( .B1(n16595), .B2(n16614), .A(n16594), .ZN(U237) );
  AOI22_X1 U19527 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16611), .ZN(n16596) );
  OAI21_X1 U19528 ( .B1(n20955), .B2(n16614), .A(n16596), .ZN(U238) );
  INV_X1 U19529 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16598) );
  AOI22_X1 U19530 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16611), .ZN(n16597) );
  OAI21_X1 U19531 ( .B1(n16598), .B2(n16614), .A(n16597), .ZN(U239) );
  INV_X1 U19532 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16600) );
  AOI22_X1 U19533 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16611), .ZN(n16599) );
  OAI21_X1 U19534 ( .B1(n16600), .B2(n16614), .A(n16599), .ZN(U240) );
  INV_X1 U19535 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16602) );
  AOI22_X1 U19536 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16611), .ZN(n16601) );
  OAI21_X1 U19537 ( .B1(n16602), .B2(n16614), .A(n16601), .ZN(U241) );
  INV_X1 U19538 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20928) );
  AOI22_X1 U19539 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16611), .ZN(n16603) );
  OAI21_X1 U19540 ( .B1(n20928), .B2(n16614), .A(n16603), .ZN(U242) );
  AOI22_X1 U19541 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16611), .ZN(n16604) );
  OAI21_X1 U19542 ( .B1(n16605), .B2(n16614), .A(n16604), .ZN(U243) );
  INV_X1 U19543 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20864) );
  AOI22_X1 U19544 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16611), .ZN(n16606) );
  OAI21_X1 U19545 ( .B1(n20864), .B2(n16614), .A(n16606), .ZN(U244) );
  INV_X1 U19546 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16608) );
  AOI22_X1 U19547 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16611), .ZN(n16607) );
  OAI21_X1 U19548 ( .B1(n16608), .B2(n16614), .A(n16607), .ZN(U245) );
  INV_X1 U19549 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16610) );
  AOI22_X1 U19550 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16611), .ZN(n16609) );
  OAI21_X1 U19551 ( .B1(n16610), .B2(n16614), .A(n16609), .ZN(U246) );
  INV_X1 U19552 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16615) );
  AOI22_X1 U19553 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16612), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16611), .ZN(n16613) );
  OAI21_X1 U19554 ( .B1(n16615), .B2(n16614), .A(n16613), .ZN(U247) );
  OAI22_X1 U19555 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16642), .ZN(n16616) );
  INV_X1 U19556 ( .A(n16616), .ZN(U251) );
  OAI22_X1 U19557 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16642), .ZN(n16617) );
  INV_X1 U19558 ( .A(n16617), .ZN(U252) );
  OAI22_X1 U19559 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16642), .ZN(n16618) );
  INV_X1 U19560 ( .A(n16618), .ZN(U253) );
  OAI22_X1 U19561 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16642), .ZN(n16619) );
  INV_X1 U19562 ( .A(n16619), .ZN(U254) );
  OAI22_X1 U19563 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16642), .ZN(n16620) );
  INV_X1 U19564 ( .A(n16620), .ZN(U255) );
  OAI22_X1 U19565 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16642), .ZN(n16621) );
  INV_X1 U19566 ( .A(n16621), .ZN(U256) );
  OAI22_X1 U19567 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16642), .ZN(n16622) );
  INV_X1 U19568 ( .A(n16622), .ZN(U257) );
  OAI22_X1 U19569 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16642), .ZN(n16623) );
  INV_X1 U19570 ( .A(n16623), .ZN(U258) );
  OAI22_X1 U19571 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16642), .ZN(n16624) );
  INV_X1 U19572 ( .A(n16624), .ZN(U259) );
  OAI22_X1 U19573 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16642), .ZN(n16625) );
  INV_X1 U19574 ( .A(n16625), .ZN(U260) );
  OAI22_X1 U19575 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16642), .ZN(n16626) );
  INV_X1 U19576 ( .A(n16626), .ZN(U261) );
  OAI22_X1 U19577 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16642), .ZN(n16627) );
  INV_X1 U19578 ( .A(n16627), .ZN(U262) );
  OAI22_X1 U19579 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16642), .ZN(n16628) );
  INV_X1 U19580 ( .A(n16628), .ZN(U263) );
  INV_X1 U19581 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U19582 ( .A1(n16642), .A2(n16629), .B1(n17424), .B2(U215), .ZN(U264) );
  OAI22_X1 U19583 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16642), .ZN(n16630) );
  INV_X1 U19584 ( .A(n16630), .ZN(U265) );
  OAI22_X1 U19585 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16642), .ZN(n16631) );
  INV_X1 U19586 ( .A(n16631), .ZN(U266) );
  INV_X1 U19587 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19271) );
  AOI22_X1 U19588 ( .A1(n16642), .A2(n21025), .B1(n19271), .B2(U215), .ZN(U267) );
  OAI22_X1 U19589 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16642), .ZN(n16632) );
  INV_X1 U19590 ( .A(n16632), .ZN(U268) );
  OAI22_X1 U19591 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16642), .ZN(n16633) );
  INV_X1 U19592 ( .A(n16633), .ZN(U269) );
  OAI22_X1 U19593 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16642), .ZN(n16634) );
  INV_X1 U19594 ( .A(n16634), .ZN(U270) );
  OAI22_X1 U19595 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16642), .ZN(n16635) );
  INV_X1 U19596 ( .A(n16635), .ZN(U271) );
  OAI22_X1 U19597 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16642), .ZN(n16636) );
  INV_X1 U19598 ( .A(n16636), .ZN(U272) );
  OAI22_X1 U19599 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16642), .ZN(n16637) );
  INV_X1 U19600 ( .A(n16637), .ZN(U273) );
  OAI22_X1 U19601 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16642), .ZN(n16638) );
  INV_X1 U19602 ( .A(n16638), .ZN(U274) );
  OAI22_X1 U19603 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16642), .ZN(n16639) );
  INV_X1 U19604 ( .A(n16639), .ZN(U275) );
  OAI22_X1 U19605 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16642), .ZN(n16640) );
  INV_X1 U19606 ( .A(n16640), .ZN(U277) );
  OAI22_X1 U19607 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16642), .ZN(n16641) );
  INV_X1 U19608 ( .A(n16641), .ZN(U278) );
  OAI22_X1 U19609 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16642), .ZN(n16643) );
  INV_X1 U19610 ( .A(n16643), .ZN(U279) );
  OAI22_X1 U19611 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16642), .ZN(n16644) );
  INV_X1 U19612 ( .A(n16644), .ZN(U280) );
  INV_X1 U19613 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18308) );
  AOI22_X1 U19614 ( .A1(n16642), .A2(n16646), .B1(n18308), .B2(U215), .ZN(U281) );
  INV_X1 U19615 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n20992) );
  AOI22_X1 U19616 ( .A1(n16642), .A2(n16645), .B1(n20992), .B2(U215), .ZN(U282) );
  INV_X1 U19617 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n20960) );
  OAI222_X1 U19618 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n21011), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n16646), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n20960), .ZN(n16648) );
  INV_X2 U19619 ( .A(n16649), .ZN(n16647) );
  INV_X1 U19620 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18827) );
  INV_X1 U19621 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U19622 ( .A1(n16647), .A2(n18827), .B1(n19881), .B2(n16649), .ZN(
        U347) );
  INV_X1 U19623 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18825) );
  INV_X1 U19624 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U19625 ( .A1(n16647), .A2(n18825), .B1(n19879), .B2(n16649), .ZN(
        U348) );
  INV_X1 U19626 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18823) );
  INV_X1 U19627 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n21144) );
  AOI22_X1 U19628 ( .A1(n16647), .A2(n18823), .B1(n21144), .B2(n16649), .ZN(
        U349) );
  INV_X1 U19629 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18822) );
  INV_X1 U19630 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U19631 ( .A1(n16647), .A2(n18822), .B1(n19877), .B2(n16649), .ZN(
        U350) );
  INV_X1 U19632 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18820) );
  INV_X1 U19633 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U19634 ( .A1(n16647), .A2(n18820), .B1(n19875), .B2(n16649), .ZN(
        U351) );
  INV_X1 U19635 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18817) );
  INV_X1 U19636 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U19637 ( .A1(n16647), .A2(n18817), .B1(n19874), .B2(n16649), .ZN(
        U352) );
  INV_X1 U19638 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18816) );
  INV_X1 U19639 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19873) );
  AOI22_X1 U19640 ( .A1(n16647), .A2(n18816), .B1(n19873), .B2(n16649), .ZN(
        U353) );
  INV_X1 U19641 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18814) );
  AOI22_X1 U19642 ( .A1(n16647), .A2(n18814), .B1(n19871), .B2(n16649), .ZN(
        U354) );
  INV_X1 U19643 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18866) );
  AOI22_X1 U19644 ( .A1(n16647), .A2(n18866), .B1(n19913), .B2(n16648), .ZN(
        U355) );
  INV_X1 U19645 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18864) );
  INV_X1 U19646 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19910) );
  AOI22_X1 U19647 ( .A1(n16647), .A2(n18864), .B1(n19910), .B2(n16649), .ZN(
        U356) );
  INV_X1 U19648 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18862) );
  INV_X1 U19649 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19908) );
  AOI22_X1 U19650 ( .A1(n16647), .A2(n18862), .B1(n19908), .B2(n16649), .ZN(
        U357) );
  INV_X1 U19651 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18859) );
  INV_X1 U19652 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19906) );
  AOI22_X1 U19653 ( .A1(n16647), .A2(n18859), .B1(n19906), .B2(n16648), .ZN(
        U358) );
  INV_X1 U19654 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18858) );
  INV_X1 U19655 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U19656 ( .A1(n16647), .A2(n18858), .B1(n19905), .B2(n16648), .ZN(
        U359) );
  INV_X1 U19657 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18856) );
  INV_X1 U19658 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19904) );
  AOI22_X1 U19659 ( .A1(n16647), .A2(n18856), .B1(n19904), .B2(n16648), .ZN(
        U360) );
  INV_X1 U19660 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18854) );
  INV_X1 U19661 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U19662 ( .A1(n16647), .A2(n18854), .B1(n19902), .B2(n16648), .ZN(
        U361) );
  INV_X1 U19663 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18851) );
  INV_X1 U19664 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19900) );
  AOI22_X1 U19665 ( .A1(n16647), .A2(n18851), .B1(n19900), .B2(n16648), .ZN(
        U362) );
  INV_X1 U19666 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18850) );
  INV_X1 U19667 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U19668 ( .A1(n16647), .A2(n18850), .B1(n19899), .B2(n16648), .ZN(
        U363) );
  INV_X1 U19669 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18848) );
  INV_X1 U19670 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19898) );
  AOI22_X1 U19671 ( .A1(n16647), .A2(n18848), .B1(n19898), .B2(n16649), .ZN(
        U364) );
  INV_X1 U19672 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18811) );
  INV_X1 U19673 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19869) );
  AOI22_X1 U19674 ( .A1(n16647), .A2(n18811), .B1(n19869), .B2(n16649), .ZN(
        U365) );
  INV_X1 U19675 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18846) );
  INV_X1 U19676 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19677 ( .A1(n16647), .A2(n18846), .B1(n19897), .B2(n16649), .ZN(
        U366) );
  INV_X1 U19678 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18845) );
  INV_X1 U19679 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19895) );
  AOI22_X1 U19680 ( .A1(n16647), .A2(n18845), .B1(n19895), .B2(n16649), .ZN(
        U367) );
  INV_X1 U19681 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18843) );
  INV_X1 U19682 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U19683 ( .A1(n16647), .A2(n18843), .B1(n19894), .B2(n16649), .ZN(
        U368) );
  INV_X1 U19684 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18840) );
  INV_X1 U19685 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U19686 ( .A1(n16647), .A2(n18840), .B1(n19892), .B2(n16649), .ZN(
        U369) );
  INV_X1 U19687 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18839) );
  INV_X1 U19688 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U19689 ( .A1(n16647), .A2(n18839), .B1(n19891), .B2(n16649), .ZN(
        U370) );
  INV_X1 U19690 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18837) );
  INV_X1 U19691 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U19692 ( .A1(n16647), .A2(n18837), .B1(n19889), .B2(n16649), .ZN(
        U371) );
  INV_X1 U19693 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18834) );
  INV_X1 U19694 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n21005) );
  AOI22_X1 U19695 ( .A1(n16647), .A2(n18834), .B1(n21005), .B2(n16649), .ZN(
        U372) );
  INV_X1 U19696 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18833) );
  INV_X1 U19697 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U19698 ( .A1(n16647), .A2(n18833), .B1(n19887), .B2(n16649), .ZN(
        U373) );
  INV_X1 U19699 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18831) );
  INV_X1 U19700 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U19701 ( .A1(n16647), .A2(n18831), .B1(n19885), .B2(n16649), .ZN(
        U374) );
  INV_X1 U19702 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18829) );
  INV_X1 U19703 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U19704 ( .A1(n16647), .A2(n18829), .B1(n19883), .B2(n16648), .ZN(
        U375) );
  INV_X1 U19705 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18808) );
  INV_X1 U19706 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U19707 ( .A1(n16647), .A2(n18808), .B1(n19868), .B2(n16649), .ZN(
        U376) );
  INV_X1 U19708 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18807) );
  NAND2_X1 U19709 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18807), .ZN(n18797) );
  AOI22_X1 U19710 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18797), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18805), .ZN(n18792) );
  AOI21_X1 U19711 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18792), .ZN(n16650) );
  INV_X1 U19712 ( .A(n16650), .ZN(P3_U2633) );
  NAND2_X1 U19713 ( .A1(n18930), .A2(n18880), .ZN(n16652) );
  OAI21_X1 U19714 ( .B1(n16656), .B2(n17484), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16651) );
  OAI21_X1 U19715 ( .B1(n16652), .B2(n18783), .A(n16651), .ZN(P3_U2634) );
  AOI21_X1 U19716 ( .B1(n18805), .B2(n18807), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16653) );
  AOI22_X1 U19717 ( .A1(n18872), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16653), 
        .B2(n18940), .ZN(P3_U2635) );
  OAI21_X1 U19718 ( .B1(n18793), .B2(BS16), .A(n18792), .ZN(n18874) );
  OAI21_X1 U19719 ( .B1(n18792), .B2(n16675), .A(n18874), .ZN(P3_U2636) );
  INV_X1 U19720 ( .A(n16654), .ZN(n16655) );
  NOR3_X1 U19721 ( .A1(n16656), .A2(n16655), .A3(n18749), .ZN(n18762) );
  NOR2_X1 U19722 ( .A1(n18762), .A2(n18925), .ZN(n18922) );
  OAI21_X1 U19723 ( .B1(n18922), .B2(n18265), .A(n16657), .ZN(P3_U2637) );
  NOR4_X1 U19724 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16661) );
  NOR4_X1 U19725 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16660) );
  NOR4_X1 U19726 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16659) );
  NOR4_X1 U19727 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16658) );
  NAND4_X1 U19728 ( .A1(n16661), .A2(n16660), .A3(n16659), .A4(n16658), .ZN(
        n16667) );
  NOR4_X1 U19729 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_2__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16665) );
  AOI211_X1 U19730 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_7__SCAN_IN), .B(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16664) );
  NOR4_X1 U19731 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16663) );
  NOR4_X1 U19732 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16662) );
  NAND4_X1 U19733 ( .A1(n16665), .A2(n16664), .A3(n16663), .A4(n16662), .ZN(
        n16666) );
  NOR2_X1 U19734 ( .A1(n16667), .A2(n16666), .ZN(n18920) );
  INV_X1 U19735 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16669) );
  NOR3_X1 U19736 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16670) );
  OAI21_X1 U19737 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16670), .A(n18920), .ZN(
        n16668) );
  OAI21_X1 U19738 ( .B1(n18920), .B2(n16669), .A(n16668), .ZN(P3_U2638) );
  INV_X1 U19739 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16672) );
  NOR2_X1 U19740 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18914) );
  OAI21_X1 U19741 ( .B1(n16670), .B2(n18914), .A(n18920), .ZN(n16671) );
  OAI21_X1 U19742 ( .B1(n18920), .B2(n16672), .A(n16671), .ZN(P3_U2639) );
  NAND2_X1 U19743 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18929), .ZN(n16674) );
  AOI211_X4 U19744 ( .C1(n18796), .C2(n16675), .A(n18945), .B(n16674), .ZN(
        n17035) );
  NOR3_X1 U19745 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17004) );
  NAND2_X1 U19746 ( .A1(n17004), .A2(n17316), .ZN(n17000) );
  NOR2_X1 U19747 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17000), .ZN(n16982) );
  NAND2_X1 U19748 ( .A1(n16982), .A2(n17311), .ZN(n16969) );
  NOR2_X1 U19749 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16969), .ZN(n16951) );
  NAND2_X1 U19750 ( .A1(n16951), .A2(n17305), .ZN(n16943) );
  NOR2_X1 U19751 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16943), .ZN(n16922) );
  NAND2_X1 U19752 ( .A1(n16922), .A2(n17265), .ZN(n16903) );
  NAND2_X1 U19753 ( .A1(n16902), .A2(n17236), .ZN(n16896) );
  INV_X1 U19754 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16873) );
  NAND2_X1 U19755 ( .A1(n16889), .A2(n16873), .ZN(n16872) );
  INV_X1 U19756 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16855) );
  NAND2_X1 U19757 ( .A1(n16858), .A2(n16855), .ZN(n16854) );
  INV_X1 U19758 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16832) );
  NAND2_X1 U19759 ( .A1(n16836), .A2(n16832), .ZN(n16831) );
  NAND2_X1 U19760 ( .A1(n16815), .A2(n16812), .ZN(n16811) );
  NOR2_X1 U19761 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16811), .ZN(n16794) );
  NAND2_X1 U19762 ( .A1(n16794), .A2(n20879), .ZN(n16789) );
  NOR2_X1 U19763 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16789), .ZN(n16775) );
  NAND2_X1 U19764 ( .A1(n16775), .A2(n17044), .ZN(n16767) );
  NOR2_X1 U19765 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16767), .ZN(n16757) );
  NAND2_X1 U19766 ( .A1(n16757), .A2(n21154), .ZN(n16747) );
  NOR2_X1 U19767 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16747), .ZN(n16740) );
  NAND2_X1 U19768 ( .A1(n16740), .A2(n21125), .ZN(n16734) );
  NOR2_X1 U19769 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16734), .ZN(n16722) );
  INV_X1 U19770 ( .A(n16722), .ZN(n16711) );
  NOR2_X1 U19771 ( .A1(n17028), .A2(n16701), .ZN(n16705) );
  INV_X1 U19772 ( .A(n16705), .ZN(n16698) );
  OAI211_X1 U19773 ( .C1(n18928), .C2(n18929), .A(n18796), .B(n16675), .ZN(
        n18773) );
  INV_X1 U19774 ( .A(n18773), .ZN(n16676) );
  AOI211_X4 U19775 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18929), .A(n16676), .B(
        n18945), .ZN(n17036) );
  INV_X1 U19776 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16678) );
  NAND2_X1 U19777 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16680), .ZN(
        n16679) );
  AOI21_X1 U19778 ( .B1(n16678), .B2(n16679), .A(n16677), .ZN(n17590) );
  OAI21_X1 U19779 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16680), .A(
        n16679), .ZN(n17610) );
  AOI21_X1 U19780 ( .B1(n20970), .B2(n17589), .A(n16680), .ZN(n17625) );
  INV_X1 U19781 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17935) );
  INV_X1 U19782 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21112) );
  NOR3_X1 U19783 ( .A1(n17935), .A2(n17633), .A3(n21112), .ZN(n16681) );
  OAI21_X1 U19784 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16681), .A(
        n17589), .ZN(n17636) );
  NOR2_X1 U19785 ( .A1(n17935), .A2(n17633), .ZN(n16683) );
  INV_X1 U19786 ( .A(n16681), .ZN(n16682) );
  OAI21_X1 U19787 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16683), .A(
        n16682), .ZN(n17646) );
  NOR2_X1 U19788 ( .A1(n17935), .A2(n17672), .ZN(n16686) );
  INV_X1 U19789 ( .A(n16686), .ZN(n16687) );
  NOR2_X1 U19790 ( .A1(n17673), .A2(n16687), .ZN(n17631) );
  OAI22_X1 U19791 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17631), .B1(
        n17935), .B2(n17633), .ZN(n17661) );
  INV_X1 U19792 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17686) );
  NOR2_X1 U19793 ( .A1(n17686), .A2(n16687), .ZN(n16685) );
  INV_X1 U19794 ( .A(n17631), .ZN(n16684) );
  OAI21_X1 U19795 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16685), .A(
        n16684), .ZN(n17676) );
  AOI22_X1 U19796 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16687), .B1(
        n16686), .B2(n17686), .ZN(n17683) );
  AND2_X1 U19797 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17695), .ZN(
        n17669) );
  OAI21_X1 U19798 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17669), .A(
        n16687), .ZN(n17693) );
  INV_X1 U19799 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17716) );
  NOR2_X1 U19800 ( .A1(n17935), .A2(n17744), .ZN(n17745) );
  INV_X1 U19801 ( .A(n17745), .ZN(n16860) );
  NOR2_X1 U19802 ( .A1(n17748), .A2(n16860), .ZN(n16824) );
  NAND2_X1 U19803 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16824), .ZN(
        n17708) );
  NAND2_X1 U19804 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17745), .ZN(
        n16846) );
  OAI21_X1 U19805 ( .B1(n16846), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n9751), .ZN(n16838) );
  INV_X1 U19806 ( .A(n16838), .ZN(n16849) );
  INV_X1 U19807 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20971) );
  XNOR2_X1 U19808 ( .A(n20971), .B(n17708), .ZN(n17724) );
  NAND2_X1 U19809 ( .A1(n16817), .A2(n17724), .ZN(n16816) );
  OAI21_X1 U19810 ( .B1(n17716), .B2(n16816), .A(n16953), .ZN(n16800) );
  NAND2_X1 U19811 ( .A1(n17693), .A2(n16800), .ZN(n16799) );
  NAND2_X1 U19812 ( .A1(n16953), .A2(n16799), .ZN(n16788) );
  NAND2_X1 U19813 ( .A1(n17683), .A2(n16788), .ZN(n16787) );
  NAND2_X1 U19814 ( .A1(n16953), .A2(n16787), .ZN(n16781) );
  NAND2_X1 U19815 ( .A1(n17676), .A2(n16781), .ZN(n16780) );
  NAND2_X1 U19816 ( .A1(n16953), .A2(n16780), .ZN(n16772) );
  NAND2_X1 U19817 ( .A1(n17661), .A2(n16772), .ZN(n16771) );
  NAND2_X1 U19818 ( .A1(n16953), .A2(n16771), .ZN(n16763) );
  NAND2_X1 U19819 ( .A1(n17646), .A2(n16763), .ZN(n16762) );
  NAND2_X1 U19820 ( .A1(n16953), .A2(n16762), .ZN(n16753) );
  NAND2_X1 U19821 ( .A1(n17636), .A2(n16753), .ZN(n16752) );
  OAI21_X1 U19822 ( .B1(n17625), .B2(n16752), .A(n16953), .ZN(n16731) );
  NOR2_X1 U19823 ( .A1(n16738), .A2(n17006), .ZN(n16724) );
  NOR2_X1 U19824 ( .A1(n17590), .A2(n16724), .ZN(n16723) );
  NOR2_X1 U19825 ( .A1(n16723), .A2(n17006), .ZN(n16713) );
  NOR2_X1 U19826 ( .A1(n16714), .A2(n16713), .ZN(n16712) );
  NOR2_X1 U19827 ( .A1(n16712), .A2(n17006), .ZN(n16699) );
  NOR4_X4 U19828 ( .A1(n18889), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n16929)
         );
  NAND2_X1 U19829 ( .A1(n18930), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18777) );
  INV_X1 U19830 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18857) );
  INV_X1 U19831 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18855) );
  INV_X1 U19832 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n21120) );
  INV_X1 U19833 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18841) );
  INV_X1 U19834 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18830) );
  INV_X1 U19835 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n21110) );
  INV_X1 U19836 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18815) );
  NAND3_X1 U19837 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16975) );
  NOR2_X1 U19838 ( .A1(n18815), .A2(n16975), .ZN(n16962) );
  NAND2_X1 U19839 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16962), .ZN(n16939) );
  NAND2_X1 U19840 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16938) );
  NOR3_X1 U19841 ( .A1(n21110), .A2(n16939), .A3(n16938), .ZN(n16909) );
  NAND4_X1 U19842 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16909), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16888) );
  NOR2_X1 U19843 ( .A1(n18830), .A2(n16888), .ZN(n16869) );
  NAND3_X1 U19844 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16869), .ZN(n16865) );
  NAND2_X1 U19845 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16843) );
  NOR3_X1 U19846 ( .A1(n18841), .A2(n16865), .A3(n16843), .ZN(n16804) );
  NAND3_X1 U19847 ( .A1(n16804), .A2(P3_REIP_REG_19__SCAN_IN), .A3(
        P3_REIP_REG_18__SCAN_IN), .ZN(n16796) );
  NOR2_X1 U19848 ( .A1(n21120), .A2(n16796), .ZN(n16786) );
  NAND4_X1 U19849 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .A4(n16786), .ZN(n16759) );
  INV_X1 U19850 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18853) );
  NAND4_X1 U19851 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16733), .ZN(n16692) );
  NAND2_X1 U19852 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18867), .ZN(n16688) );
  OAI22_X1 U19853 ( .A1(n16689), .A2(n17014), .B1(n16692), .B2(n16688), .ZN(
        n16690) );
  AOI211_X1 U19854 ( .C1(n17036), .C2(P3_EBX_REG_31__SCAN_IN), .A(n16691), .B(
        n16690), .ZN(n16697) );
  NOR2_X1 U19855 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16692), .ZN(n16704) );
  NAND2_X1 U19856 ( .A1(n17039), .A2(n17029), .ZN(n17038) );
  INV_X1 U19857 ( .A(n17038), .ZN(n16695) );
  INV_X1 U19858 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18863) );
  NAND2_X1 U19859 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16727) );
  NOR2_X1 U19860 ( .A1(n18863), .A2(n16727), .ZN(n16694) );
  NAND2_X1 U19861 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16693) );
  AOI21_X1 U19862 ( .B1(n17018), .B2(n16759), .A(n16974), .ZN(n16766) );
  OAI21_X1 U19863 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17029), .A(n16766), 
        .ZN(n16751) );
  AOI21_X1 U19864 ( .B1(n17018), .B2(n16693), .A(n16751), .ZN(n16721) );
  OAI21_X1 U19865 ( .B1(n16695), .B2(n16694), .A(n16721), .ZN(n16717) );
  OAI21_X1 U19866 ( .B1(n16704), .B2(n16717), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16696) );
  OAI211_X1 U19867 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16698), .A(n16697), .B(
        n16696), .ZN(P3_U2640) );
  XNOR2_X1 U19868 ( .A(n16700), .B(n16699), .ZN(n16708) );
  NAND2_X1 U19869 ( .A1(n17035), .A2(n16701), .ZN(n16710) );
  OAI22_X1 U19870 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16710), .B1(n16702), 
        .B2(n17014), .ZN(n16703) );
  AOI211_X1 U19871 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n16717), .A(n16704), 
        .B(n16703), .ZN(n16707) );
  OAI21_X1 U19872 ( .B1(n17036), .B2(n16705), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16706) );
  OAI211_X1 U19873 ( .C1(n18787), .C2(n16708), .A(n16707), .B(n16706), .ZN(
        P3_U2641) );
  NOR2_X1 U19874 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16727), .ZN(n16709) );
  AOI22_X1 U19875 ( .A1(n17036), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16733), 
        .B2(n16709), .ZN(n16719) );
  AOI21_X1 U19876 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16711), .A(n16710), .ZN(
        n16716) );
  AOI211_X1 U19877 ( .C1(n16714), .C2(n16713), .A(n16712), .B(n18787), .ZN(
        n16715) );
  AOI211_X1 U19878 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16717), .A(n16716), 
        .B(n16715), .ZN(n16718) );
  OAI211_X1 U19879 ( .C1(n16720), .C2(n17014), .A(n16719), .B(n16718), .ZN(
        P3_U2642) );
  AOI22_X1 U19880 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17021), .B1(
        n17036), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16730) );
  INV_X1 U19881 ( .A(n16721), .ZN(n16743) );
  AOI211_X1 U19882 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16734), .A(n16722), .B(
        n17028), .ZN(n16726) );
  AOI211_X1 U19883 ( .C1(n17590), .C2(n16724), .A(n16723), .B(n18787), .ZN(
        n16725) );
  AOI211_X1 U19884 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16743), .A(n16726), 
        .B(n16725), .ZN(n16729) );
  OAI211_X1 U19885 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16733), .B(n16727), .ZN(n16728) );
  NAND3_X1 U19886 ( .A1(n16730), .A2(n16729), .A3(n16728), .ZN(P3_U2643) );
  OAI21_X1 U19887 ( .B1(n17610), .B2(n16731), .A(n16929), .ZN(n16737) );
  INV_X1 U19888 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21014) );
  INV_X1 U19889 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17613) );
  OAI22_X1 U19890 ( .A1(n17613), .A2(n17014), .B1(n17026), .B2(n21125), .ZN(
        n16732) );
  AOI221_X1 U19891 ( .B1(n16733), .B2(n21014), .C1(n16743), .C2(
        P3_REIP_REG_27__SCAN_IN), .A(n16732), .ZN(n16736) );
  OAI211_X1 U19892 ( .C1(n16740), .C2(n21125), .A(n17035), .B(n16734), .ZN(
        n16735) );
  OAI211_X1 U19893 ( .C1(n16738), .C2(n16737), .A(n16736), .B(n16735), .ZN(
        P3_U2644) );
  NAND2_X1 U19894 ( .A1(n16953), .A2(n16752), .ZN(n16739) );
  XOR2_X1 U19895 ( .A(n17625), .B(n16739), .Z(n16746) );
  AOI22_X1 U19896 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17021), .B1(
        n17036), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16745) );
  OAI21_X1 U19897 ( .B1(n18855), .B2(n16749), .A(n18857), .ZN(n16742) );
  AOI211_X1 U19898 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16747), .A(n16740), .B(
        n17028), .ZN(n16741) );
  AOI21_X1 U19899 ( .B1(n16743), .B2(n16742), .A(n16741), .ZN(n16744) );
  OAI211_X1 U19900 ( .C1(n18787), .C2(n16746), .A(n16745), .B(n16744), .ZN(
        P3_U2645) );
  AOI22_X1 U19901 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17021), .B1(
        n17036), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16756) );
  OAI211_X1 U19902 ( .C1(n16757), .C2(n21154), .A(n17035), .B(n16747), .ZN(
        n16748) );
  OAI21_X1 U19903 ( .B1(n16749), .B2(P3_REIP_REG_25__SCAN_IN), .A(n16748), 
        .ZN(n16750) );
  AOI21_X1 U19904 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16751), .A(n16750), 
        .ZN(n16755) );
  OAI211_X1 U19905 ( .C1(n17636), .C2(n16753), .A(n16929), .B(n16752), .ZN(
        n16754) );
  NAND3_X1 U19906 ( .A1(n16756), .A2(n16755), .A3(n16754), .ZN(P3_U2646) );
  AOI211_X1 U19907 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16767), .A(n16757), .B(
        n17028), .ZN(n16761) );
  NAND2_X1 U19908 ( .A1(n17018), .A2(n18853), .ZN(n16758) );
  OAI22_X1 U19909 ( .A1(n21112), .A2(n17014), .B1(n16759), .B2(n16758), .ZN(
        n16760) );
  AOI211_X1 U19910 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17036), .A(n16761), .B(
        n16760), .ZN(n16765) );
  OAI211_X1 U19911 ( .C1(n17646), .C2(n16763), .A(n16929), .B(n16762), .ZN(
        n16764) );
  OAI211_X1 U19912 ( .C1(n16766), .C2(n18853), .A(n16765), .B(n16764), .ZN(
        P3_U2647) );
  INV_X1 U19913 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18849) );
  INV_X1 U19914 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18852) );
  NAND3_X1 U19915 ( .A1(n17018), .A2(P3_REIP_REG_21__SCAN_IN), .A3(n16786), 
        .ZN(n16784) );
  AOI221_X1 U19916 ( .B1(n18849), .B2(n18852), .C1(n16784), .C2(n18852), .A(
        n16766), .ZN(n16770) );
  OAI211_X1 U19917 ( .C1(n17044), .C2(n16775), .A(n16767), .B(n17035), .ZN(
        n16768) );
  INV_X1 U19918 ( .A(n16768), .ZN(n16769) );
  AOI211_X1 U19919 ( .C1(n17021), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16770), .B(n16769), .ZN(n16774) );
  OAI211_X1 U19920 ( .C1(n17661), .C2(n16772), .A(n16929), .B(n16771), .ZN(
        n16773) );
  OAI211_X1 U19921 ( .C1(n17044), .C2(n17026), .A(n16774), .B(n16773), .ZN(
        P3_U2648) );
  OAI221_X1 U19922 ( .B1(n17029), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n17029), 
        .C2(n16786), .A(n17039), .ZN(n16779) );
  AOI211_X1 U19923 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16789), .A(n16775), .B(
        n17028), .ZN(n16778) );
  AOI22_X1 U19924 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17021), .B1(
        n17036), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16776) );
  INV_X1 U19925 ( .A(n16776), .ZN(n16777) );
  AOI211_X1 U19926 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16779), .A(n16778), 
        .B(n16777), .ZN(n16783) );
  OAI211_X1 U19927 ( .C1(n17676), .C2(n16781), .A(n16929), .B(n16780), .ZN(
        n16782) );
  OAI211_X1 U19928 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16784), .A(n16783), 
        .B(n16782), .ZN(P3_U2649) );
  OAI21_X1 U19929 ( .B1(n16786), .B2(n17029), .A(n17039), .ZN(n16798) );
  OAI22_X1 U19930 ( .A1(n17686), .A2(n17014), .B1(n17026), .B2(n20879), .ZN(
        n16785) );
  AOI21_X1 U19931 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16798), .A(n16785), 
        .ZN(n16793) );
  INV_X1 U19932 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18847) );
  NAND3_X1 U19933 ( .A1(n17018), .A2(n16786), .A3(n18847), .ZN(n16792) );
  OAI211_X1 U19934 ( .C1(n17683), .C2(n16788), .A(n16929), .B(n16787), .ZN(
        n16791) );
  OAI211_X1 U19935 ( .C1(n16794), .C2(n20879), .A(n17035), .B(n16789), .ZN(
        n16790) );
  NAND4_X1 U19936 ( .A1(n16793), .A2(n16792), .A3(n16791), .A4(n16790), .ZN(
        P3_U2650) );
  AOI211_X1 U19937 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16811), .A(n16794), .B(
        n17028), .ZN(n16795) );
  AOI21_X1 U19938 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17036), .A(n16795), .ZN(
        n16803) );
  OAI21_X1 U19939 ( .B1(n17029), .B2(n16796), .A(n21120), .ZN(n16797) );
  AOI22_X1 U19940 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17021), .B1(
        n16798), .B2(n16797), .ZN(n16802) );
  OAI211_X1 U19941 ( .C1(n17693), .C2(n16800), .A(n16929), .B(n16799), .ZN(
        n16801) );
  NAND3_X1 U19942 ( .A1(n16803), .A2(n16802), .A3(n16801), .ZN(P3_U2651) );
  OAI21_X1 U19943 ( .B1(n16804), .B2(n17029), .A(n17039), .ZN(n16830) );
  INV_X1 U19944 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18844) );
  INV_X1 U19945 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18842) );
  NOR3_X1 U19946 ( .A1(n17029), .A2(n16865), .A3(n16843), .ZN(n16829) );
  NAND2_X1 U19947 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16829), .ZN(n16823) );
  AOI221_X1 U19948 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n18844), .C2(n18842), .A(n16823), .ZN(n16810) );
  OR2_X1 U19949 ( .A1(n20971), .A2(n17708), .ZN(n16805) );
  AOI21_X1 U19950 ( .B1(n17716), .B2(n16805), .A(n17669), .ZN(n17710) );
  AND2_X1 U19951 ( .A1(n16816), .A2(n16953), .ZN(n16807) );
  AOI21_X1 U19952 ( .B1(n17710), .B2(n16807), .A(n18787), .ZN(n16806) );
  OAI21_X1 U19953 ( .B1(n17710), .B2(n16807), .A(n16806), .ZN(n16808) );
  OAI211_X1 U19954 ( .C1(n17026), .C2(n16812), .A(n18148), .B(n16808), .ZN(
        n16809) );
  AOI211_X1 U19955 ( .C1(n16830), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16810), 
        .B(n16809), .ZN(n16814) );
  OAI211_X1 U19956 ( .C1(n16815), .C2(n16812), .A(n17035), .B(n16811), .ZN(
        n16813) );
  OAI211_X1 U19957 ( .C1(n17014), .C2(n17716), .A(n16814), .B(n16813), .ZN(
        P3_U2652) );
  INV_X1 U19958 ( .A(n16830), .ZN(n16822) );
  AOI211_X1 U19959 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16831), .A(n16815), .B(
        n17028), .ZN(n16820) );
  OAI211_X1 U19960 ( .C1(n16817), .C2(n17724), .A(n16929), .B(n16816), .ZN(
        n16818) );
  OAI211_X1 U19961 ( .C1(n17026), .C2(n17168), .A(n18148), .B(n16818), .ZN(
        n16819) );
  AOI211_X1 U19962 ( .C1(n17021), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16820), .B(n16819), .ZN(n16821) );
  OAI221_X1 U19963 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16823), .C1(n18842), 
        .C2(n16822), .A(n16821), .ZN(P3_U2653) );
  INV_X1 U19964 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16835) );
  OAI21_X1 U19965 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16824), .A(
        n17708), .ZN(n17737) );
  INV_X1 U19966 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16840) );
  AOI21_X1 U19967 ( .B1(n16840), .B2(n16846), .A(n16824), .ZN(n16837) );
  OAI21_X1 U19968 ( .B1(n16837), .B2(n16849), .A(n16953), .ZN(n16826) );
  AOI21_X1 U19969 ( .B1(n17737), .B2(n16826), .A(n18787), .ZN(n16825) );
  OAI21_X1 U19970 ( .B1(n17737), .B2(n16826), .A(n16825), .ZN(n16827) );
  OAI211_X1 U19971 ( .C1(n17026), .C2(n16832), .A(n18148), .B(n16827), .ZN(
        n16828) );
  AOI221_X1 U19972 ( .B1(n16830), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16829), 
        .C2(n18841), .A(n16828), .ZN(n16834) );
  OAI211_X1 U19973 ( .C1(n16836), .C2(n16832), .A(n17035), .B(n16831), .ZN(
        n16833) );
  OAI211_X1 U19974 ( .C1(n17014), .C2(n16835), .A(n16834), .B(n16833), .ZN(
        P3_U2654) );
  AOI21_X1 U19975 ( .B1(n17018), .B2(n16865), .A(n16974), .ZN(n16868) );
  INV_X1 U19976 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18838) );
  AOI211_X1 U19977 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16854), .A(n16836), .B(
        n17028), .ZN(n16842) );
  INV_X1 U19978 ( .A(n16837), .ZN(n17751) );
  OAI221_X1 U19979 ( .B1(n16838), .B2(n17751), .C1(n16849), .C2(n16837), .A(
        n16929), .ZN(n16839) );
  OAI211_X1 U19980 ( .C1(n16840), .C2(n17014), .A(n18148), .B(n16839), .ZN(
        n16841) );
  AOI211_X1 U19981 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17036), .A(n16842), .B(
        n16841), .ZN(n16845) );
  NOR2_X1 U19982 ( .A1(n17029), .A2(n16865), .ZN(n16853) );
  OAI211_X1 U19983 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16853), .B(n16843), .ZN(n16844) );
  OAI211_X1 U19984 ( .C1(n16868), .C2(n18838), .A(n16845), .B(n16844), .ZN(
        P3_U2655) );
  INV_X1 U19985 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17759) );
  INV_X1 U19986 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18836) );
  OAI21_X1 U19987 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17745), .A(
        n16846), .ZN(n17756) );
  NAND2_X1 U19988 ( .A1(n16953), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16847) );
  NAND2_X1 U19989 ( .A1(n16929), .A2(n16847), .ZN(n17023) );
  AOI211_X1 U19990 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16953), .A(
        n17756), .B(n17023), .ZN(n16848) );
  AOI211_X1 U19991 ( .C1(n17036), .C2(P3_EBX_REG_15__SCAN_IN), .A(n18255), .B(
        n16848), .ZN(n16851) );
  NAND3_X1 U19992 ( .A1(n16929), .A2(n16849), .A3(n17756), .ZN(n16850) );
  OAI211_X1 U19993 ( .C1(n16868), .C2(n18836), .A(n16851), .B(n16850), .ZN(
        n16852) );
  AOI21_X1 U19994 ( .B1(n16853), .B2(n18836), .A(n16852), .ZN(n16857) );
  OAI211_X1 U19995 ( .C1(n16858), .C2(n16855), .A(n17035), .B(n16854), .ZN(
        n16856) );
  OAI211_X1 U19996 ( .C1(n17014), .C2(n17759), .A(n16857), .B(n16856), .ZN(
        P3_U2656) );
  INV_X1 U19997 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18835) );
  AOI211_X1 U19998 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16872), .A(n16858), .B(
        n17028), .ZN(n16864) );
  INV_X1 U19999 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17825) );
  INV_X1 U20000 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20914) );
  INV_X1 U20001 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17883) );
  NAND2_X1 U20002 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17872), .ZN(
        n16963) );
  NOR2_X1 U20003 ( .A1(n17883), .A2(n16963), .ZN(n16952) );
  NAND2_X1 U20004 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16952), .ZN(
        n16940) );
  NOR2_X1 U20005 ( .A1(n20914), .A2(n16940), .ZN(n16925) );
  NAND2_X1 U20006 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16925), .ZN(
        n16916) );
  NOR2_X1 U20007 ( .A1(n17825), .A2(n16916), .ZN(n16905) );
  NAND2_X1 U20008 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16905), .ZN(
        n17784) );
  NOR2_X1 U20009 ( .A1(n16859), .A2(n17784), .ZN(n16870) );
  OAI21_X1 U20010 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16870), .A(
        n16860), .ZN(n17770) );
  INV_X1 U20011 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17007) );
  NAND2_X1 U20012 ( .A1(n16952), .A2(n17007), .ZN(n16941) );
  OAI21_X1 U20013 ( .B1(n17767), .B2(n16941), .A(n16953), .ZN(n16884) );
  OAI21_X1 U20014 ( .B1(n17780), .B2(n17006), .A(n16884), .ZN(n16874) );
  OAI21_X1 U20015 ( .B1(n17770), .B2(n16874), .A(n18148), .ZN(n16861) );
  AOI21_X1 U20016 ( .B1(n17770), .B2(n16874), .A(n16861), .ZN(n16862) );
  INV_X1 U20017 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n21135) );
  OAI22_X1 U20018 ( .A1(n16967), .A2(n16862), .B1(n17026), .B2(n21135), .ZN(
        n16863) );
  AOI211_X1 U20019 ( .C1(n17021), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16864), .B(n16863), .ZN(n16867) );
  NAND4_X1 U20020 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17018), .A3(n16869), 
        .A4(n16865), .ZN(n16866) );
  OAI211_X1 U20021 ( .C1(n16868), .C2(n18835), .A(n16867), .B(n16866), .ZN(
        P3_U2657) );
  NAND2_X1 U20022 ( .A1(n17018), .A2(n16869), .ZN(n16882) );
  AOI22_X1 U20023 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17021), .B1(
        n17036), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16881) );
  AOI21_X1 U20024 ( .B1(n17018), .B2(n16888), .A(n16974), .ZN(n16894) );
  OAI21_X1 U20025 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17029), .A(n16894), 
        .ZN(n16879) );
  INV_X1 U20026 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17797) );
  NOR2_X1 U20027 ( .A1(n17797), .A2(n17784), .ZN(n16883) );
  INV_X1 U20028 ( .A(n16870), .ZN(n16871) );
  OAI21_X1 U20029 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16883), .A(
        n16871), .ZN(n17785) );
  AOI211_X1 U20030 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16953), .A(
        n17785), .B(n17023), .ZN(n16878) );
  OAI211_X1 U20031 ( .C1(n16889), .C2(n16873), .A(n17035), .B(n16872), .ZN(
        n16876) );
  NAND3_X1 U20032 ( .A1(n16929), .A2(n17785), .A3(n16874), .ZN(n16875) );
  NAND3_X1 U20033 ( .A1(n18148), .A2(n16876), .A3(n16875), .ZN(n16877) );
  AOI211_X1 U20034 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16879), .A(n16878), 
        .B(n16877), .ZN(n16880) );
  OAI211_X1 U20035 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16882), .A(n16881), 
        .B(n16880), .ZN(P3_U2658) );
  AOI21_X1 U20036 ( .B1(n17797), .B2(n17784), .A(n16883), .ZN(n17800) );
  INV_X1 U20037 ( .A(n16884), .ZN(n16886) );
  INV_X1 U20038 ( .A(n17800), .ZN(n16885) );
  AOI221_X1 U20039 ( .B1(n17800), .B2(n16886), .C1(n16885), .C2(n16884), .A(
        n18787), .ZN(n16887) );
  AOI211_X1 U20040 ( .C1(n17036), .C2(P3_EBX_REG_12__SCAN_IN), .A(n18255), .B(
        n16887), .ZN(n16893) );
  NOR3_X1 U20041 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17029), .A3(n16888), 
        .ZN(n16891) );
  AOI211_X1 U20042 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16896), .A(n16889), .B(
        n17028), .ZN(n16890) );
  AOI211_X1 U20043 ( .C1(n17021), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16891), .B(n16890), .ZN(n16892) );
  OAI211_X1 U20044 ( .C1(n16894), .C2(n18830), .A(n16893), .B(n16892), .ZN(
        P3_U2659) );
  NAND2_X1 U20045 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16911) );
  INV_X1 U20046 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18828) );
  NAND2_X1 U20047 ( .A1(n17018), .A2(n16909), .ZN(n16915) );
  AOI221_X1 U20048 ( .B1(n16911), .B2(n18828), .C1(n16915), .C2(n18828), .A(
        n16894), .ZN(n16900) );
  OAI21_X1 U20049 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16905), .A(
        n17784), .ZN(n17811) );
  AOI21_X1 U20050 ( .B1(n16905), .B2(n17007), .A(n17006), .ZN(n16895) );
  XOR2_X1 U20051 ( .A(n17811), .B(n16895), .Z(n16898) );
  OAI211_X1 U20052 ( .C1(n16902), .C2(n17236), .A(n17035), .B(n16896), .ZN(
        n16897) );
  OAI211_X1 U20053 ( .C1(n16898), .C2(n18787), .A(n18148), .B(n16897), .ZN(
        n16899) );
  AOI211_X1 U20054 ( .C1(n17021), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16900), .B(n16899), .ZN(n16901) );
  OAI21_X1 U20055 ( .B1(n17026), .B2(n17236), .A(n16901), .ZN(P3_U2660) );
  AOI211_X1 U20056 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16903), .A(n16902), .B(
        n17028), .ZN(n16908) );
  OAI21_X1 U20057 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16916), .A(
        n16953), .ZN(n16904) );
  INV_X1 U20058 ( .A(n16904), .ZN(n16918) );
  AOI21_X1 U20059 ( .B1(n17825), .B2(n16916), .A(n16905), .ZN(n17820) );
  XNOR2_X1 U20060 ( .A(n16918), .B(n17820), .ZN(n16906) );
  OAI21_X1 U20061 ( .B1(n16906), .B2(n18787), .A(n18148), .ZN(n16907) );
  AOI211_X1 U20062 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17036), .A(n16908), .B(
        n16907), .ZN(n16913) );
  NAND2_X1 U20063 ( .A1(n16909), .A2(n17039), .ZN(n16914) );
  INV_X1 U20064 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18824) );
  INV_X1 U20065 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18826) );
  OAI21_X1 U20066 ( .B1(n18824), .B2(n16915), .A(n18826), .ZN(n16910) );
  OAI211_X1 U20067 ( .C1(n16911), .C2(n16914), .A(n16910), .B(n17038), .ZN(
        n16912) );
  OAI211_X1 U20068 ( .C1(n17014), .C2(n17825), .A(n16913), .B(n16912), .ZN(
        P3_U2661) );
  NAND2_X1 U20069 ( .A1(n17038), .A2(n16914), .ZN(n16931) );
  OR2_X1 U20070 ( .A1(n17028), .A2(n16922), .ZN(n16930) );
  OAI22_X1 U20071 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16915), .B1(
        P3_EBX_REG_9__SCAN_IN), .B2(n16930), .ZN(n16921) );
  OAI21_X1 U20072 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16925), .A(
        n16916), .ZN(n17838) );
  NOR3_X1 U20073 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17834), .A3(
        n16941), .ZN(n16917) );
  AOI211_X1 U20074 ( .C1(n17838), .C2(n16918), .A(n18255), .B(n16917), .ZN(
        n16919) );
  NOR2_X1 U20075 ( .A1(n18787), .A2(n16953), .ZN(n17005) );
  INV_X1 U20076 ( .A(n17005), .ZN(n16983) );
  OAI22_X1 U20077 ( .A1(n16967), .A2(n16919), .B1(n16983), .B2(n17838), .ZN(
        n16920) );
  AOI211_X1 U20078 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17021), .A(
        n16921), .B(n16920), .ZN(n16924) );
  OAI221_X1 U20079 ( .B1(n17036), .B2(n17035), .C1(n17036), .C2(n16922), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n16923) );
  OAI211_X1 U20080 ( .C1(n16931), .C2(n18824), .A(n16924), .B(n16923), .ZN(
        P3_U2662) );
  AOI21_X1 U20081 ( .B1(n20914), .B2(n16940), .A(n16925), .ZN(n17853) );
  INV_X1 U20082 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17868) );
  OR2_X1 U20083 ( .A1(n17849), .A2(n17868), .ZN(n17848) );
  NOR2_X1 U20084 ( .A1(n17935), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17011) );
  INV_X1 U20085 ( .A(n17011), .ZN(n16926) );
  OAI21_X1 U20086 ( .B1(n17848), .B2(n16926), .A(n16953), .ZN(n16927) );
  XNOR2_X1 U20087 ( .A(n17853), .B(n16927), .ZN(n16928) );
  AOI22_X1 U20088 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17021), .B1(
        n16929), .B2(n16928), .ZN(n16937) );
  AOI21_X1 U20089 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16943), .A(n16930), .ZN(
        n16935) );
  OR2_X1 U20090 ( .A1(n17029), .A2(n16939), .ZN(n16961) );
  NOR2_X1 U20091 ( .A1(n16938), .A2(n16961), .ZN(n16933) );
  INV_X1 U20092 ( .A(n16931), .ZN(n16932) );
  MUX2_X1 U20093 ( .A(n16933), .B(n16932), .S(P3_REIP_REG_8__SCAN_IN), .Z(
        n16934) );
  AOI211_X1 U20094 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17036), .A(n16935), .B(
        n16934), .ZN(n16936) );
  NAND3_X1 U20095 ( .A1(n16937), .A2(n16936), .A3(n18148), .ZN(P3_U2663) );
  OAI21_X1 U20096 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16938), .ZN(n16950) );
  AOI21_X1 U20097 ( .B1(n16939), .B2(n17018), .A(n16974), .ZN(n16972) );
  INV_X1 U20098 ( .A(n16972), .ZN(n16948) );
  OAI22_X1 U20099 ( .A1(n17868), .A2(n17014), .B1(n17026), .B2(n17305), .ZN(
        n16947) );
  OAI21_X1 U20100 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16952), .A(
        n16940), .ZN(n17864) );
  NAND2_X1 U20101 ( .A1(n16953), .A2(n16941), .ZN(n16954) );
  XNOR2_X1 U20102 ( .A(n17864), .B(n16954), .ZN(n16945) );
  OAI211_X1 U20103 ( .C1(n16951), .C2(n17305), .A(n17035), .B(n16943), .ZN(
        n16944) );
  OAI211_X1 U20104 ( .C1(n18787), .C2(n16945), .A(n18148), .B(n16944), .ZN(
        n16946) );
  AOI211_X1 U20105 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n16948), .A(n16947), .B(
        n16946), .ZN(n16949) );
  OAI21_X1 U20106 ( .B1(n16961), .B2(n16950), .A(n16949), .ZN(P3_U2664) );
  INV_X1 U20107 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18819) );
  AOI211_X1 U20108 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16969), .A(n16951), .B(
        n17028), .ZN(n16959) );
  AOI21_X1 U20109 ( .B1(n17883), .B2(n16963), .A(n16952), .ZN(n17880) );
  AOI21_X1 U20110 ( .B1(n16953), .B2(n16963), .A(n17023), .ZN(n16956) );
  NOR3_X1 U20111 ( .A1(n17880), .A2(n18787), .A3(n16954), .ZN(n16955) );
  AOI211_X1 U20112 ( .C1(n17880), .C2(n16956), .A(n18255), .B(n16955), .ZN(
        n16957) );
  OAI21_X1 U20113 ( .B1(n17026), .B2(n10029), .A(n16957), .ZN(n16958) );
  AOI211_X1 U20114 ( .C1(n17021), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16959), .B(n16958), .ZN(n16960) );
  OAI221_X1 U20115 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16961), .C1(n18819), 
        .C2(n16972), .A(n16960), .ZN(P3_U2665) );
  AOI21_X1 U20116 ( .B1(n17018), .B2(n16962), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16973) );
  NOR3_X1 U20117 ( .A1(n17935), .A2(n16976), .A3(n16978), .ZN(n16977) );
  OAI21_X1 U20118 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16977), .A(
        n16963), .ZN(n17890) );
  INV_X1 U20119 ( .A(n17890), .ZN(n16965) );
  AOI21_X1 U20120 ( .B1(n16977), .B2(n17007), .A(n17006), .ZN(n16980) );
  INV_X1 U20121 ( .A(n16980), .ZN(n16964) );
  AOI221_X1 U20122 ( .B1(n16965), .B2(n16964), .C1(n17890), .C2(n16980), .A(
        n18255), .ZN(n16966) );
  OAI22_X1 U20123 ( .A1(n16967), .A2(n16966), .B1(n17026), .B2(n17311), .ZN(
        n16968) );
  AOI21_X1 U20124 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17021), .A(
        n16968), .ZN(n16971) );
  OAI211_X1 U20125 ( .C1(n16982), .C2(n17311), .A(n17035), .B(n16969), .ZN(
        n16970) );
  OAI211_X1 U20126 ( .C1(n16973), .C2(n16972), .A(n16971), .B(n16970), .ZN(
        P3_U2666) );
  AOI21_X1 U20127 ( .B1(n17018), .B2(n16975), .A(n16974), .ZN(n16991) );
  AOI22_X1 U20128 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17021), .B1(
        n17036), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16990) );
  INV_X1 U20129 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18813) );
  NAND3_X1 U20130 ( .A1(n17018), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .ZN(n16992) );
  NOR3_X1 U20131 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18813), .A3(n16992), .ZN(
        n16988) );
  NOR2_X1 U20132 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16976), .ZN(
        n17900) );
  OR2_X1 U20133 ( .A1(n17935), .A2(n16976), .ZN(n16994) );
  AOI21_X1 U20134 ( .B1(n16978), .B2(n16994), .A(n16977), .ZN(n16979) );
  INV_X1 U20135 ( .A(n16979), .ZN(n17907) );
  AOI22_X1 U20136 ( .A1(n17011), .A2(n17900), .B1(n17907), .B2(n16980), .ZN(
        n16981) );
  OAI21_X1 U20137 ( .B1(n16981), .B2(n18787), .A(n18148), .ZN(n16987) );
  AOI211_X1 U20138 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17000), .A(n16982), .B(
        n17028), .ZN(n16986) );
  NOR2_X1 U20139 ( .A1(n17275), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16984) );
  NOR2_X1 U20140 ( .A1(n17485), .A2(n18943), .ZN(n17037) );
  INV_X1 U20141 ( .A(n17037), .ZN(n17025) );
  OAI22_X1 U20142 ( .A1(n16984), .A2(n17025), .B1(n17907), .B2(n16983), .ZN(
        n16985) );
  NOR4_X1 U20143 ( .A1(n16988), .A2(n16987), .A3(n16986), .A4(n16985), .ZN(
        n16989) );
  OAI211_X1 U20144 ( .C1(n16991), .C2(n18815), .A(n16990), .B(n16989), .ZN(
        P3_U2667) );
  INV_X1 U20145 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17003) );
  AOI21_X1 U20146 ( .B1(n18813), .B2(n16992), .A(n16991), .ZN(n16999) );
  NAND2_X1 U20147 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18735) );
  NOR2_X1 U20148 ( .A1(n18910), .A2(n18735), .ZN(n18715) );
  OAI21_X1 U20149 ( .B1(n18886), .B2(n18715), .A(n16993), .ZN(n18884) );
  INV_X1 U20150 ( .A(n18884), .ZN(n16997) );
  INV_X1 U20151 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17925) );
  NOR2_X1 U20152 ( .A1(n17935), .A2(n17925), .ZN(n17008) );
  AOI21_X1 U20153 ( .B1(n17008), .B2(n17007), .A(n17006), .ZN(n16995) );
  OAI21_X1 U20154 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17008), .A(
        n16994), .ZN(n17918) );
  XOR2_X1 U20155 ( .A(n16995), .B(n17918), .Z(n16996) );
  OAI22_X1 U20156 ( .A1(n16997), .A2(n17025), .B1(n18787), .B2(n16996), .ZN(
        n16998) );
  AOI211_X1 U20157 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n17036), .A(n16999), .B(
        n16998), .ZN(n17002) );
  OAI211_X1 U20158 ( .C1(n17004), .C2(n17316), .A(n17035), .B(n17000), .ZN(
        n17001) );
  OAI211_X1 U20159 ( .C1(n17014), .C2(n17003), .A(n17002), .B(n17001), .ZN(
        P3_U2668) );
  INV_X1 U20160 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18810) );
  INV_X1 U20161 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17042) );
  NAND2_X1 U20162 ( .A1(n17042), .A2(n17325), .ZN(n17027) );
  AOI211_X1 U20163 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17027), .A(n17004), .B(
        n17028), .ZN(n17016) );
  AOI21_X1 U20164 ( .B1(n18896), .B2(n18741), .A(n18715), .ZN(n18892) );
  AOI21_X1 U20165 ( .B1(n17935), .B2(n17925), .A(n17008), .ZN(n17928) );
  AOI22_X1 U20166 ( .A1(n18892), .A2(n17037), .B1(n17928), .B2(n17005), .ZN(
        n17013) );
  INV_X1 U20167 ( .A(n17928), .ZN(n17010) );
  NOR2_X1 U20168 ( .A1(n17006), .A2(n18787), .ZN(n17022) );
  NAND2_X1 U20169 ( .A1(n17008), .A2(n17007), .ZN(n17009) );
  OAI211_X1 U20170 ( .C1(n17011), .C2(n17010), .A(n17022), .B(n17009), .ZN(
        n17012) );
  OAI211_X1 U20171 ( .C1(n17014), .C2(n17925), .A(n17013), .B(n17012), .ZN(
        n17015) );
  AOI211_X1 U20172 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17036), .A(n17016), .B(
        n17015), .ZN(n17020) );
  NAND2_X1 U20173 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17017) );
  OAI211_X1 U20174 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17018), .B(n17017), .ZN(n17019) );
  OAI211_X1 U20175 ( .C1(n18810), .C2(n17039), .A(n17020), .B(n17019), .ZN(
        P3_U2669) );
  AOI21_X1 U20176 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17022), .A(
        n17021), .ZN(n17034) );
  INV_X1 U20177 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18809) );
  OAI22_X1 U20178 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17023), .B1(
        n18809), .B2(n17039), .ZN(n17032) );
  NAND2_X1 U20179 ( .A1(n17024), .A2(n18741), .ZN(n18897) );
  OAI22_X1 U20180 ( .A1(n17026), .A2(n17325), .B1(n18897), .B2(n17025), .ZN(
        n17031) );
  OAI21_X1 U20181 ( .B1(n17325), .B2(n17042), .A(n17027), .ZN(n17326) );
  OAI22_X1 U20182 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17029), .B1(n17028), 
        .B2(n17326), .ZN(n17030) );
  NOR3_X1 U20183 ( .A1(n17032), .A2(n17031), .A3(n17030), .ZN(n17033) );
  OAI21_X1 U20184 ( .B1(n17034), .B2(n17935), .A(n17033), .ZN(P3_U2670) );
  NOR2_X1 U20185 ( .A1(n17036), .A2(n17035), .ZN(n17043) );
  AOI22_X1 U20186 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17038), .B1(n17037), 
        .B2(n18910), .ZN(n17041) );
  NAND3_X1 U20187 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18881), .A3(
        n17039), .ZN(n17040) );
  OAI211_X1 U20188 ( .C1(n17043), .C2(n17042), .A(n17041), .B(n17040), .ZN(
        P3_U2671) );
  INV_X1 U20189 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17050) );
  NOR2_X1 U20190 ( .A1(n17044), .A2(n17106), .ZN(n17046) );
  AND4_X1 U20191 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n17045)
         );
  NAND4_X1 U20192 ( .A1(n9760), .A2(n17046), .A3(n17082), .A4(n17045), .ZN(
        n17049) );
  NAND2_X1 U20193 ( .A1(n17331), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17048) );
  NAND2_X1 U20194 ( .A1(n17077), .A2(n18316), .ZN(n17047) );
  OAI22_X1 U20195 ( .A1(n17077), .A2(n17048), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17047), .ZN(P3_U2672) );
  NAND2_X1 U20196 ( .A1(n17050), .A2(n17049), .ZN(n17051) );
  NAND2_X1 U20197 ( .A1(n17051), .A2(n17318), .ZN(n17076) );
  AOI22_X1 U20198 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17063) );
  AOI22_X1 U20199 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20200 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17052) );
  OAI21_X1 U20201 ( .B1(n9779), .B2(n20889), .A(n17052), .ZN(n17059) );
  AOI22_X1 U20202 ( .A1(n15481), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20203 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20204 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20205 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17054) );
  NAND4_X1 U20206 ( .A1(n17057), .A2(n17056), .A3(n17055), .A4(n17054), .ZN(
        n17058) );
  AOI211_X1 U20207 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n17059), .B(n17058), .ZN(n17061) );
  NAND3_X1 U20208 ( .A1(n17063), .A2(n17062), .A3(n17061), .ZN(n17075) );
  AOI22_X1 U20209 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20210 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20211 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17064) );
  OAI21_X1 U20212 ( .B1(n10254), .B2(n18313), .A(n17064), .ZN(n17070) );
  AOI22_X1 U20213 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20214 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15430), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20215 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20216 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17065) );
  NAND4_X1 U20217 ( .A1(n17068), .A2(n17067), .A3(n17066), .A4(n17065), .ZN(
        n17069) );
  AOI211_X1 U20218 ( .C1(n9738), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17070), .B(n17069), .ZN(n17071) );
  AND3_X1 U20219 ( .A1(n17073), .A2(n17072), .A3(n17071), .ZN(n17079) );
  NOR3_X1 U20220 ( .A1(n17079), .A2(n17078), .A3(n17351), .ZN(n17074) );
  XNOR2_X1 U20221 ( .A(n17075), .B(n17074), .ZN(n17341) );
  OAI22_X1 U20222 ( .A1(n17077), .A2(n17076), .B1(n17341), .B2(n17318), .ZN(
        P3_U2673) );
  NOR2_X1 U20223 ( .A1(n17351), .A2(n17078), .ZN(n17080) );
  XOR2_X1 U20224 ( .A(n17080), .B(n17079), .Z(n17345) );
  NOR2_X1 U20225 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17087), .ZN(n17081) );
  AOI22_X1 U20226 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17083), .B1(n17082), 
        .B2(n17081), .ZN(n17084) );
  OAI21_X1 U20227 ( .B1(n17331), .B2(n17345), .A(n17084), .ZN(P3_U2674) );
  OAI211_X1 U20228 ( .C1(n17353), .C2(n17352), .A(n17323), .B(n17351), .ZN(
        n17085) );
  OAI221_X1 U20229 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17087), .C1(n21125), 
        .C2(n17086), .A(n17085), .ZN(P3_U2676) );
  INV_X1 U20230 ( .A(n17087), .ZN(n17090) );
  AOI21_X1 U20231 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17331), .A(n17096), .ZN(
        n17089) );
  XNOR2_X1 U20232 ( .A(n17088), .B(n17092), .ZN(n17361) );
  OAI22_X1 U20233 ( .A1(n17090), .A2(n17089), .B1(n17331), .B2(n17361), .ZN(
        P3_U2677) );
  INV_X1 U20234 ( .A(n17091), .ZN(n17099) );
  AOI21_X1 U20235 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17331), .A(n17099), .ZN(
        n17095) );
  OAI21_X1 U20236 ( .B1(n17094), .B2(n17093), .A(n17092), .ZN(n17366) );
  OAI22_X1 U20237 ( .A1(n17096), .A2(n17095), .B1(n17318), .B2(n17366), .ZN(
        P3_U2678) );
  AOI21_X1 U20238 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17331), .A(n17104), .ZN(
        n17098) );
  XNOR2_X1 U20239 ( .A(n17097), .B(n17100), .ZN(n17371) );
  OAI22_X1 U20240 ( .A1(n17099), .A2(n17098), .B1(n17331), .B2(n17371), .ZN(
        P3_U2679) );
  NOR2_X1 U20241 ( .A1(n17106), .A2(n17105), .ZN(n17119) );
  AOI21_X1 U20242 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17331), .A(n17119), .ZN(
        n17103) );
  OAI21_X1 U20243 ( .B1(n17102), .B2(n17101), .A(n17100), .ZN(n17376) );
  OAI22_X1 U20244 ( .A1(n17104), .A2(n17103), .B1(n17318), .B2(n17376), .ZN(
        P3_U2680) );
  OAI21_X1 U20245 ( .B1(n17106), .B2(n17323), .A(n17105), .ZN(n17107) );
  INV_X1 U20246 ( .A(n17107), .ZN(n17118) );
  AOI22_X1 U20247 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17274), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20248 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9741), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20249 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17238), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20250 ( .A1(n17273), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17108) );
  NAND4_X1 U20251 ( .A1(n17111), .A2(n17110), .A3(n17109), .A4(n17108), .ZN(
        n17117) );
  AOI22_X1 U20252 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20253 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20254 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20255 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17112) );
  NAND4_X1 U20256 ( .A1(n17115), .A2(n17114), .A3(n17113), .A4(n17112), .ZN(
        n17116) );
  NOR2_X1 U20257 ( .A1(n17117), .A2(n17116), .ZN(n17379) );
  OAI22_X1 U20258 ( .A1(n17119), .A2(n17118), .B1(n17379), .B2(n17331), .ZN(
        P3_U2681) );
  AOI21_X1 U20259 ( .B1(n20879), .B2(n17142), .A(n17323), .ZN(n17120) );
  INV_X1 U20260 ( .A(n17120), .ZN(n17131) );
  AOI22_X1 U20261 ( .A1(n17273), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20262 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U20263 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20264 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17121) );
  NAND4_X1 U20265 ( .A1(n17124), .A2(n17123), .A3(n17122), .A4(n17121), .ZN(
        n17130) );
  AOI22_X1 U20266 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20267 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20268 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20269 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17125) );
  NAND4_X1 U20270 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17129) );
  NOR2_X1 U20271 ( .A1(n17130), .A2(n17129), .ZN(n17386) );
  OAI22_X1 U20272 ( .A1(n9760), .A2(n17131), .B1(n17386), .B2(n17318), .ZN(
        P3_U2682) );
  AOI22_X1 U20273 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20274 ( .A1(n15460), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20275 ( .A1(n15669), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17133) );
  AOI22_X1 U20276 ( .A1(n15653), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17132) );
  NAND4_X1 U20277 ( .A1(n17135), .A2(n17134), .A3(n17133), .A4(n17132), .ZN(
        n17141) );
  AOI22_X1 U20278 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9739), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20279 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20280 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20281 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17136) );
  NAND4_X1 U20282 ( .A1(n17139), .A2(n17138), .A3(n17137), .A4(n17136), .ZN(
        n17140) );
  NOR2_X1 U20283 ( .A1(n17141), .A2(n17140), .ZN(n17391) );
  OAI21_X1 U20284 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17156), .A(n17142), .ZN(
        n17143) );
  AOI22_X1 U20285 ( .A1(n17323), .A2(n17391), .B1(n17143), .B2(n17331), .ZN(
        P3_U2683) );
  OAI21_X1 U20286 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17144), .A(n17318), .ZN(
        n17155) );
  AOI22_X1 U20287 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20288 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20289 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20290 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17145) );
  NAND4_X1 U20291 ( .A1(n17148), .A2(n17147), .A3(n17146), .A4(n17145), .ZN(
        n17154) );
  AOI22_X1 U20292 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20293 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9738), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20294 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20295 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17149) );
  NAND4_X1 U20296 ( .A1(n17152), .A2(n17151), .A3(n17150), .A4(n17149), .ZN(
        n17153) );
  NOR2_X1 U20297 ( .A1(n17154), .A2(n17153), .ZN(n17395) );
  OAI22_X1 U20298 ( .A1(n17156), .A2(n17155), .B1(n17395), .B2(n17318), .ZN(
        P3_U2684) );
  NAND2_X1 U20299 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17157), .ZN(n17170) );
  AOI22_X1 U20300 ( .A1(n15430), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20301 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20302 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20303 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17158) );
  NAND4_X1 U20304 ( .A1(n17161), .A2(n17160), .A3(n17159), .A4(n17158), .ZN(
        n17167) );
  AOI22_X1 U20305 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20306 ( .A1(n15653), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20307 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9739), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20308 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17162) );
  NAND4_X1 U20309 ( .A1(n17165), .A2(n17164), .A3(n17163), .A4(n17162), .ZN(
        n17166) );
  NOR2_X1 U20310 ( .A1(n17167), .A2(n17166), .ZN(n17400) );
  NOR2_X1 U20311 ( .A1(n17450), .A2(n17195), .ZN(n17209) );
  NAND3_X1 U20312 ( .A1(n9850), .A2(n17209), .A3(n17168), .ZN(n17169) );
  OAI221_X1 U20313 ( .B1(n17323), .B2(n17170), .C1(n17331), .C2(n17400), .A(
        n17169), .ZN(P3_U2685) );
  NAND2_X1 U20314 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17208), .ZN(n17182) );
  AOI22_X1 U20315 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20316 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n15669), .B1(
        n15460), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20317 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17286), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17290), .ZN(n17172) );
  AOI22_X1 U20318 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17267), .ZN(n17171) );
  NAND4_X1 U20319 ( .A1(n17174), .A2(n17173), .A3(n17172), .A4(n17171), .ZN(
        n17180) );
  AOI22_X1 U20320 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17275), .ZN(n17178) );
  AOI22_X1 U20321 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9741), .ZN(n17177) );
  AOI22_X1 U20322 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17289), .ZN(n17176) );
  AOI22_X1 U20323 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17175) );
  NAND4_X1 U20324 ( .A1(n17178), .A2(n17177), .A3(n17176), .A4(n17175), .ZN(
        n17179) );
  NOR2_X1 U20325 ( .A1(n17180), .A2(n17179), .ZN(n17405) );
  NAND3_X1 U20326 ( .A1(n17182), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17331), 
        .ZN(n17181) );
  OAI221_X1 U20327 ( .B1(n17182), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17318), 
        .C2(n17405), .A(n17181), .ZN(P3_U2686) );
  INV_X1 U20328 ( .A(n17182), .ZN(n17194) );
  AOI21_X1 U20329 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17331), .A(n17208), .ZN(
        n17193) );
  AOI22_X1 U20330 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U20331 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20332 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20333 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17183) );
  NAND4_X1 U20334 ( .A1(n17186), .A2(n17185), .A3(n17184), .A4(n17183), .ZN(
        n17192) );
  AOI22_X1 U20335 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9737), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20336 ( .A1(n15669), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20337 ( .A1(n15653), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20338 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17187) );
  NAND4_X1 U20339 ( .A1(n17190), .A2(n17189), .A3(n17188), .A4(n17187), .ZN(
        n17191) );
  NOR2_X1 U20340 ( .A1(n17192), .A2(n17191), .ZN(n17411) );
  OAI22_X1 U20341 ( .A1(n17194), .A2(n17193), .B1(n17411), .B2(n17318), .ZN(
        P3_U2687) );
  NOR2_X1 U20342 ( .A1(n21135), .A2(n17195), .ZN(n17222) );
  OAI21_X1 U20343 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17222), .A(n17318), .ZN(
        n17207) );
  AOI22_X1 U20344 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U20345 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17199) );
  AOI22_X1 U20346 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20347 ( .A1(n15460), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17197) );
  NAND4_X1 U20348 ( .A1(n17200), .A2(n17199), .A3(n17198), .A4(n17197), .ZN(
        n17206) );
  AOI22_X1 U20349 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20350 ( .A1(n15669), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20351 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20352 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17201) );
  NAND4_X1 U20353 ( .A1(n17204), .A2(n17203), .A3(n17202), .A4(n17201), .ZN(
        n17205) );
  NOR2_X1 U20354 ( .A1(n17206), .A2(n17205), .ZN(n17415) );
  OAI22_X1 U20355 ( .A1(n17208), .A2(n17207), .B1(n17415), .B2(n17318), .ZN(
        P3_U2688) );
  OAI21_X1 U20356 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17209), .A(n17318), .ZN(
        n17221) );
  AOI22_X1 U20357 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20358 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20359 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20360 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17210) );
  NAND4_X1 U20361 ( .A1(n17213), .A2(n17212), .A3(n17211), .A4(n17210), .ZN(
        n17220) );
  AOI22_X1 U20362 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20363 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20364 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20365 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17215) );
  NAND4_X1 U20366 ( .A1(n17218), .A2(n17217), .A3(n17216), .A4(n17215), .ZN(
        n17219) );
  NOR2_X1 U20367 ( .A1(n17220), .A2(n17219), .ZN(n17421) );
  OAI22_X1 U20368 ( .A1(n17222), .A2(n17221), .B1(n17421), .B2(n17318), .ZN(
        P3_U2689) );
  AOI22_X1 U20369 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20370 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20371 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20372 ( .A1(n9739), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17223) );
  NAND4_X1 U20373 ( .A1(n17226), .A2(n17225), .A3(n17224), .A4(n17223), .ZN(
        n17233) );
  AOI22_X1 U20374 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20375 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20376 ( .A1(n15653), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20377 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17228) );
  NAND4_X1 U20378 ( .A1(n17231), .A2(n17230), .A3(n17229), .A4(n17228), .ZN(
        n17232) );
  NOR2_X1 U20379 ( .A1(n17233), .A2(n17232), .ZN(n17429) );
  OAI21_X1 U20380 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17251), .A(n17234), .ZN(
        n17235) );
  AOI22_X1 U20381 ( .A1(n17323), .A2(n17429), .B1(n17235), .B2(n17318), .ZN(
        P3_U2691) );
  AOI21_X1 U20382 ( .B1(n17236), .B2(n17263), .A(n17323), .ZN(n17237) );
  INV_X1 U20383 ( .A(n17237), .ZN(n17250) );
  AOI22_X1 U20384 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9741), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20385 ( .A1(n17238), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20386 ( .A1(n17053), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15669), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20387 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17239), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17240) );
  NAND4_X1 U20388 ( .A1(n17243), .A2(n17242), .A3(n17241), .A4(n17240), .ZN(
        n17249) );
  AOI22_X1 U20389 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20390 ( .A1(n17289), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U20391 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U20392 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17244) );
  NAND4_X1 U20393 ( .A1(n17247), .A2(n17246), .A3(n17245), .A4(n17244), .ZN(
        n17248) );
  NOR2_X1 U20394 ( .A1(n17249), .A2(n17248), .ZN(n17433) );
  OAI22_X1 U20395 ( .A1(n17251), .A2(n17250), .B1(n17433), .B2(n17318), .ZN(
        P3_U2692) );
  AOI22_X1 U20396 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20397 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U20398 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20399 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17267), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17253) );
  NAND4_X1 U20400 ( .A1(n17256), .A2(n17255), .A3(n17254), .A4(n17253), .ZN(
        n17262) );
  AOI22_X1 U20401 ( .A1(n17298), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20402 ( .A1(n15669), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U20403 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17273), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20404 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17257) );
  NAND4_X1 U20405 ( .A1(n17260), .A2(n17259), .A3(n17258), .A4(n17257), .ZN(
        n17261) );
  NOR2_X1 U20406 ( .A1(n17262), .A2(n17261), .ZN(n17440) );
  OAI21_X1 U20407 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17283), .A(n17263), .ZN(
        n17264) );
  AOI22_X1 U20408 ( .A1(n17323), .A2(n17440), .B1(n17264), .B2(n17331), .ZN(
        P3_U2693) );
  AOI21_X1 U20409 ( .B1(n17265), .B2(n17302), .A(n17323), .ZN(n17266) );
  INV_X1 U20410 ( .A(n17266), .ZN(n17282) );
  AOI22_X1 U20411 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17286), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20412 ( .A1(n15595), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17284), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20413 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9741), .B1(
        n17298), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20414 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17267), .ZN(n17268) );
  NAND4_X1 U20415 ( .A1(n17271), .A2(n17270), .A3(n17269), .A4(n17268), .ZN(
        n17281) );
  AOI22_X1 U20416 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17238), .ZN(n17279) );
  AOI22_X1 U20417 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17273), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17289), .ZN(n17278) );
  AOI22_X1 U20418 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17214), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20419 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17275), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17274), .ZN(n17276) );
  NAND4_X1 U20420 ( .A1(n17279), .A2(n17278), .A3(n17277), .A4(n17276), .ZN(
        n17280) );
  NOR2_X1 U20421 ( .A1(n17281), .A2(n17280), .ZN(n17441) );
  OAI22_X1 U20422 ( .A1(n17283), .A2(n17282), .B1(n17441), .B2(n17318), .ZN(
        P3_U2694) );
  AOI22_X1 U20423 ( .A1(n17284), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15460), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20424 ( .A1(n17286), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17285), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20425 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17287) );
  OAI21_X1 U20426 ( .B1(n17288), .B2(n18282), .A(n17287), .ZN(n17297) );
  AOI22_X1 U20427 ( .A1(n15669), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17289), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20428 ( .A1(n17291), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U20429 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17275), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U20430 ( .A1(n17272), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17292) );
  NAND4_X1 U20431 ( .A1(n17295), .A2(n17294), .A3(n17293), .A4(n17292), .ZN(
        n17296) );
  AOI211_X1 U20432 ( .C1(n17298), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17297), .B(n17296), .ZN(n17299) );
  NAND3_X1 U20433 ( .A1(n17301), .A2(n17300), .A3(n17299), .ZN(n17446) );
  INV_X1 U20434 ( .A(n17446), .ZN(n17304) );
  OAI21_X1 U20435 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17308), .A(n17302), .ZN(
        n17303) );
  AOI22_X1 U20436 ( .A1(n17323), .A2(n17304), .B1(n17303), .B2(n17318), .ZN(
        P3_U2695) );
  AOI21_X1 U20437 ( .B1(n17305), .B2(n17309), .A(n17323), .ZN(n17306) );
  INV_X1 U20438 ( .A(n17306), .ZN(n17307) );
  INV_X1 U20439 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18321) );
  OAI22_X1 U20440 ( .A1(n17308), .A2(n17307), .B1(n18321), .B2(n17318), .ZN(
        P3_U2696) );
  OAI21_X1 U20441 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n9767), .A(n17309), .ZN(
        n17310) );
  AOI22_X1 U20442 ( .A1(n17323), .A2(n18313), .B1(n17310), .B2(n17318), .ZN(
        P3_U2697) );
  AOI21_X1 U20443 ( .B1(n17311), .B2(n17314), .A(n17323), .ZN(n17312) );
  INV_X1 U20444 ( .A(n17312), .ZN(n17313) );
  INV_X1 U20445 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18307) );
  OAI22_X1 U20446 ( .A1(n9767), .A2(n17313), .B1(n18307), .B2(n17318), .ZN(
        P3_U2698) );
  OAI21_X1 U20447 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17320), .A(n17314), .ZN(
        n17315) );
  AOI22_X1 U20448 ( .A1(n17323), .A2(n18302), .B1(n17315), .B2(n17318), .ZN(
        P3_U2699) );
  OAI22_X1 U20449 ( .A1(n17450), .A2(n17321), .B1(n17316), .B2(n17323), .ZN(
        n17317) );
  INV_X1 U20450 ( .A(n17317), .ZN(n17319) );
  INV_X1 U20451 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n21155) );
  OAI22_X1 U20452 ( .A1(n17320), .A2(n17319), .B1(n21155), .B2(n17318), .ZN(
        P3_U2700) );
  INV_X1 U20453 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18291) );
  OAI21_X1 U20454 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n9821), .A(n17321), .ZN(
        n17322) );
  AOI22_X1 U20455 ( .A1(n17323), .A2(n18291), .B1(n17322), .B2(n17318), .ZN(
        P3_U2701) );
  OAI222_X1 U20456 ( .A1(n17326), .A2(n17327), .B1(n17325), .B2(n17324), .C1(
        n18285), .C2(n17331), .ZN(P3_U2702) );
  INV_X1 U20457 ( .A(n17327), .ZN(n17329) );
  OAI21_X1 U20458 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17329), .A(n17328), .ZN(
        n17330) );
  OAI21_X1 U20459 ( .B1(n17331), .B2(n18282), .A(n17330), .ZN(P3_U2703) );
  INV_X1 U20460 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17547) );
  INV_X1 U20461 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17543) );
  INV_X1 U20462 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17587) );
  INV_X1 U20463 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17580) );
  INV_X1 U20464 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17577) );
  INV_X1 U20465 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17575) );
  INV_X1 U20466 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17573) );
  NOR4_X1 U20467 ( .A1(n17580), .A2(n17577), .A3(n17575), .A4(n17573), .ZN(
        n17417) );
  INV_X1 U20468 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17569) );
  INV_X1 U20469 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17555) );
  NAND2_X1 U20470 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17377) );
  NAND2_X1 U20471 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17368), .ZN(n17367) );
  NAND2_X1 U20472 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17346), .ZN(n17342) );
  NAND2_X1 U20473 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17338), .ZN(n17337) );
  NAND2_X1 U20474 ( .A1(n17337), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17335) );
  NAND2_X1 U20475 ( .A1(n17333), .A2(n17470), .ZN(n17378) );
  NAND2_X1 U20476 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17406), .ZN(n17334) );
  OAI221_X1 U20477 ( .B1(n17337), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17335), 
        .C2(n17470), .A(n17334), .ZN(P3_U2704) );
  AOI22_X1 U20478 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17406), .ZN(n17340) );
  OAI211_X1 U20479 ( .C1(n17338), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17465), .B(
        n17337), .ZN(n17339) );
  OAI211_X1 U20480 ( .C1(n17341), .C2(n17473), .A(n17340), .B(n17339), .ZN(
        P3_U2705) );
  AOI22_X1 U20481 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17406), .ZN(n17344) );
  OAI211_X1 U20482 ( .C1(n17346), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17465), .B(
        n17342), .ZN(n17343) );
  OAI211_X1 U20483 ( .C1(n17473), .C2(n17345), .A(n17344), .B(n17343), .ZN(
        P3_U2706) );
  AOI22_X1 U20484 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17406), .ZN(n17349) );
  AOI211_X1 U20485 ( .C1(n17547), .C2(n17354), .A(n17346), .B(n17470), .ZN(
        n17347) );
  INV_X1 U20486 ( .A(n17347), .ZN(n17348) );
  OAI211_X1 U20487 ( .C1(n17473), .C2(n17350), .A(n17349), .B(n17348), .ZN(
        P3_U2707) );
  OAI21_X1 U20488 ( .B1(n17353), .B2(n17352), .A(n17351), .ZN(n17357) );
  AOI22_X1 U20489 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17406), .ZN(n17356) );
  OAI211_X1 U20490 ( .C1(n9784), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17465), .B(
        n17354), .ZN(n17355) );
  OAI211_X1 U20491 ( .C1(n17473), .C2(n17357), .A(n17356), .B(n17355), .ZN(
        P3_U2708) );
  AOI22_X1 U20492 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17406), .ZN(n17360) );
  AOI211_X1 U20493 ( .C1(n17543), .C2(n17362), .A(n9784), .B(n17470), .ZN(
        n17358) );
  INV_X1 U20494 ( .A(n17358), .ZN(n17359) );
  OAI211_X1 U20495 ( .C1(n17473), .C2(n17361), .A(n17360), .B(n17359), .ZN(
        P3_U2709) );
  AOI22_X1 U20496 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17406), .ZN(n17365) );
  OAI211_X1 U20497 ( .C1(n17363), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17465), .B(
        n17362), .ZN(n17364) );
  OAI211_X1 U20498 ( .C1(n17473), .C2(n17366), .A(n17365), .B(n17364), .ZN(
        P3_U2710) );
  AOI22_X1 U20499 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17406), .ZN(n17370) );
  OAI211_X1 U20500 ( .C1(n17368), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17465), .B(
        n17367), .ZN(n17369) );
  OAI211_X1 U20501 ( .C1(n17371), .C2(n17473), .A(n17370), .B(n17369), .ZN(
        P3_U2711) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17406), .ZN(n17375) );
  OAI211_X1 U20503 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17373), .A(n17465), .B(
        n17372), .ZN(n17374) );
  OAI211_X1 U20504 ( .C1(n17376), .C2(n17473), .A(n17375), .B(n17374), .ZN(
        P3_U2712) );
  INV_X1 U20505 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17535) );
  INV_X1 U20506 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17533) );
  NAND2_X1 U20507 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17396), .ZN(n17392) );
  NAND2_X1 U20508 ( .A1(n17383), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17382) );
  INV_X1 U20509 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19306) );
  OAI22_X1 U20510 ( .A1(n17379), .A2(n17473), .B1(n19306), .B2(n17378), .ZN(
        n17380) );
  AOI21_X1 U20511 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17407), .A(n17380), .ZN(
        n17381) );
  OAI221_X1 U20512 ( .B1(n17383), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17382), 
        .C2(n17470), .A(n17381), .ZN(P3_U2713) );
  AOI22_X1 U20513 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17406), .ZN(n17385) );
  NOR2_X1 U20514 ( .A1(n17533), .A2(n17392), .ZN(n17387) );
  OAI211_X1 U20515 ( .C1(n17387), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17465), .B(
        n17383), .ZN(n17384) );
  OAI211_X1 U20516 ( .C1(n17386), .C2(n17473), .A(n17385), .B(n17384), .ZN(
        P3_U2714) );
  AOI22_X1 U20517 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17406), .ZN(n17390) );
  AOI211_X1 U20518 ( .C1(n17533), .C2(n17392), .A(n17387), .B(n17470), .ZN(
        n17388) );
  INV_X1 U20519 ( .A(n17388), .ZN(n17389) );
  OAI211_X1 U20520 ( .C1(n17391), .C2(n17473), .A(n17390), .B(n17389), .ZN(
        P3_U2715) );
  AOI22_X1 U20521 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17406), .ZN(n17394) );
  OAI211_X1 U20522 ( .C1(n17396), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17465), .B(
        n17392), .ZN(n17393) );
  OAI211_X1 U20523 ( .C1(n17395), .C2(n17473), .A(n17394), .B(n17393), .ZN(
        P3_U2716) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17406), .ZN(n17399) );
  INV_X1 U20525 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17529) );
  INV_X1 U20526 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17527) );
  OR2_X1 U20527 ( .A1(n17527), .A2(n17408), .ZN(n17401) );
  AOI211_X1 U20528 ( .C1(n17529), .C2(n17401), .A(n17396), .B(n17470), .ZN(
        n17397) );
  INV_X1 U20529 ( .A(n17397), .ZN(n17398) );
  OAI211_X1 U20530 ( .C1(n17400), .C2(n17473), .A(n17399), .B(n17398), .ZN(
        P3_U2717) );
  AOI22_X1 U20531 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17406), .ZN(n17404) );
  INV_X1 U20532 ( .A(n17408), .ZN(n17402) );
  OAI211_X1 U20533 ( .C1(n17402), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17465), .B(
        n17401), .ZN(n17403) );
  OAI211_X1 U20534 ( .C1(n17405), .C2(n17473), .A(n17404), .B(n17403), .ZN(
        P3_U2718) );
  AOI22_X1 U20535 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17407), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17406), .ZN(n17410) );
  OAI211_X1 U20536 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17412), .A(n17465), .B(
        n17408), .ZN(n17409) );
  OAI211_X1 U20537 ( .C1(n17411), .C2(n17473), .A(n17410), .B(n17409), .ZN(
        P3_U2719) );
  AOI211_X1 U20538 ( .C1(n17587), .C2(n17418), .A(n17470), .B(n17412), .ZN(
        n17413) );
  AOI21_X1 U20539 ( .B1(n17478), .B2(BUF2_REG_15__SCAN_IN), .A(n17413), .ZN(
        n17414) );
  OAI21_X1 U20540 ( .B1(n17415), .B2(n17473), .A(n17414), .ZN(P3_U2720) );
  NAND3_X1 U20541 ( .A1(n18316), .A2(P3_EAX_REG_9__SCAN_IN), .A3(n9754), .ZN(
        n17437) );
  NOR2_X1 U20542 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17437), .ZN(n17416) );
  AOI22_X1 U20543 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17478), .B1(n17417), .B2(
        n17416), .ZN(n17420) );
  NAND3_X1 U20544 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17465), .A3(n17418), 
        .ZN(n17419) );
  OAI211_X1 U20545 ( .C1(n17421), .C2(n17473), .A(n17420), .B(n17419), .ZN(
        P3_U2721) );
  NAND2_X1 U20546 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n17422) );
  NOR2_X1 U20547 ( .A1(n17422), .A2(n17437), .ZN(n17435) );
  NAND2_X1 U20548 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17435), .ZN(n17428) );
  NAND2_X1 U20549 ( .A1(n17428), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17427) );
  OAI22_X1 U20550 ( .A1(n17424), .A2(n17476), .B1(n17473), .B2(n17423), .ZN(
        n17425) );
  INV_X1 U20551 ( .A(n17425), .ZN(n17426) );
  OAI221_X1 U20552 ( .B1(n17428), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17427), 
        .C2(n17470), .A(n17426), .ZN(P3_U2722) );
  INV_X1 U20553 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17432) );
  INV_X1 U20554 ( .A(n17428), .ZN(n17431) );
  AOI21_X1 U20555 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17465), .A(n17435), .ZN(
        n17430) );
  OAI222_X1 U20556 ( .A1(n17476), .A2(n17432), .B1(n17431), .B2(n17430), .C1(
        n17473), .C2(n17429), .ZN(P3_U2723) );
  INV_X1 U20557 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17436) );
  INV_X1 U20558 ( .A(n17437), .ZN(n17443) );
  AOI22_X1 U20559 ( .A1(n17443), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n17465), .ZN(n17434) );
  OAI222_X1 U20560 ( .A1(n17476), .A2(n17436), .B1(n17435), .B2(n17434), .C1(
        n17473), .C2(n17433), .ZN(P3_U2724) );
  AOI221_X1 U20561 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n17443), .C1(n17573), 
        .C2(n17437), .A(n17470), .ZN(n17438) );
  AOI21_X1 U20562 ( .B1(n17478), .B2(BUF2_REG_10__SCAN_IN), .A(n17438), .ZN(
        n17439) );
  OAI21_X1 U20563 ( .B1(n17440), .B2(n17473), .A(n17439), .ZN(P3_U2725) );
  INV_X1 U20564 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20565 ( .A1(n18316), .A2(n9754), .B1(P3_EAX_REG_9__SCAN_IN), .B2(
        n17465), .ZN(n17442) );
  OAI222_X1 U20566 ( .A1(n17476), .A2(n17444), .B1(n17443), .B2(n17442), .C1(
        n17473), .C2(n17441), .ZN(P3_U2726) );
  NOR2_X1 U20567 ( .A1(n17450), .A2(n17445), .ZN(n17453) );
  AOI21_X1 U20568 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17465), .A(n17453), .ZN(
        n17449) );
  AOI22_X1 U20569 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17478), .B1(n17447), .B2(
        n17446), .ZN(n17448) );
  OAI21_X1 U20570 ( .B1(n9754), .B2(n17449), .A(n17448), .ZN(P3_U2727) );
  INV_X1 U20571 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20954) );
  INV_X1 U20572 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17565) );
  INV_X1 U20573 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17561) );
  INV_X1 U20574 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17557) );
  NOR3_X1 U20575 ( .A1(n17450), .A2(n17479), .A3(n17553), .ZN(n17477) );
  NAND2_X1 U20576 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17477), .ZN(n17469) );
  NAND2_X1 U20577 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17475), .ZN(n17461) );
  NAND2_X1 U20578 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17464), .ZN(n17454) );
  NOR2_X1 U20579 ( .A1(n17565), .A2(n17454), .ZN(n17457) );
  AOI21_X1 U20580 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17465), .A(n17457), .ZN(
        n17452) );
  OAI222_X1 U20581 ( .A1(n17476), .A2(n20954), .B1(n17453), .B2(n17452), .C1(
        n17473), .C2(n17451), .ZN(P3_U2728) );
  INV_X1 U20582 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18309) );
  INV_X1 U20583 ( .A(n17454), .ZN(n17460) );
  AOI21_X1 U20584 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17465), .A(n17460), .ZN(
        n17456) );
  OAI222_X1 U20585 ( .A1(n18309), .A2(n17476), .B1(n17457), .B2(n17456), .C1(
        n17473), .C2(n17455), .ZN(P3_U2729) );
  INV_X1 U20586 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21139) );
  AOI21_X1 U20587 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17465), .A(n17464), .ZN(
        n17459) );
  OAI222_X1 U20588 ( .A1(n21139), .A2(n17476), .B1(n17460), .B2(n17459), .C1(
        n17473), .C2(n17458), .ZN(P3_U2730) );
  INV_X1 U20589 ( .A(n17461), .ZN(n17468) );
  AOI21_X1 U20590 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17465), .A(n17468), .ZN(
        n17463) );
  OAI222_X1 U20591 ( .A1(n18297), .A2(n17476), .B1(n17464), .B2(n17463), .C1(
        n17473), .C2(n17462), .ZN(P3_U2731) );
  INV_X1 U20592 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18293) );
  AOI21_X1 U20593 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17465), .A(n17475), .ZN(
        n17467) );
  OAI222_X1 U20594 ( .A1(n18293), .A2(n17476), .B1(n17468), .B2(n17467), .C1(
        n17473), .C2(n17466), .ZN(P3_U2732) );
  INV_X1 U20595 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18286) );
  OAI21_X1 U20596 ( .B1(n17557), .B2(n17470), .A(n17469), .ZN(n17471) );
  INV_X1 U20597 ( .A(n17471), .ZN(n17474) );
  OAI222_X1 U20598 ( .A1(n18286), .A2(n17476), .B1(n17475), .B2(n17474), .C1(
        n17473), .C2(n17472), .ZN(P3_U2733) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17478), .B1(n17477), .B2(
        n17555), .ZN(n17481) );
  OAI221_X1 U20600 ( .B1(n17479), .B2(n18316), .C1(n17479), .C2(n17553), .A(
        P3_EAX_REG_1__SCAN_IN), .ZN(n17480) );
  OAI211_X1 U20601 ( .C1(n17482), .C2(n17473), .A(n17481), .B(n17480), .ZN(
        P3_U2734) );
  NAND2_X1 U20602 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17709), .ZN(n18927) );
  INV_X2 U20603 ( .A(n18927), .ZN(n17519) );
  NOR2_X4 U20604 ( .A1(n17519), .A2(n17503), .ZN(n17500) );
  AND2_X1 U20605 ( .A1(n17500), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20606 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17551) );
  NAND2_X1 U20607 ( .A1(n17503), .A2(n17485), .ZN(n17502) );
  AOI22_X1 U20608 ( .A1(n17519), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17500), .ZN(n17486) );
  OAI21_X1 U20609 ( .B1(n17551), .B2(n17502), .A(n17486), .ZN(P3_U2737) );
  INV_X1 U20610 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17549) );
  AOI22_X1 U20611 ( .A1(n17519), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17487) );
  OAI21_X1 U20612 ( .B1(n17549), .B2(n17502), .A(n17487), .ZN(P3_U2738) );
  AOI22_X1 U20613 ( .A1(n17519), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17488) );
  OAI21_X1 U20614 ( .B1(n17547), .B2(n17502), .A(n17488), .ZN(P3_U2739) );
  INV_X1 U20615 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n21119) );
  AOI22_X1 U20616 ( .A1(n17519), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17489) );
  OAI21_X1 U20617 ( .B1(n21119), .B2(n17502), .A(n17489), .ZN(P3_U2740) );
  AOI22_X1 U20618 ( .A1(n17519), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17490) );
  OAI21_X1 U20619 ( .B1(n17543), .B2(n17502), .A(n17490), .ZN(P3_U2741) );
  AOI22_X1 U20620 ( .A1(n17519), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17491) );
  OAI21_X1 U20621 ( .B1(n9999), .B2(n17502), .A(n17491), .ZN(P3_U2742) );
  INV_X1 U20622 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17540) );
  AOI22_X1 U20623 ( .A1(n17519), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17492) );
  OAI21_X1 U20624 ( .B1(n17540), .B2(n17502), .A(n17492), .ZN(P3_U2743) );
  INV_X1 U20625 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20861) );
  AOI22_X1 U20626 ( .A1(n17519), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17493) );
  OAI21_X1 U20627 ( .B1(n20861), .B2(n17502), .A(n17493), .ZN(P3_U2744) );
  INV_X1 U20628 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U20629 ( .A1(n17519), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17494) );
  OAI21_X1 U20630 ( .B1(n17537), .B2(n17502), .A(n17494), .ZN(P3_U2745) );
  AOI22_X1 U20631 ( .A1(n17519), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17495) );
  OAI21_X1 U20632 ( .B1(n17535), .B2(n17502), .A(n17495), .ZN(P3_U2746) );
  AOI22_X1 U20633 ( .A1(n17519), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17496) );
  OAI21_X1 U20634 ( .B1(n17533), .B2(n17502), .A(n17496), .ZN(P3_U2747) );
  INV_X1 U20635 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20636 ( .A1(n17519), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17497) );
  OAI21_X1 U20637 ( .B1(n17531), .B2(n17502), .A(n17497), .ZN(P3_U2748) );
  AOI22_X1 U20638 ( .A1(n17519), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17498) );
  OAI21_X1 U20639 ( .B1(n17529), .B2(n17502), .A(n17498), .ZN(P3_U2749) );
  AOI22_X1 U20640 ( .A1(n17519), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17499) );
  OAI21_X1 U20641 ( .B1(n17527), .B2(n17502), .A(n17499), .ZN(P3_U2750) );
  INV_X1 U20642 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20643 ( .A1(n17519), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17501) );
  OAI21_X1 U20644 ( .B1(n17525), .B2(n17502), .A(n17501), .ZN(P3_U2751) );
  AOI22_X1 U20645 ( .A1(n17519), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17504) );
  OAI21_X1 U20646 ( .B1(n17587), .B2(n17521), .A(n17504), .ZN(P3_U2752) );
  INV_X1 U20647 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17582) );
  AOI22_X1 U20648 ( .A1(n17519), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17505) );
  OAI21_X1 U20649 ( .B1(n17582), .B2(n17521), .A(n17505), .ZN(P3_U2753) );
  AOI22_X1 U20650 ( .A1(n17519), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17506) );
  OAI21_X1 U20651 ( .B1(n17580), .B2(n17521), .A(n17506), .ZN(P3_U2754) );
  AOI22_X1 U20652 ( .A1(n17519), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17507) );
  OAI21_X1 U20653 ( .B1(n17577), .B2(n17521), .A(n17507), .ZN(P3_U2755) );
  AOI22_X1 U20654 ( .A1(n17519), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17508) );
  OAI21_X1 U20655 ( .B1(n17575), .B2(n17521), .A(n17508), .ZN(P3_U2756) );
  AOI22_X1 U20656 ( .A1(n17519), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17509) );
  OAI21_X1 U20657 ( .B1(n17573), .B2(n17521), .A(n17509), .ZN(P3_U2757) );
  INV_X1 U20658 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17571) );
  AOI22_X1 U20659 ( .A1(n17519), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17510) );
  OAI21_X1 U20660 ( .B1(n17571), .B2(n17521), .A(n17510), .ZN(P3_U2758) );
  AOI22_X1 U20661 ( .A1(n17519), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17511) );
  OAI21_X1 U20662 ( .B1(n17569), .B2(n17521), .A(n17511), .ZN(P3_U2759) );
  INV_X1 U20663 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17567) );
  AOI22_X1 U20664 ( .A1(n17519), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17512) );
  OAI21_X1 U20665 ( .B1(n17567), .B2(n17521), .A(n17512), .ZN(P3_U2760) );
  AOI22_X1 U20666 ( .A1(n17519), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17513) );
  OAI21_X1 U20667 ( .B1(n17565), .B2(n17521), .A(n17513), .ZN(P3_U2761) );
  INV_X1 U20668 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17563) );
  AOI22_X1 U20669 ( .A1(n17519), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17514) );
  OAI21_X1 U20670 ( .B1(n17563), .B2(n17521), .A(n17514), .ZN(P3_U2762) );
  AOI22_X1 U20671 ( .A1(n17519), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17515) );
  OAI21_X1 U20672 ( .B1(n17561), .B2(n17521), .A(n17515), .ZN(P3_U2763) );
  INV_X1 U20673 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17559) );
  AOI22_X1 U20674 ( .A1(n17519), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17516) );
  OAI21_X1 U20675 ( .B1(n17559), .B2(n17521), .A(n17516), .ZN(P3_U2764) );
  AOI22_X1 U20676 ( .A1(n17519), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17517) );
  OAI21_X1 U20677 ( .B1(n17557), .B2(n17521), .A(n17517), .ZN(P3_U2765) );
  AOI22_X1 U20678 ( .A1(n17519), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17518) );
  OAI21_X1 U20679 ( .B1(n17555), .B2(n17521), .A(n17518), .ZN(P3_U2766) );
  AOI22_X1 U20680 ( .A1(n17519), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17500), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17520) );
  OAI21_X1 U20681 ( .B1(n17553), .B2(n17521), .A(n17520), .ZN(P3_U2767) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17584), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17583), .ZN(n17524) );
  OAI21_X1 U20683 ( .B1(n17525), .B2(n17586), .A(n17524), .ZN(P3_U2768) );
  AOI22_X1 U20684 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17583), .ZN(n17526) );
  OAI21_X1 U20685 ( .B1(n17527), .B2(n17586), .A(n17526), .ZN(P3_U2769) );
  AOI22_X1 U20686 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17583), .ZN(n17528) );
  OAI21_X1 U20687 ( .B1(n17529), .B2(n17586), .A(n17528), .ZN(P3_U2770) );
  AOI22_X1 U20688 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17583), .ZN(n17530) );
  OAI21_X1 U20689 ( .B1(n17531), .B2(n17586), .A(n17530), .ZN(P3_U2771) );
  AOI22_X1 U20690 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17583), .ZN(n17532) );
  OAI21_X1 U20691 ( .B1(n17533), .B2(n17586), .A(n17532), .ZN(P3_U2772) );
  AOI22_X1 U20692 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17583), .ZN(n17534) );
  OAI21_X1 U20693 ( .B1(n17535), .B2(n17586), .A(n17534), .ZN(P3_U2773) );
  AOI22_X1 U20694 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17583), .ZN(n17536) );
  OAI21_X1 U20695 ( .B1(n17537), .B2(n17586), .A(n17536), .ZN(P3_U2774) );
  AOI22_X1 U20696 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17583), .ZN(n17538) );
  OAI21_X1 U20697 ( .B1(n20861), .B2(n17586), .A(n17538), .ZN(P3_U2775) );
  AOI22_X1 U20698 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17583), .ZN(n17539) );
  OAI21_X1 U20699 ( .B1(n17540), .B2(n17586), .A(n17539), .ZN(P3_U2776) );
  AOI22_X1 U20700 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17583), .ZN(n17541) );
  OAI21_X1 U20701 ( .B1(n9999), .B2(n17586), .A(n17541), .ZN(P3_U2777) );
  AOI22_X1 U20702 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17583), .ZN(n17542) );
  OAI21_X1 U20703 ( .B1(n17543), .B2(n17586), .A(n17542), .ZN(P3_U2778) );
  AOI22_X1 U20704 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17544), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17583), .ZN(n17545) );
  OAI21_X1 U20705 ( .B1(n21119), .B2(n17586), .A(n17545), .ZN(P3_U2779) );
  AOI22_X1 U20706 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17584), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17583), .ZN(n17546) );
  OAI21_X1 U20707 ( .B1(n17547), .B2(n17586), .A(n17546), .ZN(P3_U2780) );
  AOI22_X1 U20708 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17584), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17583), .ZN(n17548) );
  OAI21_X1 U20709 ( .B1(n17549), .B2(n17586), .A(n17548), .ZN(P3_U2781) );
  AOI22_X1 U20710 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17584), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17583), .ZN(n17550) );
  OAI21_X1 U20711 ( .B1(n17551), .B2(n17586), .A(n17550), .ZN(P3_U2782) );
  AOI22_X1 U20712 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17583), .ZN(n17552) );
  OAI21_X1 U20713 ( .B1(n17553), .B2(n17586), .A(n17552), .ZN(P3_U2783) );
  AOI22_X1 U20714 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17583), .ZN(n17554) );
  OAI21_X1 U20715 ( .B1(n17555), .B2(n17586), .A(n17554), .ZN(P3_U2784) );
  AOI22_X1 U20716 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17583), .ZN(n17556) );
  OAI21_X1 U20717 ( .B1(n17557), .B2(n17586), .A(n17556), .ZN(P3_U2785) );
  AOI22_X1 U20718 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17583), .ZN(n17558) );
  OAI21_X1 U20719 ( .B1(n17559), .B2(n17586), .A(n17558), .ZN(P3_U2786) );
  AOI22_X1 U20720 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17578), .ZN(n17560) );
  OAI21_X1 U20721 ( .B1(n17561), .B2(n17586), .A(n17560), .ZN(P3_U2787) );
  AOI22_X1 U20722 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17578), .ZN(n17562) );
  OAI21_X1 U20723 ( .B1(n17563), .B2(n17586), .A(n17562), .ZN(P3_U2788) );
  AOI22_X1 U20724 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17578), .ZN(n17564) );
  OAI21_X1 U20725 ( .B1(n17565), .B2(n17586), .A(n17564), .ZN(P3_U2789) );
  AOI22_X1 U20726 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17578), .ZN(n17566) );
  OAI21_X1 U20727 ( .B1(n17567), .B2(n17586), .A(n17566), .ZN(P3_U2790) );
  AOI22_X1 U20728 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17578), .ZN(n17568) );
  OAI21_X1 U20729 ( .B1(n17569), .B2(n17586), .A(n17568), .ZN(P3_U2791) );
  AOI22_X1 U20730 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17578), .ZN(n17570) );
  OAI21_X1 U20731 ( .B1(n17571), .B2(n17586), .A(n17570), .ZN(P3_U2792) );
  AOI22_X1 U20732 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17578), .ZN(n17572) );
  OAI21_X1 U20733 ( .B1(n17573), .B2(n17586), .A(n17572), .ZN(P3_U2793) );
  AOI22_X1 U20734 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17578), .ZN(n17574) );
  OAI21_X1 U20735 ( .B1(n17575), .B2(n17586), .A(n17574), .ZN(P3_U2794) );
  AOI22_X1 U20736 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17578), .ZN(n17576) );
  OAI21_X1 U20737 ( .B1(n17577), .B2(n17586), .A(n17576), .ZN(P3_U2795) );
  AOI22_X1 U20738 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17578), .ZN(n17579) );
  OAI21_X1 U20739 ( .B1(n17580), .B2(n17586), .A(n17579), .ZN(P3_U2796) );
  AOI22_X1 U20740 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17583), .ZN(n17581) );
  OAI21_X1 U20741 ( .B1(n17582), .B2(n17586), .A(n17581), .ZN(P3_U2797) );
  AOI22_X1 U20742 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17584), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17583), .ZN(n17585) );
  OAI21_X1 U20743 ( .B1(n17587), .B2(n17586), .A(n17585), .ZN(P3_U2798) );
  OAI21_X1 U20744 ( .B1(n17602), .B2(n17781), .A(n17940), .ZN(n17588) );
  AOI21_X1 U20745 ( .B1(n17709), .B2(n17589), .A(n17588), .ZN(n17622) );
  OAI21_X1 U20746 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17694), .A(
        n17622), .ZN(n17612) );
  AOI22_X1 U20747 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17612), .B1(
        n17801), .B2(n17590), .ZN(n17607) );
  AOI21_X1 U20748 ( .B1(n17593), .B2(n17592), .A(n17591), .ZN(n17601) );
  INV_X1 U20749 ( .A(n17594), .ZN(n17595) );
  NAND2_X1 U20750 ( .A1(n17595), .A2(n17719), .ZN(n17665) );
  NOR4_X1 U20751 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17596), .A3(
        n17953), .A4(n17665), .ZN(n17600) );
  NOR2_X1 U20752 ( .A1(n9734), .A2(n17777), .ZN(n17701) );
  OAI22_X1 U20753 ( .A1(n17945), .A2(n16499), .B1(n17946), .B2(n17944), .ZN(
        n17627) );
  NOR2_X1 U20754 ( .A1(n17953), .A2(n17627), .ZN(n17598) );
  NOR3_X1 U20755 ( .A1(n17701), .A2(n17598), .A3(n17597), .ZN(n17599) );
  AOI211_X1 U20756 ( .C1(n17857), .C2(n17601), .A(n17600), .B(n17599), .ZN(
        n17606) );
  NAND2_X1 U20757 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18255), .ZN(n17605) );
  AND2_X1 U20758 ( .A1(n17602), .A2(n17746), .ZN(n17614) );
  NAND2_X1 U20759 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17603) );
  OAI211_X1 U20760 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17614), .B(n17603), .ZN(n17604) );
  NAND4_X1 U20761 ( .A1(n17607), .A2(n17606), .A3(n17605), .A4(n17604), .ZN(
        P3_U2802) );
  AOI21_X1 U20762 ( .B1(n17792), .B2(n17609), .A(n17608), .ZN(n17958) );
  OAI22_X1 U20763 ( .A1(n18148), .A2(n21014), .B1(n17786), .B2(n17610), .ZN(
        n17611) );
  AOI221_X1 U20764 ( .B1(n17614), .B2(n17613), .C1(n17612), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17611), .ZN(n17618) );
  NOR2_X1 U20765 ( .A1(n17615), .A2(n17755), .ZN(n17616) );
  AOI22_X1 U20766 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17627), .B1(
        n17616), .B2(n17953), .ZN(n17617) );
  OAI211_X1 U20767 ( .C1(n17958), .C2(n17844), .A(n17618), .B(n17617), .ZN(
        P3_U2803) );
  INV_X1 U20768 ( .A(n17619), .ZN(n17620) );
  AOI21_X1 U20769 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17621), .A(
        n17620), .ZN(n17965) );
  NAND2_X1 U20770 ( .A1(n17786), .A2(n17694), .ZN(n17934) );
  NOR2_X1 U20771 ( .A1(n18148), .A2(n18857), .ZN(n17960) );
  AOI221_X1 U20772 ( .B1(n18365), .B2(n20970), .C1(n17623), .C2(n20970), .A(
        n17622), .ZN(n17624) );
  AOI211_X1 U20773 ( .C1(n17625), .C2(n17934), .A(n17960), .B(n17624), .ZN(
        n17629) );
  NOR3_X1 U20774 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17626), .A3(
        n17986), .ZN(n17961) );
  NOR2_X1 U20775 ( .A1(n17959), .A2(n17755), .ZN(n17652) );
  AOI22_X1 U20776 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17627), .B1(
        n17961), .B2(n17652), .ZN(n17628) );
  OAI211_X1 U20777 ( .C1(n17965), .C2(n17844), .A(n17629), .B(n17628), .ZN(
        P3_U2804) );
  NOR2_X1 U20778 ( .A1(n17986), .A2(n17959), .ZN(n17969) );
  NAND2_X1 U20779 ( .A1(n18001), .A2(n17969), .ZN(n17630) );
  XOR2_X1 U20780 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17630), .Z(
        n17973) );
  OAI21_X1 U20781 ( .B1(n17631), .B2(n18791), .A(n17940), .ZN(n17632) );
  AOI21_X1 U20782 ( .B1(n18662), .B2(n17633), .A(n17632), .ZN(n17660) );
  OAI21_X1 U20783 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17694), .A(
        n17660), .ZN(n17648) );
  NOR2_X1 U20784 ( .A1(n17712), .A2(n17633), .ZN(n17649) );
  OAI211_X1 U20785 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17649), .B(n17634), .ZN(n17635) );
  NAND2_X1 U20786 ( .A1(n18255), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17971) );
  OAI211_X1 U20787 ( .C1(n17786), .C2(n17636), .A(n17635), .B(n17971), .ZN(
        n17642) );
  INV_X1 U20788 ( .A(n18079), .ZN(n18000) );
  NAND2_X1 U20789 ( .A1(n18000), .A2(n17969), .ZN(n17637) );
  XOR2_X1 U20790 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17637), .Z(
        n17978) );
  OAI21_X1 U20791 ( .B1(n17792), .B2(n17639), .A(n17638), .ZN(n17640) );
  XOR2_X1 U20792 ( .A(n17640), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17974) );
  OAI22_X1 U20793 ( .A1(n16499), .A2(n17978), .B1(n17844), .B2(n17974), .ZN(
        n17641) );
  AOI211_X1 U20794 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17648), .A(
        n17642), .B(n17641), .ZN(n17643) );
  OAI21_X1 U20795 ( .B1(n17944), .B2(n17973), .A(n17643), .ZN(P3_U2805) );
  NAND2_X1 U20796 ( .A1(n18001), .A2(n17644), .ZN(n17980) );
  NOR2_X1 U20797 ( .A1(n18079), .A2(n17959), .ZN(n17982) );
  INV_X1 U20798 ( .A(n17982), .ZN(n17645) );
  AOI22_X1 U20799 ( .A1(n9734), .A2(n17980), .B1(n17777), .B2(n17645), .ZN(
        n17664) );
  OAI22_X1 U20800 ( .A1(n18148), .A2(n18853), .B1(n17786), .B2(n17646), .ZN(
        n17647) );
  AOI221_X1 U20801 ( .B1(n17649), .B2(n21112), .C1(n17648), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17647), .ZN(n17654) );
  OAI21_X1 U20802 ( .B1(n17651), .B2(n17986), .A(n17650), .ZN(n17988) );
  AOI22_X1 U20803 ( .A1(n17857), .A2(n17988), .B1(n17652), .B2(n17986), .ZN(
        n17653) );
  OAI211_X1 U20804 ( .C1(n17664), .C2(n17986), .A(n17654), .B(n17653), .ZN(
        P3_U2806) );
  OAI22_X1 U20805 ( .A1(n17856), .A2(n17950), .B1(n17666), .B2(n17655), .ZN(
        n17656) );
  NOR2_X1 U20806 ( .A1(n17656), .A2(n17691), .ZN(n17657) );
  XOR2_X1 U20807 ( .A(n17657), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n17995) );
  NOR2_X1 U20808 ( .A1(n18148), .A2(n18852), .ZN(n17994) );
  AOI21_X1 U20809 ( .B1(n17658), .B2(n18662), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17659) );
  OAI22_X1 U20810 ( .A1(n17919), .A2(n17661), .B1(n17660), .B2(n17659), .ZN(
        n17662) );
  AOI211_X1 U20811 ( .C1(n17995), .C2(n17857), .A(n17994), .B(n17662), .ZN(
        n17663) );
  OAI221_X1 U20812 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17665), 
        .C1(n17998), .C2(n17664), .A(n17663), .ZN(P3_U2807) );
  INV_X1 U20813 ( .A(n17666), .ZN(n17667) );
  AOI221_X1 U20814 ( .B1(n17742), .B2(n17667), .C1(n18005), .C2(n17667), .A(
        n17691), .ZN(n17668) );
  XOR2_X1 U20815 ( .A(n17950), .B(n17668), .Z(n18017) );
  NOR2_X1 U20816 ( .A1(n18005), .A2(n17755), .ZN(n17678) );
  AOI22_X1 U20817 ( .A1(n17777), .A2(n18079), .B1(n9734), .B2(n18090), .ZN(
        n17754) );
  OAI21_X1 U20818 ( .B1(n18010), .B2(n17701), .A(n17754), .ZN(n17688) );
  INV_X1 U20819 ( .A(n17672), .ZN(n17670) );
  OAI22_X1 U20820 ( .A1(n17670), .A2(n17781), .B1(n17669), .B2(n18791), .ZN(
        n17671) );
  NOR2_X1 U20821 ( .A1(n17889), .A2(n17671), .ZN(n17697) );
  OAI21_X1 U20822 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17694), .A(
        n17697), .ZN(n17685) );
  AOI22_X1 U20823 ( .A1(n18255), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17685), .ZN(n17675) );
  NOR2_X1 U20824 ( .A1(n17712), .A2(n17672), .ZN(n17687) );
  OAI211_X1 U20825 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17687), .B(n17673), .ZN(n17674) );
  OAI211_X1 U20826 ( .C1(n17676), .C2(n17786), .A(n17675), .B(n17674), .ZN(
        n17677) );
  AOI221_X1 U20827 ( .B1(n17678), .B2(n17950), .C1(n17688), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17677), .ZN(n17679) );
  OAI21_X1 U20828 ( .B1(n17844), .B2(n18017), .A(n17679), .ZN(P3_U2808) );
  NAND3_X1 U20829 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17856), .A3(
        n17680), .ZN(n17704) );
  INV_X1 U20830 ( .A(n17722), .ZN(n17705) );
  OAI22_X1 U20831 ( .A1(n18023), .A2(n17704), .B1(n17681), .B2(n17705), .ZN(
        n17682) );
  XOR2_X1 U20832 ( .A(n18024), .B(n17682), .Z(n18031) );
  OAI22_X1 U20833 ( .A1(n18148), .A2(n18847), .B1(n17786), .B2(n17683), .ZN(
        n17684) );
  AOI221_X1 U20834 ( .B1(n17687), .B2(n17686), .C1(n17685), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17684), .ZN(n17690) );
  NOR2_X1 U20835 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18023), .ZN(
        n18028) );
  AOI22_X1 U20836 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17688), .B1(
        n17719), .B2(n18028), .ZN(n17689) );
  OAI211_X1 U20837 ( .C1(n18031), .C2(n17844), .A(n17690), .B(n17689), .ZN(
        P3_U2809) );
  INV_X1 U20838 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18046) );
  AOI221_X1 U20839 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17704), 
        .C1(n18046), .C2(n17721), .A(n17691), .ZN(n17692) );
  XOR2_X1 U20840 ( .A(n18006), .B(n17692), .Z(n18039) );
  INV_X1 U20841 ( .A(n17693), .ZN(n17699) );
  AOI21_X1 U20842 ( .B1(n17695), .B2(n18662), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17696) );
  OAI22_X1 U20843 ( .A1(n17697), .A2(n17696), .B1(n18148), .B2(n21120), .ZN(
        n17698) );
  AOI221_X1 U20844 ( .B1(n17801), .B2(n17699), .C1(n16488), .C2(n17699), .A(
        n17698), .ZN(n17703) );
  NAND2_X1 U20845 ( .A1(n17700), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18032) );
  INV_X1 U20846 ( .A(n18032), .ZN(n18002) );
  OAI21_X1 U20847 ( .B1(n17701), .B2(n18002), .A(n17754), .ZN(n17718) );
  NOR2_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18046), .ZN(
        n18035) );
  AOI22_X1 U20849 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17718), .B1(
        n17719), .B2(n18035), .ZN(n17702) );
  OAI211_X1 U20850 ( .C1(n17844), .C2(n18039), .A(n17703), .B(n17702), .ZN(
        P3_U2810) );
  OAI21_X1 U20851 ( .B1(n17705), .B2(n17721), .A(n17704), .ZN(n17706) );
  XOR2_X1 U20852 ( .A(n17706), .B(n18046), .Z(n18040) );
  AOI21_X1 U20853 ( .B1(n17711), .B2(n17850), .A(n17889), .ZN(n17707) );
  INV_X1 U20854 ( .A(n17707), .ZN(n17734) );
  AOI21_X1 U20855 ( .B1(n17709), .B2(n17708), .A(n17734), .ZN(n17725) );
  AOI22_X1 U20856 ( .A1(n18255), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n17801), 
        .B2(n17710), .ZN(n17715) );
  NOR2_X1 U20857 ( .A1(n17712), .A2(n17711), .ZN(n17727) );
  OAI211_X1 U20858 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17727), .B(n17713), .ZN(n17714) );
  OAI211_X1 U20859 ( .C1(n17725), .C2(n17716), .A(n17715), .B(n17714), .ZN(
        n17717) );
  AOI221_X1 U20860 ( .B1(n17719), .B2(n18046), .C1(n17718), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17717), .ZN(n17720) );
  OAI21_X1 U20861 ( .B1(n18040), .B2(n17844), .A(n17720), .ZN(P3_U2811) );
  OAI21_X1 U20862 ( .B1(n17792), .B2(n21129), .A(n17721), .ZN(n17723) );
  XOR2_X1 U20863 ( .A(n17723), .B(n17722), .Z(n18061) );
  NOR2_X1 U20864 ( .A1(n18148), .A2(n18842), .ZN(n18049) );
  OAI22_X1 U20865 ( .A1(n17725), .A2(n20971), .B1(n17786), .B2(n17724), .ZN(
        n17726) );
  AOI211_X1 U20866 ( .C1(n17727), .C2(n20971), .A(n18049), .B(n17726), .ZN(
        n17731) );
  OAI21_X1 U20867 ( .B1(n17728), .B2(n17755), .A(n17754), .ZN(n17740) );
  NOR2_X1 U20868 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18054), .ZN(
        n18050) );
  AOI22_X1 U20869 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17740), .B1(
        n17729), .B2(n18050), .ZN(n17730) );
  OAI211_X1 U20870 ( .C1(n17844), .C2(n18061), .A(n17731), .B(n17730), .ZN(
        P3_U2812) );
  AOI21_X1 U20871 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17733), .A(
        n17732), .ZN(n18067) );
  NOR3_X1 U20872 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18074), .A3(
        n17755), .ZN(n17739) );
  NAND2_X1 U20873 ( .A1(n18255), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18065) );
  OAI221_X1 U20874 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18662), .C1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n17735), .A(n17734), .ZN(
        n17736) );
  OAI211_X1 U20875 ( .C1(n17919), .C2(n17737), .A(n18065), .B(n17736), .ZN(
        n17738) );
  AOI211_X1 U20876 ( .C1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17740), .A(
        n17739), .B(n17738), .ZN(n17741) );
  OAI21_X1 U20877 ( .B1(n18067), .B2(n17844), .A(n17741), .ZN(P3_U2813) );
  INV_X1 U20878 ( .A(n17845), .ZN(n17790) );
  NAND2_X1 U20879 ( .A1(n17856), .A2(n17790), .ZN(n17822) );
  INV_X1 U20880 ( .A(n17822), .ZN(n17832) );
  AOI22_X1 U20881 ( .A1(n18048), .A2(n17832), .B1(n17742), .B2(n17792), .ZN(
        n17743) );
  XOR2_X1 U20882 ( .A(n18074), .B(n17743), .Z(n18076) );
  AOI21_X1 U20883 ( .B1(n17850), .B2(n17744), .A(n17889), .ZN(n17769) );
  OAI21_X1 U20884 ( .B1(n17745), .B2(n18791), .A(n17769), .ZN(n17758) );
  AOI22_X1 U20885 ( .A1(n18255), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17758), .ZN(n17750) );
  NAND2_X1 U20886 ( .A1(n17780), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17747) );
  NAND2_X1 U20887 ( .A1(n17782), .A2(n17746), .ZN(n17798) );
  NOR2_X1 U20888 ( .A1(n17747), .A2(n17798), .ZN(n17760) );
  OAI211_X1 U20889 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17760), .B(n17748), .ZN(n17749) );
  OAI211_X1 U20890 ( .C1(n17786), .C2(n17751), .A(n17750), .B(n17749), .ZN(
        n17752) );
  AOI21_X1 U20891 ( .B1(n17857), .B2(n18076), .A(n17752), .ZN(n17753) );
  OAI221_X1 U20892 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17755), 
        .C1(n18074), .C2(n17754), .A(n17753), .ZN(P3_U2814) );
  NOR2_X1 U20893 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17772), .ZN(
        n18086) );
  NAND2_X1 U20894 ( .A1(n17777), .A2(n18079), .ZN(n17765) );
  OAI22_X1 U20895 ( .A1(n18148), .A2(n18836), .B1(n17786), .B2(n17756), .ZN(
        n17757) );
  AOI221_X1 U20896 ( .B1(n17760), .B2(n17759), .C1(n17758), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17757), .ZN(n17764) );
  NOR2_X1 U20897 ( .A1(n18099), .A2(n17822), .ZN(n17774) );
  NAND2_X1 U20898 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18095), .ZN(
        n18124) );
  OAI221_X1 U20899 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17775), 
        .C1(n18098), .C2(n17774), .A(n18124), .ZN(n17761) );
  XOR2_X1 U20900 ( .A(n15698), .B(n17761), .Z(n18087) );
  NOR2_X1 U20901 ( .A1(n18001), .A2(n17944), .ZN(n17762) );
  NAND2_X1 U20902 ( .A1(n18083), .A2(n17808), .ZN(n17766) );
  NAND2_X1 U20903 ( .A1(n15698), .A2(n17766), .ZN(n18089) );
  AOI22_X1 U20904 ( .A1(n17857), .A2(n18087), .B1(n17762), .B2(n18089), .ZN(
        n17763) );
  OAI211_X1 U20905 ( .C1(n18086), .C2(n17765), .A(n17764), .B(n17763), .ZN(
        P3_U2815) );
  NOR2_X1 U20906 ( .A1(n18135), .A2(n18099), .ZN(n18118) );
  OAI221_X1 U20907 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18118), .A(n17766), .ZN(
        n18111) );
  NAND3_X1 U20908 ( .A1(n18662), .A2(n17872), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17863) );
  NOR2_X1 U20909 ( .A1(n17767), .A2(n17863), .ZN(n17813) );
  AOI21_X1 U20910 ( .B1(n17780), .B2(n17813), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17768) );
  OAI22_X1 U20911 ( .A1(n17919), .A2(n17770), .B1(n17769), .B2(n17768), .ZN(
        n17771) );
  AOI21_X1 U20912 ( .B1(n18255), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17771), 
        .ZN(n17779) );
  AOI21_X1 U20913 ( .B1(n18098), .B2(n17773), .A(n17772), .ZN(n18106) );
  OAI21_X1 U20914 ( .B1(n17775), .B2(n17774), .A(n18124), .ZN(n17776) );
  XOR2_X1 U20915 ( .A(n17776), .B(n18098), .Z(n18108) );
  AOI22_X1 U20916 ( .A1(n17777), .A2(n18106), .B1(n17857), .B2(n18108), .ZN(
        n17778) );
  OAI211_X1 U20917 ( .C1(n17944), .C2(n18111), .A(n17779), .B(n17778), .ZN(
        P3_U2816) );
  NAND2_X1 U20918 ( .A1(n18113), .A2(n17840), .ZN(n17807) );
  INV_X1 U20919 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17787) );
  AOI211_X1 U20920 ( .C1(n17797), .C2(n17787), .A(n17780), .B(n17798), .ZN(
        n17789) );
  OAI21_X1 U20921 ( .B1(n17782), .B2(n17781), .A(n18791), .ZN(n17783) );
  AOI21_X1 U20922 ( .B1(n17784), .B2(n17783), .A(n17889), .ZN(n17796) );
  OAI22_X1 U20923 ( .A1(n17796), .A2(n17787), .B1(n17786), .B2(n17785), .ZN(
        n17788) );
  AOI211_X1 U20924 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18255), .A(n17789), 
        .B(n17788), .ZN(n17795) );
  NOR2_X1 U20925 ( .A1(n18099), .A2(n18133), .ZN(n18116) );
  OAI22_X1 U20926 ( .A1(n18118), .A2(n17944), .B1(n18116), .B2(n16499), .ZN(
        n17804) );
  INV_X1 U20927 ( .A(n18099), .ZN(n18094) );
  AOI22_X1 U20928 ( .A1(n17790), .A2(n18094), .B1(n18132), .B2(n17792), .ZN(
        n17791) );
  AOI21_X1 U20929 ( .B1(n17802), .B2(n17792), .A(n17791), .ZN(n17793) );
  XOR2_X1 U20930 ( .A(n17793), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18112) );
  AOI22_X1 U20931 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17804), .B1(
        n17857), .B2(n18112), .ZN(n17794) );
  OAI211_X1 U20932 ( .C1(n18124), .C2(n17807), .A(n17795), .B(n17794), .ZN(
        P3_U2817) );
  NAND2_X1 U20933 ( .A1(n18255), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18130) );
  OAI221_X1 U20934 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17798), .C1(
        n17797), .C2(n17796), .A(n18130), .ZN(n17799) );
  AOI21_X1 U20935 ( .B1(n17801), .B2(n17800), .A(n17799), .ZN(n17806) );
  OR2_X1 U20936 ( .A1(n18142), .A2(n17822), .ZN(n17815) );
  OAI21_X1 U20937 ( .B1(n17819), .B2(n17815), .A(n17802), .ZN(n17803) );
  XOR2_X1 U20938 ( .A(n17803), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18129) );
  AOI22_X1 U20939 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17804), .B1(
        n17857), .B2(n18129), .ZN(n17805) );
  OAI211_X1 U20940 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17807), .A(
        n17806), .B(n17805), .ZN(P3_U2818) );
  OAI22_X1 U20941 ( .A1(n17809), .A2(n16499), .B1(n17808), .B2(n17944), .ZN(
        n17842) );
  AOI21_X1 U20942 ( .B1(n18142), .B2(n17840), .A(n17842), .ZN(n17830) );
  NOR2_X1 U20943 ( .A1(n17889), .A2(n17850), .ZN(n17904) );
  INV_X1 U20944 ( .A(n17904), .ZN(n17936) );
  INV_X1 U20945 ( .A(n17863), .ZN(n17810) );
  NAND3_X1 U20946 ( .A1(n17847), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17810), .ZN(n17835) );
  NOR2_X1 U20947 ( .A1(n17825), .A2(n17835), .ZN(n17824) );
  AOI21_X1 U20948 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17936), .A(
        n17824), .ZN(n17812) );
  OAI22_X1 U20949 ( .A1(n17813), .A2(n17812), .B1(n17919), .B2(n17811), .ZN(
        n17814) );
  AOI21_X1 U20950 ( .B1(n18255), .B2(P3_REIP_REG_11__SCAN_IN), .A(n17814), 
        .ZN(n17818) );
  OAI21_X1 U20951 ( .B1(n17821), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17815), .ZN(n17816) );
  XOR2_X1 U20952 ( .A(n17816), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18146) );
  NOR2_X1 U20953 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18142), .ZN(
        n18145) );
  AOI22_X1 U20954 ( .A1(n17857), .A2(n18146), .B1(n18145), .B2(n17840), .ZN(
        n17817) );
  OAI211_X1 U20955 ( .C1(n17830), .C2(n17819), .A(n17818), .B(n17817), .ZN(
        P3_U2819) );
  AOI21_X1 U20956 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17840), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17829) );
  AOI22_X1 U20957 ( .A1(n18255), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17820), 
        .B2(n17934), .ZN(n17828) );
  OAI21_X1 U20958 ( .B1(n17841), .B2(n17822), .A(n17821), .ZN(n17823) );
  XNOR2_X1 U20959 ( .A(n10101), .B(n17823), .ZN(n18152) );
  AOI211_X1 U20960 ( .C1(n17835), .C2(n17825), .A(n17904), .B(n17824), .ZN(
        n17826) );
  AOI21_X1 U20961 ( .B1(n17857), .B2(n18152), .A(n17826), .ZN(n17827) );
  OAI211_X1 U20962 ( .C1(n17830), .C2(n17829), .A(n17828), .B(n17827), .ZN(
        P3_U2820) );
  NOR2_X1 U20963 ( .A1(n17832), .A2(n17831), .ZN(n17833) );
  XOR2_X1 U20964 ( .A(n17833), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18163) );
  NOR2_X1 U20965 ( .A1(n17834), .A2(n17863), .ZN(n17836) );
  OAI211_X1 U20966 ( .C1(n17836), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17936), .B(n17835), .ZN(n17837) );
  NAND2_X1 U20967 ( .A1(n18255), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18160) );
  OAI211_X1 U20968 ( .C1(n17919), .C2(n17838), .A(n17837), .B(n18160), .ZN(
        n17839) );
  AOI221_X1 U20969 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17842), .C1(
        n17841), .C2(n17840), .A(n17839), .ZN(n17843) );
  OAI21_X1 U20970 ( .B1(n18163), .B2(n17844), .A(n17843), .ZN(P3_U2821) );
  OAI21_X1 U20971 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17846), .A(
        n17845), .ZN(n18178) );
  AOI211_X1 U20972 ( .C1(n20914), .C2(n17848), .A(n17847), .B(n18365), .ZN(
        n17852) );
  AOI21_X1 U20973 ( .B1(n17850), .B2(n17849), .A(n17889), .ZN(n17867) );
  OAI22_X1 U20974 ( .A1(n18148), .A2(n21110), .B1(n20914), .B2(n17867), .ZN(
        n17851) );
  AOI211_X1 U20975 ( .C1(n17853), .C2(n17934), .A(n17852), .B(n17851), .ZN(
        n17859) );
  AOI21_X1 U20976 ( .B1(n17855), .B2(n18171), .A(n17854), .ZN(n18173) );
  XOR2_X1 U20977 ( .A(n17856), .B(n18178), .Z(n18174) );
  AOI22_X1 U20978 ( .A1(n9734), .A2(n18173), .B1(n17857), .B2(n18174), .ZN(
        n17858) );
  OAI211_X1 U20979 ( .C1(n16499), .C2(n18178), .A(n17859), .B(n17858), .ZN(
        P3_U2822) );
  NAND2_X1 U20980 ( .A1(n17861), .A2(n17860), .ZN(n17862) );
  XOR2_X1 U20981 ( .A(n17862), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18184) );
  OAI22_X1 U20982 ( .A1(n17919), .A2(n17864), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17863), .ZN(n17870) );
  OAI21_X1 U20983 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17866), .A(
        n17865), .ZN(n18183) );
  OAI22_X1 U20984 ( .A1(n17943), .A2(n18183), .B1(n17868), .B2(n17867), .ZN(
        n17869) );
  AOI211_X1 U20985 ( .C1(n18255), .C2(P3_REIP_REG_7__SCAN_IN), .A(n17870), .B(
        n17869), .ZN(n17871) );
  OAI21_X1 U20986 ( .B1(n17944), .B2(n18184), .A(n17871), .ZN(P3_U2823) );
  NAND2_X1 U20987 ( .A1(n18662), .A2(n17872), .ZN(n17876) );
  NAND2_X1 U20988 ( .A1(n17936), .A2(n17876), .ZN(n17891) );
  OAI21_X1 U20989 ( .B1(n17875), .B2(n17874), .A(n17873), .ZN(n18191) );
  OAI22_X1 U20990 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17876), .B1(
        n17943), .B2(n18191), .ZN(n17877) );
  AOI21_X1 U20991 ( .B1(n18255), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17877), .ZN(
        n17882) );
  AOI21_X1 U20992 ( .B1(n17879), .B2(n18195), .A(n17878), .ZN(n18193) );
  AOI22_X1 U20993 ( .A1(n9734), .A2(n18193), .B1(n17880), .B2(n17934), .ZN(
        n17881) );
  OAI211_X1 U20994 ( .C1(n17883), .C2(n17891), .A(n17882), .B(n17881), .ZN(
        P3_U2824) );
  OAI21_X1 U20995 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17885), .A(
        n17884), .ZN(n18206) );
  AOI21_X1 U20996 ( .B1(n17888), .B2(n17887), .A(n17886), .ZN(n18204) );
  NOR2_X1 U20997 ( .A1(n17925), .A2(n17889), .ZN(n17924) );
  AND2_X1 U20998 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17924), .ZN(
        n17903) );
  AOI21_X1 U20999 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17903), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17892) );
  OAI22_X1 U21000 ( .A1(n17892), .A2(n17891), .B1(n17919), .B2(n17890), .ZN(
        n17893) );
  AOI21_X1 U21001 ( .B1(n9734), .B2(n18204), .A(n17893), .ZN(n17895) );
  INV_X1 U21002 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18818) );
  NOR2_X1 U21003 ( .A1(n18148), .A2(n18818), .ZN(n18203) );
  INV_X1 U21004 ( .A(n18203), .ZN(n17894) );
  OAI211_X1 U21005 ( .C1(n17943), .C2(n18206), .A(n17895), .B(n17894), .ZN(
        P3_U2825) );
  OAI21_X1 U21006 ( .B1(n17898), .B2(n17897), .A(n17896), .ZN(n18216) );
  OAI22_X1 U21007 ( .A1(n18148), .A2(n18815), .B1(n17943), .B2(n18216), .ZN(
        n17899) );
  AOI21_X1 U21008 ( .B1(n18662), .B2(n17900), .A(n17899), .ZN(n17906) );
  AOI21_X1 U21009 ( .B1(n18210), .B2(n17902), .A(n17901), .ZN(n18213) );
  NOR2_X1 U21010 ( .A1(n17904), .A2(n17903), .ZN(n17915) );
  AOI22_X1 U21011 ( .A1(n9734), .A2(n18213), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17915), .ZN(n17905) );
  OAI211_X1 U21012 ( .C1(n17919), .C2(n17907), .A(n17906), .B(n17905), .ZN(
        P3_U2826) );
  AOI21_X1 U21013 ( .B1(n17910), .B2(n17909), .A(n17908), .ZN(n18223) );
  OAI21_X1 U21014 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17912), .A(
        n17911), .ZN(n18225) );
  OAI22_X1 U21015 ( .A1(n18148), .A2(n18813), .B1(n17943), .B2(n18225), .ZN(
        n17913) );
  AOI21_X1 U21016 ( .B1(n9734), .B2(n18223), .A(n17913), .ZN(n17917) );
  OAI21_X1 U21017 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17924), .A(
        n17915), .ZN(n17916) );
  OAI211_X1 U21018 ( .C1(n17919), .C2(n17918), .A(n17917), .B(n17916), .ZN(
        P3_U2827) );
  OAI21_X1 U21019 ( .B1(n17922), .B2(n17921), .A(n17920), .ZN(n18241) );
  AOI211_X1 U21020 ( .C1(n18234), .C2(n18233), .A(n17923), .B(n17944), .ZN(
        n17927) );
  AOI21_X1 U21021 ( .B1(n18365), .B2(n17925), .A(n17924), .ZN(n17926) );
  AOI211_X1 U21022 ( .C1(n17928), .C2(n17934), .A(n17927), .B(n17926), .ZN(
        n17929) );
  NAND2_X1 U21023 ( .A1(n18255), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18239) );
  OAI211_X1 U21024 ( .C1(n17943), .C2(n18241), .A(n17929), .B(n18239), .ZN(
        P3_U2828) );
  AND2_X1 U21025 ( .A1(n17939), .A2(n18907), .ZN(n17930) );
  XNOR2_X1 U21026 ( .A(n17930), .B(n17932), .ZN(n18252) );
  OAI21_X1 U21027 ( .B1(n17932), .B2(n17938), .A(n17931), .ZN(n18246) );
  OAI22_X1 U21028 ( .A1(n18148), .A2(n18809), .B1(n17943), .B2(n18246), .ZN(
        n17933) );
  AOI221_X1 U21029 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17936), .C1(
        n17935), .C2(n17934), .A(n17933), .ZN(n17937) );
  OAI21_X1 U21030 ( .B1(n18252), .B2(n17944), .A(n17937), .ZN(P3_U2829) );
  AOI21_X1 U21031 ( .B1(n17939), .B2(n18907), .A(n17938), .ZN(n18259) );
  INV_X1 U21032 ( .A(n18259), .ZN(n18257) );
  NAND3_X1 U21033 ( .A1(n18889), .A2(n18791), .A3(n17940), .ZN(n17941) );
  AOI22_X1 U21034 ( .A1(n18255), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17941), .ZN(n17942) );
  OAI221_X1 U21035 ( .B1(n18259), .B2(n17944), .C1(n18257), .C2(n17943), .A(
        n17942), .ZN(P3_U2830) );
  AOI22_X1 U21036 ( .A1(n18255), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18189), .ZN(n17957) );
  NOR2_X1 U21037 ( .A1(n18217), .A2(n17953), .ZN(n17954) );
  OAI22_X1 U21038 ( .A1(n17946), .A2(n18117), .B1(n17945), .B2(n18115), .ZN(
        n17947) );
  AOI211_X1 U21039 ( .C1(n17949), .C2(n18226), .A(n17948), .B(n17947), .ZN(
        n17952) );
  NAND2_X1 U21040 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17951) );
  OAI22_X1 U21041 ( .A1(n18721), .A2(n17950), .B1(n17992), .B2(n18071), .ZN(
        n18012) );
  NAND3_X1 U21042 ( .A1(n18051), .A2(n18010), .A3(n18012), .ZN(n17979) );
  OAI21_X1 U21043 ( .B1(n17951), .B2(n17979), .A(n18226), .ZN(n17966) );
  NAND2_X1 U21044 ( .A1(n17952), .A2(n17966), .ZN(n17962) );
  OAI22_X1 U21045 ( .A1(n17955), .A2(n17954), .B1(n17962), .B2(n17953), .ZN(
        n17956) );
  OAI211_X1 U21046 ( .C1(n17958), .C2(n18162), .A(n17957), .B(n17956), .ZN(
        P3_U2835) );
  NOR2_X1 U21047 ( .A1(n17959), .A2(n18018), .ZN(n17987) );
  AOI21_X1 U21048 ( .B1(n17961), .B2(n17987), .A(n17960), .ZN(n17964) );
  OAI221_X1 U21049 ( .B1(n18189), .B2(n18254), .C1(n18189), .C2(n17962), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17963) );
  OAI211_X1 U21050 ( .C1(n17965), .C2(n18162), .A(n17964), .B(n17963), .ZN(
        P3_U2836) );
  OAI221_X1 U21051 ( .B1(n18739), .B2(n18053), .C1(n18739), .C2(n17969), .A(
        n17966), .ZN(n17970) );
  NOR2_X1 U21052 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17967), .ZN(
        n17968) );
  AOI22_X1 U21053 ( .A1(n17970), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n17969), .B2(n17968), .ZN(n17972) );
  OAI21_X1 U21054 ( .B1(n18217), .B2(n17972), .A(n17971), .ZN(n17976) );
  OAI22_X1 U21055 ( .A1(n18162), .A2(n17974), .B1(n18251), .B2(n17973), .ZN(
        n17975) );
  AOI211_X1 U21056 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18189), .A(
        n17976), .B(n17975), .ZN(n17977) );
  OAI21_X1 U21057 ( .B1(n18179), .B2(n17978), .A(n17977), .ZN(P3_U2837) );
  AOI22_X1 U21058 ( .A1(n18750), .A2(n17980), .B1(n18226), .B2(n17979), .ZN(
        n17981) );
  OAI211_X1 U21059 ( .C1(n17982), .C2(n18115), .A(n17981), .B(n18245), .ZN(
        n17985) );
  AOI211_X1 U21060 ( .C1(n18751), .C2(n17983), .A(n17998), .B(n17985), .ZN(
        n17984) );
  OR2_X1 U21061 ( .A1(n18255), .A2(n17984), .ZN(n17999) );
  OAI21_X1 U21062 ( .B1(n18168), .B2(n17985), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17991) );
  AOI22_X1 U21063 ( .A1(n18175), .A2(n17988), .B1(n17987), .B2(n17986), .ZN(
        n17990) );
  NAND2_X1 U21064 ( .A1(n18255), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17989) );
  OAI211_X1 U21065 ( .C1(n17999), .C2(n17991), .A(n17990), .B(n17989), .ZN(
        P3_U2838) );
  INV_X1 U21066 ( .A(n17992), .ZN(n17993) );
  NAND3_X1 U21067 ( .A1(n17993), .A2(n18009), .A3(n18245), .ZN(n17997) );
  AOI21_X1 U21068 ( .B1(n17995), .B2(n18175), .A(n17994), .ZN(n17996) );
  OAI221_X1 U21069 ( .B1(n17999), .B2(n17998), .C1(n17999), .C2(n17997), .A(
        n17996), .ZN(P3_U2839) );
  OAI22_X1 U21070 ( .A1(n18001), .A2(n18117), .B1(n18000), .B2(n18115), .ZN(
        n18019) );
  AOI21_X1 U21071 ( .B1(n18051), .B2(n18002), .A(n18722), .ZN(n18003) );
  AOI21_X1 U21072 ( .B1(n18751), .B2(n18004), .A(n18003), .ZN(n18022) );
  NAND2_X1 U21073 ( .A1(n18117), .A2(n18115), .ZN(n18141) );
  AOI22_X1 U21074 ( .A1(n18716), .A2(n18006), .B1(n18005), .B2(n18141), .ZN(
        n18026) );
  OAI211_X1 U21075 ( .C1(n18151), .C2(n18007), .A(n18022), .B(n18026), .ZN(
        n18008) );
  NOR2_X1 U21076 ( .A1(n18019), .A2(n18008), .ZN(n18013) );
  AOI21_X1 U21077 ( .B1(n18010), .B2(n18009), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18011) );
  AOI21_X1 U21078 ( .B1(n18013), .B2(n18012), .A(n18011), .ZN(n18014) );
  AOI22_X1 U21079 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18189), .B1(
        n18254), .B2(n18014), .ZN(n18016) );
  NAND2_X1 U21080 ( .A1(n18255), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18015) );
  OAI211_X1 U21081 ( .C1(n18017), .C2(n18162), .A(n18016), .B(n18015), .ZN(
        P3_U2840) );
  NOR2_X1 U21082 ( .A1(n18020), .A2(n18018), .ZN(n18041) );
  NAND2_X1 U21083 ( .A1(n18732), .A2(n18739), .ZN(n18244) );
  NOR2_X1 U21084 ( .A1(n18217), .A2(n18019), .ZN(n18068) );
  OAI21_X1 U21085 ( .B1(n18020), .B2(n18071), .A(n18721), .ZN(n18021) );
  NAND3_X1 U21086 ( .A1(n18068), .A2(n18022), .A3(n18021), .ZN(n18033) );
  AOI21_X1 U21087 ( .B1(n18023), .B2(n18244), .A(n18033), .ZN(n18025) );
  AOI211_X1 U21088 ( .C1(n18026), .C2(n18025), .A(n18255), .B(n18024), .ZN(
        n18027) );
  AOI21_X1 U21089 ( .B1(n18041), .B2(n18028), .A(n18027), .ZN(n18030) );
  NAND2_X1 U21090 ( .A1(n18255), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18029) );
  OAI211_X1 U21091 ( .C1(n18031), .C2(n18162), .A(n18030), .B(n18029), .ZN(
        P3_U2841) );
  NAND3_X1 U21092 ( .A1(n18046), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18244), 
        .ZN(n18034) );
  OAI221_X1 U21093 ( .B1(n18033), .B2(n18032), .C1(n18033), .C2(n18141), .A(
        n18148), .ZN(n18045) );
  NAND2_X1 U21094 ( .A1(n18034), .A2(n18045), .ZN(n18036) );
  AOI22_X1 U21095 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18036), .B1(
        n18035), .B2(n18041), .ZN(n18038) );
  NAND2_X1 U21096 ( .A1(n18255), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18037) );
  OAI211_X1 U21097 ( .C1(n18039), .C2(n18162), .A(n18038), .B(n18037), .ZN(
        P3_U2842) );
  INV_X1 U21098 ( .A(n18040), .ZN(n18042) );
  AOI22_X1 U21099 ( .A1(n18175), .A2(n18042), .B1(n18041), .B2(n18046), .ZN(
        n18044) );
  NAND2_X1 U21100 ( .A1(n18255), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18043) );
  OAI211_X1 U21101 ( .C1(n18046), .C2(n18045), .A(n18044), .B(n18043), .ZN(
        P3_U2843) );
  INV_X1 U21102 ( .A(n18228), .ZN(n18047) );
  OAI22_X1 U21103 ( .A1(n18207), .A2(n18739), .B1(n18209), .B2(n18047), .ZN(
        n18080) );
  NAND2_X1 U21104 ( .A1(n18254), .A2(n18080), .ZN(n18197) );
  OAI222_X1 U21105 ( .A1(n18135), .A2(n18251), .B1(n18081), .B2(n18196), .C1(
        n18179), .C2(n18133), .ZN(n18159) );
  AND2_X1 U21106 ( .A1(n18159), .A2(n18048), .ZN(n18075) );
  AOI21_X1 U21107 ( .B1(n18050), .B2(n18075), .A(n18049), .ZN(n18060) );
  NOR2_X1 U21108 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18164), .ZN(
        n18058) );
  NOR2_X1 U21109 ( .A1(n18732), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18227) );
  INV_X1 U21110 ( .A(n18051), .ZN(n18052) );
  NOR3_X1 U21111 ( .A1(n18227), .A2(n18052), .A3(n18074), .ZN(n18057) );
  NOR2_X1 U21112 ( .A1(n18053), .A2(n18739), .ZN(n18055) );
  OAI22_X1 U21113 ( .A1(n18751), .A2(n18141), .B1(n18055), .B2(n18054), .ZN(
        n18056) );
  OAI211_X1 U21114 ( .C1(n18164), .C2(n18057), .A(n18068), .B(n18056), .ZN(
        n18062) );
  OAI211_X1 U21115 ( .C1(n18058), .C2(n18062), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n18148), .ZN(n18059) );
  OAI211_X1 U21116 ( .C1(n18061), .C2(n18162), .A(n18060), .B(n18059), .ZN(
        P3_U2844) );
  NOR2_X1 U21117 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18074), .ZN(
        n18064) );
  AND2_X1 U21118 ( .A1(n18148), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18063) );
  AOI22_X1 U21119 ( .A1(n18075), .A2(n18064), .B1(n18063), .B2(n18062), .ZN(
        n18066) );
  OAI211_X1 U21120 ( .C1(n18067), .C2(n18162), .A(n18066), .B(n18065), .ZN(
        P3_U2845) );
  INV_X1 U21121 ( .A(n18068), .ZN(n18073) );
  AOI22_X1 U21122 ( .A1(n18751), .A2(n18070), .B1(n18716), .B2(n18069), .ZN(
        n18114) );
  OAI21_X1 U21123 ( .B1(n15698), .B2(n18721), .A(n18071), .ZN(n18072) );
  OAI211_X1 U21124 ( .C1(n18151), .C2(n18083), .A(n18114), .B(n18072), .ZN(
        n18082) );
  OAI221_X1 U21125 ( .B1(n18073), .B2(n18168), .C1(n18073), .C2(n18082), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U21126 ( .A1(n18175), .A2(n18076), .B1(n18075), .B2(n18074), .ZN(
        n18077) );
  OAI221_X1 U21127 ( .B1(n18255), .B2(n18078), .C1(n18148), .C2(n18838), .A(
        n18077), .ZN(P3_U2846) );
  AOI22_X1 U21128 ( .A1(n18255), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18189), .ZN(n18093) );
  NAND2_X1 U21129 ( .A1(n18134), .A2(n18079), .ZN(n18085) );
  INV_X1 U21130 ( .A(n18080), .ZN(n18219) );
  NOR3_X1 U21131 ( .A1(n18219), .A2(n18081), .A3(n18180), .ZN(n18100) );
  OAI221_X1 U21132 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18083), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18100), .A(n18082), .ZN(
        n18084) );
  OAI21_X1 U21133 ( .B1(n18086), .B2(n18085), .A(n18084), .ZN(n18088) );
  AOI22_X1 U21134 ( .A1(n18254), .A2(n18088), .B1(n18175), .B2(n18087), .ZN(
        n18092) );
  NAND3_X1 U21135 ( .A1(n18258), .A2(n18090), .A3(n18089), .ZN(n18091) );
  NAND3_X1 U21136 ( .A1(n18093), .A2(n18092), .A3(n18091), .ZN(P3_U2847) );
  NOR2_X1 U21137 ( .A1(n18148), .A2(n18835), .ZN(n18105) );
  AOI21_X1 U21138 ( .B1(n18094), .B2(n18137), .A(n18732), .ZN(n18120) );
  OAI21_X1 U21139 ( .B1(n18120), .B2(n18095), .A(n18244), .ZN(n18096) );
  OAI211_X1 U21140 ( .C1(n18722), .C2(n18101), .A(n18114), .B(n18096), .ZN(
        n18097) );
  AOI211_X1 U21141 ( .C1(n18751), .C2(n18099), .A(n18098), .B(n18097), .ZN(
        n18103) );
  AOI21_X1 U21142 ( .B1(n18101), .B2(n18100), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18102) );
  NOR3_X1 U21143 ( .A1(n18103), .A2(n18102), .A3(n18217), .ZN(n18104) );
  AOI211_X1 U21144 ( .C1(n18189), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18105), .B(n18104), .ZN(n18110) );
  AOI22_X1 U21145 ( .A1(n18175), .A2(n18108), .B1(n18107), .B2(n18106), .ZN(
        n18109) );
  OAI211_X1 U21146 ( .C1(n18251), .C2(n18111), .A(n18110), .B(n18109), .ZN(
        P3_U2848) );
  NAND2_X1 U21147 ( .A1(n18113), .A2(n18159), .ZN(n18126) );
  AOI22_X1 U21148 ( .A1(n18255), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18175), 
        .B2(n18112), .ZN(n18123) );
  NOR2_X1 U21149 ( .A1(n18151), .A2(n18113), .ZN(n18144) );
  INV_X1 U21150 ( .A(n18114), .ZN(n18139) );
  OAI22_X1 U21151 ( .A1(n18118), .A2(n18117), .B1(n18116), .B2(n18115), .ZN(
        n18119) );
  NOR4_X1 U21152 ( .A1(n18144), .A2(n18120), .A3(n18139), .A4(n18119), .ZN(
        n18127) );
  OAI211_X1 U21153 ( .C1(n18151), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18254), .B(n18127), .ZN(n18121) );
  NAND3_X1 U21154 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18148), .A3(
        n18121), .ZN(n18122) );
  OAI211_X1 U21155 ( .C1(n18126), .C2(n18124), .A(n18123), .B(n18122), .ZN(
        P3_U2849) );
  NAND2_X1 U21156 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18254), .ZN(
        n18125) );
  AOI22_X1 U21157 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18127), .B1(
        n18126), .B2(n18125), .ZN(n18128) );
  AOI21_X1 U21158 ( .B1(n18175), .B2(n18129), .A(n18128), .ZN(n18131) );
  OAI211_X1 U21159 ( .C1(n18245), .C2(n18132), .A(n18131), .B(n18130), .ZN(
        P3_U2850) );
  AOI22_X1 U21160 ( .A1(n18750), .A2(n18135), .B1(n18134), .B2(n18133), .ZN(
        n18136) );
  OAI211_X1 U21161 ( .C1(n18732), .C2(n18137), .A(n18254), .B(n18136), .ZN(
        n18138) );
  NOR2_X1 U21162 ( .A1(n18139), .A2(n18138), .ZN(n18157) );
  OAI21_X1 U21163 ( .B1(n18732), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18157), .ZN(n18140) );
  AOI21_X1 U21164 ( .B1(n18142), .B2(n18141), .A(n18140), .ZN(n18150) );
  OAI21_X1 U21165 ( .B1(n18732), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18150), .ZN(n18143) );
  OAI21_X1 U21166 ( .B1(n18144), .B2(n18143), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18149) );
  AOI22_X1 U21167 ( .A1(n18175), .A2(n18146), .B1(n18145), .B2(n18159), .ZN(
        n18147) );
  OAI221_X1 U21168 ( .B1(n18255), .B2(n18149), .C1(n18148), .C2(n18828), .A(
        n18147), .ZN(P3_U2851) );
  NAND2_X1 U21169 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18159), .ZN(
        n18156) );
  AOI221_X1 U21170 ( .B1(n18151), .B2(n18150), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18150), .A(n18255), .ZN(
        n18153) );
  AOI22_X1 U21171 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18153), .B1(
        n18175), .B2(n18152), .ZN(n18155) );
  NAND2_X1 U21172 ( .A1(n18255), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18154) );
  OAI211_X1 U21173 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n18156), .A(
        n18155), .B(n18154), .ZN(P3_U2852) );
  OAI21_X1 U21174 ( .B1(n18255), .B2(n18157), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18158) );
  OAI21_X1 U21175 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18159), .A(
        n18158), .ZN(n18161) );
  OAI211_X1 U21176 ( .C1(n18163), .C2(n18162), .A(n18161), .B(n18160), .ZN(
        P3_U2853) );
  INV_X1 U21177 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21107) );
  NOR3_X1 U21178 ( .A1(n21107), .A2(n18195), .A3(n18196), .ZN(n18172) );
  OAI22_X1 U21179 ( .A1(n18166), .A2(n18739), .B1(n18165), .B2(n18164), .ZN(
        n18167) );
  OR2_X1 U21180 ( .A1(n18227), .A2(n18167), .ZN(n18190) );
  AOI211_X1 U21181 ( .C1(n18168), .C2(n18195), .A(n21107), .B(n18190), .ZN(
        n18181) );
  OAI21_X1 U21182 ( .B1(n18181), .B2(n18242), .A(n18245), .ZN(n18170) );
  NOR2_X1 U21183 ( .A1(n18148), .A2(n21110), .ZN(n18169) );
  AOI221_X1 U21184 ( .B1(n18172), .B2(n18171), .C1(n18170), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18169), .ZN(n18177) );
  AOI22_X1 U21185 ( .A1(n18175), .A2(n18174), .B1(n18258), .B2(n18173), .ZN(
        n18176) );
  OAI211_X1 U21186 ( .C1(n18179), .C2(n18178), .A(n18177), .B(n18176), .ZN(
        P3_U2854) );
  OR2_X1 U21187 ( .A1(n18180), .A2(n18219), .ZN(n18182) );
  AOI221_X1 U21188 ( .B1(n18195), .B2(n21107), .C1(n18182), .C2(n21107), .A(
        n18181), .ZN(n18186) );
  OAI22_X1 U21189 ( .A1(n18251), .A2(n18184), .B1(n18247), .B2(n18183), .ZN(
        n18185) );
  AOI21_X1 U21190 ( .B1(n18254), .B2(n18186), .A(n18185), .ZN(n18188) );
  NAND2_X1 U21191 ( .A1(n18255), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n18187) );
  OAI211_X1 U21192 ( .C1(n18245), .C2(n21107), .A(n18188), .B(n18187), .ZN(
        P3_U2855) );
  AOI21_X1 U21193 ( .B1(n18254), .B2(n18190), .A(n18189), .ZN(n18199) );
  OAI22_X1 U21194 ( .A1(n18148), .A2(n18819), .B1(n18247), .B2(n18191), .ZN(
        n18192) );
  AOI21_X1 U21195 ( .B1(n18258), .B2(n18193), .A(n18192), .ZN(n18194) );
  OAI221_X1 U21196 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18196), .C1(
        n18195), .C2(n18199), .A(n18194), .ZN(P3_U2856) );
  NAND2_X1 U21197 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18198) );
  NOR2_X1 U21198 ( .A1(n18198), .A2(n18197), .ZN(n18201) );
  INV_X1 U21199 ( .A(n18199), .ZN(n18200) );
  MUX2_X1 U21200 ( .A(n18201), .B(n18200), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18202) );
  AOI211_X1 U21201 ( .C1(n18204), .C2(n18258), .A(n18203), .B(n18202), .ZN(
        n18205) );
  OAI21_X1 U21202 ( .B1(n18247), .B2(n18206), .A(n18205), .ZN(P3_U2857) );
  NAND2_X1 U21203 ( .A1(n18751), .A2(n18207), .ZN(n18232) );
  NAND2_X1 U21204 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18232), .ZN(
        n18208) );
  AOI211_X1 U21205 ( .C1(n18209), .C2(n18226), .A(n18227), .B(n18208), .ZN(
        n18218) );
  AOI221_X1 U21206 ( .B1(n18218), .B2(n18245), .C1(n18242), .C2(n18245), .A(
        n18210), .ZN(n18212) );
  NOR4_X1 U21207 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18219), .A3(
        n18220), .A4(n18217), .ZN(n18211) );
  AOI211_X1 U21208 ( .C1(n18213), .C2(n18258), .A(n18212), .B(n18211), .ZN(
        n18215) );
  NAND2_X1 U21209 ( .A1(n18255), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18214) );
  OAI211_X1 U21210 ( .C1(n18247), .C2(n18216), .A(n18215), .B(n18214), .ZN(
        P3_U2858) );
  AOI211_X1 U21211 ( .C1(n18219), .C2(n18220), .A(n18218), .B(n18217), .ZN(
        n18222) );
  OAI22_X1 U21212 ( .A1(n18148), .A2(n18813), .B1(n18220), .B2(n18245), .ZN(
        n18221) );
  AOI211_X1 U21213 ( .C1(n18223), .C2(n18258), .A(n18222), .B(n18221), .ZN(
        n18224) );
  OAI21_X1 U21214 ( .B1(n18247), .B2(n18225), .A(n18224), .ZN(P3_U2859) );
  INV_X1 U21215 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18891) );
  OAI211_X1 U21216 ( .C1(n18227), .C2(n18891), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n18226), .ZN(n18231) );
  NAND3_X1 U21217 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18228), .A3(
        n18236), .ZN(n18230) );
  NAND4_X1 U21218 ( .A1(n18751), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18229) );
  NAND4_X1 U21219 ( .A1(n18232), .A2(n18231), .A3(n18230), .A4(n18229), .ZN(
        n18238) );
  XNOR2_X1 U21220 ( .A(n18234), .B(n18233), .ZN(n18235) );
  OAI22_X1 U21221 ( .A1(n18236), .A2(n18245), .B1(n18251), .B2(n18235), .ZN(
        n18237) );
  AOI21_X1 U21222 ( .B1(n18254), .B2(n18238), .A(n18237), .ZN(n18240) );
  OAI211_X1 U21223 ( .C1(n18247), .C2(n18241), .A(n18240), .B(n18239), .ZN(
        P3_U2860) );
  NOR2_X1 U21224 ( .A1(n18243), .A2(n18242), .ZN(n18249) );
  NAND3_X1 U21225 ( .A1(n18254), .A2(n18907), .A3(n18244), .ZN(n18262) );
  NAND2_X1 U21226 ( .A1(n18245), .A2(n18262), .ZN(n18253) );
  OAI22_X1 U21227 ( .A1(n18148), .A2(n18809), .B1(n18247), .B2(n18246), .ZN(
        n18248) );
  AOI221_X1 U21228 ( .B1(n18249), .B2(n18891), .C1(n18253), .C2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n18248), .ZN(n18250) );
  OAI21_X1 U21229 ( .B1(n18252), .B2(n18251), .A(n18250), .ZN(P3_U2861) );
  AOI21_X1 U21230 ( .B1(n18254), .B2(n18716), .A(n18253), .ZN(n18263) );
  AND2_X1 U21231 ( .A1(n18255), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18256) );
  AOI221_X1 U21232 ( .B1(n18260), .B2(n18259), .C1(n18258), .C2(n18257), .A(
        n18256), .ZN(n18261) );
  OAI211_X1 U21233 ( .C1(n18263), .C2(n18907), .A(n18262), .B(n18261), .ZN(
        P3_U2862) );
  AOI211_X1 U21234 ( .C1(n18265), .C2(n18264), .A(n18889), .B(n18930), .ZN(
        n18774) );
  OAI21_X1 U21235 ( .B1(n18774), .B2(n18322), .A(n18271), .ZN(n18266) );
  OAI221_X1 U21236 ( .B1(n18273), .B2(n18267), .C1(n18273), .C2(n18271), .A(
        n18266), .ZN(P3_U2863) );
  INV_X1 U21237 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18758) );
  NAND2_X1 U21238 ( .A1(n18746), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18550) );
  INV_X1 U21239 ( .A(n18550), .ZN(n18571) );
  NAND2_X1 U21240 ( .A1(n18758), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18453) );
  INV_X1 U21241 ( .A(n18453), .ZN(n18455) );
  NOR2_X1 U21242 ( .A1(n18571), .A2(n18455), .ZN(n18268) );
  OAI22_X1 U21243 ( .A1(n18270), .A2(n18758), .B1(n18269), .B2(n18268), .ZN(
        P3_U2866) );
  NOR2_X1 U21244 ( .A1(n21010), .A2(n18271), .ZN(P3_U2867) );
  NAND2_X1 U21245 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18548) );
  INV_X1 U21246 ( .A(n18548), .ZN(n18729) );
  NOR2_X1 U21247 ( .A1(n18746), .A2(n18758), .ZN(n18274) );
  NAND2_X1 U21248 ( .A1(n18729), .A2(n18274), .ZN(n18713) );
  NAND2_X1 U21249 ( .A1(n18725), .A2(n18273), .ZN(n18727) );
  NOR2_X1 U21250 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18368) );
  INV_X1 U21251 ( .A(n18368), .ZN(n18409) );
  NOR2_X1 U21252 ( .A1(n18727), .A2(n18409), .ZN(n18356) );
  NOR2_X1 U21253 ( .A1(n18360), .A2(n18384), .ZN(n18342) );
  NAND2_X1 U21254 ( .A1(n18576), .A2(n18272), .ZN(n18619) );
  INV_X1 U21255 ( .A(n18274), .ZN(n18278) );
  NOR2_X1 U21256 ( .A1(n18725), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18525) );
  NOR2_X1 U21257 ( .A1(n18273), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18501) );
  NOR2_X1 U21258 ( .A1(n18525), .A2(n18501), .ZN(n18574) );
  OR2_X1 U21259 ( .A1(n18278), .A2(n18574), .ZN(n18622) );
  OAI22_X1 U21260 ( .A1(n18342), .A2(n18619), .B1(n18365), .B2(n18622), .ZN(
        n18320) );
  NOR2_X2 U21261 ( .A1(n18365), .A2(n19271), .ZN(n18658) );
  AND2_X1 U21262 ( .A1(n18274), .A2(n18525), .ZN(n18652) );
  AND2_X1 U21263 ( .A1(n18576), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18657) );
  INV_X1 U21264 ( .A(n18777), .ZN(n18781) );
  NOR2_X1 U21265 ( .A1(n18781), .A2(n18342), .ZN(n18314) );
  AOI22_X1 U21266 ( .A1(n18658), .A2(n18652), .B1(n18657), .B2(n18314), .ZN(
        n18281) );
  NAND2_X1 U21267 ( .A1(n18276), .A2(n18275), .ZN(n18315) );
  NOR2_X1 U21268 ( .A1(n18277), .A2(n18315), .ZN(n18623) );
  NOR2_X1 U21269 ( .A1(n18278), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18661) );
  NAND2_X1 U21270 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18661), .ZN(
        n18618) );
  INV_X1 U21271 ( .A(n18618), .ZN(n18706) );
  INV_X1 U21272 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18279) );
  NOR2_X2 U21273 ( .A1(n18279), .A2(n18365), .ZN(n18663) );
  AOI22_X1 U21274 ( .A1(n18384), .A2(n18623), .B1(n18706), .B2(n18663), .ZN(
        n18280) );
  OAI211_X1 U21275 ( .C1(n18282), .C2(n18320), .A(n18281), .B(n18280), .ZN(
        P3_U2868) );
  AND2_X1 U21276 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18662), .ZN(n18668) );
  AND2_X1 U21277 ( .A1(n18576), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18667) );
  AOI22_X1 U21278 ( .A1(n18706), .A2(n18668), .B1(n18314), .B2(n18667), .ZN(
        n18284) );
  NOR2_X1 U21279 ( .A1(n9961), .A2(n18315), .ZN(n18626) );
  AND2_X1 U21280 ( .A1(n18662), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18669) );
  AOI22_X1 U21281 ( .A1(n18356), .A2(n18626), .B1(n18652), .B2(n18669), .ZN(
        n18283) );
  OAI211_X1 U21282 ( .C1(n18285), .C2(n18320), .A(n18284), .B(n18283), .ZN(
        P3_U2869) );
  AND2_X1 U21283 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18662), .ZN(n18675) );
  NOR2_X2 U21284 ( .A1(n18367), .A2(n18286), .ZN(n18673) );
  AOI22_X1 U21285 ( .A1(n18706), .A2(n18675), .B1(n18314), .B2(n18673), .ZN(
        n18290) );
  NOR2_X1 U21286 ( .A1(n18287), .A2(n18315), .ZN(n18630) );
  INV_X1 U21287 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18288) );
  NOR2_X2 U21288 ( .A1(n18365), .A2(n18288), .ZN(n18674) );
  AOI22_X1 U21289 ( .A1(n18356), .A2(n18630), .B1(n18652), .B2(n18674), .ZN(
        n18289) );
  OAI211_X1 U21290 ( .C1(n18291), .C2(n18320), .A(n18290), .B(n18289), .ZN(
        P3_U2870) );
  INV_X1 U21291 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18292) );
  NOR2_X2 U21292 ( .A1(n18365), .A2(n18292), .ZN(n18680) );
  NOR2_X2 U21293 ( .A1(n18367), .A2(n18293), .ZN(n18679) );
  AOI22_X1 U21294 ( .A1(n18652), .A2(n18680), .B1(n18314), .B2(n18679), .ZN(
        n18296) );
  NOR2_X1 U21295 ( .A1(n18294), .A2(n18315), .ZN(n18633) );
  AOI22_X1 U21296 ( .A1(n18356), .A2(n18633), .B1(n18706), .B2(n18681), .ZN(
        n18295) );
  OAI211_X1 U21297 ( .C1(n21155), .C2(n18320), .A(n18296), .B(n18295), .ZN(
        P3_U2871) );
  AND2_X1 U21298 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18662), .ZN(n18685) );
  NOR2_X2 U21299 ( .A1(n18367), .A2(n18297), .ZN(n18686) );
  AOI22_X1 U21300 ( .A1(n18706), .A2(n18685), .B1(n18314), .B2(n18686), .ZN(
        n18301) );
  NOR2_X1 U21301 ( .A1(n18298), .A2(n18315), .ZN(n18637) );
  INV_X1 U21302 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18299) );
  NOR2_X2 U21303 ( .A1(n18365), .A2(n18299), .ZN(n18687) );
  AOI22_X1 U21304 ( .A1(n18356), .A2(n18637), .B1(n18652), .B2(n18687), .ZN(
        n18300) );
  OAI211_X1 U21305 ( .C1(n18302), .C2(n18320), .A(n18301), .B(n18300), .ZN(
        P3_U2872) );
  AND2_X1 U21306 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18662), .ZN(n18691) );
  NOR2_X2 U21307 ( .A1(n18367), .A2(n21139), .ZN(n18692) );
  AOI22_X1 U21308 ( .A1(n18706), .A2(n18691), .B1(n18314), .B2(n18692), .ZN(
        n18306) );
  NOR2_X1 U21309 ( .A1(n18303), .A2(n18315), .ZN(n18641) );
  INV_X1 U21310 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18304) );
  NOR2_X2 U21311 ( .A1(n18365), .A2(n18304), .ZN(n18693) );
  AOI22_X1 U21312 ( .A1(n18356), .A2(n18641), .B1(n18652), .B2(n18693), .ZN(
        n18305) );
  OAI211_X1 U21313 ( .C1(n18307), .C2(n18320), .A(n18306), .B(n18305), .ZN(
        P3_U2873) );
  NOR2_X2 U21314 ( .A1(n18308), .A2(n18365), .ZN(n18697) );
  NOR2_X2 U21315 ( .A1(n18367), .A2(n18309), .ZN(n18698) );
  AOI22_X1 U21316 ( .A1(n18706), .A2(n18697), .B1(n18314), .B2(n18698), .ZN(
        n18312) );
  NOR2_X1 U21317 ( .A1(n18310), .A2(n18315), .ZN(n18645) );
  NOR2_X2 U21318 ( .A1(n18365), .A2(n19306), .ZN(n18699) );
  AOI22_X1 U21319 ( .A1(n18384), .A2(n18645), .B1(n18652), .B2(n18699), .ZN(
        n18311) );
  OAI211_X1 U21320 ( .C1(n18313), .C2(n18320), .A(n18312), .B(n18311), .ZN(
        P3_U2874) );
  NOR2_X2 U21321 ( .A1(n18365), .A2(n20992), .ZN(n18708) );
  NOR2_X2 U21322 ( .A1(n20954), .A2(n18367), .ZN(n18704) );
  AOI22_X1 U21323 ( .A1(n18706), .A2(n18708), .B1(n18314), .B2(n18704), .ZN(
        n18319) );
  NOR2_X1 U21324 ( .A1(n18316), .A2(n18315), .ZN(n18651) );
  INV_X1 U21325 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18317) );
  NOR2_X2 U21326 ( .A1(n18317), .A2(n18365), .ZN(n18705) );
  AOI22_X1 U21327 ( .A1(n18384), .A2(n18651), .B1(n18652), .B2(n18705), .ZN(
        n18318) );
  OAI211_X1 U21328 ( .C1(n18321), .C2(n18320), .A(n18319), .B(n18318), .ZN(
        P3_U2875) );
  NAND2_X1 U21329 ( .A1(n18368), .A2(n18501), .ZN(n18341) );
  NAND2_X1 U21330 ( .A1(n18725), .A2(n18777), .ZN(n18502) );
  NOR2_X1 U21331 ( .A1(n18409), .A2(n18502), .ZN(n18337) );
  AOI22_X1 U21332 ( .A1(n18663), .A2(n18652), .B1(n18657), .B2(n18337), .ZN(
        n18324) );
  NOR2_X1 U21333 ( .A1(n18758), .A2(n18503), .ZN(n18659) );
  NOR2_X1 U21334 ( .A1(n18367), .A2(n18322), .ZN(n18660) );
  AND2_X1 U21335 ( .A1(n18725), .A2(n18660), .ZN(n18410) );
  AOI22_X1 U21336 ( .A1(n18662), .A2(n18659), .B1(n18368), .B2(n18410), .ZN(
        n18338) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18338), .B1(
        n18360), .B2(n18658), .ZN(n18323) );
  OAI211_X1 U21338 ( .C1(n18666), .C2(n18341), .A(n18324), .B(n18323), .ZN(
        P3_U2876) );
  AOI22_X1 U21339 ( .A1(n18652), .A2(n18668), .B1(n18667), .B2(n18337), .ZN(
        n18326) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18338), .B1(
        n18360), .B2(n18669), .ZN(n18325) );
  OAI211_X1 U21341 ( .C1(n18672), .C2(n18341), .A(n18326), .B(n18325), .ZN(
        P3_U2877) );
  INV_X1 U21342 ( .A(n18630), .ZN(n18678) );
  AOI22_X1 U21343 ( .A1(n18360), .A2(n18674), .B1(n18673), .B2(n18337), .ZN(
        n18328) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18338), .B1(
        n18652), .B2(n18675), .ZN(n18327) );
  OAI211_X1 U21345 ( .C1(n18678), .C2(n18341), .A(n18328), .B(n18327), .ZN(
        P3_U2878) );
  INV_X1 U21346 ( .A(n18633), .ZN(n18684) );
  AOI22_X1 U21347 ( .A1(n18652), .A2(n18681), .B1(n18679), .B2(n18337), .ZN(
        n18330) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18338), .B1(
        n18360), .B2(n18680), .ZN(n18329) );
  OAI211_X1 U21349 ( .C1(n18684), .C2(n18341), .A(n18330), .B(n18329), .ZN(
        P3_U2879) );
  INV_X1 U21350 ( .A(n18637), .ZN(n18690) );
  AOI22_X1 U21351 ( .A1(n18652), .A2(n18685), .B1(n18686), .B2(n18337), .ZN(
        n18332) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18338), .B1(
        n18360), .B2(n18687), .ZN(n18331) );
  OAI211_X1 U21353 ( .C1(n18690), .C2(n18341), .A(n18332), .B(n18331), .ZN(
        P3_U2880) );
  INV_X1 U21354 ( .A(n18641), .ZN(n18696) );
  AOI22_X1 U21355 ( .A1(n18652), .A2(n18691), .B1(n18692), .B2(n18337), .ZN(
        n18334) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18338), .B1(
        n18360), .B2(n18693), .ZN(n18333) );
  OAI211_X1 U21357 ( .C1(n18696), .C2(n18341), .A(n18334), .B(n18333), .ZN(
        P3_U2881) );
  AOI22_X1 U21358 ( .A1(n18360), .A2(n18699), .B1(n18698), .B2(n18337), .ZN(
        n18336) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18338), .B1(
        n18652), .B2(n18697), .ZN(n18335) );
  OAI211_X1 U21360 ( .C1(n18702), .C2(n18341), .A(n18336), .B(n18335), .ZN(
        P3_U2882) );
  INV_X1 U21361 ( .A(n18651), .ZN(n18712) );
  AOI22_X1 U21362 ( .A1(n18652), .A2(n18708), .B1(n18704), .B2(n18337), .ZN(
        n18340) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18338), .B1(
        n18360), .B2(n18705), .ZN(n18339) );
  OAI211_X1 U21364 ( .C1(n18712), .C2(n18341), .A(n18340), .B(n18339), .ZN(
        P3_U2883) );
  NAND2_X1 U21365 ( .A1(n18368), .A2(n18525), .ZN(n18364) );
  INV_X1 U21366 ( .A(n18341), .ZN(n18404) );
  NOR2_X1 U21367 ( .A1(n18404), .A2(n18426), .ZN(n18388) );
  NOR2_X1 U21368 ( .A1(n18781), .A2(n18388), .ZN(n18359) );
  AOI22_X1 U21369 ( .A1(n18360), .A2(n18663), .B1(n18657), .B2(n18359), .ZN(
        n18345) );
  AOI221_X1 U21370 ( .B1(n18388), .B2(n18620), .C1(n18388), .C2(n18342), .A(
        n18619), .ZN(n18343) );
  INV_X1 U21371 ( .A(n18343), .ZN(n18361) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18361), .B1(
        n18356), .B2(n18658), .ZN(n18344) );
  OAI211_X1 U21373 ( .C1(n18666), .C2(n18364), .A(n18345), .B(n18344), .ZN(
        P3_U2884) );
  AOI22_X1 U21374 ( .A1(n18384), .A2(n18669), .B1(n18667), .B2(n18359), .ZN(
        n18347) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18361), .B1(
        n18360), .B2(n18668), .ZN(n18346) );
  OAI211_X1 U21376 ( .C1(n18672), .C2(n18364), .A(n18347), .B(n18346), .ZN(
        P3_U2885) );
  AOI22_X1 U21377 ( .A1(n18360), .A2(n18675), .B1(n18673), .B2(n18359), .ZN(
        n18349) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18361), .B1(
        n18356), .B2(n18674), .ZN(n18348) );
  OAI211_X1 U21379 ( .C1(n18678), .C2(n18364), .A(n18349), .B(n18348), .ZN(
        P3_U2886) );
  AOI22_X1 U21380 ( .A1(n18384), .A2(n18680), .B1(n18679), .B2(n18359), .ZN(
        n18351) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18361), .B1(
        n18360), .B2(n18681), .ZN(n18350) );
  OAI211_X1 U21382 ( .C1(n18684), .C2(n18364), .A(n18351), .B(n18350), .ZN(
        P3_U2887) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18361), .B1(
        n18686), .B2(n18359), .ZN(n18353) );
  AOI22_X1 U21384 ( .A1(n18360), .A2(n18685), .B1(n18356), .B2(n18687), .ZN(
        n18352) );
  OAI211_X1 U21385 ( .C1(n18690), .C2(n18364), .A(n18353), .B(n18352), .ZN(
        P3_U2888) );
  AOI22_X1 U21386 ( .A1(n18384), .A2(n18693), .B1(n18692), .B2(n18359), .ZN(
        n18355) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18361), .B1(
        n18360), .B2(n18691), .ZN(n18354) );
  OAI211_X1 U21388 ( .C1(n18696), .C2(n18364), .A(n18355), .B(n18354), .ZN(
        P3_U2889) );
  AOI22_X1 U21389 ( .A1(n18360), .A2(n18697), .B1(n18698), .B2(n18359), .ZN(
        n18358) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18361), .B1(
        n18356), .B2(n18699), .ZN(n18357) );
  OAI211_X1 U21391 ( .C1(n18702), .C2(n18364), .A(n18358), .B(n18357), .ZN(
        P3_U2890) );
  AOI22_X1 U21392 ( .A1(n18384), .A2(n18705), .B1(n18704), .B2(n18359), .ZN(
        n18363) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18361), .B1(
        n18360), .B2(n18708), .ZN(n18362) );
  OAI211_X1 U21394 ( .C1(n18712), .C2(n18364), .A(n18363), .B(n18362), .ZN(
        P3_U2891) );
  NOR2_X2 U21395 ( .A1(n18548), .A2(n18409), .ZN(n18449) );
  AOI22_X1 U21396 ( .A1(n18384), .A2(n18663), .B1(n18657), .B2(n18383), .ZN(
        n18370) );
  OAI21_X1 U21397 ( .B1(n18367), .B2(n18366), .A(n18365), .ZN(n18454) );
  NAND2_X1 U21398 ( .A1(n18368), .A2(n18454), .ZN(n18385) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18385), .B1(
        n18658), .B2(n18404), .ZN(n18369) );
  OAI211_X1 U21400 ( .C1(n18666), .C2(n18432), .A(n18370), .B(n18369), .ZN(
        P3_U2892) );
  AOI22_X1 U21401 ( .A1(n18384), .A2(n18668), .B1(n18667), .B2(n18383), .ZN(
        n18372) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18385), .B1(
        n18669), .B2(n18404), .ZN(n18371) );
  OAI211_X1 U21403 ( .C1(n18672), .C2(n18432), .A(n18372), .B(n18371), .ZN(
        P3_U2893) );
  AOI22_X1 U21404 ( .A1(n18384), .A2(n18675), .B1(n18673), .B2(n18383), .ZN(
        n18374) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18385), .B1(
        n18674), .B2(n18404), .ZN(n18373) );
  OAI211_X1 U21406 ( .C1(n18678), .C2(n18432), .A(n18374), .B(n18373), .ZN(
        P3_U2894) );
  AOI22_X1 U21407 ( .A1(n18680), .A2(n18404), .B1(n18679), .B2(n18383), .ZN(
        n18376) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18385), .B1(
        n18384), .B2(n18681), .ZN(n18375) );
  OAI211_X1 U21409 ( .C1(n18684), .C2(n18432), .A(n18376), .B(n18375), .ZN(
        P3_U2895) );
  AOI22_X1 U21410 ( .A1(n18384), .A2(n18685), .B1(n18686), .B2(n18383), .ZN(
        n18378) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18385), .B1(
        n18687), .B2(n18404), .ZN(n18377) );
  OAI211_X1 U21412 ( .C1(n18690), .C2(n18432), .A(n18378), .B(n18377), .ZN(
        P3_U2896) );
  AOI22_X1 U21413 ( .A1(n18693), .A2(n18404), .B1(n18692), .B2(n18383), .ZN(
        n18380) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18385), .B1(
        n18384), .B2(n18691), .ZN(n18379) );
  OAI211_X1 U21415 ( .C1(n18696), .C2(n18432), .A(n18380), .B(n18379), .ZN(
        P3_U2897) );
  AOI22_X1 U21416 ( .A1(n18699), .A2(n18404), .B1(n18698), .B2(n18383), .ZN(
        n18382) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18385), .B1(
        n18384), .B2(n18697), .ZN(n18381) );
  OAI211_X1 U21418 ( .C1(n18702), .C2(n18432), .A(n18382), .B(n18381), .ZN(
        P3_U2898) );
  AOI22_X1 U21419 ( .A1(n18705), .A2(n18404), .B1(n18704), .B2(n18383), .ZN(
        n18387) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18385), .B1(
        n18384), .B2(n18708), .ZN(n18386) );
  OAI211_X1 U21421 ( .C1(n18712), .C2(n18432), .A(n18387), .B(n18386), .ZN(
        P3_U2899) );
  NOR2_X2 U21422 ( .A1(n18727), .A2(n18453), .ZN(n18471) );
  AOI21_X1 U21423 ( .B1(n18432), .B2(n18431), .A(n18781), .ZN(n18405) );
  AOI22_X1 U21424 ( .A1(n18658), .A2(n18426), .B1(n18657), .B2(n18405), .ZN(
        n18391) );
  AOI221_X1 U21425 ( .B1(n18388), .B2(n18432), .C1(n18620), .C2(n18432), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18389) );
  OAI21_X1 U21426 ( .B1(n18471), .B2(n18389), .A(n18576), .ZN(n18406) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18406), .B1(
        n18663), .B2(n18404), .ZN(n18390) );
  OAI211_X1 U21428 ( .C1(n18666), .C2(n18431), .A(n18391), .B(n18390), .ZN(
        P3_U2900) );
  AOI22_X1 U21429 ( .A1(n18669), .A2(n18426), .B1(n18667), .B2(n18405), .ZN(
        n18393) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18406), .B1(
        n18668), .B2(n18404), .ZN(n18392) );
  OAI211_X1 U21431 ( .C1(n18672), .C2(n18431), .A(n18393), .B(n18392), .ZN(
        P3_U2901) );
  AOI22_X1 U21432 ( .A1(n18675), .A2(n18404), .B1(n18673), .B2(n18405), .ZN(
        n18395) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18406), .B1(
        n18674), .B2(n18426), .ZN(n18394) );
  OAI211_X1 U21434 ( .C1(n18678), .C2(n18431), .A(n18395), .B(n18394), .ZN(
        P3_U2902) );
  AOI22_X1 U21435 ( .A1(n18680), .A2(n18426), .B1(n18679), .B2(n18405), .ZN(
        n18397) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18406), .B1(
        n18681), .B2(n18404), .ZN(n18396) );
  OAI211_X1 U21437 ( .C1(n18684), .C2(n18431), .A(n18397), .B(n18396), .ZN(
        P3_U2903) );
  AOI22_X1 U21438 ( .A1(n18686), .A2(n18405), .B1(n18685), .B2(n18404), .ZN(
        n18399) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18406), .B1(
        n18687), .B2(n18426), .ZN(n18398) );
  OAI211_X1 U21440 ( .C1(n18690), .C2(n18431), .A(n18399), .B(n18398), .ZN(
        P3_U2904) );
  AOI22_X1 U21441 ( .A1(n18692), .A2(n18405), .B1(n18691), .B2(n18404), .ZN(
        n18401) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18406), .B1(
        n18693), .B2(n18426), .ZN(n18400) );
  OAI211_X1 U21443 ( .C1(n18696), .C2(n18431), .A(n18401), .B(n18400), .ZN(
        P3_U2905) );
  AOI22_X1 U21444 ( .A1(n18699), .A2(n18426), .B1(n18698), .B2(n18405), .ZN(
        n18403) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18406), .B1(
        n18697), .B2(n18404), .ZN(n18402) );
  OAI211_X1 U21446 ( .C1(n18702), .C2(n18431), .A(n18403), .B(n18402), .ZN(
        P3_U2906) );
  AOI22_X1 U21447 ( .A1(n18704), .A2(n18405), .B1(n18708), .B2(n18404), .ZN(
        n18408) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18406), .B1(
        n18705), .B2(n18426), .ZN(n18407) );
  OAI211_X1 U21449 ( .C1(n18712), .C2(n18431), .A(n18408), .B(n18407), .ZN(
        P3_U2907) );
  NAND2_X1 U21450 ( .A1(n18455), .A2(n18501), .ZN(n18456) );
  NOR2_X1 U21451 ( .A1(n18453), .A2(n18502), .ZN(n18427) );
  AOI22_X1 U21452 ( .A1(n18663), .A2(n18426), .B1(n18657), .B2(n18427), .ZN(
        n18413) );
  NOR2_X1 U21453 ( .A1(n18725), .A2(n18409), .ZN(n18411) );
  AOI22_X1 U21454 ( .A1(n18662), .A2(n18411), .B1(n18455), .B2(n18410), .ZN(
        n18428) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18428), .B1(
        n18658), .B2(n18449), .ZN(n18412) );
  OAI211_X1 U21456 ( .C1(n18666), .C2(n18456), .A(n18413), .B(n18412), .ZN(
        P3_U2908) );
  AOI22_X1 U21457 ( .A1(n18668), .A2(n18426), .B1(n18667), .B2(n18427), .ZN(
        n18415) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18428), .B1(
        n18669), .B2(n18449), .ZN(n18414) );
  OAI211_X1 U21459 ( .C1(n18672), .C2(n18456), .A(n18415), .B(n18414), .ZN(
        P3_U2909) );
  AOI22_X1 U21460 ( .A1(n18674), .A2(n18449), .B1(n18673), .B2(n18427), .ZN(
        n18417) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18428), .B1(
        n18675), .B2(n18426), .ZN(n18416) );
  OAI211_X1 U21462 ( .C1(n18678), .C2(n18456), .A(n18417), .B(n18416), .ZN(
        P3_U2910) );
  AOI22_X1 U21463 ( .A1(n18681), .A2(n18426), .B1(n18679), .B2(n18427), .ZN(
        n18419) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18428), .B1(
        n18680), .B2(n18449), .ZN(n18418) );
  OAI211_X1 U21465 ( .C1(n18684), .C2(n18456), .A(n18419), .B(n18418), .ZN(
        P3_U2911) );
  AOI22_X1 U21466 ( .A1(n18687), .A2(n18449), .B1(n18686), .B2(n18427), .ZN(
        n18421) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18428), .B1(
        n18685), .B2(n18426), .ZN(n18420) );
  OAI211_X1 U21468 ( .C1(n18690), .C2(n18456), .A(n18421), .B(n18420), .ZN(
        P3_U2912) );
  AOI22_X1 U21469 ( .A1(n18693), .A2(n18449), .B1(n18692), .B2(n18427), .ZN(
        n18423) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18428), .B1(
        n18691), .B2(n18426), .ZN(n18422) );
  OAI211_X1 U21471 ( .C1(n18696), .C2(n18456), .A(n18423), .B(n18422), .ZN(
        P3_U2913) );
  AOI22_X1 U21472 ( .A1(n18698), .A2(n18427), .B1(n18697), .B2(n18426), .ZN(
        n18425) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18428), .B1(
        n18699), .B2(n18449), .ZN(n18424) );
  OAI211_X1 U21474 ( .C1(n18702), .C2(n18456), .A(n18425), .B(n18424), .ZN(
        P3_U2914) );
  AOI22_X1 U21475 ( .A1(n18704), .A2(n18427), .B1(n18708), .B2(n18426), .ZN(
        n18430) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18428), .B1(
        n18705), .B2(n18449), .ZN(n18429) );
  OAI211_X1 U21477 ( .C1(n18712), .C2(n18456), .A(n18430), .B(n18429), .ZN(
        P3_U2915) );
  NAND2_X1 U21478 ( .A1(n18455), .A2(n18525), .ZN(n18480) );
  NAND2_X1 U21479 ( .A1(n18456), .A2(n18480), .ZN(n18478) );
  AND2_X1 U21480 ( .A1(n18777), .A2(n18478), .ZN(n18448) );
  AOI22_X1 U21481 ( .A1(n18663), .A2(n18449), .B1(n18657), .B2(n18448), .ZN(
        n18435) );
  NAND2_X1 U21482 ( .A1(n18432), .A2(n18431), .ZN(n18433) );
  INV_X1 U21483 ( .A(n18619), .ZN(n18477) );
  OAI221_X1 U21484 ( .B1(n18478), .B2(n18572), .C1(n18478), .C2(n18433), .A(
        n18477), .ZN(n18450) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18450), .B1(
        n18658), .B2(n18471), .ZN(n18434) );
  OAI211_X1 U21486 ( .C1(n18666), .C2(n18480), .A(n18435), .B(n18434), .ZN(
        P3_U2916) );
  AOI22_X1 U21487 ( .A1(n18669), .A2(n18471), .B1(n18667), .B2(n18448), .ZN(
        n18437) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18450), .B1(
        n18668), .B2(n18449), .ZN(n18436) );
  OAI211_X1 U21489 ( .C1(n18672), .C2(n18480), .A(n18437), .B(n18436), .ZN(
        P3_U2917) );
  AOI22_X1 U21490 ( .A1(n18674), .A2(n18471), .B1(n18673), .B2(n18448), .ZN(
        n18439) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18450), .B1(
        n18675), .B2(n18449), .ZN(n18438) );
  OAI211_X1 U21492 ( .C1(n18678), .C2(n18480), .A(n18439), .B(n18438), .ZN(
        P3_U2918) );
  AOI22_X1 U21493 ( .A1(n18680), .A2(n18471), .B1(n18679), .B2(n18448), .ZN(
        n18441) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18450), .B1(
        n18681), .B2(n18449), .ZN(n18440) );
  OAI211_X1 U21495 ( .C1(n18684), .C2(n18480), .A(n18441), .B(n18440), .ZN(
        P3_U2919) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18450), .B1(
        n18686), .B2(n18448), .ZN(n18443) );
  AOI22_X1 U21497 ( .A1(n18687), .A2(n18471), .B1(n18685), .B2(n18449), .ZN(
        n18442) );
  OAI211_X1 U21498 ( .C1(n18690), .C2(n18480), .A(n18443), .B(n18442), .ZN(
        P3_U2920) );
  AOI22_X1 U21499 ( .A1(n18692), .A2(n18448), .B1(n18691), .B2(n18449), .ZN(
        n18445) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18450), .B1(
        n18693), .B2(n18471), .ZN(n18444) );
  OAI211_X1 U21501 ( .C1(n18696), .C2(n18480), .A(n18445), .B(n18444), .ZN(
        P3_U2921) );
  AOI22_X1 U21502 ( .A1(n18698), .A2(n18448), .B1(n18697), .B2(n18449), .ZN(
        n18447) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18450), .B1(
        n18699), .B2(n18471), .ZN(n18446) );
  OAI211_X1 U21504 ( .C1(n18702), .C2(n18480), .A(n18447), .B(n18446), .ZN(
        P3_U2922) );
  AOI22_X1 U21505 ( .A1(n18705), .A2(n18471), .B1(n18704), .B2(n18448), .ZN(
        n18452) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18450), .B1(
        n18708), .B2(n18449), .ZN(n18451) );
  OAI211_X1 U21507 ( .C1(n18712), .C2(n18480), .A(n18452), .B(n18451), .ZN(
        P3_U2923) );
  NOR2_X2 U21508 ( .A1(n18548), .A2(n18453), .ZN(n18542) );
  AOI22_X1 U21509 ( .A1(n18663), .A2(n18471), .B1(n18657), .B2(n18472), .ZN(
        n18458) );
  NAND2_X1 U21510 ( .A1(n18455), .A2(n18454), .ZN(n18473) );
  INV_X1 U21511 ( .A(n18456), .ZN(n18495) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18473), .B1(
        n18658), .B2(n18495), .ZN(n18457) );
  OAI211_X1 U21513 ( .C1(n18666), .C2(n18476), .A(n18458), .B(n18457), .ZN(
        P3_U2924) );
  AOI22_X1 U21514 ( .A1(n18669), .A2(n18495), .B1(n18667), .B2(n18472), .ZN(
        n18460) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18473), .B1(
        n18668), .B2(n18471), .ZN(n18459) );
  OAI211_X1 U21516 ( .C1(n18672), .C2(n18476), .A(n18460), .B(n18459), .ZN(
        P3_U2925) );
  AOI22_X1 U21517 ( .A1(n18674), .A2(n18495), .B1(n18673), .B2(n18472), .ZN(
        n18462) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18473), .B1(
        n18675), .B2(n18471), .ZN(n18461) );
  OAI211_X1 U21519 ( .C1(n18678), .C2(n18476), .A(n18462), .B(n18461), .ZN(
        P3_U2926) );
  AOI22_X1 U21520 ( .A1(n18680), .A2(n18495), .B1(n18679), .B2(n18472), .ZN(
        n18464) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18473), .B1(
        n18681), .B2(n18471), .ZN(n18463) );
  OAI211_X1 U21522 ( .C1(n18684), .C2(n18476), .A(n18464), .B(n18463), .ZN(
        P3_U2927) );
  AOI22_X1 U21523 ( .A1(n18686), .A2(n18472), .B1(n18685), .B2(n18471), .ZN(
        n18466) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18473), .B1(
        n18687), .B2(n18495), .ZN(n18465) );
  OAI211_X1 U21525 ( .C1(n18690), .C2(n18476), .A(n18466), .B(n18465), .ZN(
        P3_U2928) );
  AOI22_X1 U21526 ( .A1(n18693), .A2(n18495), .B1(n18692), .B2(n18472), .ZN(
        n18468) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18473), .B1(
        n18691), .B2(n18471), .ZN(n18467) );
  OAI211_X1 U21528 ( .C1(n18696), .C2(n18476), .A(n18468), .B(n18467), .ZN(
        P3_U2929) );
  AOI22_X1 U21529 ( .A1(n18699), .A2(n18495), .B1(n18698), .B2(n18472), .ZN(
        n18470) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18473), .B1(
        n18697), .B2(n18471), .ZN(n18469) );
  OAI211_X1 U21531 ( .C1(n18702), .C2(n18476), .A(n18470), .B(n18469), .ZN(
        P3_U2930) );
  AOI22_X1 U21532 ( .A1(n18704), .A2(n18472), .B1(n18708), .B2(n18471), .ZN(
        n18475) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18473), .B1(
        n18705), .B2(n18495), .ZN(n18474) );
  OAI211_X1 U21534 ( .C1(n18712), .C2(n18476), .A(n18475), .B(n18474), .ZN(
        P3_U2931) );
  NOR2_X2 U21535 ( .A1(n18727), .A2(n18550), .ZN(n18566) );
  NAND2_X1 U21536 ( .A1(n18476), .A2(n18500), .ZN(n18479) );
  OAI221_X1 U21537 ( .B1(n18479), .B2(n18572), .C1(n18479), .C2(n18478), .A(
        n18477), .ZN(n18497) );
  INV_X1 U21538 ( .A(n18479), .ZN(n18526) );
  NOR2_X1 U21539 ( .A1(n18781), .A2(n18526), .ZN(n18496) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18497), .B1(
        n18657), .B2(n18496), .ZN(n18482) );
  AOI22_X1 U21541 ( .A1(n18663), .A2(n18495), .B1(n18658), .B2(n18520), .ZN(
        n18481) );
  OAI211_X1 U21542 ( .C1(n18666), .C2(n18500), .A(n18482), .B(n18481), .ZN(
        P3_U2932) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18497), .B1(
        n18667), .B2(n18496), .ZN(n18484) );
  AOI22_X1 U21544 ( .A1(n18669), .A2(n18520), .B1(n18668), .B2(n18495), .ZN(
        n18483) );
  OAI211_X1 U21545 ( .C1(n18672), .C2(n18500), .A(n18484), .B(n18483), .ZN(
        P3_U2933) );
  AOI22_X1 U21546 ( .A1(n18675), .A2(n18495), .B1(n18673), .B2(n18496), .ZN(
        n18486) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18497), .B1(
        n18674), .B2(n18520), .ZN(n18485) );
  OAI211_X1 U21548 ( .C1(n18678), .C2(n18500), .A(n18486), .B(n18485), .ZN(
        P3_U2934) );
  AOI22_X1 U21549 ( .A1(n18680), .A2(n18520), .B1(n18679), .B2(n18496), .ZN(
        n18488) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18497), .B1(
        n18681), .B2(n18495), .ZN(n18487) );
  OAI211_X1 U21551 ( .C1(n18684), .C2(n18500), .A(n18488), .B(n18487), .ZN(
        P3_U2935) );
  AOI22_X1 U21552 ( .A1(n18686), .A2(n18496), .B1(n18685), .B2(n18495), .ZN(
        n18490) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18497), .B1(
        n18687), .B2(n18520), .ZN(n18489) );
  OAI211_X1 U21554 ( .C1(n18690), .C2(n18500), .A(n18490), .B(n18489), .ZN(
        P3_U2936) );
  AOI22_X1 U21555 ( .A1(n18692), .A2(n18496), .B1(n18691), .B2(n18495), .ZN(
        n18492) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18497), .B1(
        n18693), .B2(n18520), .ZN(n18491) );
  OAI211_X1 U21557 ( .C1(n18696), .C2(n18500), .A(n18492), .B(n18491), .ZN(
        P3_U2937) );
  AOI22_X1 U21558 ( .A1(n18698), .A2(n18496), .B1(n18697), .B2(n18495), .ZN(
        n18494) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18497), .B1(
        n18699), .B2(n18520), .ZN(n18493) );
  OAI211_X1 U21560 ( .C1(n18702), .C2(n18500), .A(n18494), .B(n18493), .ZN(
        P3_U2938) );
  AOI22_X1 U21561 ( .A1(n18704), .A2(n18496), .B1(n18708), .B2(n18495), .ZN(
        n18499) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18497), .B1(
        n18705), .B2(n18520), .ZN(n18498) );
  OAI211_X1 U21563 ( .C1(n18712), .C2(n18500), .A(n18499), .B(n18498), .ZN(
        P3_U2939) );
  NAND2_X1 U21564 ( .A1(n18571), .A2(n18501), .ZN(n18549) );
  NOR2_X1 U21565 ( .A1(n18550), .A2(n18502), .ZN(n18521) );
  AOI22_X1 U21566 ( .A1(n18663), .A2(n18520), .B1(n18657), .B2(n18521), .ZN(
        n18507) );
  NOR2_X1 U21567 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18503), .ZN(
        n18505) );
  NOR2_X1 U21568 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18550), .ZN(
        n18504) );
  AOI22_X1 U21569 ( .A1(n18662), .A2(n18505), .B1(n18660), .B2(n18504), .ZN(
        n18522) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18522), .B1(
        n18658), .B2(n18542), .ZN(n18506) );
  OAI211_X1 U21571 ( .C1(n18666), .C2(n18549), .A(n18507), .B(n18506), .ZN(
        P3_U2940) );
  AOI22_X1 U21572 ( .A1(n18668), .A2(n18520), .B1(n18667), .B2(n18521), .ZN(
        n18509) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18522), .B1(
        n18669), .B2(n18542), .ZN(n18508) );
  OAI211_X1 U21574 ( .C1(n18672), .C2(n18549), .A(n18509), .B(n18508), .ZN(
        P3_U2941) );
  AOI22_X1 U21575 ( .A1(n18675), .A2(n18520), .B1(n18673), .B2(n18521), .ZN(
        n18511) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18522), .B1(
        n18674), .B2(n18542), .ZN(n18510) );
  OAI211_X1 U21577 ( .C1(n18678), .C2(n18549), .A(n18511), .B(n18510), .ZN(
        P3_U2942) );
  AOI22_X1 U21578 ( .A1(n18681), .A2(n18520), .B1(n18679), .B2(n18521), .ZN(
        n18513) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18522), .B1(
        n18680), .B2(n18542), .ZN(n18512) );
  OAI211_X1 U21580 ( .C1(n18684), .C2(n18549), .A(n18513), .B(n18512), .ZN(
        P3_U2943) );
  AOI22_X1 U21581 ( .A1(n18686), .A2(n18521), .B1(n18685), .B2(n18520), .ZN(
        n18515) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18522), .B1(
        n18687), .B2(n18542), .ZN(n18514) );
  OAI211_X1 U21583 ( .C1(n18690), .C2(n18549), .A(n18515), .B(n18514), .ZN(
        P3_U2944) );
  AOI22_X1 U21584 ( .A1(n18692), .A2(n18521), .B1(n18691), .B2(n18520), .ZN(
        n18517) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18522), .B1(
        n18693), .B2(n18542), .ZN(n18516) );
  OAI211_X1 U21586 ( .C1(n18696), .C2(n18549), .A(n18517), .B(n18516), .ZN(
        P3_U2945) );
  AOI22_X1 U21587 ( .A1(n18698), .A2(n18521), .B1(n18697), .B2(n18520), .ZN(
        n18519) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18522), .B1(
        n18699), .B2(n18542), .ZN(n18518) );
  OAI211_X1 U21589 ( .C1(n18702), .C2(n18549), .A(n18519), .B(n18518), .ZN(
        P3_U2946) );
  AOI22_X1 U21590 ( .A1(n18704), .A2(n18521), .B1(n18708), .B2(n18520), .ZN(
        n18524) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18522), .B1(
        n18705), .B2(n18542), .ZN(n18523) );
  OAI211_X1 U21592 ( .C1(n18712), .C2(n18549), .A(n18524), .B(n18523), .ZN(
        P3_U2947) );
  NAND2_X1 U21593 ( .A1(n18571), .A2(n18525), .ZN(n18547) );
  AOI22_X1 U21594 ( .A1(n18663), .A2(n18542), .B1(n18657), .B2(n18543), .ZN(
        n18529) );
  AOI221_X1 U21595 ( .B1(n18526), .B2(n18549), .C1(n18620), .C2(n18549), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18527) );
  OAI21_X1 U21596 ( .B1(n18614), .B2(n18527), .A(n18576), .ZN(n18544) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18544), .B1(
        n18658), .B2(n18566), .ZN(n18528) );
  OAI211_X1 U21598 ( .C1(n18666), .C2(n18547), .A(n18529), .B(n18528), .ZN(
        P3_U2948) );
  AOI22_X1 U21599 ( .A1(n18669), .A2(n18566), .B1(n18667), .B2(n18543), .ZN(
        n18531) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18544), .B1(
        n18668), .B2(n18542), .ZN(n18530) );
  OAI211_X1 U21601 ( .C1(n18672), .C2(n18547), .A(n18531), .B(n18530), .ZN(
        P3_U2949) );
  AOI22_X1 U21602 ( .A1(n18674), .A2(n18566), .B1(n18673), .B2(n18543), .ZN(
        n18533) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18544), .B1(
        n18675), .B2(n18542), .ZN(n18532) );
  OAI211_X1 U21604 ( .C1(n18678), .C2(n18547), .A(n18533), .B(n18532), .ZN(
        P3_U2950) );
  AOI22_X1 U21605 ( .A1(n18681), .A2(n18542), .B1(n18679), .B2(n18543), .ZN(
        n18535) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18544), .B1(
        n18680), .B2(n18566), .ZN(n18534) );
  OAI211_X1 U21607 ( .C1(n18684), .C2(n18547), .A(n18535), .B(n18534), .ZN(
        P3_U2951) );
  AOI22_X1 U21608 ( .A1(n18687), .A2(n18566), .B1(n18686), .B2(n18543), .ZN(
        n18537) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18544), .B1(
        n18685), .B2(n18542), .ZN(n18536) );
  OAI211_X1 U21610 ( .C1(n18690), .C2(n18547), .A(n18537), .B(n18536), .ZN(
        P3_U2952) );
  AOI22_X1 U21611 ( .A1(n18692), .A2(n18543), .B1(n18691), .B2(n18542), .ZN(
        n18539) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18544), .B1(
        n18693), .B2(n18566), .ZN(n18538) );
  OAI211_X1 U21613 ( .C1(n18696), .C2(n18547), .A(n18539), .B(n18538), .ZN(
        P3_U2953) );
  AOI22_X1 U21614 ( .A1(n18698), .A2(n18543), .B1(n18697), .B2(n18542), .ZN(
        n18541) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18544), .B1(
        n18699), .B2(n18566), .ZN(n18540) );
  OAI211_X1 U21616 ( .C1(n18702), .C2(n18547), .A(n18541), .B(n18540), .ZN(
        P3_U2954) );
  AOI22_X1 U21617 ( .A1(n18704), .A2(n18543), .B1(n18708), .B2(n18542), .ZN(
        n18546) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18544), .B1(
        n18705), .B2(n18566), .ZN(n18545) );
  OAI211_X1 U21619 ( .C1(n18712), .C2(n18547), .A(n18546), .B(n18545), .ZN(
        P3_U2955) );
  NOR2_X2 U21620 ( .A1(n18548), .A2(n18550), .ZN(n18650) );
  INV_X1 U21621 ( .A(n18650), .ZN(n18570) );
  INV_X1 U21622 ( .A(n18549), .ZN(n18592) );
  NOR2_X1 U21623 ( .A1(n18725), .A2(n18550), .ZN(n18598) );
  AND2_X1 U21624 ( .A1(n18777), .A2(n18598), .ZN(n18565) );
  AOI22_X1 U21625 ( .A1(n18658), .A2(n18592), .B1(n18657), .B2(n18565), .ZN(
        n18552) );
  OAI211_X1 U21626 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18662), .A(
        n18660), .B(n18571), .ZN(n18567) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18567), .B1(
        n18663), .B2(n18566), .ZN(n18551) );
  OAI211_X1 U21628 ( .C1(n18666), .C2(n18570), .A(n18552), .B(n18551), .ZN(
        P3_U2956) );
  AOI22_X1 U21629 ( .A1(n18669), .A2(n18592), .B1(n18667), .B2(n18565), .ZN(
        n18554) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18567), .B1(
        n18668), .B2(n18566), .ZN(n18553) );
  OAI211_X1 U21631 ( .C1(n18672), .C2(n18570), .A(n18554), .B(n18553), .ZN(
        P3_U2957) );
  AOI22_X1 U21632 ( .A1(n18675), .A2(n18566), .B1(n18673), .B2(n18565), .ZN(
        n18556) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18567), .B1(
        n18674), .B2(n18592), .ZN(n18555) );
  OAI211_X1 U21634 ( .C1(n18678), .C2(n18570), .A(n18556), .B(n18555), .ZN(
        P3_U2958) );
  AOI22_X1 U21635 ( .A1(n18680), .A2(n18592), .B1(n18679), .B2(n18565), .ZN(
        n18558) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18567), .B1(
        n18681), .B2(n18566), .ZN(n18557) );
  OAI211_X1 U21637 ( .C1(n18684), .C2(n18570), .A(n18558), .B(n18557), .ZN(
        P3_U2959) );
  AOI22_X1 U21638 ( .A1(n18686), .A2(n18565), .B1(n18685), .B2(n18566), .ZN(
        n18560) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18567), .B1(
        n18687), .B2(n18592), .ZN(n18559) );
  OAI211_X1 U21640 ( .C1(n18690), .C2(n18570), .A(n18560), .B(n18559), .ZN(
        P3_U2960) );
  AOI22_X1 U21641 ( .A1(n18692), .A2(n18565), .B1(n18691), .B2(n18566), .ZN(
        n18562) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18567), .B1(
        n18693), .B2(n18592), .ZN(n18561) );
  OAI211_X1 U21643 ( .C1(n18696), .C2(n18570), .A(n18562), .B(n18561), .ZN(
        P3_U2961) );
  AOI22_X1 U21644 ( .A1(n18699), .A2(n18592), .B1(n18698), .B2(n18565), .ZN(
        n18564) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18567), .B1(
        n18697), .B2(n18566), .ZN(n18563) );
  OAI211_X1 U21646 ( .C1(n18702), .C2(n18570), .A(n18564), .B(n18563), .ZN(
        P3_U2962) );
  AOI22_X1 U21647 ( .A1(n18705), .A2(n18592), .B1(n18704), .B2(n18565), .ZN(
        n18569) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18567), .B1(
        n18708), .B2(n18566), .ZN(n18568) );
  OAI211_X1 U21649 ( .C1(n18712), .C2(n18570), .A(n18569), .B(n18568), .ZN(
        P3_U2963) );
  INV_X1 U21650 ( .A(n18661), .ZN(n18597) );
  NOR2_X2 U21651 ( .A1(n18597), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18707) );
  INV_X1 U21652 ( .A(n18707), .ZN(n18596) );
  NAND2_X1 U21653 ( .A1(n18572), .A2(n18571), .ZN(n18573) );
  NOR2_X1 U21654 ( .A1(n18650), .A2(n18707), .ZN(n18621) );
  OAI21_X1 U21655 ( .B1(n18574), .B2(n18573), .A(n18621), .ZN(n18575) );
  OAI211_X1 U21656 ( .C1(n18707), .C2(n18880), .A(n18576), .B(n18575), .ZN(
        n18593) );
  NOR2_X1 U21657 ( .A1(n18781), .A2(n18621), .ZN(n18591) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18593), .B1(
        n18657), .B2(n18591), .ZN(n18578) );
  AOI22_X1 U21659 ( .A1(n18663), .A2(n18592), .B1(n18658), .B2(n18614), .ZN(
        n18577) );
  OAI211_X1 U21660 ( .C1(n18666), .C2(n18596), .A(n18578), .B(n18577), .ZN(
        P3_U2964) );
  AOI22_X1 U21661 ( .A1(n18669), .A2(n18614), .B1(n18667), .B2(n18591), .ZN(
        n18580) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18593), .B1(
        n18668), .B2(n18592), .ZN(n18579) );
  OAI211_X1 U21663 ( .C1(n18672), .C2(n18596), .A(n18580), .B(n18579), .ZN(
        P3_U2965) );
  AOI22_X1 U21664 ( .A1(n18674), .A2(n18614), .B1(n18673), .B2(n18591), .ZN(
        n18582) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18593), .B1(
        n18675), .B2(n18592), .ZN(n18581) );
  OAI211_X1 U21666 ( .C1(n18678), .C2(n18596), .A(n18582), .B(n18581), .ZN(
        P3_U2966) );
  AOI22_X1 U21667 ( .A1(n18681), .A2(n18592), .B1(n18679), .B2(n18591), .ZN(
        n18584) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18593), .B1(
        n18680), .B2(n18614), .ZN(n18583) );
  OAI211_X1 U21669 ( .C1(n18684), .C2(n18596), .A(n18584), .B(n18583), .ZN(
        P3_U2967) );
  AOI22_X1 U21670 ( .A1(n18686), .A2(n18591), .B1(n18685), .B2(n18592), .ZN(
        n18586) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18593), .B1(
        n18687), .B2(n18614), .ZN(n18585) );
  OAI211_X1 U21672 ( .C1(n18690), .C2(n18596), .A(n18586), .B(n18585), .ZN(
        P3_U2968) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18593), .B1(
        n18692), .B2(n18591), .ZN(n18588) );
  AOI22_X1 U21674 ( .A1(n18693), .A2(n18614), .B1(n18691), .B2(n18592), .ZN(
        n18587) );
  OAI211_X1 U21675 ( .C1(n18696), .C2(n18596), .A(n18588), .B(n18587), .ZN(
        P3_U2969) );
  AOI22_X1 U21676 ( .A1(n18699), .A2(n18614), .B1(n18698), .B2(n18591), .ZN(
        n18590) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18593), .B1(
        n18697), .B2(n18592), .ZN(n18589) );
  OAI211_X1 U21678 ( .C1(n18702), .C2(n18596), .A(n18590), .B(n18589), .ZN(
        P3_U2970) );
  AOI22_X1 U21679 ( .A1(n18705), .A2(n18614), .B1(n18704), .B2(n18591), .ZN(
        n18595) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18593), .B1(
        n18708), .B2(n18592), .ZN(n18594) );
  OAI211_X1 U21681 ( .C1(n18712), .C2(n18596), .A(n18595), .B(n18594), .ZN(
        P3_U2971) );
  NOR2_X1 U21682 ( .A1(n18781), .A2(n18597), .ZN(n18613) );
  AOI22_X1 U21683 ( .A1(n18658), .A2(n18650), .B1(n18657), .B2(n18613), .ZN(
        n18600) );
  AOI22_X1 U21684 ( .A1(n18662), .A2(n18598), .B1(n18661), .B2(n18660), .ZN(
        n18615) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18615), .B1(
        n18663), .B2(n18614), .ZN(n18599) );
  OAI211_X1 U21686 ( .C1(n18618), .C2(n18666), .A(n18600), .B(n18599), .ZN(
        P3_U2972) );
  AOI22_X1 U21687 ( .A1(n18669), .A2(n18650), .B1(n18667), .B2(n18613), .ZN(
        n18602) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18615), .B1(
        n18668), .B2(n18614), .ZN(n18601) );
  OAI211_X1 U21689 ( .C1(n18618), .C2(n18672), .A(n18602), .B(n18601), .ZN(
        P3_U2973) );
  AOI22_X1 U21690 ( .A1(n18675), .A2(n18614), .B1(n18673), .B2(n18613), .ZN(
        n18604) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18615), .B1(
        n18674), .B2(n18650), .ZN(n18603) );
  OAI211_X1 U21692 ( .C1(n18618), .C2(n18678), .A(n18604), .B(n18603), .ZN(
        P3_U2974) );
  AOI22_X1 U21693 ( .A1(n18681), .A2(n18614), .B1(n18679), .B2(n18613), .ZN(
        n18606) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18615), .B1(
        n18680), .B2(n18650), .ZN(n18605) );
  OAI211_X1 U21695 ( .C1(n18618), .C2(n18684), .A(n18606), .B(n18605), .ZN(
        P3_U2975) );
  AOI22_X1 U21696 ( .A1(n18687), .A2(n18650), .B1(n18686), .B2(n18613), .ZN(
        n18608) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18615), .B1(
        n18685), .B2(n18614), .ZN(n18607) );
  OAI211_X1 U21698 ( .C1(n18618), .C2(n18690), .A(n18608), .B(n18607), .ZN(
        P3_U2976) );
  AOI22_X1 U21699 ( .A1(n18693), .A2(n18650), .B1(n18692), .B2(n18613), .ZN(
        n18610) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18615), .B1(
        n18691), .B2(n18614), .ZN(n18609) );
  OAI211_X1 U21701 ( .C1(n18618), .C2(n18696), .A(n18610), .B(n18609), .ZN(
        P3_U2977) );
  AOI22_X1 U21702 ( .A1(n18699), .A2(n18650), .B1(n18698), .B2(n18613), .ZN(
        n18612) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18615), .B1(
        n18697), .B2(n18614), .ZN(n18611) );
  OAI211_X1 U21704 ( .C1(n18618), .C2(n18702), .A(n18612), .B(n18611), .ZN(
        P3_U2978) );
  AOI22_X1 U21705 ( .A1(n18705), .A2(n18650), .B1(n18704), .B2(n18613), .ZN(
        n18617) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18615), .B1(
        n18708), .B2(n18614), .ZN(n18616) );
  OAI211_X1 U21707 ( .C1(n18618), .C2(n18712), .A(n18617), .B(n18616), .ZN(
        P3_U2979) );
  INV_X1 U21708 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20925) );
  NOR2_X1 U21709 ( .A1(n18781), .A2(n18622), .ZN(n18649) );
  AOI22_X1 U21710 ( .A1(n18663), .A2(n18650), .B1(n18657), .B2(n18649), .ZN(
        n18625) );
  AOI22_X1 U21711 ( .A1(n18623), .A2(n18652), .B1(n18658), .B2(n18707), .ZN(
        n18624) );
  OAI211_X1 U21712 ( .C1(n18656), .C2(n20925), .A(n18625), .B(n18624), .ZN(
        P3_U2980) );
  INV_X1 U21713 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18629) );
  AOI22_X1 U21714 ( .A1(n18668), .A2(n18650), .B1(n18667), .B2(n18649), .ZN(
        n18628) );
  AOI22_X1 U21715 ( .A1(n18652), .A2(n18626), .B1(n18669), .B2(n18707), .ZN(
        n18627) );
  OAI211_X1 U21716 ( .C1(n18656), .C2(n18629), .A(n18628), .B(n18627), .ZN(
        P3_U2981) );
  INV_X1 U21717 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20877) );
  AOI22_X1 U21718 ( .A1(n18675), .A2(n18650), .B1(n18673), .B2(n18649), .ZN(
        n18632) );
  AOI22_X1 U21719 ( .A1(n18652), .A2(n18630), .B1(n18674), .B2(n18707), .ZN(
        n18631) );
  OAI211_X1 U21720 ( .C1(n18656), .C2(n20877), .A(n18632), .B(n18631), .ZN(
        P3_U2982) );
  INV_X1 U21721 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18636) );
  AOI22_X1 U21722 ( .A1(n18681), .A2(n18650), .B1(n18679), .B2(n18649), .ZN(
        n18635) );
  AOI22_X1 U21723 ( .A1(n18652), .A2(n18633), .B1(n18680), .B2(n18707), .ZN(
        n18634) );
  OAI211_X1 U21724 ( .C1(n18656), .C2(n18636), .A(n18635), .B(n18634), .ZN(
        P3_U2983) );
  INV_X1 U21725 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18640) );
  AOI22_X1 U21726 ( .A1(n18687), .A2(n18707), .B1(n18686), .B2(n18649), .ZN(
        n18639) );
  AOI22_X1 U21727 ( .A1(n18652), .A2(n18637), .B1(n18685), .B2(n18650), .ZN(
        n18638) );
  OAI211_X1 U21728 ( .C1(n18656), .C2(n18640), .A(n18639), .B(n18638), .ZN(
        P3_U2984) );
  INV_X1 U21729 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18644) );
  AOI22_X1 U21730 ( .A1(n18692), .A2(n18649), .B1(n18691), .B2(n18650), .ZN(
        n18643) );
  AOI22_X1 U21731 ( .A1(n18652), .A2(n18641), .B1(n18693), .B2(n18707), .ZN(
        n18642) );
  OAI211_X1 U21732 ( .C1(n18656), .C2(n18644), .A(n18643), .B(n18642), .ZN(
        P3_U2985) );
  INV_X1 U21733 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18648) );
  AOI22_X1 U21734 ( .A1(n18698), .A2(n18649), .B1(n18697), .B2(n18650), .ZN(
        n18647) );
  AOI22_X1 U21735 ( .A1(n18652), .A2(n18645), .B1(n18699), .B2(n18707), .ZN(
        n18646) );
  OAI211_X1 U21736 ( .C1(n18656), .C2(n18648), .A(n18647), .B(n18646), .ZN(
        P3_U2986) );
  INV_X1 U21737 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18655) );
  AOI22_X1 U21738 ( .A1(n18705), .A2(n18707), .B1(n18704), .B2(n18649), .ZN(
        n18654) );
  AOI22_X1 U21739 ( .A1(n18652), .A2(n18651), .B1(n18708), .B2(n18650), .ZN(
        n18653) );
  OAI211_X1 U21740 ( .C1(n18656), .C2(n18655), .A(n18654), .B(n18653), .ZN(
        P3_U2987) );
  AND2_X1 U21741 ( .A1(n18777), .A2(n18659), .ZN(n18703) );
  AOI22_X1 U21742 ( .A1(n18706), .A2(n18658), .B1(n18657), .B2(n18703), .ZN(
        n18665) );
  AOI22_X1 U21743 ( .A1(n18662), .A2(n18661), .B1(n18660), .B2(n18659), .ZN(
        n18709) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18709), .B1(
        n18663), .B2(n18707), .ZN(n18664) );
  OAI211_X1 U21745 ( .C1(n18713), .C2(n18666), .A(n18665), .B(n18664), .ZN(
        P3_U2988) );
  AOI22_X1 U21746 ( .A1(n18668), .A2(n18707), .B1(n18667), .B2(n18703), .ZN(
        n18671) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18709), .B1(
        n18706), .B2(n18669), .ZN(n18670) );
  OAI211_X1 U21748 ( .C1(n18713), .C2(n18672), .A(n18671), .B(n18670), .ZN(
        P3_U2989) );
  AOI22_X1 U21749 ( .A1(n18706), .A2(n18674), .B1(n18673), .B2(n18703), .ZN(
        n18677) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18709), .B1(
        n18675), .B2(n18707), .ZN(n18676) );
  OAI211_X1 U21751 ( .C1(n18713), .C2(n18678), .A(n18677), .B(n18676), .ZN(
        P3_U2990) );
  AOI22_X1 U21752 ( .A1(n18706), .A2(n18680), .B1(n18679), .B2(n18703), .ZN(
        n18683) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18709), .B1(
        n18681), .B2(n18707), .ZN(n18682) );
  OAI211_X1 U21754 ( .C1(n18713), .C2(n18684), .A(n18683), .B(n18682), .ZN(
        P3_U2991) );
  AOI22_X1 U21755 ( .A1(n18686), .A2(n18703), .B1(n18685), .B2(n18707), .ZN(
        n18689) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18709), .B1(
        n18706), .B2(n18687), .ZN(n18688) );
  OAI211_X1 U21757 ( .C1(n18713), .C2(n18690), .A(n18689), .B(n18688), .ZN(
        P3_U2992) );
  AOI22_X1 U21758 ( .A1(n18692), .A2(n18703), .B1(n18691), .B2(n18707), .ZN(
        n18695) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18709), .B1(
        n18706), .B2(n18693), .ZN(n18694) );
  OAI211_X1 U21760 ( .C1(n18713), .C2(n18696), .A(n18695), .B(n18694), .ZN(
        P3_U2993) );
  AOI22_X1 U21761 ( .A1(n18698), .A2(n18703), .B1(n18697), .B2(n18707), .ZN(
        n18701) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18709), .B1(
        n18706), .B2(n18699), .ZN(n18700) );
  OAI211_X1 U21763 ( .C1(n18713), .C2(n18702), .A(n18701), .B(n18700), .ZN(
        P3_U2994) );
  AOI22_X1 U21764 ( .A1(n18706), .A2(n18705), .B1(n18704), .B2(n18703), .ZN(
        n18711) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18709), .B1(
        n18708), .B2(n18707), .ZN(n18710) );
  OAI211_X1 U21766 ( .C1(n18713), .C2(n18712), .A(n18711), .B(n18710), .ZN(
        P3_U2995) );
  AOI22_X1 U21767 ( .A1(n18896), .A2(n18741), .B1(n18716), .B2(n18735), .ZN(
        n18714) );
  OAI21_X1 U21768 ( .B1(n18731), .B2(n18715), .A(n18714), .ZN(n18885) );
  NOR2_X1 U21769 ( .A1(n18761), .A2(n18885), .ZN(n18719) );
  AND2_X1 U21770 ( .A1(n18896), .A2(n18741), .ZN(n18717) );
  NOR2_X1 U21771 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18716), .ZN(
        n18723) );
  OAI22_X1 U21772 ( .A1(n18717), .A2(n18739), .B1(n18723), .B2(n18735), .ZN(
        n18882) );
  NAND2_X1 U21773 ( .A1(n18886), .A2(n18882), .ZN(n18718) );
  OAI22_X1 U21774 ( .A1(n18719), .A2(n18886), .B1(n18761), .B2(n18718), .ZN(
        n18769) );
  NOR2_X1 U21775 ( .A1(n18721), .A2(n18720), .ZN(n18724) );
  OAI22_X1 U21776 ( .A1(n18910), .A2(n18722), .B1(n18724), .B2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18905) );
  INV_X1 U21777 ( .A(n18905), .ZN(n18728) );
  OAI22_X1 U21778 ( .A1(n18724), .A2(n18897), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18723), .ZN(n18901) );
  OAI221_X1 U21779 ( .B1(n18901), .B2(n18905), .C1(n18901), .C2(n18725), .A(
        n18744), .ZN(n18726) );
  AOI22_X1 U21780 ( .A1(n18729), .A2(n18728), .B1(n18727), .B2(n18726), .ZN(
        n18747) );
  AOI221_X1 U21781 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18731), 
        .C1(n18730), .C2(n18731), .A(n18896), .ZN(n18742) );
  NOR2_X1 U21782 ( .A1(n18732), .A2(n18910), .ZN(n18734) );
  OAI211_X1 U21783 ( .C1(n18734), .C2(n18733), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18896), .ZN(n18738) );
  OAI211_X1 U21784 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18736), .B(n18735), .ZN(
        n18737) );
  OAI211_X1 U21785 ( .C1(n18892), .C2(n18739), .A(n18738), .B(n18737), .ZN(
        n18740) );
  AOI21_X1 U21786 ( .B1(n18742), .B2(n18741), .A(n18740), .ZN(n18743) );
  INV_X1 U21787 ( .A(n18743), .ZN(n18894) );
  OAI22_X1 U21788 ( .A1(n18744), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18894), .B2(n18761), .ZN(n18748) );
  INV_X1 U21789 ( .A(n18748), .ZN(n18745) );
  AOI222_X1 U21790 ( .A1(n18747), .A2(n18746), .B1(n18747), .B2(n18745), .C1(
        n18746), .C2(n18745), .ZN(n18765) );
  OAI221_X1 U21791 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n18765), .A(n18748), .ZN(
        n18768) );
  INV_X1 U21792 ( .A(n18749), .ZN(n18755) );
  NOR2_X1 U21793 ( .A1(n18751), .A2(n18750), .ZN(n18753) );
  OAI222_X1 U21794 ( .A1(n18757), .A2(n18756), .B1(n18755), .B2(n18754), .C1(
        n18753), .C2(n9960), .ZN(n18923) );
  NAND2_X1 U21795 ( .A1(n21010), .A2(n18758), .ZN(n18766) );
  AOI211_X1 U21796 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18761), .A(
        n18760), .B(n18759), .ZN(n18764) );
  OAI21_X1 U21797 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18762), .ZN(n18763) );
  OAI211_X1 U21798 ( .C1(n18766), .C2(n18765), .A(n18764), .B(n18763), .ZN(
        n18767) );
  AOI211_X1 U21799 ( .C1(n18769), .C2(n18768), .A(n18923), .B(n18767), .ZN(
        n18780) );
  AOI22_X1 U21800 ( .A1(n18931), .A2(n17519), .B1(n18904), .B2(n18936), .ZN(
        n18770) );
  INV_X1 U21801 ( .A(n18770), .ZN(n18776) );
  OAI211_X1 U21802 ( .C1(n18773), .C2(n18772), .A(n18771), .B(n18780), .ZN(
        n18879) );
  OAI21_X1 U21803 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18796), .A(n18879), 
        .ZN(n18782) );
  NOR2_X1 U21804 ( .A1(n18774), .A2(n18782), .ZN(n18775) );
  MUX2_X1 U21805 ( .A(n18776), .B(n18775), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18779) );
  OR2_X1 U21806 ( .A1(n18783), .A2(n18777), .ZN(n18778) );
  OAI211_X1 U21807 ( .C1(n18780), .C2(n18925), .A(n18779), .B(n18778), .ZN(
        P3_U2996) );
  NAND2_X1 U21808 ( .A1(n18931), .A2(n17519), .ZN(n18786) );
  NOR4_X1 U21809 ( .A1(n18933), .A2(n18889), .A3(n18796), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18789) );
  INV_X1 U21810 ( .A(n18789), .ZN(n18785) );
  OR3_X1 U21811 ( .A1(n18783), .A2(n18782), .A3(n18781), .ZN(n18784) );
  NAND4_X1 U21812 ( .A1(n18787), .A2(n18786), .A3(n18785), .A4(n18784), .ZN(
        P3_U2997) );
  OAI21_X1 U21813 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18788), .ZN(n18790) );
  AOI21_X1 U21814 ( .B1(n18791), .B2(n18790), .A(n18789), .ZN(P3_U2998) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18876), .ZN(
        P3_U2999) );
  AND2_X1 U21816 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18876), .ZN(
        P3_U3000) );
  AND2_X1 U21817 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18876), .ZN(
        P3_U3001) );
  AND2_X1 U21818 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18876), .ZN(
        P3_U3002) );
  AND2_X1 U21819 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18876), .ZN(
        P3_U3003) );
  AND2_X1 U21820 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18876), .ZN(
        P3_U3004) );
  AND2_X1 U21821 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18876), .ZN(
        P3_U3005) );
  AND2_X1 U21822 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18876), .ZN(
        P3_U3006) );
  AND2_X1 U21823 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18876), .ZN(
        P3_U3007) );
  AND2_X1 U21824 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18876), .ZN(
        P3_U3008) );
  AND2_X1 U21825 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18876), .ZN(
        P3_U3009) );
  AND2_X1 U21826 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18876), .ZN(
        P3_U3010) );
  AND2_X1 U21827 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18876), .ZN(
        P3_U3011) );
  AND2_X1 U21828 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18876), .ZN(
        P3_U3012) );
  AND2_X1 U21829 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18876), .ZN(
        P3_U3013) );
  AND2_X1 U21830 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18876), .ZN(
        P3_U3014) );
  AND2_X1 U21831 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18876), .ZN(
        P3_U3015) );
  AND2_X1 U21832 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18876), .ZN(
        P3_U3016) );
  AND2_X1 U21833 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18876), .ZN(
        P3_U3017) );
  AND2_X1 U21834 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18876), .ZN(
        P3_U3018) );
  AND2_X1 U21835 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18876), .ZN(
        P3_U3019) );
  AND2_X1 U21836 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18876), .ZN(
        P3_U3020) );
  AND2_X1 U21837 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18876), .ZN(P3_U3021) );
  AND2_X1 U21838 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18876), .ZN(P3_U3022) );
  AND2_X1 U21839 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18876), .ZN(P3_U3023) );
  AND2_X1 U21840 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18876), .ZN(P3_U3024) );
  AND2_X1 U21841 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18876), .ZN(P3_U3025) );
  AND2_X1 U21842 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18876), .ZN(P3_U3026) );
  AND2_X1 U21843 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18876), .ZN(P3_U3027) );
  AND2_X1 U21844 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18876), .ZN(P3_U3028) );
  OAI21_X1 U21845 ( .B1(n18793), .B2(n19855), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18794) );
  AOI22_X1 U21846 ( .A1(n18805), .A2(n18807), .B1(n18940), .B2(n18794), .ZN(
        n18795) );
  INV_X1 U21847 ( .A(NA), .ZN(n20759) );
  OR3_X1 U21848 ( .A1(n20759), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18800) );
  OAI211_X1 U21849 ( .C1(n18796), .C2(n18797), .A(n18795), .B(n18800), .ZN(
        P3_U3029) );
  NOR2_X1 U21850 ( .A1(n18807), .A2(n19855), .ZN(n18803) );
  INV_X1 U21851 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18938) );
  OAI22_X1 U21852 ( .A1(n18803), .A2(n18938), .B1(n19855), .B2(n18797), .ZN(
        n18798) );
  AOI21_X1 U21853 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n18798), .A(n18928), 
        .ZN(n18799) );
  NAND2_X1 U21854 ( .A1(n18931), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18801) );
  NAND2_X1 U21855 ( .A1(n18799), .A2(n18801), .ZN(P3_U3030) );
  AOI22_X1 U21856 ( .A1(n18931), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18805), 
        .B2(n18800), .ZN(n18806) );
  OAI22_X1 U21857 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18801), .ZN(n18802) );
  OAI22_X1 U21858 ( .A1(n18803), .A2(n18802), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18804) );
  OAI22_X1 U21859 ( .A1(n18806), .A2(n18807), .B1(n18805), .B2(n18804), .ZN(
        P3_U3031) );
  INV_X2 U21860 ( .A(n18812), .ZN(n18860) );
  OAI222_X1 U21861 ( .A1(n18809), .A2(n18860), .B1(n18808), .B2(n18872), .C1(
        n18810), .C2(n18868), .ZN(P3_U3032) );
  OAI222_X1 U21862 ( .A1(n18868), .A2(n18813), .B1(n18811), .B2(n18872), .C1(
        n18810), .C2(n18860), .ZN(P3_U3033) );
  OAI222_X1 U21863 ( .A1(n18868), .A2(n18815), .B1(n18814), .B2(n18872), .C1(
        n18813), .C2(n18860), .ZN(P3_U3034) );
  OAI222_X1 U21864 ( .A1(n18868), .A2(n18818), .B1(n18816), .B2(n18872), .C1(
        n18815), .C2(n18860), .ZN(P3_U3035) );
  OAI222_X1 U21865 ( .A1(n18818), .A2(n18860), .B1(n18817), .B2(n18872), .C1(
        n18819), .C2(n18868), .ZN(P3_U3036) );
  INV_X1 U21866 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18821) );
  OAI222_X1 U21867 ( .A1(n18868), .A2(n18821), .B1(n18820), .B2(n18872), .C1(
        n18819), .C2(n18860), .ZN(P3_U3037) );
  OAI222_X1 U21868 ( .A1(n18868), .A2(n21110), .B1(n18822), .B2(n18872), .C1(
        n18821), .C2(n18860), .ZN(P3_U3038) );
  OAI222_X1 U21869 ( .A1(n21110), .A2(n18860), .B1(n18823), .B2(n18872), .C1(
        n18824), .C2(n18868), .ZN(P3_U3039) );
  OAI222_X1 U21870 ( .A1(n18868), .A2(n18826), .B1(n18825), .B2(n18872), .C1(
        n18824), .C2(n18860), .ZN(P3_U3040) );
  OAI222_X1 U21871 ( .A1(n18868), .A2(n18828), .B1(n18827), .B2(n18872), .C1(
        n18826), .C2(n18860), .ZN(P3_U3041) );
  OAI222_X1 U21872 ( .A1(n18868), .A2(n18830), .B1(n18829), .B2(n18872), .C1(
        n18828), .C2(n18860), .ZN(P3_U3042) );
  INV_X1 U21873 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18832) );
  OAI222_X1 U21874 ( .A1(n18868), .A2(n18832), .B1(n18831), .B2(n18872), .C1(
        n18830), .C2(n18860), .ZN(P3_U3043) );
  OAI222_X1 U21875 ( .A1(n18868), .A2(n18835), .B1(n18833), .B2(n18872), .C1(
        n18832), .C2(n18860), .ZN(P3_U3044) );
  OAI222_X1 U21876 ( .A1(n18835), .A2(n18860), .B1(n18834), .B2(n18872), .C1(
        n18836), .C2(n18868), .ZN(P3_U3045) );
  OAI222_X1 U21877 ( .A1(n18868), .A2(n18838), .B1(n18837), .B2(n18872), .C1(
        n18836), .C2(n18860), .ZN(P3_U3046) );
  OAI222_X1 U21878 ( .A1(n18868), .A2(n18841), .B1(n18839), .B2(n18872), .C1(
        n18838), .C2(n18860), .ZN(P3_U3047) );
  OAI222_X1 U21879 ( .A1(n18841), .A2(n18860), .B1(n18840), .B2(n18872), .C1(
        n18842), .C2(n18868), .ZN(P3_U3048) );
  OAI222_X1 U21880 ( .A1(n18868), .A2(n18844), .B1(n18843), .B2(n18872), .C1(
        n18842), .C2(n18860), .ZN(P3_U3049) );
  OAI222_X1 U21881 ( .A1(n18868), .A2(n21120), .B1(n18845), .B2(n18872), .C1(
        n18844), .C2(n18860), .ZN(P3_U3050) );
  OAI222_X1 U21882 ( .A1(n18868), .A2(n18847), .B1(n18846), .B2(n18872), .C1(
        n21120), .C2(n18860), .ZN(P3_U3051) );
  OAI222_X1 U21883 ( .A1(n18868), .A2(n18849), .B1(n18848), .B2(n18872), .C1(
        n18847), .C2(n18860), .ZN(P3_U3052) );
  OAI222_X1 U21884 ( .A1(n18868), .A2(n18852), .B1(n18850), .B2(n18872), .C1(
        n18849), .C2(n18860), .ZN(P3_U3053) );
  OAI222_X1 U21885 ( .A1(n18852), .A2(n18860), .B1(n18851), .B2(n18872), .C1(
        n18853), .C2(n18868), .ZN(P3_U3054) );
  OAI222_X1 U21886 ( .A1(n18868), .A2(n18855), .B1(n18854), .B2(n18872), .C1(
        n18853), .C2(n18860), .ZN(P3_U3055) );
  OAI222_X1 U21887 ( .A1(n18868), .A2(n18857), .B1(n18856), .B2(n18872), .C1(
        n18855), .C2(n18860), .ZN(P3_U3056) );
  OAI222_X1 U21888 ( .A1(n18868), .A2(n21014), .B1(n18858), .B2(n18872), .C1(
        n18857), .C2(n18860), .ZN(P3_U3057) );
  INV_X1 U21889 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18861) );
  OAI222_X1 U21890 ( .A1(n18860), .A2(n21014), .B1(n18859), .B2(n18872), .C1(
        n18861), .C2(n18868), .ZN(P3_U3058) );
  OAI222_X1 U21891 ( .A1(n18868), .A2(n18863), .B1(n18862), .B2(n18872), .C1(
        n18861), .C2(n18860), .ZN(P3_U3059) );
  INV_X1 U21892 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18865) );
  OAI222_X1 U21893 ( .A1(n18868), .A2(n18865), .B1(n18864), .B2(n18872), .C1(
        n18863), .C2(n18860), .ZN(P3_U3060) );
  OAI222_X1 U21894 ( .A1(n18868), .A2(n18867), .B1(n18866), .B2(n18872), .C1(
        n18865), .C2(n18860), .ZN(P3_U3061) );
  OAI22_X1 U21895 ( .A1(n18940), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18872), .ZN(n18869) );
  INV_X1 U21896 ( .A(n18869), .ZN(P3_U3274) );
  OAI22_X1 U21897 ( .A1(n18940), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18872), .ZN(n18870) );
  INV_X1 U21898 ( .A(n18870), .ZN(P3_U3275) );
  OAI22_X1 U21899 ( .A1(n18940), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18872), .ZN(n18871) );
  INV_X1 U21900 ( .A(n18871), .ZN(P3_U3276) );
  OAI22_X1 U21901 ( .A1(n18940), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18872), .ZN(n18873) );
  INV_X1 U21902 ( .A(n18873), .ZN(P3_U3277) );
  INV_X1 U21903 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18913) );
  INV_X1 U21904 ( .A(n18874), .ZN(n18875) );
  AOI21_X1 U21905 ( .B1(n18876), .B2(n18913), .A(n18875), .ZN(P3_U3280) );
  AOI21_X1 U21906 ( .B1(n18876), .B2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n18875), 
        .ZN(n18877) );
  INV_X1 U21907 ( .A(n18877), .ZN(P3_U3281) );
  OAI221_X1 U21908 ( .B1(n18880), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18880), 
        .C2(n18879), .A(n18878), .ZN(P3_U3282) );
  NOR2_X1 U21909 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18881), .ZN(
        n18883) );
  AOI22_X1 U21910 ( .A1(n18904), .A2(n18884), .B1(n18883), .B2(n18882), .ZN(
        n18888) );
  AOI21_X1 U21911 ( .B1(n18906), .B2(n18885), .A(n18911), .ZN(n18887) );
  OAI22_X1 U21912 ( .A1(n18911), .A2(n18888), .B1(n18887), .B2(n18886), .ZN(
        P3_U3285) );
  NOR2_X1 U21913 ( .A1(n18889), .A2(n18907), .ZN(n18898) );
  OAI22_X1 U21914 ( .A1(n18891), .A2(n18890), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18899) );
  INV_X1 U21915 ( .A(n18899), .ZN(n18893) );
  AOI222_X1 U21916 ( .A1(n18894), .A2(n18906), .B1(n18898), .B2(n18893), .C1(
        n18904), .C2(n18892), .ZN(n18895) );
  AOI22_X1 U21917 ( .A1(n18911), .A2(n18896), .B1(n18895), .B2(n18908), .ZN(
        P3_U3288) );
  INV_X1 U21918 ( .A(n18897), .ZN(n18900) );
  AOI222_X1 U21919 ( .A1(n18901), .A2(n18906), .B1(n18904), .B2(n18900), .C1(
        n18899), .C2(n18898), .ZN(n18902) );
  AOI22_X1 U21920 ( .A1(n18911), .A2(n18903), .B1(n18902), .B2(n18908), .ZN(
        P3_U3289) );
  AOI222_X1 U21921 ( .A1(n18907), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18906), 
        .B2(n18905), .C1(n18910), .C2(n18904), .ZN(n18909) );
  AOI22_X1 U21922 ( .A1(n18911), .A2(n18910), .B1(n18909), .B2(n18908), .ZN(
        P3_U3290) );
  NOR3_X1 U21923 ( .A1(n18913), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18912) );
  AOI221_X1 U21924 ( .B1(n18914), .B2(n18913), .C1(P3_REIP_REG_1__SCAN_IN), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18912), .ZN(n18916) );
  INV_X1 U21925 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18915) );
  INV_X1 U21926 ( .A(n18920), .ZN(n18917) );
  AOI22_X1 U21927 ( .A1(n18920), .A2(n18916), .B1(n18915), .B2(n18917), .ZN(
        P3_U3292) );
  NOR2_X1 U21928 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18919) );
  INV_X1 U21929 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18918) );
  AOI22_X1 U21930 ( .A1(n18920), .A2(n18919), .B1(n18918), .B2(n18917), .ZN(
        P3_U3293) );
  INV_X1 U21931 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18921) );
  AOI22_X1 U21932 ( .A1(n18872), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18921), 
        .B2(n18940), .ZN(P3_U3294) );
  MUX2_X1 U21933 ( .A(P3_MORE_REG_SCAN_IN), .B(n18923), .S(n18922), .Z(
        P3_U3295) );
  AOI21_X1 U21934 ( .B1(n18925), .B2(n18924), .A(n18947), .ZN(n18926) );
  OAI21_X1 U21935 ( .B1(n18931), .B2(n18927), .A(n18926), .ZN(n18939) );
  OAI21_X1 U21936 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18929), .A(n18928), 
        .ZN(n18932) );
  AOI211_X1 U21937 ( .C1(n18942), .C2(n18932), .A(n18931), .B(n18930), .ZN(
        n18934) );
  NOR2_X1 U21938 ( .A1(n18934), .A2(n18933), .ZN(n18935) );
  OAI21_X1 U21939 ( .B1(n18936), .B2(n18935), .A(n18939), .ZN(n18937) );
  OAI21_X1 U21940 ( .B1(n18939), .B2(n18938), .A(n18937), .ZN(P3_U3296) );
  MUX2_X1 U21941 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n18940), .Z(P3_U3297) );
  OAI21_X1 U21942 ( .B1(n18944), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n18943), 
        .ZN(n18941) );
  OAI21_X1 U21943 ( .B1(n18943), .B2(n18942), .A(n18941), .ZN(P3_U3298) );
  NOR2_X1 U21944 ( .A1(n18944), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18946)
         );
  OAI21_X1 U21945 ( .B1(n18947), .B2(n18946), .A(n18945), .ZN(P3_U3299) );
  INV_X1 U21946 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19845) );
  NAND2_X1 U21947 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19866), .ZN(n19854) );
  NAND2_X1 U21948 ( .A1(n19845), .A2(n18948), .ZN(n19851) );
  OAI21_X1 U21949 ( .B1(n19845), .B2(n19854), .A(n19851), .ZN(n19922) );
  AOI21_X1 U21950 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19922), .ZN(n18949) );
  INV_X1 U21951 ( .A(n18949), .ZN(P2_U2815) );
  INV_X1 U21952 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18952) );
  OAI22_X1 U21953 ( .A1(n18951), .A2(n18952), .B1(n19924), .B2(n18950), .ZN(
        P2_U2816) );
  INV_X2 U21954 ( .A(n19970), .ZN(n19969) );
  AOI22_X1 U21955 ( .A1(n19969), .A2(n18952), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19970), .ZN(n18953) );
  OAI21_X1 U21956 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19851), .A(n18953), 
        .ZN(P2_U2817) );
  OAI21_X1 U21957 ( .B1(n19859), .B2(BS16), .A(n19922), .ZN(n19920) );
  OAI21_X1 U21958 ( .B1(n19922), .B2(n19661), .A(n19920), .ZN(P2_U2818) );
  NOR4_X1 U21959 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n18957) );
  NOR4_X1 U21960 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_14__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n18956) );
  NOR4_X1 U21961 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18955) );
  NOR4_X1 U21962 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18954) );
  NAND4_X1 U21963 ( .A1(n18957), .A2(n18956), .A3(n18955), .A4(n18954), .ZN(
        n18963) );
  NOR4_X1 U21964 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_2__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18961) );
  AOI211_X1 U21965 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_17__SCAN_IN), .B(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18960) );
  NOR4_X1 U21966 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18959) );
  NOR4_X1 U21967 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18958) );
  NAND4_X1 U21968 ( .A1(n18961), .A2(n18960), .A3(n18959), .A4(n18958), .ZN(
        n18962) );
  NOR2_X1 U21969 ( .A1(n18963), .A2(n18962), .ZN(n18973) );
  INV_X1 U21970 ( .A(n18973), .ZN(n18971) );
  NOR2_X1 U21971 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18971), .ZN(n18966) );
  NOR2_X1 U21972 ( .A1(n18973), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18964)
         );
  OAI22_X1 U21973 ( .A1(n18966), .A2(n18964), .B1(n12290), .B2(n18971), .ZN(
        P2_U2820) );
  OR3_X1 U21974 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18970) );
  INV_X1 U21975 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18965) );
  AOI22_X1 U21976 ( .A1(n18966), .A2(n18970), .B1(n18971), .B2(n18965), .ZN(
        P2_U2821) );
  INV_X1 U21977 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19921) );
  NAND2_X1 U21978 ( .A1(n18966), .A2(n19921), .ZN(n18969) );
  OAI21_X1 U21979 ( .B1(n12290), .B2(n19867), .A(n18973), .ZN(n18967) );
  OAI21_X1 U21980 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18973), .A(n18967), 
        .ZN(n18968) );
  OAI221_X1 U21981 ( .B1(n18969), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18969), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18968), .ZN(P2_U2822) );
  INV_X1 U21982 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18972) );
  OAI221_X1 U21983 ( .B1(n18973), .B2(n18972), .C1(n18971), .C2(n18970), .A(
        n18969), .ZN(P2_U2823) );
  OAI22_X1 U21984 ( .A1(n19101), .A2(n12544), .B1(n19896), .B2(n19059), .ZN(
        n18975) );
  NOR2_X1 U21985 ( .A1(n19024), .A2(n12957), .ZN(n18974) );
  AOI211_X1 U21986 ( .C1(n18976), .C2(n19119), .A(n18975), .B(n18974), .ZN(
        n18977) );
  OAI21_X1 U21987 ( .B1(n18978), .B2(n19090), .A(n18977), .ZN(n18979) );
  INV_X1 U21988 ( .A(n18979), .ZN(n18984) );
  OAI211_X1 U21989 ( .C1(n18982), .C2(n18981), .A(n19080), .B(n18980), .ZN(
        n18983) );
  OAI211_X1 U21990 ( .C1(n19100), .C2(n18985), .A(n18984), .B(n18983), .ZN(
        P2_U2835) );
  AOI22_X1 U21991 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19130), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n19117), .ZN(n18986) );
  OAI21_X1 U21992 ( .B1(n18987), .B2(n19090), .A(n18986), .ZN(n18988) );
  AOI211_X1 U21993 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19122), .A(n19255), 
        .B(n18988), .ZN(n18997) );
  INV_X1 U21994 ( .A(n18989), .ZN(n18990) );
  AOI22_X1 U21995 ( .A1(n19119), .A2(n18991), .B1(n18990), .B2(n19121), .ZN(
        n18996) );
  OAI211_X1 U21996 ( .C1(n18994), .C2(n18993), .A(n19080), .B(n18992), .ZN(
        n18995) );
  NAND3_X1 U21997 ( .A1(n18997), .A2(n18996), .A3(n18995), .ZN(P2_U2836) );
  NOR2_X1 U21998 ( .A1(n19105), .A2(n18998), .ZN(n19001) );
  AOI22_X1 U21999 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19130), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19117), .ZN(n18999) );
  OAI211_X1 U22000 ( .C1(n19059), .C2(n19893), .A(n18999), .B(n19058), .ZN(
        n19000) );
  AOI211_X1 U22001 ( .C1(n19002), .C2(n19125), .A(n19001), .B(n19000), .ZN(
        n19007) );
  OAI211_X1 U22002 ( .C1(n19005), .C2(n19004), .A(n19080), .B(n19003), .ZN(
        n19006) );
  OAI211_X1 U22003 ( .C1(n19100), .C2(n19008), .A(n19007), .B(n19006), .ZN(
        P2_U2837) );
  NOR2_X1 U22004 ( .A1(n19108), .A2(n19009), .ZN(n19033) );
  XOR2_X1 U22005 ( .A(n19010), .B(n19033), .Z(n19019) );
  INV_X1 U22006 ( .A(n19011), .ZN(n19012) );
  AOI22_X1 U22007 ( .A1(n19012), .A2(n19125), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19130), .ZN(n19013) );
  OAI211_X1 U22008 ( .C1(n19890), .C2(n19059), .A(n19013), .B(n19058), .ZN(
        n19017) );
  OAI22_X1 U22009 ( .A1(n19100), .A2(n19015), .B1(n19105), .B2(n19014), .ZN(
        n19016) );
  AOI211_X1 U22010 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19117), .A(n19017), .B(
        n19016), .ZN(n19018) );
  OAI21_X1 U22011 ( .B1(n19841), .B2(n19019), .A(n19018), .ZN(P2_U2839) );
  AOI21_X1 U22012 ( .B1(n19021), .B2(n19020), .A(n19841), .ZN(n19032) );
  NAND2_X1 U22013 ( .A1(n19022), .A2(n19021), .ZN(n19029) );
  OAI21_X1 U22014 ( .B1(n19105), .B2(n19023), .A(n19058), .ZN(n19027) );
  OAI22_X1 U22015 ( .A1(n19025), .A2(n19024), .B1(n19888), .B2(n19059), .ZN(
        n19026) );
  AOI211_X1 U22016 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19117), .A(n19027), .B(
        n19026), .ZN(n19028) );
  OAI211_X1 U22017 ( .C1(n19090), .C2(n19030), .A(n19029), .B(n19028), .ZN(
        n19031) );
  AOI21_X1 U22018 ( .B1(n19033), .B2(n19032), .A(n19031), .ZN(n19034) );
  OAI21_X1 U22019 ( .B1(n19035), .B2(n19100), .A(n19034), .ZN(P2_U2840) );
  AOI22_X1 U22020 ( .A1(n19036), .A2(n19125), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19117), .ZN(n19037) );
  OAI211_X1 U22021 ( .C1(n12408), .C2(n19059), .A(n19037), .B(n19058), .ZN(
        n19038) );
  AOI21_X1 U22022 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19130), .A(
        n19038), .ZN(n19044) );
  XOR2_X1 U22023 ( .A(n19040), .B(n19039), .Z(n19042) );
  AOI22_X1 U22024 ( .A1(n19042), .A2(n19080), .B1(n19119), .B2(n19041), .ZN(
        n19043) );
  OAI211_X1 U22025 ( .C1(n19045), .C2(n19100), .A(n19044), .B(n19043), .ZN(
        P2_U2841) );
  NOR2_X1 U22026 ( .A1(n19108), .A2(n19046), .ZN(n19048) );
  XOR2_X1 U22027 ( .A(n19048), .B(n19047), .Z(n19057) );
  AOI22_X1 U22028 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n19117), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19130), .ZN(n19049) );
  OAI21_X1 U22029 ( .B1(n19050), .B2(n19090), .A(n19049), .ZN(n19051) );
  AOI211_X1 U22030 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19122), .A(n19255), 
        .B(n19051), .ZN(n19056) );
  INV_X1 U22031 ( .A(n19052), .ZN(n19054) );
  INV_X1 U22032 ( .A(n19053), .ZN(n19139) );
  AOI22_X1 U22033 ( .A1(n19054), .A2(n19119), .B1(n19121), .B2(n19139), .ZN(
        n19055) );
  OAI211_X1 U22034 ( .C1(n19841), .C2(n19057), .A(n19056), .B(n19055), .ZN(
        P2_U2843) );
  OAI21_X1 U22035 ( .B1(n19880), .B2(n19059), .A(n19058), .ZN(n19062) );
  OAI22_X1 U22036 ( .A1(n19060), .A2(n19090), .B1(n19101), .B2(n12516), .ZN(
        n19061) );
  AOI211_X1 U22037 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19130), .A(
        n19062), .B(n19061), .ZN(n19070) );
  NOR2_X1 U22038 ( .A1(n19108), .A2(n19063), .ZN(n19065) );
  XNOR2_X1 U22039 ( .A(n19065), .B(n19064), .ZN(n19068) );
  INV_X1 U22040 ( .A(n19066), .ZN(n19067) );
  AOI22_X1 U22041 ( .A1(n19068), .A2(n19080), .B1(n19119), .B2(n19067), .ZN(
        n19069) );
  OAI211_X1 U22042 ( .C1(n19100), .C2(n19071), .A(n19070), .B(n19069), .ZN(
        P2_U2845) );
  AOI22_X1 U22043 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19117), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19130), .ZN(n19072) );
  OAI21_X1 U22044 ( .B1(n19073), .B2(n19090), .A(n19072), .ZN(n19074) );
  AOI211_X1 U22045 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19122), .A(n19255), .B(
        n19074), .ZN(n19083) );
  NOR2_X1 U22046 ( .A1(n19108), .A2(n19075), .ZN(n19077) );
  XNOR2_X1 U22047 ( .A(n19077), .B(n19076), .ZN(n19081) );
  INV_X1 U22048 ( .A(n19078), .ZN(n19079) );
  AOI22_X1 U22049 ( .A1(n19081), .A2(n19080), .B1(n19119), .B2(n19079), .ZN(
        n19082) );
  OAI211_X1 U22050 ( .C1(n19100), .C2(n19084), .A(n19083), .B(n19082), .ZN(
        P2_U2847) );
  NOR2_X1 U22051 ( .A1(n19108), .A2(n19085), .ZN(n19087) );
  XOR2_X1 U22052 ( .A(n19087), .B(n19086), .Z(n19097) );
  AOI22_X1 U22053 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19130), .B1(
        P2_EBX_REG_6__SCAN_IN), .B2(n19117), .ZN(n19088) );
  OAI21_X1 U22054 ( .B1(n19090), .B2(n19089), .A(n19088), .ZN(n19091) );
  AOI211_X1 U22055 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19122), .A(n19255), .B(
        n19091), .ZN(n19096) );
  INV_X1 U22056 ( .A(n19092), .ZN(n19094) );
  INV_X1 U22057 ( .A(n19093), .ZN(n19144) );
  AOI22_X1 U22058 ( .A1(n19119), .A2(n19094), .B1(n19121), .B2(n19144), .ZN(
        n19095) );
  OAI211_X1 U22059 ( .C1(n19841), .C2(n19097), .A(n19096), .B(n19095), .ZN(
        P2_U2849) );
  AOI22_X1 U22060 ( .A1(n19125), .A2(n19098), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19130), .ZN(n19115) );
  OAI22_X1 U22061 ( .A1(n19101), .A2(n12495), .B1(n19100), .B2(n19099), .ZN(
        n19102) );
  AOI211_X1 U22062 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19122), .A(n19103), .B(
        n19102), .ZN(n19114) );
  OAI22_X1 U22063 ( .A1(n19148), .A2(n19123), .B1(n19105), .B2(n19104), .ZN(
        n19106) );
  INV_X1 U22064 ( .A(n19106), .ZN(n19113) );
  INV_X1 U22065 ( .A(n19266), .ZN(n19111) );
  NOR2_X1 U22066 ( .A1(n19108), .A2(n19107), .ZN(n19110) );
  AOI21_X1 U22067 ( .B1(n19111), .B2(n19110), .A(n19841), .ZN(n19109) );
  OAI21_X1 U22068 ( .B1(n19111), .B2(n19110), .A(n19109), .ZN(n19112) );
  NAND4_X1 U22069 ( .A1(n19115), .A2(n19114), .A3(n19113), .A4(n19112), .ZN(
        P2_U2851) );
  AOI22_X1 U22070 ( .A1(n19119), .A2(n19118), .B1(P2_EBX_REG_0__SCAN_IN), .B2(
        n19117), .ZN(n19129) );
  INV_X1 U22071 ( .A(n19120), .ZN(n19177) );
  AOI22_X1 U22072 ( .A1(n19122), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19121), 
        .B2(n19177), .ZN(n19128) );
  OR2_X1 U22073 ( .A1(n19953), .A2(n19123), .ZN(n19127) );
  NAND2_X1 U22074 ( .A1(n19125), .A2(n19124), .ZN(n19126) );
  AND4_X1 U22075 ( .A1(n19129), .A2(n19128), .A3(n19127), .A4(n19126), .ZN(
        n19132) );
  NAND2_X1 U22076 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19130), .ZN(
        n19131) );
  OAI211_X1 U22077 ( .C1(n13758), .C2(n19841), .A(n19132), .B(n19131), .ZN(
        P2_U2855) );
  AOI22_X1 U22078 ( .A1(n19134), .A2(BUF2_REG_31__SCAN_IN), .B1(n19173), .B2(
        n10154), .ZN(n19137) );
  AOI22_X1 U22079 ( .A1(n19135), .A2(BUF1_REG_31__SCAN_IN), .B1(n19172), .B2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n19136) );
  NAND2_X1 U22080 ( .A1(n19137), .A2(n19136), .ZN(P2_U2888) );
  INV_X1 U22081 ( .A(n19138), .ZN(n19147) );
  AOI22_X1 U22082 ( .A1(n19147), .A2(n19139), .B1(n19172), .B2(
        P2_EAX_REG_12__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U22083 ( .B1(n19141), .B2(n19180), .A(n19140), .ZN(P2_U2907) );
  AOI22_X1 U22084 ( .A1(n19147), .A2(n19142), .B1(n19172), .B2(
        P2_EAX_REG_7__SCAN_IN), .ZN(n19143) );
  OAI21_X1 U22085 ( .B1(n19318), .B2(n19180), .A(n19143), .ZN(P2_U2912) );
  AOI22_X1 U22086 ( .A1(n19147), .A2(n19144), .B1(n19172), .B2(
        P2_EAX_REG_6__SCAN_IN), .ZN(n19145) );
  OAI21_X1 U22087 ( .B1(n19308), .B2(n19180), .A(n19145), .ZN(P2_U2913) );
  AOI22_X1 U22088 ( .A1(n19147), .A2(n19146), .B1(n19172), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n19152) );
  INV_X1 U22089 ( .A(n19148), .ZN(n19149) );
  NAND3_X1 U22090 ( .A1(n19150), .A2(n19149), .A3(n19175), .ZN(n19151) );
  OAI211_X1 U22091 ( .C1(n19303), .C2(n19180), .A(n19152), .B(n19151), .ZN(
        P2_U2914) );
  AOI22_X1 U22092 ( .A1(n19173), .A2(n19929), .B1(n19172), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19158) );
  AOI21_X1 U22093 ( .B1(n19155), .B2(n19154), .A(n19153), .ZN(n19156) );
  OR2_X1 U22094 ( .A1(n19156), .A2(n19168), .ZN(n19157) );
  OAI211_X1 U22095 ( .C1(n19294), .C2(n19180), .A(n19158), .B(n19157), .ZN(
        P2_U2916) );
  AOI22_X1 U22096 ( .A1(n19173), .A2(n19938), .B1(n19172), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19164) );
  AOI21_X1 U22097 ( .B1(n19161), .B2(n19160), .A(n19159), .ZN(n19162) );
  OR2_X1 U22098 ( .A1(n19162), .A2(n19168), .ZN(n19163) );
  OAI211_X1 U22099 ( .C1(n19291), .C2(n19180), .A(n19164), .B(n19163), .ZN(
        P2_U2917) );
  INV_X1 U22100 ( .A(n19165), .ZN(n19947) );
  AOI22_X1 U22101 ( .A1(n19173), .A2(n19947), .B1(n19172), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19171) );
  AOI21_X1 U22102 ( .B1(n19174), .B2(n19167), .A(n19166), .ZN(n19169) );
  OR2_X1 U22103 ( .A1(n19169), .A2(n19168), .ZN(n19170) );
  OAI211_X1 U22104 ( .C1(n19287), .C2(n19180), .A(n19171), .B(n19170), .ZN(
        P2_U2918) );
  AOI22_X1 U22105 ( .A1(n19173), .A2(n19177), .B1(n19172), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19179) );
  INV_X1 U22106 ( .A(n19174), .ZN(n19176) );
  OAI211_X1 U22107 ( .C1(n19534), .C2(n19177), .A(n19176), .B(n19175), .ZN(
        n19178) );
  OAI211_X1 U22108 ( .C1(n19280), .C2(n19180), .A(n19179), .B(n19178), .ZN(
        P2_U2919) );
  INV_X1 U22109 ( .A(n19181), .ZN(n19182) );
  NAND2_X1 U22110 ( .A1(n19183), .A2(n19182), .ZN(n19184) );
  NAND2_X1 U22111 ( .A1(n19185), .A2(n19184), .ZN(n19186) );
  NOR2_X4 U22112 ( .A1(n19218), .A2(n19251), .ZN(n19237) );
  AND2_X1 U22113 ( .A1(n19237), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22114 ( .A1(n19251), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n19188) );
  OAI21_X1 U22115 ( .B1(n19189), .B2(n19216), .A(n19188), .ZN(P2_U2921) );
  AOI22_X1 U22116 ( .A1(n19251), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19190) );
  OAI21_X1 U22117 ( .B1(n19191), .B2(n19216), .A(n19190), .ZN(P2_U2922) );
  AOI22_X1 U22118 ( .A1(n19251), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19192) );
  OAI21_X1 U22119 ( .B1(n19193), .B2(n19216), .A(n19192), .ZN(P2_U2923) );
  AOI22_X1 U22120 ( .A1(n19251), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U22121 ( .B1(n19195), .B2(n19216), .A(n19194), .ZN(P2_U2924) );
  AOI22_X1 U22122 ( .A1(n19251), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U22123 ( .B1(n19197), .B2(n19216), .A(n19196), .ZN(P2_U2925) );
  AOI22_X1 U22124 ( .A1(n19251), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22125 ( .B1(n19199), .B2(n19216), .A(n19198), .ZN(P2_U2926) );
  INV_X1 U22126 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19201) );
  AOI22_X1 U22127 ( .A1(n19251), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U22128 ( .B1(n19201), .B2(n19216), .A(n19200), .ZN(P2_U2927) );
  INV_X1 U22129 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19203) );
  AOI22_X1 U22130 ( .A1(n19251), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19202) );
  OAI21_X1 U22131 ( .B1(n19203), .B2(n19216), .A(n19202), .ZN(P2_U2928) );
  INV_X1 U22132 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19205) );
  AOI22_X1 U22133 ( .A1(n19251), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U22134 ( .B1(n19205), .B2(n19216), .A(n19204), .ZN(P2_U2929) );
  INV_X1 U22135 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19207) );
  AOI22_X1 U22136 ( .A1(n19251), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19206) );
  OAI21_X1 U22137 ( .B1(n19207), .B2(n19216), .A(n19206), .ZN(P2_U2930) );
  INV_X1 U22138 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19209) );
  AOI22_X1 U22139 ( .A1(n19251), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19208) );
  OAI21_X1 U22140 ( .B1(n19209), .B2(n19216), .A(n19208), .ZN(P2_U2931) );
  INV_X1 U22141 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19211) );
  AOI22_X1 U22142 ( .A1(n19251), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19210) );
  OAI21_X1 U22143 ( .B1(n19211), .B2(n19216), .A(n19210), .ZN(P2_U2932) );
  INV_X1 U22144 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19213) );
  AOI22_X1 U22145 ( .A1(n19251), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19212) );
  OAI21_X1 U22146 ( .B1(n19213), .B2(n19216), .A(n19212), .ZN(P2_U2933) );
  INV_X1 U22147 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n20998) );
  AOI22_X1 U22148 ( .A1(n19251), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19214) );
  OAI21_X1 U22149 ( .B1(n20998), .B2(n19216), .A(n19214), .ZN(P2_U2934) );
  INV_X1 U22150 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19217) );
  AOI22_X1 U22151 ( .A1(n19251), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19215) );
  OAI21_X1 U22152 ( .B1(n19217), .B2(n19216), .A(n19215), .ZN(P2_U2935) );
  AOI22_X1 U22153 ( .A1(n19251), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19219) );
  OAI21_X1 U22154 ( .B1(n19220), .B2(n19253), .A(n19219), .ZN(P2_U2936) );
  AOI22_X1 U22155 ( .A1(n19251), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19221) );
  OAI21_X1 U22156 ( .B1(n19222), .B2(n19253), .A(n19221), .ZN(P2_U2937) );
  AOI22_X1 U22157 ( .A1(n19251), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19223) );
  OAI21_X1 U22158 ( .B1(n19224), .B2(n19253), .A(n19223), .ZN(P2_U2938) );
  INV_X1 U22159 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19226) );
  AOI22_X1 U22160 ( .A1(n19244), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19225) );
  OAI21_X1 U22161 ( .B1(n19226), .B2(n19253), .A(n19225), .ZN(P2_U2939) );
  AOI22_X1 U22162 ( .A1(n19244), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19227) );
  OAI21_X1 U22163 ( .B1(n19228), .B2(n19253), .A(n19227), .ZN(P2_U2940) );
  AOI22_X1 U22164 ( .A1(n19244), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19229) );
  OAI21_X1 U22165 ( .B1(n19230), .B2(n19253), .A(n19229), .ZN(P2_U2941) );
  AOI22_X1 U22166 ( .A1(n19244), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19231) );
  OAI21_X1 U22167 ( .B1(n19232), .B2(n19253), .A(n19231), .ZN(P2_U2942) );
  AOI22_X1 U22168 ( .A1(n19244), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19233) );
  OAI21_X1 U22169 ( .B1(n19234), .B2(n19253), .A(n19233), .ZN(P2_U2943) );
  INV_X1 U22170 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19236) );
  AOI22_X1 U22171 ( .A1(n19244), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19235) );
  OAI21_X1 U22172 ( .B1(n19236), .B2(n19253), .A(n19235), .ZN(P2_U2944) );
  INV_X1 U22173 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19239) );
  AOI22_X1 U22174 ( .A1(n19244), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19238) );
  OAI21_X1 U22175 ( .B1(n19239), .B2(n19253), .A(n19238), .ZN(P2_U2945) );
  INV_X1 U22176 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19241) );
  AOI22_X1 U22177 ( .A1(n19244), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19240) );
  OAI21_X1 U22178 ( .B1(n19241), .B2(n19253), .A(n19240), .ZN(P2_U2946) );
  INV_X1 U22179 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19243) );
  AOI22_X1 U22180 ( .A1(n19244), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19242) );
  OAI21_X1 U22181 ( .B1(n19243), .B2(n19253), .A(n19242), .ZN(P2_U2947) );
  INV_X1 U22182 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19246) );
  AOI22_X1 U22183 ( .A1(n19244), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19245) );
  OAI21_X1 U22184 ( .B1(n19246), .B2(n19253), .A(n19245), .ZN(P2_U2948) );
  INV_X1 U22185 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19248) );
  AOI22_X1 U22186 ( .A1(n19251), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19247) );
  OAI21_X1 U22187 ( .B1(n19248), .B2(n19253), .A(n19247), .ZN(P2_U2949) );
  INV_X1 U22188 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19250) );
  AOI22_X1 U22189 ( .A1(n19251), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19249) );
  OAI21_X1 U22190 ( .B1(n19250), .B2(n19253), .A(n19249), .ZN(P2_U2950) );
  AOI22_X1 U22191 ( .A1(n19251), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19237), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19252) );
  OAI21_X1 U22192 ( .B1(n19254), .B2(n19253), .A(n19252), .ZN(P2_U2951) );
  AOI22_X1 U22193 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19256), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19255), .ZN(n19265) );
  OAI22_X1 U22194 ( .A1(n19260), .A2(n19259), .B1(n19258), .B2(n19257), .ZN(
        n19261) );
  AOI21_X1 U22195 ( .B1(n19263), .B2(n19262), .A(n19261), .ZN(n19264) );
  OAI211_X1 U22196 ( .C1(n19267), .C2(n19266), .A(n19265), .B(n19264), .ZN(
        P2_U3010) );
  AOI22_X1 U22197 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19311), .ZN(n19740) );
  NOR2_X2 U22198 ( .A1(n11750), .A2(n19315), .ZN(n19774) );
  NAND2_X1 U22199 ( .A1(n19933), .A2(n19940), .ZN(n19380) );
  OR2_X1 U22200 ( .A1(n19380), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19326) );
  NOR2_X1 U22201 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19326), .ZN(
        n19317) );
  AOI22_X1 U22202 ( .A1(n19784), .A2(n19831), .B1(n19774), .B2(n19317), .ZN(
        n19286) );
  INV_X1 U22203 ( .A(n19349), .ZN(n19272) );
  OAI21_X1 U22204 ( .B1(n19831), .B2(n19272), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19273) );
  NAND2_X1 U22205 ( .A1(n19273), .A2(n19928), .ZN(n19284) );
  NOR2_X1 U22206 ( .A1(n19933), .A2(n19274), .ZN(n19826) );
  NOR2_X1 U22207 ( .A1(n19826), .A2(n19317), .ZN(n19283) );
  INV_X1 U22208 ( .A(n19283), .ZN(n19279) );
  INV_X1 U22209 ( .A(n19275), .ZN(n19281) );
  OAI21_X1 U22210 ( .B1(n19281), .B2(n19951), .A(n19509), .ZN(n19277) );
  INV_X1 U22211 ( .A(n19317), .ZN(n19276) );
  AOI21_X1 U22212 ( .B1(n19277), .B2(n19276), .A(n19778), .ZN(n19278) );
  NOR2_X2 U22213 ( .A1(n19280), .A2(n19778), .ZN(n19775) );
  OAI21_X1 U22214 ( .B1(n19281), .B2(n19317), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19282) );
  AOI22_X1 U22215 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19320), .B1(
        n19775), .B2(n19319), .ZN(n19285) );
  OAI211_X1 U22216 ( .C1(n19787), .C2(n19349), .A(n19286), .B(n19285), .ZN(
        P2_U3048) );
  AOI22_X2 U22217 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19311), .ZN(n19793) );
  AOI22_X1 U22218 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19311), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19312), .ZN(n19704) );
  NOR2_X2 U22219 ( .A1(n11776), .A2(n19315), .ZN(n19788) );
  AOI22_X1 U22220 ( .A1(n19790), .A2(n19831), .B1(n19788), .B2(n19317), .ZN(
        n19289) );
  NOR2_X2 U22221 ( .A1(n19287), .A2(n19778), .ZN(n19789) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19320), .B1(
        n19789), .B2(n19319), .ZN(n19288) );
  OAI211_X1 U22223 ( .C1(n19793), .C2(n19349), .A(n19289), .B(n19288), .ZN(
        P2_U3049) );
  AOI22_X2 U22224 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19311), .ZN(n19746) );
  AOI22_X1 U22225 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19311), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19312), .ZN(n19799) );
  AOI22_X1 U22226 ( .A1(n19743), .A2(n19831), .B1(n9852), .B2(n19317), .ZN(
        n19293) );
  NOR2_X2 U22227 ( .A1(n19291), .A2(n19778), .ZN(n19795) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19320), .B1(
        n19795), .B2(n19319), .ZN(n19292) );
  OAI211_X1 U22229 ( .C1(n19746), .C2(n19349), .A(n19293), .B(n19292), .ZN(
        P2_U3050) );
  AOI22_X2 U22230 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19311), .ZN(n19750) );
  AOI22_X1 U22231 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19311), .ZN(n19805) );
  NOR2_X2 U22232 ( .A1(n11751), .A2(n19315), .ZN(n19800) );
  AOI22_X1 U22233 ( .A1(n19747), .A2(n19831), .B1(n19800), .B2(n19317), .ZN(
        n19296) );
  NOR2_X2 U22234 ( .A1(n19294), .A2(n19778), .ZN(n19801) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19320), .B1(
        n19801), .B2(n19319), .ZN(n19295) );
  OAI211_X1 U22236 ( .C1(n19750), .C2(n19349), .A(n19296), .B(n19295), .ZN(
        P2_U3051) );
  AOI22_X1 U22237 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19311), .ZN(n19712) );
  AOI22_X1 U22238 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19311), .ZN(n19811) );
  INV_X1 U22239 ( .A(n19811), .ZN(n19709) );
  NOR2_X2 U22240 ( .A1(n19297), .A2(n19315), .ZN(n19806) );
  AOI22_X1 U22241 ( .A1(n19709), .A2(n19831), .B1(n19806), .B2(n19317), .ZN(
        n19301) );
  INV_X1 U22242 ( .A(n19298), .ZN(n19299) );
  NOR2_X2 U22243 ( .A1(n19299), .A2(n19778), .ZN(n19807) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19320), .B1(
        n19807), .B2(n19319), .ZN(n19300) );
  OAI211_X1 U22245 ( .C1(n19712), .C2(n19349), .A(n19301), .B(n19300), .ZN(
        P2_U3052) );
  AOI22_X1 U22246 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19311), .ZN(n19756) );
  AOI22_X1 U22247 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19311), .ZN(n19817) );
  INV_X1 U22248 ( .A(n19817), .ZN(n19753) );
  NOR2_X2 U22249 ( .A1(n19302), .A2(n19315), .ZN(n19812) );
  AOI22_X1 U22250 ( .A1(n19753), .A2(n19831), .B1(n19812), .B2(n19317), .ZN(
        n19305) );
  NOR2_X2 U22251 ( .A1(n19303), .A2(n19778), .ZN(n19813) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19320), .B1(
        n19813), .B2(n19319), .ZN(n19304) );
  OAI211_X1 U22253 ( .C1(n19756), .C2(n19349), .A(n19305), .B(n19304), .ZN(
        P2_U3053) );
  AOI22_X1 U22254 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19311), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19312), .ZN(n19761) );
  INV_X1 U22255 ( .A(n19761), .ZN(n19820) );
  NOR2_X2 U22256 ( .A1(n19307), .A2(n19315), .ZN(n19818) );
  AOI22_X1 U22257 ( .A1(n19820), .A2(n19831), .B1(n19818), .B2(n19317), .ZN(
        n19310) );
  NOR2_X2 U22258 ( .A1(n19308), .A2(n19778), .ZN(n19819) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19320), .B1(
        n19819), .B2(n19319), .ZN(n19309) );
  OAI211_X1 U22260 ( .C1(n19825), .C2(n19349), .A(n19310), .B(n19309), .ZN(
        P2_U3054) );
  AOI22_X1 U22261 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19312), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19311), .ZN(n19769) );
  NOR2_X2 U22262 ( .A1(n19316), .A2(n19315), .ZN(n19827) );
  AOI22_X1 U22263 ( .A1(n19764), .A2(n19831), .B1(n19827), .B2(n19317), .ZN(
        n19322) );
  NOR2_X2 U22264 ( .A1(n19318), .A2(n19778), .ZN(n19828) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19320), .B1(
        n19828), .B2(n19319), .ZN(n19321) );
  OAI211_X1 U22266 ( .C1(n19769), .C2(n19349), .A(n19322), .B(n19321), .ZN(
        P2_U3055) );
  INV_X1 U22267 ( .A(n19325), .ZN(n19323) );
  NOR2_X1 U22268 ( .A1(n19564), .A2(n19380), .ZN(n19344) );
  OAI21_X1 U22269 ( .B1(n19323), .B2(n19344), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19324) );
  OAI21_X1 U22270 ( .B1(n19326), .B2(n19728), .A(n19324), .ZN(n19345) );
  AOI22_X1 U22271 ( .A1(n19345), .A2(n19775), .B1(n19774), .B2(n19344), .ZN(
        n19331) );
  AOI21_X1 U22272 ( .B1(n19325), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19328) );
  NAND2_X1 U22273 ( .A1(n19565), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19507) );
  OAI21_X1 U22274 ( .B1(n19507), .B2(n19566), .A(n19326), .ZN(n19327) );
  OAI211_X1 U22275 ( .C1(n19344), .C2(n19328), .A(n19327), .B(n19731), .ZN(
        n19346) );
  NAND2_X1 U22276 ( .A1(n19329), .A2(n19513), .ZN(n19354) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19346), .B1(
        n19376), .B2(n19725), .ZN(n19330) );
  OAI211_X1 U22278 ( .C1(n19740), .C2(n19349), .A(n19331), .B(n19330), .ZN(
        P2_U3056) );
  AOI22_X1 U22279 ( .A1(n19345), .A2(n19789), .B1(n19788), .B2(n19344), .ZN(
        n19333) );
  INV_X1 U22280 ( .A(n19793), .ZN(n19701) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19346), .B1(
        n19376), .B2(n19701), .ZN(n19332) );
  OAI211_X1 U22282 ( .C1(n19704), .C2(n19349), .A(n19333), .B(n19332), .ZN(
        P2_U3057) );
  AOI22_X1 U22283 ( .A1(n19345), .A2(n19795), .B1(n9852), .B2(n19344), .ZN(
        n19335) );
  INV_X1 U22284 ( .A(n19746), .ZN(n19796) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19346), .B1(
        n19376), .B2(n19796), .ZN(n19334) );
  OAI211_X1 U22286 ( .C1(n19799), .C2(n19349), .A(n19335), .B(n19334), .ZN(
        P2_U3058) );
  AOI22_X1 U22287 ( .A1(n19345), .A2(n19801), .B1(n19800), .B2(n19344), .ZN(
        n19337) );
  INV_X1 U22288 ( .A(n19750), .ZN(n19802) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19346), .B1(
        n19376), .B2(n19802), .ZN(n19336) );
  OAI211_X1 U22290 ( .C1(n19805), .C2(n19349), .A(n19337), .B(n19336), .ZN(
        P2_U3059) );
  AOI22_X1 U22291 ( .A1(n19345), .A2(n19807), .B1(n19806), .B2(n19344), .ZN(
        n19339) );
  INV_X1 U22292 ( .A(n19712), .ZN(n19808) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19346), .B1(
        n19376), .B2(n19808), .ZN(n19338) );
  OAI211_X1 U22294 ( .C1(n19811), .C2(n19349), .A(n19339), .B(n19338), .ZN(
        P2_U3060) );
  AOI22_X1 U22295 ( .A1(n19345), .A2(n19813), .B1(n19812), .B2(n19344), .ZN(
        n19341) );
  INV_X1 U22296 ( .A(n19756), .ZN(n19814) );
  AOI22_X1 U22297 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19346), .B1(
        n19376), .B2(n19814), .ZN(n19340) );
  OAI211_X1 U22298 ( .C1(n19817), .C2(n19349), .A(n19341), .B(n19340), .ZN(
        P2_U3061) );
  AOI22_X1 U22299 ( .A1(n19345), .A2(n19819), .B1(n19818), .B2(n19344), .ZN(
        n19343) );
  AOI22_X1 U22300 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19346), .B1(
        n19376), .B2(n19757), .ZN(n19342) );
  OAI211_X1 U22301 ( .C1(n19761), .C2(n19349), .A(n19343), .B(n19342), .ZN(
        P2_U3062) );
  AOI22_X1 U22302 ( .A1(n19345), .A2(n19828), .B1(n19827), .B2(n19344), .ZN(
        n19348) );
  AOI22_X1 U22303 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19346), .B1(
        n19376), .B2(n19830), .ZN(n19347) );
  OAI211_X1 U22304 ( .C1(n19836), .C2(n19349), .A(n19348), .B(n19347), .ZN(
        P2_U3063) );
  INV_X1 U22305 ( .A(n19350), .ZN(n19353) );
  NOR2_X1 U22306 ( .A1(n19597), .A2(n19380), .ZN(n19374) );
  OAI21_X1 U22307 ( .B1(n19353), .B2(n19374), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19352) );
  NOR2_X1 U22308 ( .A1(n19600), .A2(n19380), .ZN(n19355) );
  INV_X1 U22309 ( .A(n19355), .ZN(n19351) );
  NAND2_X1 U22310 ( .A1(n19352), .A2(n19351), .ZN(n19375) );
  AOI22_X1 U22311 ( .A1(n19375), .A2(n19775), .B1(n19774), .B2(n19374), .ZN(
        n19361) );
  AOI21_X1 U22312 ( .B1(n19353), .B2(n19509), .A(n19374), .ZN(n19358) );
  AOI21_X1 U22313 ( .B1(n19409), .B2(n19354), .A(n19661), .ZN(n19356) );
  NOR2_X1 U22314 ( .A1(n19356), .A2(n19355), .ZN(n19357) );
  MUX2_X1 U22315 ( .A(n19358), .B(n19357), .S(n19928), .Z(n19359) );
  OR2_X1 U22316 ( .A1(n19359), .A2(n19778), .ZN(n19377) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19377), .B1(
        n19376), .B2(n19784), .ZN(n19360) );
  OAI211_X1 U22318 ( .C1(n19787), .C2(n19409), .A(n19361), .B(n19360), .ZN(
        P2_U3064) );
  AOI22_X1 U22319 ( .A1(n19375), .A2(n19789), .B1(n19788), .B2(n19374), .ZN(
        n19363) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19377), .B1(
        n19376), .B2(n19790), .ZN(n19362) );
  OAI211_X1 U22321 ( .C1(n19793), .C2(n19409), .A(n19363), .B(n19362), .ZN(
        P2_U3065) );
  AOI22_X1 U22322 ( .A1(n19375), .A2(n19795), .B1(n9852), .B2(n19374), .ZN(
        n19365) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19377), .B1(
        n19376), .B2(n19743), .ZN(n19364) );
  OAI211_X1 U22324 ( .C1(n19746), .C2(n19409), .A(n19365), .B(n19364), .ZN(
        P2_U3066) );
  AOI22_X1 U22325 ( .A1(n19375), .A2(n19801), .B1(n19800), .B2(n19374), .ZN(
        n19367) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19377), .B1(
        n19376), .B2(n19747), .ZN(n19366) );
  OAI211_X1 U22327 ( .C1(n19750), .C2(n19409), .A(n19367), .B(n19366), .ZN(
        P2_U3067) );
  AOI22_X1 U22328 ( .A1(n19375), .A2(n19807), .B1(n19806), .B2(n19374), .ZN(
        n19369) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19377), .B1(
        n19376), .B2(n19709), .ZN(n19368) );
  OAI211_X1 U22330 ( .C1(n19712), .C2(n19409), .A(n19369), .B(n19368), .ZN(
        P2_U3068) );
  AOI22_X1 U22331 ( .A1(n19375), .A2(n19813), .B1(n19812), .B2(n19374), .ZN(
        n19371) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19377), .B1(
        n19376), .B2(n19753), .ZN(n19370) );
  OAI211_X1 U22333 ( .C1(n19756), .C2(n19409), .A(n19371), .B(n19370), .ZN(
        P2_U3069) );
  AOI22_X1 U22334 ( .A1(n19375), .A2(n19819), .B1(n19818), .B2(n19374), .ZN(
        n19373) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19377), .B1(
        n19376), .B2(n19820), .ZN(n19372) );
  OAI211_X1 U22336 ( .C1(n19825), .C2(n19409), .A(n19373), .B(n19372), .ZN(
        P2_U3070) );
  AOI22_X1 U22337 ( .A1(n19375), .A2(n19828), .B1(n19827), .B2(n19374), .ZN(
        n19379) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19377), .B1(
        n19376), .B2(n19764), .ZN(n19378) );
  OAI211_X1 U22339 ( .C1(n19769), .C2(n19409), .A(n19379), .B(n19378), .ZN(
        P2_U3071) );
  INV_X1 U22340 ( .A(n19409), .ZN(n19399) );
  NOR2_X1 U22341 ( .A1(n19629), .A2(n19380), .ZN(n19404) );
  AOI22_X1 U22342 ( .A1(n19784), .A2(n19399), .B1(n19404), .B2(n19774), .ZN(
        n19390) );
  OAI21_X1 U22343 ( .B1(n19507), .B2(n19635), .A(n19928), .ZN(n19388) );
  NOR2_X1 U22344 ( .A1(n19949), .A2(n19380), .ZN(n19383) );
  INV_X1 U22345 ( .A(n19404), .ZN(n19381) );
  OAI211_X1 U22346 ( .C1(n19384), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19381), 
        .B(n19728), .ZN(n19382) );
  OAI211_X1 U22347 ( .C1(n19388), .C2(n19383), .A(n19731), .B(n19382), .ZN(
        n19406) );
  INV_X1 U22348 ( .A(n19383), .ZN(n19387) );
  INV_X1 U22349 ( .A(n19384), .ZN(n19385) );
  OAI21_X1 U22350 ( .B1(n19385), .B2(n19404), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19386) );
  OAI21_X1 U22351 ( .B1(n19388), .B2(n19387), .A(n19386), .ZN(n19405) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19406), .B1(
        n19775), .B2(n19405), .ZN(n19389) );
  OAI211_X1 U22353 ( .C1(n19787), .C2(n19441), .A(n19390), .B(n19389), .ZN(
        P2_U3072) );
  AOI22_X1 U22354 ( .A1(n19399), .A2(n19790), .B1(n19404), .B2(n19788), .ZN(
        n19392) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19406), .B1(
        n19789), .B2(n19405), .ZN(n19391) );
  OAI211_X1 U22356 ( .C1(n19793), .C2(n19441), .A(n19392), .B(n19391), .ZN(
        P2_U3073) );
  AOI22_X1 U22357 ( .A1(n19399), .A2(n19743), .B1(n19404), .B2(n9852), .ZN(
        n19394) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19406), .B1(
        n19795), .B2(n19405), .ZN(n19393) );
  OAI211_X1 U22359 ( .C1(n19746), .C2(n19441), .A(n19394), .B(n19393), .ZN(
        P2_U3074) );
  AOI22_X1 U22360 ( .A1(n19399), .A2(n19747), .B1(n19404), .B2(n19800), .ZN(
        n19396) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19406), .B1(
        n19801), .B2(n19405), .ZN(n19395) );
  OAI211_X1 U22362 ( .C1(n19750), .C2(n19441), .A(n19396), .B(n19395), .ZN(
        P2_U3075) );
  AOI22_X1 U22363 ( .A1(n19808), .A2(n19431), .B1(n19404), .B2(n19806), .ZN(
        n19398) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19406), .B1(
        n19807), .B2(n19405), .ZN(n19397) );
  OAI211_X1 U22365 ( .C1(n19811), .C2(n19409), .A(n19398), .B(n19397), .ZN(
        P2_U3076) );
  AOI22_X1 U22366 ( .A1(n19753), .A2(n19399), .B1(n19404), .B2(n19812), .ZN(
        n19401) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19406), .B1(
        n19813), .B2(n19405), .ZN(n19400) );
  OAI211_X1 U22368 ( .C1(n19756), .C2(n19441), .A(n19401), .B(n19400), .ZN(
        P2_U3077) );
  AOI22_X1 U22369 ( .A1(n19757), .A2(n19431), .B1(n19404), .B2(n19818), .ZN(
        n19403) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19406), .B1(
        n19819), .B2(n19405), .ZN(n19402) );
  OAI211_X1 U22371 ( .C1(n19761), .C2(n19409), .A(n19403), .B(n19402), .ZN(
        P2_U3078) );
  AOI22_X1 U22372 ( .A1(n19830), .A2(n19431), .B1(n19404), .B2(n19827), .ZN(
        n19408) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19406), .B1(
        n19828), .B2(n19405), .ZN(n19407) );
  OAI211_X1 U22374 ( .C1(n19836), .C2(n19409), .A(n19408), .B(n19407), .ZN(
        P2_U3079) );
  NOR3_X1 U22375 ( .A1(n19940), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19443) );
  INV_X1 U22376 ( .A(n19443), .ZN(n19447) );
  NOR2_X1 U22377 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19447), .ZN(
        n19436) );
  AOI22_X1 U22378 ( .A1(n19725), .A2(n19459), .B1(n19774), .B2(n19436), .ZN(
        n19422) );
  OAI21_X1 U22379 ( .B1(n19459), .B2(n19431), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19410) );
  NAND2_X1 U22380 ( .A1(n19410), .A2(n19928), .ZN(n19420) );
  NAND2_X1 U22381 ( .A1(n19412), .A2(n19411), .ZN(n19659) );
  NOR2_X1 U22382 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19659), .ZN(
        n19415) );
  INV_X1 U22383 ( .A(n19436), .ZN(n19413) );
  OAI211_X1 U22384 ( .C1(n19416), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19413), 
        .B(n19728), .ZN(n19414) );
  OAI211_X1 U22385 ( .C1(n19420), .C2(n19415), .A(n19731), .B(n19414), .ZN(
        n19438) );
  INV_X1 U22386 ( .A(n19415), .ZN(n19419) );
  INV_X1 U22387 ( .A(n19416), .ZN(n19417) );
  OAI21_X1 U22388 ( .B1(n19417), .B2(n19436), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19418) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19438), .B1(
        n19775), .B2(n19437), .ZN(n19421) );
  OAI211_X1 U22390 ( .C1(n19740), .C2(n19441), .A(n19422), .B(n19421), .ZN(
        P2_U3080) );
  AOI22_X1 U22391 ( .A1(n19701), .A2(n19459), .B1(n19788), .B2(n19436), .ZN(
        n19424) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19438), .B1(
        n19789), .B2(n19437), .ZN(n19423) );
  OAI211_X1 U22393 ( .C1(n19704), .C2(n19441), .A(n19424), .B(n19423), .ZN(
        P2_U3081) );
  AOI22_X1 U22394 ( .A1(n19431), .A2(n19743), .B1(n9852), .B2(n19436), .ZN(
        n19426) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19438), .B1(
        n19795), .B2(n19437), .ZN(n19425) );
  OAI211_X1 U22396 ( .C1(n19746), .C2(n19470), .A(n19426), .B(n19425), .ZN(
        P2_U3082) );
  AOI22_X1 U22397 ( .A1(n19431), .A2(n19747), .B1(n19800), .B2(n19436), .ZN(
        n19428) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19438), .B1(
        n19801), .B2(n19437), .ZN(n19427) );
  OAI211_X1 U22399 ( .C1(n19750), .C2(n19470), .A(n19428), .B(n19427), .ZN(
        P2_U3083) );
  AOI22_X1 U22400 ( .A1(n19808), .A2(n19459), .B1(n19806), .B2(n19436), .ZN(
        n19430) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19438), .B1(
        n19807), .B2(n19437), .ZN(n19429) );
  OAI211_X1 U22402 ( .C1(n19811), .C2(n19441), .A(n19430), .B(n19429), .ZN(
        P2_U3084) );
  AOI22_X1 U22403 ( .A1(n19753), .A2(n19431), .B1(n19812), .B2(n19436), .ZN(
        n19433) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19438), .B1(
        n19813), .B2(n19437), .ZN(n19432) );
  OAI211_X1 U22405 ( .C1(n19756), .C2(n19470), .A(n19433), .B(n19432), .ZN(
        P2_U3085) );
  AOI22_X1 U22406 ( .A1(n19757), .A2(n19459), .B1(n19818), .B2(n19436), .ZN(
        n19435) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19438), .B1(
        n19819), .B2(n19437), .ZN(n19434) );
  OAI211_X1 U22408 ( .C1(n19761), .C2(n19441), .A(n19435), .B(n19434), .ZN(
        P2_U3086) );
  AOI22_X1 U22409 ( .A1(n19830), .A2(n19459), .B1(n19827), .B2(n19436), .ZN(
        n19440) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19438), .B1(
        n19828), .B2(n19437), .ZN(n19439) );
  OAI211_X1 U22411 ( .C1(n19836), .C2(n19441), .A(n19440), .B(n19439), .ZN(
        P2_U3087) );
  NAND2_X1 U22412 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19443), .ZN(
        n19478) );
  INV_X1 U22413 ( .A(n19478), .ZN(n19465) );
  AOI22_X1 U22414 ( .A1(n19725), .A2(n19497), .B1(n19774), .B2(n19465), .ZN(
        n19450) );
  OAI21_X1 U22415 ( .B1(n19507), .B2(n19687), .A(n19928), .ZN(n19448) );
  OAI211_X1 U22416 ( .C1(n19444), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19478), 
        .B(n19728), .ZN(n19442) );
  OAI211_X1 U22417 ( .C1(n19448), .C2(n19443), .A(n19731), .B(n19442), .ZN(
        n19467) );
  INV_X1 U22418 ( .A(n19444), .ZN(n19445) );
  OAI21_X1 U22419 ( .B1(n19445), .B2(n19465), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19446) );
  OAI21_X1 U22420 ( .B1(n19448), .B2(n19447), .A(n19446), .ZN(n19466) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19467), .B1(
        n19775), .B2(n19466), .ZN(n19449) );
  OAI211_X1 U22422 ( .C1(n19740), .C2(n19470), .A(n19450), .B(n19449), .ZN(
        P2_U3088) );
  AOI22_X1 U22423 ( .A1(n19701), .A2(n19497), .B1(n19788), .B2(n19465), .ZN(
        n19452) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19467), .B1(
        n19789), .B2(n19466), .ZN(n19451) );
  OAI211_X1 U22425 ( .C1(n19704), .C2(n19470), .A(n19452), .B(n19451), .ZN(
        P2_U3089) );
  AOI22_X1 U22426 ( .A1(n19796), .A2(n19497), .B1(n9852), .B2(n19465), .ZN(
        n19454) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19467), .B1(
        n19795), .B2(n19466), .ZN(n19453) );
  OAI211_X1 U22428 ( .C1(n19799), .C2(n19470), .A(n19454), .B(n19453), .ZN(
        P2_U3090) );
  INV_X1 U22429 ( .A(n19497), .ZN(n19462) );
  AOI22_X1 U22430 ( .A1(n19459), .A2(n19747), .B1(n19800), .B2(n19465), .ZN(
        n19456) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19467), .B1(
        n19801), .B2(n19466), .ZN(n19455) );
  OAI211_X1 U22432 ( .C1(n19750), .C2(n19462), .A(n19456), .B(n19455), .ZN(
        P2_U3091) );
  AOI22_X1 U22433 ( .A1(n19808), .A2(n19497), .B1(n19806), .B2(n19465), .ZN(
        n19458) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19467), .B1(
        n19807), .B2(n19466), .ZN(n19457) );
  OAI211_X1 U22435 ( .C1(n19811), .C2(n19470), .A(n19458), .B(n19457), .ZN(
        P2_U3092) );
  AOI22_X1 U22436 ( .A1(n19753), .A2(n19459), .B1(n19812), .B2(n19465), .ZN(
        n19461) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19467), .B1(
        n19813), .B2(n19466), .ZN(n19460) );
  OAI211_X1 U22438 ( .C1(n19756), .C2(n19462), .A(n19461), .B(n19460), .ZN(
        P2_U3093) );
  AOI22_X1 U22439 ( .A1(n19757), .A2(n19497), .B1(n19818), .B2(n19465), .ZN(
        n19464) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19467), .B1(
        n19819), .B2(n19466), .ZN(n19463) );
  OAI211_X1 U22441 ( .C1(n19761), .C2(n19470), .A(n19464), .B(n19463), .ZN(
        P2_U3094) );
  AOI22_X1 U22442 ( .A1(n19830), .A2(n19497), .B1(n19827), .B2(n19465), .ZN(
        n19469) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19467), .B1(
        n19828), .B2(n19466), .ZN(n19468) );
  OAI211_X1 U22444 ( .C1(n19836), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U3095) );
  INV_X1 U22445 ( .A(n19471), .ZN(n19472) );
  MUX2_X1 U22446 ( .A(n19478), .B(n19475), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19474) );
  INV_X1 U22447 ( .A(n19512), .ZN(n19505) );
  NOR2_X1 U22448 ( .A1(n19505), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19495) );
  INV_X1 U22449 ( .A(n19495), .ZN(n19473) );
  AOI21_X1 U22450 ( .B1(n19474), .B2(n19473), .A(n19504), .ZN(n19496) );
  AOI22_X1 U22451 ( .A1(n19496), .A2(n19775), .B1(n19774), .B2(n19495), .ZN(
        n19482) );
  OAI21_X1 U22452 ( .B1(n19522), .B2(n19497), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19479) );
  INV_X1 U22453 ( .A(n19475), .ZN(n19476) );
  OAI21_X1 U22454 ( .B1(n19476), .B2(n19951), .A(n19509), .ZN(n19477) );
  AOI21_X1 U22455 ( .B1(n19479), .B2(n19478), .A(n19477), .ZN(n19480) );
  OAI21_X1 U22456 ( .B1(n19495), .B2(n19480), .A(n19731), .ZN(n19498) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19784), .ZN(n19481) );
  OAI211_X1 U22458 ( .C1(n19787), .C2(n19533), .A(n19482), .B(n19481), .ZN(
        P2_U3096) );
  AOI22_X1 U22459 ( .A1(n19496), .A2(n19789), .B1(n19788), .B2(n19495), .ZN(
        n19484) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19790), .ZN(n19483) );
  OAI211_X1 U22461 ( .C1(n19793), .C2(n19533), .A(n19484), .B(n19483), .ZN(
        P2_U3097) );
  AOI22_X1 U22462 ( .A1(n19496), .A2(n19795), .B1(n9852), .B2(n19495), .ZN(
        n19486) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19743), .ZN(n19485) );
  OAI211_X1 U22464 ( .C1(n19746), .C2(n19533), .A(n19486), .B(n19485), .ZN(
        P2_U3098) );
  AOI22_X1 U22465 ( .A1(n19496), .A2(n19801), .B1(n19800), .B2(n19495), .ZN(
        n19488) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19747), .ZN(n19487) );
  OAI211_X1 U22467 ( .C1(n19750), .C2(n19533), .A(n19488), .B(n19487), .ZN(
        P2_U3099) );
  AOI22_X1 U22468 ( .A1(n19496), .A2(n19807), .B1(n19806), .B2(n19495), .ZN(
        n19490) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19709), .ZN(n19489) );
  OAI211_X1 U22470 ( .C1(n19712), .C2(n19533), .A(n19490), .B(n19489), .ZN(
        P2_U3100) );
  AOI22_X1 U22471 ( .A1(n19496), .A2(n19813), .B1(n19812), .B2(n19495), .ZN(
        n19492) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19753), .ZN(n19491) );
  OAI211_X1 U22473 ( .C1(n19756), .C2(n19533), .A(n19492), .B(n19491), .ZN(
        P2_U3101) );
  AOI22_X1 U22474 ( .A1(n19496), .A2(n19819), .B1(n19818), .B2(n19495), .ZN(
        n19494) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19820), .ZN(n19493) );
  OAI211_X1 U22476 ( .C1(n19825), .C2(n19533), .A(n19494), .B(n19493), .ZN(
        P2_U3102) );
  AOI22_X1 U22477 ( .A1(n19496), .A2(n19828), .B1(n19827), .B2(n19495), .ZN(
        n19500) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19764), .ZN(n19499) );
  OAI211_X1 U22479 ( .C1(n19769), .C2(n19533), .A(n19500), .B(n19499), .ZN(
        P2_U3103) );
  AND2_X1 U22480 ( .A1(n19506), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19501) );
  NAND2_X1 U22481 ( .A1(n19502), .A2(n19501), .ZN(n19508) );
  INV_X1 U22482 ( .A(n19508), .ZN(n19503) );
  AOI211_X2 U22483 ( .C1(n19951), .C2(n19505), .A(n19504), .B(n19503), .ZN(
        n19529) );
  INV_X1 U22484 ( .A(n19506), .ZN(n19538) );
  AOI22_X1 U22485 ( .A1(n19529), .A2(n19775), .B1(n19538), .B2(n19774), .ZN(
        n19515) );
  NOR2_X1 U22486 ( .A1(n19507), .A2(n19723), .ZN(n19927) );
  OAI211_X1 U22487 ( .C1(n19538), .C2(n19509), .A(n19508), .B(n19731), .ZN(
        n19510) );
  INV_X1 U22488 ( .A(n19510), .ZN(n19511) );
  OAI21_X1 U22489 ( .B1(n19927), .B2(n19512), .A(n19511), .ZN(n19530) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19530), .B1(
        n19555), .B2(n19725), .ZN(n19514) );
  OAI211_X1 U22491 ( .C1(n19740), .C2(n19533), .A(n19515), .B(n19514), .ZN(
        P2_U3104) );
  AOI22_X1 U22492 ( .A1(n19529), .A2(n19789), .B1(n19538), .B2(n19788), .ZN(
        n19517) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19530), .B1(
        n19522), .B2(n19790), .ZN(n19516) );
  OAI211_X1 U22494 ( .C1(n19793), .C2(n19563), .A(n19517), .B(n19516), .ZN(
        P2_U3105) );
  AOI22_X1 U22495 ( .A1(n19529), .A2(n19795), .B1(n19538), .B2(n9852), .ZN(
        n19519) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19530), .B1(
        n19522), .B2(n19743), .ZN(n19518) );
  OAI211_X1 U22497 ( .C1(n19746), .C2(n19563), .A(n19519), .B(n19518), .ZN(
        P2_U3106) );
  AOI22_X1 U22498 ( .A1(n19529), .A2(n19801), .B1(n19538), .B2(n19800), .ZN(
        n19521) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19530), .B1(
        n19522), .B2(n19747), .ZN(n19520) );
  OAI211_X1 U22500 ( .C1(n19750), .C2(n19563), .A(n19521), .B(n19520), .ZN(
        P2_U3107) );
  AOI22_X1 U22501 ( .A1(n19529), .A2(n19807), .B1(n19538), .B2(n19806), .ZN(
        n19524) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19530), .B1(
        n19522), .B2(n19709), .ZN(n19523) );
  OAI211_X1 U22503 ( .C1(n19712), .C2(n19563), .A(n19524), .B(n19523), .ZN(
        P2_U3108) );
  AOI22_X1 U22504 ( .A1(n19529), .A2(n19813), .B1(n19538), .B2(n19812), .ZN(
        n19526) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19530), .B1(
        n19555), .B2(n19814), .ZN(n19525) );
  OAI211_X1 U22506 ( .C1(n19817), .C2(n19533), .A(n19526), .B(n19525), .ZN(
        P2_U3109) );
  AOI22_X1 U22507 ( .A1(n19529), .A2(n19819), .B1(n19538), .B2(n19818), .ZN(
        n19528) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19530), .B1(
        n19555), .B2(n19757), .ZN(n19527) );
  OAI211_X1 U22509 ( .C1(n19761), .C2(n19533), .A(n19528), .B(n19527), .ZN(
        P2_U3110) );
  AOI22_X1 U22510 ( .A1(n19529), .A2(n19828), .B1(n19538), .B2(n19827), .ZN(
        n19532) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19530), .B1(
        n19555), .B2(n19830), .ZN(n19531) );
  OAI211_X1 U22512 ( .C1(n19836), .C2(n19533), .A(n19532), .B(n19531), .ZN(
        P2_U3111) );
  NAND2_X1 U22513 ( .A1(n19940), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19634) );
  INV_X1 U22514 ( .A(n19634), .ZN(n19628) );
  NAND2_X1 U22515 ( .A1(n19628), .A2(n19949), .ZN(n19574) );
  NOR2_X1 U22516 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19574), .ZN(
        n19558) );
  AOI22_X1 U22517 ( .A1(n19784), .A2(n19555), .B1(n19558), .B2(n19774), .ZN(
        n19544) );
  OAI21_X1 U22518 ( .B1(n19555), .B2(n19588), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19535) );
  NAND2_X1 U22519 ( .A1(n19535), .A2(n19928), .ZN(n19542) );
  NOR2_X1 U22520 ( .A1(n19542), .A2(n19538), .ZN(n19536) );
  AOI211_X1 U22521 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n11934), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19536), .ZN(n19537) );
  OAI21_X1 U22522 ( .B1(n19558), .B2(n19537), .A(n19731), .ZN(n19560) );
  NOR2_X1 U22523 ( .A1(n19538), .A2(n19558), .ZN(n19541) );
  INV_X1 U22524 ( .A(n11934), .ZN(n19539) );
  OAI21_X1 U22525 ( .B1(n19539), .B2(n19558), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19540) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19560), .B1(
        n19775), .B2(n19559), .ZN(n19543) );
  OAI211_X1 U22527 ( .C1(n19787), .C2(n19596), .A(n19544), .B(n19543), .ZN(
        P2_U3112) );
  AOI22_X1 U22528 ( .A1(n19555), .A2(n19790), .B1(n19558), .B2(n19788), .ZN(
        n19546) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19560), .B1(
        n19559), .B2(n19789), .ZN(n19545) );
  OAI211_X1 U22530 ( .C1(n19793), .C2(n19596), .A(n19546), .B(n19545), .ZN(
        P2_U3113) );
  AOI22_X1 U22531 ( .A1(n19796), .A2(n19588), .B1(n19558), .B2(n9852), .ZN(
        n19548) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19560), .B1(
        n19559), .B2(n19795), .ZN(n19547) );
  OAI211_X1 U22533 ( .C1(n19799), .C2(n19563), .A(n19548), .B(n19547), .ZN(
        P2_U3114) );
  AOI22_X1 U22534 ( .A1(n19802), .A2(n19588), .B1(n19558), .B2(n19800), .ZN(
        n19550) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19560), .B1(
        n19559), .B2(n19801), .ZN(n19549) );
  OAI211_X1 U22536 ( .C1(n19805), .C2(n19563), .A(n19550), .B(n19549), .ZN(
        P2_U3115) );
  AOI22_X1 U22537 ( .A1(n19808), .A2(n19588), .B1(n19558), .B2(n19806), .ZN(
        n19552) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19560), .B1(
        n19559), .B2(n19807), .ZN(n19551) );
  OAI211_X1 U22539 ( .C1(n19811), .C2(n19563), .A(n19552), .B(n19551), .ZN(
        P2_U3116) );
  AOI22_X1 U22540 ( .A1(n19814), .A2(n19588), .B1(n19558), .B2(n19812), .ZN(
        n19554) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19560), .B1(
        n19559), .B2(n19813), .ZN(n19553) );
  OAI211_X1 U22542 ( .C1(n19817), .C2(n19563), .A(n19554), .B(n19553), .ZN(
        P2_U3117) );
  AOI22_X1 U22543 ( .A1(n19820), .A2(n19555), .B1(n19558), .B2(n19818), .ZN(
        n19557) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19560), .B1(
        n19559), .B2(n19819), .ZN(n19556) );
  OAI211_X1 U22545 ( .C1(n19825), .C2(n19596), .A(n19557), .B(n19556), .ZN(
        P2_U3118) );
  AOI22_X1 U22546 ( .A1(n19830), .A2(n19588), .B1(n19558), .B2(n19827), .ZN(
        n19562) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19560), .B1(
        n19559), .B2(n19828), .ZN(n19561) );
  OAI211_X1 U22548 ( .C1(n19836), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P2_U3119) );
  NOR2_X1 U22549 ( .A1(n19564), .A2(n19634), .ZN(n19601) );
  AOI22_X1 U22550 ( .A1(n19784), .A2(n19588), .B1(n19774), .B2(n19601), .ZN(
        n19577) );
  OR2_X1 U22551 ( .A1(n19565), .A2(n19661), .ZN(n19693) );
  OR2_X1 U22552 ( .A1(n19693), .A2(n19566), .ZN(n19567) );
  AND2_X1 U22553 ( .A1(n19567), .A2(n19928), .ZN(n19571) );
  INV_X1 U22554 ( .A(n19601), .ZN(n19568) );
  NAND2_X1 U22555 ( .A1(n11921), .A2(n19568), .ZN(n19572) );
  NOR2_X1 U22556 ( .A1(n19572), .A2(n19951), .ZN(n19569) );
  AOI21_X1 U22557 ( .B1(n19571), .B2(n19574), .A(n19569), .ZN(n19570) );
  OAI211_X1 U22558 ( .C1(n19601), .C2(n19509), .A(n19570), .B(n19731), .ZN(
        n19593) );
  INV_X1 U22559 ( .A(n19571), .ZN(n19575) );
  INV_X1 U22560 ( .A(n19572), .ZN(n19573) );
  OAI22_X1 U22561 ( .A1(n19575), .A2(n19574), .B1(n19573), .B2(n19951), .ZN(
        n19592) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19593), .B1(
        n19775), .B2(n19592), .ZN(n19576) );
  OAI211_X1 U22563 ( .C1(n19787), .C2(n19591), .A(n19577), .B(n19576), .ZN(
        P2_U3120) );
  AOI22_X1 U22564 ( .A1(n19790), .A2(n19588), .B1(n19601), .B2(n19788), .ZN(
        n19579) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19593), .B1(
        n19789), .B2(n19592), .ZN(n19578) );
  OAI211_X1 U22566 ( .C1(n19793), .C2(n19591), .A(n19579), .B(n19578), .ZN(
        P2_U3121) );
  AOI22_X1 U22567 ( .A1(n19743), .A2(n19588), .B1(n9852), .B2(n19601), .ZN(
        n19581) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19593), .B1(
        n19795), .B2(n19592), .ZN(n19580) );
  OAI211_X1 U22569 ( .C1(n19746), .C2(n19591), .A(n19581), .B(n19580), .ZN(
        P2_U3122) );
  AOI22_X1 U22570 ( .A1(n19802), .A2(n19622), .B1(n19800), .B2(n19601), .ZN(
        n19583) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19593), .B1(
        n19801), .B2(n19592), .ZN(n19582) );
  OAI211_X1 U22572 ( .C1(n19805), .C2(n19596), .A(n19583), .B(n19582), .ZN(
        P2_U3123) );
  AOI22_X1 U22573 ( .A1(n19709), .A2(n19588), .B1(n19806), .B2(n19601), .ZN(
        n19585) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19593), .B1(
        n19807), .B2(n19592), .ZN(n19584) );
  OAI211_X1 U22575 ( .C1(n19712), .C2(n19591), .A(n19585), .B(n19584), .ZN(
        P2_U3124) );
  AOI22_X1 U22576 ( .A1(n19814), .A2(n19622), .B1(n19812), .B2(n19601), .ZN(
        n19587) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19593), .B1(
        n19813), .B2(n19592), .ZN(n19586) );
  OAI211_X1 U22578 ( .C1(n19817), .C2(n19596), .A(n19587), .B(n19586), .ZN(
        P2_U3125) );
  AOI22_X1 U22579 ( .A1(n19820), .A2(n19588), .B1(n19601), .B2(n19818), .ZN(
        n19590) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19593), .B1(
        n19819), .B2(n19592), .ZN(n19589) );
  OAI211_X1 U22581 ( .C1(n19825), .C2(n19591), .A(n19590), .B(n19589), .ZN(
        P2_U3126) );
  AOI22_X1 U22582 ( .A1(n19830), .A2(n19622), .B1(n19827), .B2(n19601), .ZN(
        n19595) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19593), .B1(
        n19828), .B2(n19592), .ZN(n19594) );
  OAI211_X1 U22584 ( .C1(n19836), .C2(n19596), .A(n19595), .B(n19594), .ZN(
        P2_U3127) );
  INV_X1 U22585 ( .A(n19602), .ZN(n19598) );
  NOR2_X1 U22586 ( .A1(n19597), .A2(n19634), .ZN(n19620) );
  OAI21_X1 U22587 ( .B1(n19598), .B2(n19620), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19599) );
  OAI21_X1 U22588 ( .B1(n19634), .B2(n19600), .A(n19599), .ZN(n19621) );
  AOI22_X1 U22589 ( .A1(n19621), .A2(n19775), .B1(n19774), .B2(n19620), .ZN(
        n19607) );
  AOI221_X1 U22590 ( .B1(n19622), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19654), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19601), .ZN(n19603) );
  MUX2_X1 U22591 ( .A(n19603), .B(n19602), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19604) );
  NOR2_X1 U22592 ( .A1(n19604), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19605) );
  OAI21_X1 U22593 ( .B1(n19605), .B2(n19620), .A(n19731), .ZN(n19623) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19784), .ZN(n19606) );
  OAI211_X1 U22595 ( .C1(n19787), .C2(n19626), .A(n19607), .B(n19606), .ZN(
        P2_U3128) );
  AOI22_X1 U22596 ( .A1(n19621), .A2(n19789), .B1(n19788), .B2(n19620), .ZN(
        n19609) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19790), .ZN(n19608) );
  OAI211_X1 U22598 ( .C1(n19793), .C2(n19626), .A(n19609), .B(n19608), .ZN(
        P2_U3129) );
  AOI22_X1 U22599 ( .A1(n19621), .A2(n19795), .B1(n9852), .B2(n19620), .ZN(
        n19611) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19743), .ZN(n19610) );
  OAI211_X1 U22601 ( .C1(n19746), .C2(n19626), .A(n19611), .B(n19610), .ZN(
        P2_U3130) );
  AOI22_X1 U22602 ( .A1(n19621), .A2(n19801), .B1(n19800), .B2(n19620), .ZN(
        n19613) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19747), .ZN(n19612) );
  OAI211_X1 U22604 ( .C1(n19750), .C2(n19626), .A(n19613), .B(n19612), .ZN(
        P2_U3131) );
  AOI22_X1 U22605 ( .A1(n19621), .A2(n19807), .B1(n19806), .B2(n19620), .ZN(
        n19615) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19709), .ZN(n19614) );
  OAI211_X1 U22607 ( .C1(n19712), .C2(n19626), .A(n19615), .B(n19614), .ZN(
        P2_U3132) );
  AOI22_X1 U22608 ( .A1(n19621), .A2(n19813), .B1(n19812), .B2(n19620), .ZN(
        n19617) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19753), .ZN(n19616) );
  OAI211_X1 U22610 ( .C1(n19756), .C2(n19626), .A(n19617), .B(n19616), .ZN(
        P2_U3133) );
  AOI22_X1 U22611 ( .A1(n19621), .A2(n19819), .B1(n19818), .B2(n19620), .ZN(
        n19619) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19820), .ZN(n19618) );
  OAI211_X1 U22613 ( .C1(n19825), .C2(n19626), .A(n19619), .B(n19618), .ZN(
        P2_U3134) );
  AOI22_X1 U22614 ( .A1(n19621), .A2(n19828), .B1(n19827), .B2(n19620), .ZN(
        n19625) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19764), .ZN(n19624) );
  OAI211_X1 U22616 ( .C1(n19769), .C2(n19626), .A(n19625), .B(n19624), .ZN(
        P2_U3135) );
  INV_X1 U22617 ( .A(n19688), .ZN(n19627) );
  NAND2_X1 U22618 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19628), .ZN(
        n19632) );
  INV_X1 U22619 ( .A(n19633), .ZN(n19630) );
  NOR2_X1 U22620 ( .A1(n19629), .A2(n19634), .ZN(n19652) );
  OAI21_X1 U22621 ( .B1(n19630), .B2(n19652), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19631) );
  OAI21_X1 U22622 ( .B1(n19632), .B2(n19728), .A(n19631), .ZN(n19653) );
  AOI22_X1 U22623 ( .A1(n19653), .A2(n19775), .B1(n19774), .B2(n19652), .ZN(
        n19639) );
  AOI21_X1 U22624 ( .B1(n19633), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19637) );
  OAI22_X1 U22625 ( .A1(n19693), .A2(n19635), .B1(n19949), .B2(n19634), .ZN(
        n19636) );
  OAI211_X1 U22626 ( .C1(n19652), .C2(n19637), .A(n19636), .B(n19731), .ZN(
        n19655) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19784), .ZN(n19638) );
  OAI211_X1 U22628 ( .C1(n19787), .C2(n19686), .A(n19639), .B(n19638), .ZN(
        P2_U3136) );
  AOI22_X1 U22629 ( .A1(n19653), .A2(n19789), .B1(n19788), .B2(n19652), .ZN(
        n19641) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19790), .ZN(n19640) );
  OAI211_X1 U22631 ( .C1(n19793), .C2(n19686), .A(n19641), .B(n19640), .ZN(
        P2_U3137) );
  AOI22_X1 U22632 ( .A1(n19653), .A2(n19795), .B1(n9852), .B2(n19652), .ZN(
        n19643) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19743), .ZN(n19642) );
  OAI211_X1 U22634 ( .C1(n19746), .C2(n19686), .A(n19643), .B(n19642), .ZN(
        P2_U3138) );
  AOI22_X1 U22635 ( .A1(n19653), .A2(n19801), .B1(n19800), .B2(n19652), .ZN(
        n19645) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19747), .ZN(n19644) );
  OAI211_X1 U22637 ( .C1(n19750), .C2(n19686), .A(n19645), .B(n19644), .ZN(
        P2_U3139) );
  AOI22_X1 U22638 ( .A1(n19653), .A2(n19807), .B1(n19806), .B2(n19652), .ZN(
        n19647) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19709), .ZN(n19646) );
  OAI211_X1 U22640 ( .C1(n19712), .C2(n19686), .A(n19647), .B(n19646), .ZN(
        P2_U3140) );
  AOI22_X1 U22641 ( .A1(n19653), .A2(n19813), .B1(n19812), .B2(n19652), .ZN(
        n19649) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19753), .ZN(n19648) );
  OAI211_X1 U22643 ( .C1(n19756), .C2(n19686), .A(n19649), .B(n19648), .ZN(
        P2_U3141) );
  AOI22_X1 U22644 ( .A1(n19653), .A2(n19819), .B1(n19818), .B2(n19652), .ZN(
        n19651) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19820), .ZN(n19650) );
  OAI211_X1 U22646 ( .C1(n19825), .C2(n19686), .A(n19651), .B(n19650), .ZN(
        P2_U3142) );
  AOI22_X1 U22647 ( .A1(n19653), .A2(n19828), .B1(n19827), .B2(n19652), .ZN(
        n19657) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19655), .B1(
        n19654), .B2(n19764), .ZN(n19656) );
  OAI211_X1 U22649 ( .C1(n19769), .C2(n19686), .A(n19657), .B(n19656), .ZN(
        P2_U3143) );
  INV_X1 U22650 ( .A(n11917), .ZN(n19658) );
  NAND3_X1 U22651 ( .A1(n19949), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19690) );
  INV_X1 U22652 ( .A(n19690), .ZN(n19698) );
  NAND2_X1 U22653 ( .A1(n19958), .A2(n19698), .ZN(n19663) );
  INV_X1 U22654 ( .A(n19663), .ZN(n19681) );
  NOR3_X1 U22655 ( .A1(n19658), .A2(n19681), .A3(n19951), .ZN(n19662) );
  NOR2_X1 U22656 ( .A1(n19933), .A2(n19659), .ZN(n19666) );
  AOI21_X1 U22657 ( .B1(n19666), .B2(n19509), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19660) );
  AOI22_X1 U22658 ( .A1(n19682), .A2(n19775), .B1(n19774), .B2(n19681), .ZN(
        n19668) );
  NOR2_X2 U22659 ( .A1(n19724), .A2(n19687), .ZN(n19715) );
  INV_X1 U22660 ( .A(n19715), .ZN(n19722) );
  AOI21_X1 U22661 ( .B1(n19686), .B2(n19722), .A(n19661), .ZN(n19665) );
  AOI211_X1 U22662 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19663), .A(n19778), 
        .B(n19662), .ZN(n19664) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19683), .B1(
        n19715), .B2(n19725), .ZN(n19667) );
  OAI211_X1 U22664 ( .C1(n19740), .C2(n19686), .A(n19668), .B(n19667), .ZN(
        P2_U3144) );
  AOI22_X1 U22665 ( .A1(n19682), .A2(n19789), .B1(n19788), .B2(n19681), .ZN(
        n19670) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19683), .B1(
        n19715), .B2(n19701), .ZN(n19669) );
  OAI211_X1 U22667 ( .C1(n19704), .C2(n19686), .A(n19670), .B(n19669), .ZN(
        P2_U3145) );
  AOI22_X1 U22668 ( .A1(n19682), .A2(n19795), .B1(n9852), .B2(n19681), .ZN(
        n19672) );
  AOI22_X1 U22669 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19683), .B1(
        n19715), .B2(n19796), .ZN(n19671) );
  OAI211_X1 U22670 ( .C1(n19799), .C2(n19686), .A(n19672), .B(n19671), .ZN(
        P2_U3146) );
  AOI22_X1 U22671 ( .A1(n19682), .A2(n19801), .B1(n19800), .B2(n19681), .ZN(
        n19674) );
  AOI22_X1 U22672 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19683), .B1(
        n19715), .B2(n19802), .ZN(n19673) );
  OAI211_X1 U22673 ( .C1(n19805), .C2(n19686), .A(n19674), .B(n19673), .ZN(
        P2_U3147) );
  AOI22_X1 U22674 ( .A1(n19682), .A2(n19807), .B1(n19806), .B2(n19681), .ZN(
        n19676) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19683), .B1(
        n19715), .B2(n19808), .ZN(n19675) );
  OAI211_X1 U22676 ( .C1(n19811), .C2(n19686), .A(n19676), .B(n19675), .ZN(
        P2_U3148) );
  AOI22_X1 U22677 ( .A1(n19682), .A2(n19813), .B1(n19812), .B2(n19681), .ZN(
        n19678) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19683), .B1(
        n19715), .B2(n19814), .ZN(n19677) );
  OAI211_X1 U22679 ( .C1(n19817), .C2(n19686), .A(n19678), .B(n19677), .ZN(
        P2_U3149) );
  AOI22_X1 U22680 ( .A1(n19682), .A2(n19819), .B1(n19818), .B2(n19681), .ZN(
        n19680) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19683), .B1(
        n19715), .B2(n19757), .ZN(n19679) );
  OAI211_X1 U22682 ( .C1(n19761), .C2(n19686), .A(n19680), .B(n19679), .ZN(
        P2_U3150) );
  AOI22_X1 U22683 ( .A1(n19682), .A2(n19828), .B1(n19827), .B2(n19681), .ZN(
        n19685) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19683), .B1(
        n19715), .B2(n19830), .ZN(n19684) );
  OAI211_X1 U22685 ( .C1(n19836), .C2(n19686), .A(n19685), .B(n19684), .ZN(
        P2_U3151) );
  INV_X1 U22686 ( .A(n19689), .ZN(n19691) );
  NOR2_X1 U22687 ( .A1(n19958), .A2(n19690), .ZN(n19727) );
  NOR3_X1 U22688 ( .A1(n19691), .A2(n19727), .A3(n19951), .ZN(n19694) );
  AOI21_X1 U22689 ( .B1(n19509), .B2(n19698), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19692) );
  NOR2_X1 U22690 ( .A1(n19694), .A2(n19692), .ZN(n19718) );
  AOI22_X1 U22691 ( .A1(n19718), .A2(n19775), .B1(n19774), .B2(n19727), .ZN(
        n19700) );
  INV_X1 U22692 ( .A(n19693), .ZN(n19781) );
  INV_X1 U22693 ( .A(n19727), .ZN(n19695) );
  AOI211_X1 U22694 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19695), .A(n19778), 
        .B(n19694), .ZN(n19696) );
  OAI221_X1 U22695 ( .B1(n19698), .B2(n19697), .C1(n19698), .C2(n19781), .A(
        n19696), .ZN(n19719) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19719), .B1(
        n19715), .B2(n19784), .ZN(n19699) );
  OAI211_X1 U22697 ( .C1(n19787), .C2(n19760), .A(n19700), .B(n19699), .ZN(
        P2_U3152) );
  AOI22_X1 U22698 ( .A1(n19718), .A2(n19789), .B1(n19788), .B2(n19727), .ZN(
        n19703) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19719), .B1(
        n19763), .B2(n19701), .ZN(n19702) );
  OAI211_X1 U22700 ( .C1(n19704), .C2(n19722), .A(n19703), .B(n19702), .ZN(
        P2_U3153) );
  AOI22_X1 U22701 ( .A1(n19718), .A2(n19795), .B1(n9852), .B2(n19727), .ZN(
        n19706) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19719), .B1(
        n19715), .B2(n19743), .ZN(n19705) );
  OAI211_X1 U22703 ( .C1(n19746), .C2(n19760), .A(n19706), .B(n19705), .ZN(
        P2_U3154) );
  AOI22_X1 U22704 ( .A1(n19718), .A2(n19801), .B1(n19800), .B2(n19727), .ZN(
        n19708) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19719), .B1(
        n19715), .B2(n19747), .ZN(n19707) );
  OAI211_X1 U22706 ( .C1(n19750), .C2(n19760), .A(n19708), .B(n19707), .ZN(
        P2_U3155) );
  AOI22_X1 U22707 ( .A1(n19718), .A2(n19807), .B1(n19806), .B2(n19727), .ZN(
        n19711) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19719), .B1(
        n19715), .B2(n19709), .ZN(n19710) );
  OAI211_X1 U22709 ( .C1(n19712), .C2(n19760), .A(n19711), .B(n19710), .ZN(
        P2_U3156) );
  AOI22_X1 U22710 ( .A1(n19718), .A2(n19813), .B1(n19812), .B2(n19727), .ZN(
        n19714) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19719), .B1(
        n19763), .B2(n19814), .ZN(n19713) );
  OAI211_X1 U22712 ( .C1(n19817), .C2(n19722), .A(n19714), .B(n19713), .ZN(
        P2_U3157) );
  AOI22_X1 U22713 ( .A1(n19718), .A2(n19819), .B1(n19818), .B2(n19727), .ZN(
        n19717) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19719), .B1(
        n19715), .B2(n19820), .ZN(n19716) );
  OAI211_X1 U22715 ( .C1(n19825), .C2(n19760), .A(n19717), .B(n19716), .ZN(
        P2_U3158) );
  AOI22_X1 U22716 ( .A1(n19718), .A2(n19828), .B1(n19827), .B2(n19727), .ZN(
        n19721) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19719), .B1(
        n19763), .B2(n19830), .ZN(n19720) );
  OAI211_X1 U22718 ( .C1(n19836), .C2(n19722), .A(n19721), .B(n19720), .ZN(
        P2_U3159) );
  NOR3_X2 U22719 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19933), .A3(
        n19771), .ZN(n19762) );
  AOI22_X1 U22720 ( .A1(n19725), .A2(n19821), .B1(n19774), .B2(n19762), .ZN(
        n19739) );
  OAI21_X1 U22721 ( .B1(n19821), .B2(n19763), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19726) );
  NAND2_X1 U22722 ( .A1(n19726), .A2(n19928), .ZN(n19737) );
  NOR2_X1 U22723 ( .A1(n19762), .A2(n19727), .ZN(n19736) );
  INV_X1 U22724 ( .A(n19736), .ZN(n19732) );
  INV_X1 U22725 ( .A(n19762), .ZN(n19729) );
  OAI211_X1 U22726 ( .C1(n19733), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19729), 
        .B(n19728), .ZN(n19730) );
  OAI211_X1 U22727 ( .C1(n19737), .C2(n19732), .A(n19731), .B(n19730), .ZN(
        n19766) );
  INV_X1 U22728 ( .A(n19733), .ZN(n19734) );
  OAI21_X1 U22729 ( .B1(n19734), .B2(n19762), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19735) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19766), .B1(
        n19775), .B2(n19765), .ZN(n19738) );
  OAI211_X1 U22731 ( .C1(n19740), .C2(n19760), .A(n19739), .B(n19738), .ZN(
        P2_U3160) );
  AOI22_X1 U22732 ( .A1(n19790), .A2(n19763), .B1(n19788), .B2(n19762), .ZN(
        n19742) );
  AOI22_X1 U22733 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19766), .B1(
        n19789), .B2(n19765), .ZN(n19741) );
  OAI211_X1 U22734 ( .C1(n19793), .C2(n19835), .A(n19742), .B(n19741), .ZN(
        P2_U3161) );
  AOI22_X1 U22735 ( .A1(n19743), .A2(n19763), .B1(n9852), .B2(n19762), .ZN(
        n19745) );
  AOI22_X1 U22736 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19766), .B1(
        n19795), .B2(n19765), .ZN(n19744) );
  OAI211_X1 U22737 ( .C1(n19746), .C2(n19835), .A(n19745), .B(n19744), .ZN(
        P2_U3162) );
  AOI22_X1 U22738 ( .A1(n19747), .A2(n19763), .B1(n19800), .B2(n19762), .ZN(
        n19749) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19766), .B1(
        n19801), .B2(n19765), .ZN(n19748) );
  OAI211_X1 U22740 ( .C1(n19750), .C2(n19835), .A(n19749), .B(n19748), .ZN(
        P2_U3163) );
  AOI22_X1 U22741 ( .A1(n19808), .A2(n19821), .B1(n19806), .B2(n19762), .ZN(
        n19752) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19766), .B1(
        n19807), .B2(n19765), .ZN(n19751) );
  OAI211_X1 U22743 ( .C1(n19811), .C2(n19760), .A(n19752), .B(n19751), .ZN(
        P2_U3164) );
  AOI22_X1 U22744 ( .A1(n19753), .A2(n19763), .B1(n19812), .B2(n19762), .ZN(
        n19755) );
  AOI22_X1 U22745 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19766), .B1(
        n19813), .B2(n19765), .ZN(n19754) );
  OAI211_X1 U22746 ( .C1(n19756), .C2(n19835), .A(n19755), .B(n19754), .ZN(
        P2_U3165) );
  AOI22_X1 U22747 ( .A1(n19757), .A2(n19821), .B1(n19818), .B2(n19762), .ZN(
        n19759) );
  AOI22_X1 U22748 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19766), .B1(
        n19819), .B2(n19765), .ZN(n19758) );
  OAI211_X1 U22749 ( .C1(n19761), .C2(n19760), .A(n19759), .B(n19758), .ZN(
        P2_U3166) );
  AOI22_X1 U22750 ( .A1(n19764), .A2(n19763), .B1(n19827), .B2(n19762), .ZN(
        n19768) );
  AOI22_X1 U22751 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19766), .B1(
        n19828), .B2(n19765), .ZN(n19767) );
  OAI211_X1 U22752 ( .C1(n19769), .C2(n19835), .A(n19768), .B(n19767), .ZN(
        P2_U3167) );
  INV_X1 U22753 ( .A(n19826), .ZN(n19779) );
  NAND3_X1 U22754 ( .A1(n19770), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19779), 
        .ZN(n19776) );
  NOR2_X1 U22755 ( .A1(n19933), .A2(n19771), .ZN(n19783) );
  INV_X1 U22756 ( .A(n19783), .ZN(n19772) );
  OAI21_X1 U22757 ( .B1(n19772), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19951), 
        .ZN(n19773) );
  AND2_X1 U22758 ( .A1(n19776), .A2(n19773), .ZN(n19829) );
  AOI22_X1 U22759 ( .A1(n19829), .A2(n19775), .B1(n19774), .B2(n19826), .ZN(
        n19786) );
  INV_X1 U22760 ( .A(n19776), .ZN(n19777) );
  AOI211_X1 U22761 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19779), .A(n19778), 
        .B(n19777), .ZN(n19780) );
  OAI221_X1 U22762 ( .B1(n19783), .B2(n19782), .C1(n19783), .C2(n19781), .A(
        n19780), .ZN(n19832) );
  AOI22_X1 U22763 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19832), .B1(
        n19821), .B2(n19784), .ZN(n19785) );
  OAI211_X1 U22764 ( .C1(n19787), .C2(n19824), .A(n19786), .B(n19785), .ZN(
        P2_U3168) );
  AOI22_X1 U22765 ( .A1(n19829), .A2(n19789), .B1(n19788), .B2(n19826), .ZN(
        n19792) );
  AOI22_X1 U22766 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19832), .B1(
        n19821), .B2(n19790), .ZN(n19791) );
  OAI211_X1 U22767 ( .C1(n19793), .C2(n19824), .A(n19792), .B(n19791), .ZN(
        P2_U3169) );
  AOI22_X1 U22768 ( .A1(n19829), .A2(n19795), .B1(n9852), .B2(n19826), .ZN(
        n19798) );
  AOI22_X1 U22769 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19832), .B1(
        n19831), .B2(n19796), .ZN(n19797) );
  OAI211_X1 U22770 ( .C1(n19799), .C2(n19835), .A(n19798), .B(n19797), .ZN(
        P2_U3170) );
  AOI22_X1 U22771 ( .A1(n19829), .A2(n19801), .B1(n19800), .B2(n19826), .ZN(
        n19804) );
  AOI22_X1 U22772 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19832), .B1(
        n19831), .B2(n19802), .ZN(n19803) );
  OAI211_X1 U22773 ( .C1(n19805), .C2(n19835), .A(n19804), .B(n19803), .ZN(
        P2_U3171) );
  AOI22_X1 U22774 ( .A1(n19829), .A2(n19807), .B1(n19806), .B2(n19826), .ZN(
        n19810) );
  AOI22_X1 U22775 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19832), .B1(
        n19831), .B2(n19808), .ZN(n19809) );
  OAI211_X1 U22776 ( .C1(n19811), .C2(n19835), .A(n19810), .B(n19809), .ZN(
        P2_U3172) );
  AOI22_X1 U22777 ( .A1(n19829), .A2(n19813), .B1(n19812), .B2(n19826), .ZN(
        n19816) );
  AOI22_X1 U22778 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19832), .B1(
        n19831), .B2(n19814), .ZN(n19815) );
  OAI211_X1 U22779 ( .C1(n19817), .C2(n19835), .A(n19816), .B(n19815), .ZN(
        P2_U3173) );
  AOI22_X1 U22780 ( .A1(n19829), .A2(n19819), .B1(n19818), .B2(n19826), .ZN(
        n19823) );
  AOI22_X1 U22781 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19832), .B1(
        n19821), .B2(n19820), .ZN(n19822) );
  OAI211_X1 U22782 ( .C1(n19825), .C2(n19824), .A(n19823), .B(n19822), .ZN(
        P2_U3174) );
  AOI22_X1 U22783 ( .A1(n19829), .A2(n19828), .B1(n19827), .B2(n19826), .ZN(
        n19834) );
  AOI22_X1 U22784 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19832), .B1(
        n19831), .B2(n19830), .ZN(n19833) );
  OAI211_X1 U22785 ( .C1(n19836), .C2(n19835), .A(n19834), .B(n19833), .ZN(
        P2_U3175) );
  NOR4_X1 U22786 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n19857), .A4(n21158), .ZN(n19837) );
  NOR2_X1 U22787 ( .A1(n19838), .A2(n19837), .ZN(n19842) );
  OAI211_X1 U22788 ( .C1(n19843), .C2(n19839), .A(n19857), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19840) );
  OAI211_X1 U22789 ( .C1(n19843), .C2(n19842), .A(n19841), .B(n19840), .ZN(
        P2_U3177) );
  AND2_X1 U22790 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19844), .ZN(
        P2_U3179) );
  AND2_X1 U22791 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19844), .ZN(
        P2_U3180) );
  AND2_X1 U22792 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19844), .ZN(
        P2_U3181) );
  AND2_X1 U22793 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19844), .ZN(
        P2_U3182) );
  AND2_X1 U22794 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19844), .ZN(
        P2_U3183) );
  AND2_X1 U22795 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19844), .ZN(
        P2_U3184) );
  AND2_X1 U22796 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19844), .ZN(
        P2_U3185) );
  AND2_X1 U22797 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19844), .ZN(
        P2_U3186) );
  AND2_X1 U22798 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19844), .ZN(
        P2_U3187) );
  AND2_X1 U22799 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19844), .ZN(
        P2_U3188) );
  AND2_X1 U22800 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19844), .ZN(
        P2_U3189) );
  AND2_X1 U22801 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19844), .ZN(
        P2_U3190) );
  AND2_X1 U22802 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19844), .ZN(
        P2_U3191) );
  AND2_X1 U22803 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19844), .ZN(
        P2_U3192) );
  AND2_X1 U22804 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19844), .ZN(
        P2_U3193) );
  AND2_X1 U22805 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19844), .ZN(
        P2_U3194) );
  AND2_X1 U22806 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19844), .ZN(
        P2_U3195) );
  AND2_X1 U22807 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19844), .ZN(
        P2_U3196) );
  AND2_X1 U22808 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19844), .ZN(
        P2_U3197) );
  AND2_X1 U22809 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19844), .ZN(
        P2_U3198) );
  AND2_X1 U22810 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19844), .ZN(
        P2_U3199) );
  AND2_X1 U22811 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19844), .ZN(
        P2_U3200) );
  AND2_X1 U22812 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19844), .ZN(P2_U3201) );
  AND2_X1 U22813 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19844), .ZN(P2_U3202) );
  AND2_X1 U22814 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19844), .ZN(P2_U3203) );
  AND2_X1 U22815 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19844), .ZN(P2_U3204) );
  AND2_X1 U22816 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19844), .ZN(P2_U3205) );
  AND2_X1 U22817 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19844), .ZN(P2_U3206) );
  AND2_X1 U22818 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19844), .ZN(P2_U3207) );
  AND2_X1 U22819 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19844), .ZN(P2_U3208) );
  NOR2_X1 U22820 ( .A1(n20759), .A2(n19851), .ZN(n19865) );
  INV_X1 U22821 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19849) );
  NOR2_X1 U22822 ( .A1(n19845), .A2(n19849), .ZN(n19846) );
  NAND2_X1 U22823 ( .A1(n19857), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19860) );
  AOI21_X1 U22824 ( .B1(n19846), .B2(n19860), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19848) );
  AOI211_X1 U22825 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n19855), .A(
        n19859), .B(n19969), .ZN(n19847) );
  OR3_X1 U22826 ( .A1(n19865), .A2(n19848), .A3(n19847), .ZN(P2_U3209) );
  AOI21_X1 U22827 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19855), .A(n19866), 
        .ZN(n19856) );
  NOR2_X1 U22828 ( .A1(n19849), .A2(n19856), .ZN(n19852) );
  AOI21_X1 U22829 ( .B1(n19852), .B2(n19851), .A(n19850), .ZN(n19853) );
  OAI211_X1 U22830 ( .C1(n19855), .C2(n19854), .A(n19853), .B(n19860), .ZN(
        P2_U3210) );
  AOI21_X1 U22831 ( .B1(n19858), .B2(n19857), .A(n19856), .ZN(n19864) );
  INV_X1 U22832 ( .A(n19859), .ZN(n19861) );
  OAI22_X1 U22833 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19861), .B1(NA), 
        .B2(n19860), .ZN(n19862) );
  OAI211_X1 U22834 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19862), .ZN(n19863) );
  OAI21_X1 U22835 ( .B1(n19865), .B2(n19864), .A(n19863), .ZN(P2_U3211) );
  INV_X1 U22836 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19870) );
  NAND2_X2 U22837 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19969), .ZN(n19911) );
  OAI222_X1 U22838 ( .A1(n19915), .A2(n19870), .B1(n19868), .B2(n19969), .C1(
        n19867), .C2(n19911), .ZN(P2_U3212) );
  OAI222_X1 U22839 ( .A1(n19911), .A2(n19870), .B1(n19869), .B2(n19969), .C1(
        n19872), .C2(n19915), .ZN(P2_U3213) );
  OAI222_X1 U22840 ( .A1(n19911), .A2(n19872), .B1(n19871), .B2(n19969), .C1(
        n12321), .C2(n19915), .ZN(P2_U3214) );
  OAI222_X1 U22841 ( .A1(n19915), .A2(n12325), .B1(n19873), .B2(n19969), .C1(
        n12321), .C2(n19911), .ZN(P2_U3215) );
  OAI222_X1 U22842 ( .A1(n19915), .A2(n12329), .B1(n19874), .B2(n19969), .C1(
        n12325), .C2(n19911), .ZN(P2_U3216) );
  INV_X1 U22843 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19876) );
  OAI222_X1 U22844 ( .A1(n19915), .A2(n19876), .B1(n19875), .B2(n19969), .C1(
        n12329), .C2(n19911), .ZN(P2_U3217) );
  OAI222_X1 U22845 ( .A1(n19915), .A2(n12345), .B1(n19877), .B2(n19969), .C1(
        n19876), .C2(n19911), .ZN(P2_U3218) );
  OAI222_X1 U22846 ( .A1(n19915), .A2(n19878), .B1(n21144), .B2(n19969), .C1(
        n12345), .C2(n19911), .ZN(P2_U3219) );
  OAI222_X1 U22847 ( .A1(n19915), .A2(n19880), .B1(n19879), .B2(n19969), .C1(
        n19878), .C2(n19911), .ZN(P2_U3220) );
  INV_X1 U22848 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19882) );
  OAI222_X1 U22849 ( .A1(n19915), .A2(n19882), .B1(n19881), .B2(n19969), .C1(
        n19880), .C2(n19911), .ZN(P2_U3221) );
  OAI222_X1 U22850 ( .A1(n19915), .A2(n19884), .B1(n19883), .B2(n19969), .C1(
        n19882), .C2(n19911), .ZN(P2_U3222) );
  OAI222_X1 U22851 ( .A1(n19915), .A2(n19886), .B1(n19885), .B2(n19969), .C1(
        n19884), .C2(n19911), .ZN(P2_U3223) );
  OAI222_X1 U22852 ( .A1(n19915), .A2(n12408), .B1(n19887), .B2(n19969), .C1(
        n19886), .C2(n19911), .ZN(P2_U3224) );
  OAI222_X1 U22853 ( .A1(n19915), .A2(n19888), .B1(n21005), .B2(n19969), .C1(
        n12408), .C2(n19911), .ZN(P2_U3225) );
  OAI222_X1 U22854 ( .A1(n19915), .A2(n19890), .B1(n19889), .B2(n19969), .C1(
        n19888), .C2(n19911), .ZN(P2_U3226) );
  OAI222_X1 U22855 ( .A1(n19915), .A2(n12432), .B1(n19891), .B2(n19969), .C1(
        n19890), .C2(n19911), .ZN(P2_U3227) );
  OAI222_X1 U22856 ( .A1(n19915), .A2(n19893), .B1(n19892), .B2(n19969), .C1(
        n12432), .C2(n19911), .ZN(P2_U3228) );
  OAI222_X1 U22857 ( .A1(n19915), .A2(n15005), .B1(n19894), .B2(n19969), .C1(
        n19893), .C2(n19911), .ZN(P2_U3229) );
  OAI222_X1 U22858 ( .A1(n19915), .A2(n19896), .B1(n19895), .B2(n19969), .C1(
        n15005), .C2(n19911), .ZN(P2_U3230) );
  OAI222_X1 U22859 ( .A1(n19915), .A2(n12438), .B1(n19897), .B2(n19969), .C1(
        n19896), .C2(n19911), .ZN(P2_U3231) );
  OAI222_X1 U22860 ( .A1(n19915), .A2(n20948), .B1(n19898), .B2(n19969), .C1(
        n12438), .C2(n19911), .ZN(P2_U3232) );
  OAI222_X1 U22861 ( .A1(n19915), .A2(n13979), .B1(n19899), .B2(n19969), .C1(
        n20948), .C2(n19911), .ZN(P2_U3233) );
  OAI222_X1 U22862 ( .A1(n19915), .A2(n19901), .B1(n19900), .B2(n19969), .C1(
        n13979), .C2(n19911), .ZN(P2_U3234) );
  INV_X1 U22863 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19903) );
  OAI222_X1 U22864 ( .A1(n19915), .A2(n19903), .B1(n19902), .B2(n19969), .C1(
        n19901), .C2(n19911), .ZN(P2_U3235) );
  INV_X1 U22865 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20942) );
  OAI222_X1 U22866 ( .A1(n19915), .A2(n20942), .B1(n19904), .B2(n19969), .C1(
        n19903), .C2(n19911), .ZN(P2_U3236) );
  OAI222_X1 U22867 ( .A1(n19915), .A2(n12449), .B1(n19905), .B2(n19969), .C1(
        n20942), .C2(n19911), .ZN(P2_U3237) );
  OAI222_X1 U22868 ( .A1(n19911), .A2(n12449), .B1(n19906), .B2(n19969), .C1(
        n19907), .C2(n19915), .ZN(P2_U3238) );
  INV_X1 U22869 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19909) );
  OAI222_X1 U22870 ( .A1(n19915), .A2(n19909), .B1(n19908), .B2(n19969), .C1(
        n19907), .C2(n19911), .ZN(P2_U3239) );
  INV_X1 U22871 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19912) );
  OAI222_X1 U22872 ( .A1(n19915), .A2(n19912), .B1(n19910), .B2(n19969), .C1(
        n19909), .C2(n19911), .ZN(P2_U3240) );
  OAI222_X1 U22873 ( .A1(n19915), .A2(n19914), .B1(n19913), .B2(n19969), .C1(
        n19912), .C2(n19911), .ZN(P2_U3241) );
  OAI22_X1 U22874 ( .A1(n19970), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19969), .ZN(n19916) );
  INV_X1 U22875 ( .A(n19916), .ZN(P2_U3585) );
  OAI22_X1 U22876 ( .A1(n19970), .A2(P2_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P2_BE_N_REG_2__SCAN_IN), .B2(n19969), .ZN(n19917) );
  INV_X1 U22877 ( .A(n19917), .ZN(P2_U3586) );
  OAI22_X1 U22878 ( .A1(n19970), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19969), .ZN(n19918) );
  INV_X1 U22879 ( .A(n19918), .ZN(P2_U3587) );
  MUX2_X1 U22880 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .B(P2_BE_N_REG_0__SCAN_IN), .S(n19970), .Z(P2_U3588) );
  OAI21_X1 U22881 ( .B1(n19922), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19920), 
        .ZN(n19919) );
  INV_X1 U22882 ( .A(n19919), .ZN(P2_U3591) );
  OAI21_X1 U22883 ( .B1(n19922), .B2(n19921), .A(n19920), .ZN(P2_U3592) );
  AND2_X1 U22884 ( .A1(n19928), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19944) );
  NAND2_X1 U22885 ( .A1(n19923), .A2(n19944), .ZN(n19934) );
  NAND3_X1 U22886 ( .A1(n19925), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19924), 
        .ZN(n19926) );
  NAND2_X1 U22887 ( .A1(n19926), .A2(n19941), .ZN(n19935) );
  NAND2_X1 U22888 ( .A1(n19934), .A2(n19935), .ZN(n19931) );
  AOI222_X1 U22889 ( .A1(n19931), .A2(n19930), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19929), .C1(n19928), .C2(n19927), .ZN(n19932) );
  AOI22_X1 U22890 ( .A1(n19956), .A2(n19933), .B1(n19932), .B2(n19957), .ZN(
        P2_U3602) );
  OAI21_X1 U22891 ( .B1(n19936), .B2(n19935), .A(n19934), .ZN(n19937) );
  AOI21_X1 U22892 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19938), .A(n19937), 
        .ZN(n19939) );
  AOI22_X1 U22893 ( .A1(n19956), .A2(n19940), .B1(n19939), .B2(n19957), .ZN(
        P2_U3603) );
  INV_X1 U22894 ( .A(n19941), .ZN(n19952) );
  NOR2_X1 U22895 ( .A1(n19952), .A2(n19942), .ZN(n19945) );
  MUX2_X1 U22896 ( .A(n19945), .B(n19944), .S(n19943), .Z(n19946) );
  AOI21_X1 U22897 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19947), .A(n19946), 
        .ZN(n19948) );
  AOI22_X1 U22898 ( .A1(n19956), .A2(n19949), .B1(n19948), .B2(n19957), .ZN(
        P2_U3604) );
  OAI22_X1 U22899 ( .A1(n19953), .A2(n19952), .B1(n19951), .B2(n19950), .ZN(
        n19954) );
  AOI21_X1 U22900 ( .B1(n19958), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19954), 
        .ZN(n19955) );
  OAI22_X1 U22901 ( .A1(n19958), .A2(n19957), .B1(n19956), .B2(n19955), .ZN(
        P2_U3605) );
  INV_X1 U22902 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19959) );
  AOI22_X1 U22903 ( .A1(n19969), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19959), 
        .B2(n19970), .ZN(P2_U3608) );
  INV_X1 U22904 ( .A(n19960), .ZN(n19966) );
  AOI22_X1 U22905 ( .A1(n19964), .A2(n19963), .B1(n19962), .B2(n19961), .ZN(
        n19965) );
  NAND2_X1 U22906 ( .A1(n19966), .A2(n19965), .ZN(n19968) );
  MUX2_X1 U22907 ( .A(P2_MORE_REG_SCAN_IN), .B(n19968), .S(n19967), .Z(
        P2_U3609) );
  OAI22_X1 U22908 ( .A1(n19970), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19969), .ZN(n19971) );
  INV_X1 U22909 ( .A(n19971), .ZN(P2_U3611) );
  AND2_X1 U22910 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20753), .ZN(n19974) );
  INV_X1 U22911 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19973) );
  NOR2_X2 U22912 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n19972), .ZN(n20845) );
  AOI21_X1 U22913 ( .B1(n19974), .B2(n19973), .A(n20845), .ZN(P1_U2802) );
  NAND2_X1 U22914 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n19975), .ZN(n19979) );
  OAI21_X1 U22915 ( .B1(n19977), .B2(n19976), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19978) );
  OAI21_X1 U22916 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19979), .A(n19978), 
        .ZN(P1_U2803) );
  NOR2_X1 U22917 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20750) );
  OAI21_X1 U22918 ( .B1(n20750), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20799), .ZN(
        n19980) );
  OAI21_X1 U22919 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20799), .A(n19980), 
        .ZN(P1_U2804) );
  AOI21_X1 U22920 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20753), .A(n20845), 
        .ZN(n20811) );
  OAI21_X1 U22921 ( .B1(BS16), .B2(n20750), .A(n20811), .ZN(n20809) );
  OAI21_X1 U22922 ( .B1(n20811), .B2(n20814), .A(n20809), .ZN(P1_U2805) );
  OAI21_X1 U22923 ( .B1(n19983), .B2(n19982), .A(n19981), .ZN(P1_U2806) );
  NOR4_X1 U22924 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_18__SCAN_IN), .A3(P1_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19987) );
  NOR4_X1 U22925 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n19986) );
  NOR4_X1 U22926 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19985) );
  NOR4_X1 U22927 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_23__SCAN_IN), .A3(P1_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_25__SCAN_IN), .ZN(n19984) );
  NAND4_X1 U22928 ( .A1(n19987), .A2(n19986), .A3(n19985), .A4(n19984), .ZN(
        n19993) );
  NOR4_X1 U22929 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_29__SCAN_IN), .ZN(n19991) );
  AOI211_X1 U22930 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_3__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19990) );
  NOR4_X1 U22931 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19989) );
  NOR4_X1 U22932 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19988) );
  NAND4_X1 U22933 ( .A1(n19991), .A2(n19990), .A3(n19989), .A4(n19988), .ZN(
        n19992) );
  NOR2_X1 U22934 ( .A1(n19993), .A2(n19992), .ZN(n20843) );
  INV_X1 U22935 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19995) );
  NOR3_X1 U22936 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19996) );
  OAI21_X1 U22937 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19996), .A(n20843), .ZN(
        n19994) );
  OAI21_X1 U22938 ( .B1(n20843), .B2(n19995), .A(n19994), .ZN(P1_U2807) );
  INV_X1 U22939 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20810) );
  AOI21_X1 U22940 ( .B1(n20836), .B2(n20810), .A(n19996), .ZN(n19998) );
  INV_X1 U22941 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19997) );
  INV_X1 U22942 ( .A(n20843), .ZN(n20838) );
  AOI22_X1 U22943 ( .A1(n20843), .A2(n19998), .B1(n19997), .B2(n20838), .ZN(
        P1_U2808) );
  AOI22_X1 U22944 ( .A1(n19999), .A2(n20027), .B1(n20046), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n20009) );
  NAND2_X1 U22945 ( .A1(n20019), .A2(n20000), .ZN(n20002) );
  OAI22_X1 U22946 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20002), .B1(n20001), 
        .B2(n20044), .ZN(n20003) );
  AOI211_X1 U22947 ( .C1(n20040), .C2(n20004), .A(n20135), .B(n20003), .ZN(
        n20008) );
  AOI22_X1 U22948 ( .A1(n20006), .A2(n20031), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20005), .ZN(n20007) );
  NAND3_X1 U22949 ( .A1(n20009), .A2(n20008), .A3(n20007), .ZN(P1_U2831) );
  OAI22_X1 U22950 ( .A1(n20060), .A2(n20011), .B1(n20054), .B2(n20010), .ZN(
        n20015) );
  INV_X1 U22951 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20012) );
  NAND4_X1 U22952 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20038), .A4(n20012), .ZN(n20013) );
  OAI211_X1 U22953 ( .C1(n20044), .C2(n20883), .A(n20042), .B(n20013), .ZN(
        n20014) );
  AOI211_X1 U22954 ( .C1(n20027), .C2(n20016), .A(n20015), .B(n20014), .ZN(
        n20024) );
  AND2_X1 U22955 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20020) );
  AOI21_X1 U22956 ( .B1(n20019), .B2(n20018), .A(n20017), .ZN(n20071) );
  OAI21_X1 U22957 ( .B1(n20021), .B2(n20020), .A(n20071), .ZN(n20030) );
  AOI22_X1 U22958 ( .A1(n20022), .A2(n20031), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20030), .ZN(n20023) );
  NAND2_X1 U22959 ( .A1(n20024), .A2(n20023), .ZN(P1_U2833) );
  INV_X1 U22960 ( .A(n20025), .ZN(n20028) );
  AOI22_X1 U22961 ( .A1(n20028), .A2(n20040), .B1(n20027), .B2(n20026), .ZN(
        n20036) );
  NOR2_X1 U22962 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20053), .ZN(n20029) );
  AOI22_X1 U22963 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20059), .B1(
        n20038), .B2(n20029), .ZN(n20035) );
  AOI21_X1 U22964 ( .B1(n20046), .B2(P1_EBX_REG_6__SCAN_IN), .A(n20135), .ZN(
        n20034) );
  AOI22_X1 U22965 ( .A1(n20032), .A2(n20031), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20030), .ZN(n20033) );
  NAND4_X1 U22966 ( .A1(n20036), .A2(n20035), .A3(n20034), .A4(n20033), .ZN(
        P1_U2834) );
  INV_X1 U22967 ( .A(n20037), .ZN(n20049) );
  NAND2_X1 U22968 ( .A1(n20038), .A2(n20053), .ZN(n20048) );
  NAND2_X1 U22969 ( .A1(n20040), .A2(n20039), .ZN(n20041) );
  OAI211_X1 U22970 ( .C1(n20044), .C2(n20043), .A(n20042), .B(n20041), .ZN(
        n20045) );
  AOI21_X1 U22971 ( .B1(n20046), .B2(P1_EBX_REG_5__SCAN_IN), .A(n20045), .ZN(
        n20047) );
  OAI211_X1 U22972 ( .C1(n20049), .C2(n20062), .A(n20048), .B(n20047), .ZN(
        n20050) );
  AOI21_X1 U22973 ( .B1(n20051), .B2(n20067), .A(n20050), .ZN(n20052) );
  OAI21_X1 U22974 ( .B1(n20071), .B2(n20053), .A(n20052), .ZN(P1_U2835) );
  OAI22_X1 U22975 ( .A1(n20057), .A2(n20056), .B1(n20055), .B2(n20054), .ZN(
        n20058) );
  AOI211_X1 U22976 ( .C1(n20059), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20135), .B(n20058), .ZN(n20070) );
  OAI22_X1 U22977 ( .A1(n20062), .A2(n20061), .B1(n20060), .B2(n11301), .ZN(
        n20066) );
  NAND2_X1 U22978 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20064) );
  NOR3_X1 U22979 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20064), .A3(n20063), .ZN(
        n20065) );
  AOI211_X1 U22980 ( .C1(n20068), .C2(n20067), .A(n20066), .B(n20065), .ZN(
        n20069) );
  OAI211_X1 U22981 ( .C1(n20071), .C2(n20765), .A(n20070), .B(n20069), .ZN(
        P1_U2836) );
  AOI22_X1 U22982 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20073) );
  OAI21_X1 U22983 ( .B1(n13631), .B2(n20095), .A(n20073), .ZN(P1_U2921) );
  AOI22_X1 U22984 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20074) );
  OAI21_X1 U22985 ( .B1(n20908), .B2(n20095), .A(n20074), .ZN(P1_U2922) );
  INV_X1 U22986 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20076) );
  AOI22_X1 U22987 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20075) );
  OAI21_X1 U22988 ( .B1(n20076), .B2(n20095), .A(n20075), .ZN(P1_U2923) );
  INV_X1 U22989 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20078) );
  AOI22_X1 U22990 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20077) );
  OAI21_X1 U22991 ( .B1(n20078), .B2(n20095), .A(n20077), .ZN(P1_U2924) );
  AOI22_X1 U22992 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20079) );
  OAI21_X1 U22993 ( .B1(n14351), .B2(n20095), .A(n20079), .ZN(P1_U2925) );
  AOI22_X1 U22994 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20080) );
  OAI21_X1 U22995 ( .B1(n13972), .B2(n20095), .A(n20080), .ZN(P1_U2926) );
  INV_X1 U22996 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20082) );
  AOI22_X1 U22997 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20081) );
  OAI21_X1 U22998 ( .B1(n20082), .B2(n20095), .A(n20081), .ZN(P1_U2927) );
  AOI22_X1 U22999 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20849), .B1(n15844), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20083) );
  OAI21_X1 U23000 ( .B1(n13887), .B2(n20095), .A(n20083), .ZN(P1_U2928) );
  AOI22_X1 U23001 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20084) );
  OAI21_X1 U23002 ( .B1(n13772), .B2(n20095), .A(n20084), .ZN(P1_U2929) );
  AOI22_X1 U23003 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20085) );
  OAI21_X1 U23004 ( .B1(n10690), .B2(n20095), .A(n20085), .ZN(P1_U2930) );
  AOI22_X1 U23005 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20086) );
  OAI21_X1 U23006 ( .B1(n20087), .B2(n20095), .A(n20086), .ZN(P1_U2931) );
  AOI22_X1 U23007 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20088) );
  OAI21_X1 U23008 ( .B1(n20089), .B2(n20095), .A(n20088), .ZN(P1_U2932) );
  AOI22_X1 U23009 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20090) );
  OAI21_X1 U23010 ( .B1(n10613), .B2(n20095), .A(n20090), .ZN(P1_U2933) );
  AOI22_X1 U23011 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20091) );
  OAI21_X1 U23012 ( .B1(n10554), .B2(n20095), .A(n20091), .ZN(P1_U2934) );
  AOI22_X1 U23013 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20092) );
  OAI21_X1 U23014 ( .B1(n10562), .B2(n20095), .A(n20092), .ZN(P1_U2935) );
  AOI22_X1 U23015 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20093), .B1(n15844), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20094) );
  OAI21_X1 U23016 ( .B1(n20096), .B2(n20095), .A(n20094), .ZN(P1_U2936) );
  AOI22_X1 U23017 ( .A1(n20119), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20118), .ZN(n20098) );
  NAND2_X1 U23018 ( .A1(n20110), .A2(n20097), .ZN(n20112) );
  NAND2_X1 U23019 ( .A1(n20098), .A2(n20112), .ZN(P1_U2945) );
  AOI22_X1 U23020 ( .A1(n20119), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20118), .ZN(n20100) );
  NAND2_X1 U23021 ( .A1(n20110), .A2(n20099), .ZN(n20114) );
  NAND2_X1 U23022 ( .A1(n20100), .A2(n20114), .ZN(P1_U2946) );
  AOI22_X1 U23023 ( .A1(n20119), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20118), .ZN(n20102) );
  NAND2_X1 U23024 ( .A1(n20110), .A2(n20101), .ZN(n20116) );
  NAND2_X1 U23025 ( .A1(n20102), .A2(n20116), .ZN(P1_U2947) );
  AOI22_X1 U23026 ( .A1(n20119), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20118), .ZN(n20104) );
  NAND2_X1 U23027 ( .A1(n20110), .A2(n20103), .ZN(n20120) );
  NAND2_X1 U23028 ( .A1(n20104), .A2(n20120), .ZN(P1_U2948) );
  AOI22_X1 U23029 ( .A1(n20119), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20118), .ZN(n20106) );
  NAND2_X1 U23030 ( .A1(n20110), .A2(n20105), .ZN(n20122) );
  NAND2_X1 U23031 ( .A1(n20106), .A2(n20122), .ZN(P1_U2949) );
  AOI22_X1 U23032 ( .A1(n20119), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20118), .ZN(n20108) );
  NAND2_X1 U23033 ( .A1(n20110), .A2(n20107), .ZN(n20124) );
  NAND2_X1 U23034 ( .A1(n20108), .A2(n20124), .ZN(P1_U2950) );
  AOI22_X1 U23035 ( .A1(n20119), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20118), .ZN(n20111) );
  NAND2_X1 U23036 ( .A1(n20110), .A2(n20109), .ZN(n20126) );
  NAND2_X1 U23037 ( .A1(n20111), .A2(n20126), .ZN(P1_U2951) );
  AOI22_X1 U23038 ( .A1(n20119), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20118), .ZN(n20113) );
  NAND2_X1 U23039 ( .A1(n20113), .A2(n20112), .ZN(P1_U2960) );
  AOI22_X1 U23040 ( .A1(n20119), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20118), .ZN(n20115) );
  NAND2_X1 U23041 ( .A1(n20115), .A2(n20114), .ZN(P1_U2961) );
  AOI22_X1 U23042 ( .A1(n20119), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20118), .ZN(n20117) );
  NAND2_X1 U23043 ( .A1(n20117), .A2(n20116), .ZN(P1_U2962) );
  AOI22_X1 U23044 ( .A1(n20119), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20118), .ZN(n20121) );
  NAND2_X1 U23045 ( .A1(n20121), .A2(n20120), .ZN(P1_U2963) );
  AOI22_X1 U23046 ( .A1(n20119), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20118), .ZN(n20123) );
  NAND2_X1 U23047 ( .A1(n20123), .A2(n20122), .ZN(P1_U2964) );
  AOI22_X1 U23048 ( .A1(n20119), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20118), .ZN(n20125) );
  NAND2_X1 U23049 ( .A1(n20125), .A2(n20124), .ZN(P1_U2965) );
  AOI22_X1 U23050 ( .A1(n20119), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20118), .ZN(n20127) );
  NAND2_X1 U23051 ( .A1(n20127), .A2(n20126), .ZN(P1_U2966) );
  INV_X1 U23052 ( .A(n20128), .ZN(n20130) );
  AOI21_X1 U23053 ( .B1(n20130), .B2(n9916), .A(n20129), .ZN(n20141) );
  OR2_X1 U23054 ( .A1(n20132), .A2(n20131), .ZN(n20133) );
  AOI22_X1 U23055 ( .A1(n20141), .A2(n20134), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20133), .ZN(n20136) );
  NAND2_X1 U23056 ( .A1(n20135), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20148) );
  OAI211_X1 U23057 ( .C1(n20138), .C2(n20137), .A(n20136), .B(n20148), .ZN(
        P1_U2999) );
  AOI22_X1 U23058 ( .A1(n20141), .A2(n20140), .B1(n9916), .B2(n20139), .ZN(
        n20149) );
  OAI21_X1 U23059 ( .B1(n20143), .B2(n20142), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20147) );
  NAND2_X1 U23060 ( .A1(n20145), .A2(n20144), .ZN(n20146) );
  NAND4_X1 U23061 ( .A1(n20149), .A2(n20148), .A3(n20147), .A4(n20146), .ZN(
        P1_U3031) );
  NOR2_X1 U23062 ( .A1(n20150), .A2(n20835), .ZN(P1_U3032) );
  NAND2_X1 U23063 ( .A1(n20433), .A2(n20487), .ZN(n20324) );
  NOR2_X1 U23064 ( .A1(n20164), .A2(n20260), .ZN(n20561) );
  NOR2_X1 U23065 ( .A1(n20328), .A2(n20561), .ZN(n20492) );
  INV_X1 U23066 ( .A(n20492), .ZN(n20261) );
  INV_X1 U23067 ( .A(n20830), .ZN(n20151) );
  NAND2_X1 U23068 ( .A1(n20606), .A2(n20151), .ZN(n20533) );
  OAI21_X1 U23069 ( .B1(n20253), .B2(n20738), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20152) );
  NAND2_X1 U23070 ( .A1(n20152), .A2(n20682), .ZN(n20167) );
  INV_X1 U23071 ( .A(n13446), .ZN(n20153) );
  OR2_X1 U23072 ( .A1(n20817), .A2(n20153), .ZN(n20258) );
  OR2_X1 U23073 ( .A1(n20258), .A2(n20647), .ZN(n20166) );
  INV_X1 U23074 ( .A(n20166), .ZN(n20154) );
  NOR3_X1 U23075 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20236) );
  INV_X1 U23076 ( .A(n20236), .ZN(n20233) );
  NOR2_X1 U23077 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20233), .ZN(
        n20226) );
  OAI22_X1 U23078 ( .A1(n20167), .A2(n20154), .B1(n20226), .B2(n20568), .ZN(
        n20155) );
  AOI211_X1 U23079 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20324), .A(n20261), 
        .B(n20155), .ZN(n20178) );
  INV_X1 U23080 ( .A(DATAI_24_), .ZN(n20159) );
  OAI22_X2 U23081 ( .A1(n20160), .A2(n20220), .B1(n20159), .B2(n20222), .ZN(
        n20691) );
  NOR2_X2 U23082 ( .A1(n20225), .A2(n20162), .ZN(n20686) );
  AOI22_X1 U23083 ( .A1(n20738), .A2(n20691), .B1(n20686), .B2(n20226), .ZN(
        n20171) );
  INV_X1 U23084 ( .A(n20164), .ZN(n20165) );
  NOR2_X1 U23085 ( .A1(n20165), .A2(n20260), .ZN(n20489) );
  INV_X1 U23086 ( .A(n20489), .ZN(n20435) );
  INV_X1 U23087 ( .A(DATAI_16_), .ZN(n20168) );
  OAI22_X2 U23088 ( .A1(n20169), .A2(n20220), .B1(n20168), .B2(n20222), .ZN(
        n20610) );
  AOI22_X1 U23089 ( .A1(n20685), .A2(n20228), .B1(n20253), .B2(n20610), .ZN(
        n20170) );
  OAI211_X1 U23090 ( .C1(n20178), .C2(n20172), .A(n20171), .B(n20170), .ZN(
        P1_U3033) );
  INV_X1 U23091 ( .A(DATAI_17_), .ZN(n20173) );
  OAI22_X1 U23092 ( .A1(n20174), .A2(n20220), .B1(n20173), .B2(n20222), .ZN(
        n20614) );
  INV_X1 U23093 ( .A(n20614), .ZN(n20700) );
  INV_X1 U23094 ( .A(DATAI_25_), .ZN(n20175) );
  OAI22_X2 U23095 ( .A1(n20176), .A2(n20220), .B1(n20175), .B2(n20222), .ZN(
        n20697) );
  NOR2_X2 U23096 ( .A1(n20225), .A2(n20177), .ZN(n20696) );
  AOI22_X1 U23097 ( .A1(n20738), .A2(n20697), .B1(n20696), .B2(n20226), .ZN(
        n20181) );
  INV_X1 U23098 ( .A(n20178), .ZN(n20229) );
  AOI22_X1 U23099 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20229), .B1(
        n20695), .B2(n20228), .ZN(n20180) );
  OAI211_X1 U23100 ( .C1(n20700), .C2(n20232), .A(n20181), .B(n20180), .ZN(
        P1_U3034) );
  INV_X1 U23101 ( .A(DATAI_18_), .ZN(n20183) );
  OAI22_X1 U23102 ( .A1(n20183), .A2(n20222), .B1(n20182), .B2(n20220), .ZN(
        n20618) );
  INV_X1 U23103 ( .A(n20618), .ZN(n20706) );
  INV_X1 U23104 ( .A(DATAI_26_), .ZN(n20184) );
  OAI22_X2 U23105 ( .A1(n14305), .A2(n20220), .B1(n20184), .B2(n20222), .ZN(
        n20703) );
  AOI22_X1 U23106 ( .A1(n20738), .A2(n20703), .B1(n20702), .B2(n20226), .ZN(
        n20187) );
  AOI22_X1 U23107 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20229), .B1(
        n20701), .B2(n20228), .ZN(n20186) );
  OAI211_X1 U23108 ( .C1(n20706), .C2(n20232), .A(n20187), .B(n20186), .ZN(
        P1_U3035) );
  INV_X1 U23109 ( .A(DATAI_19_), .ZN(n20188) );
  OAI22_X2 U23110 ( .A1(n20189), .A2(n20220), .B1(n20188), .B2(n20222), .ZN(
        n20709) );
  INV_X1 U23111 ( .A(n20709), .ZN(n20662) );
  INV_X1 U23112 ( .A(DATAI_27_), .ZN(n20190) );
  OAI22_X2 U23113 ( .A1(n20191), .A2(n20220), .B1(n20190), .B2(n20222), .ZN(
        n20659) );
  NOR2_X2 U23114 ( .A1(n20225), .A2(n20192), .ZN(n20708) );
  AOI22_X1 U23115 ( .A1(n20738), .A2(n20659), .B1(n20708), .B2(n20226), .ZN(
        n20195) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20229), .B1(
        n20707), .B2(n20228), .ZN(n20194) );
  OAI211_X1 U23117 ( .C1(n20662), .C2(n20232), .A(n20195), .B(n20194), .ZN(
        P1_U3036) );
  INV_X1 U23118 ( .A(DATAI_20_), .ZN(n20197) );
  OAI22_X1 U23119 ( .A1(n20197), .A2(n20222), .B1(n20196), .B2(n20220), .ZN(
        n20624) );
  INV_X1 U23120 ( .A(n20624), .ZN(n20718) );
  INV_X1 U23121 ( .A(DATAI_28_), .ZN(n20198) );
  OAI22_X2 U23122 ( .A1(n14292), .A2(n20220), .B1(n20198), .B2(n20222), .ZN(
        n20715) );
  NOR2_X2 U23123 ( .A1(n20225), .A2(n20199), .ZN(n20714) );
  AOI22_X1 U23124 ( .A1(n20738), .A2(n20715), .B1(n20714), .B2(n20226), .ZN(
        n20202) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20229), .B1(
        n20713), .B2(n20228), .ZN(n20201) );
  OAI211_X1 U23126 ( .C1(n20718), .C2(n20232), .A(n20202), .B(n20201), .ZN(
        P1_U3037) );
  INV_X1 U23127 ( .A(DATAI_21_), .ZN(n20204) );
  OAI22_X1 U23128 ( .A1(n20204), .A2(n20222), .B1(n20203), .B2(n20220), .ZN(
        n20628) );
  INV_X1 U23129 ( .A(n20628), .ZN(n20724) );
  INV_X1 U23130 ( .A(DATAI_29_), .ZN(n20205) );
  OAI22_X2 U23131 ( .A1(n20206), .A2(n20220), .B1(n20205), .B2(n20222), .ZN(
        n20721) );
  NOR2_X2 U23132 ( .A1(n20225), .A2(n20207), .ZN(n20720) );
  AOI22_X1 U23133 ( .A1(n20738), .A2(n20721), .B1(n20720), .B2(n20226), .ZN(
        n20210) );
  AOI22_X1 U23134 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20229), .B1(
        n20719), .B2(n20228), .ZN(n20209) );
  OAI211_X1 U23135 ( .C1(n20724), .C2(n20232), .A(n20210), .B(n20209), .ZN(
        P1_U3038) );
  INV_X1 U23136 ( .A(DATAI_22_), .ZN(n20211) );
  OAI22_X1 U23137 ( .A1(n20211), .A2(n20222), .B1(n21037), .B2(n20220), .ZN(
        n20632) );
  INV_X1 U23138 ( .A(n20632), .ZN(n20732) );
  INV_X1 U23139 ( .A(DATAI_30_), .ZN(n20212) );
  OAI22_X2 U23140 ( .A1(n20213), .A2(n20220), .B1(n20212), .B2(n20222), .ZN(
        n20727) );
  NOR2_X2 U23141 ( .A1(n20225), .A2(n20214), .ZN(n20726) );
  AOI22_X1 U23142 ( .A1(n20738), .A2(n20727), .B1(n20726), .B2(n20226), .ZN(
        n20217) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20229), .B1(
        n20725), .B2(n20228), .ZN(n20216) );
  OAI211_X1 U23144 ( .C1(n20732), .C2(n20232), .A(n20217), .B(n20216), .ZN(
        P1_U3039) );
  INV_X1 U23145 ( .A(DATAI_23_), .ZN(n20219) );
  OAI22_X2 U23146 ( .A1(n20219), .A2(n20222), .B1(n20218), .B2(n20220), .ZN(
        n20737) );
  INV_X1 U23147 ( .A(DATAI_31_), .ZN(n20223) );
  OAI22_X2 U23148 ( .A1(n20223), .A2(n20222), .B1(n20221), .B2(n20220), .ZN(
        n20671) );
  NOR2_X2 U23149 ( .A1(n20225), .A2(n20224), .ZN(n20736) );
  AOI22_X1 U23150 ( .A1(n20738), .A2(n20671), .B1(n20736), .B2(n20226), .ZN(
        n20231) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20229), .B1(
        n20734), .B2(n20228), .ZN(n20230) );
  OAI211_X1 U23152 ( .C1(n20676), .C2(n20232), .A(n20231), .B(n20230), .ZN(
        P1_U3040) );
  INV_X1 U23153 ( .A(n20610), .ZN(n20694) );
  NOR2_X1 U23154 ( .A1(n20834), .A2(n20233), .ZN(n20252) );
  INV_X1 U23155 ( .A(n20258), .ZN(n20290) );
  INV_X1 U23156 ( .A(n20599), .ZN(n20461) );
  AOI21_X1 U23157 ( .B1(n20290), .B2(n20461), .A(n20252), .ZN(n20234) );
  OAI22_X1 U23158 ( .A1(n20234), .A2(n20829), .B1(n20233), .B2(n20260), .ZN(
        n20251) );
  AOI22_X1 U23159 ( .A1(n20686), .A2(n20252), .B1(n20251), .B2(n20685), .ZN(
        n20238) );
  OAI211_X1 U23160 ( .C1(n20294), .C2(n20814), .A(n20682), .B(n20234), .ZN(
        n20235) );
  OAI211_X1 U23161 ( .C1(n20813), .C2(n20236), .A(n20689), .B(n20235), .ZN(
        n20254) );
  AOI22_X1 U23162 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20691), .ZN(n20237) );
  OAI211_X1 U23163 ( .C1(n20694), .C2(n20279), .A(n20238), .B(n20237), .ZN(
        P1_U3041) );
  AOI22_X1 U23164 ( .A1(n20696), .A2(n20252), .B1(n20251), .B2(n20695), .ZN(
        n20240) );
  AOI22_X1 U23165 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20697), .ZN(n20239) );
  OAI211_X1 U23166 ( .C1(n20700), .C2(n20279), .A(n20240), .B(n20239), .ZN(
        P1_U3042) );
  AOI22_X1 U23167 ( .A1(n20702), .A2(n20252), .B1(n20251), .B2(n20701), .ZN(
        n20242) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20703), .ZN(n20241) );
  OAI211_X1 U23169 ( .C1(n20706), .C2(n20279), .A(n20242), .B(n20241), .ZN(
        P1_U3043) );
  AOI22_X1 U23170 ( .A1(n20708), .A2(n20252), .B1(n20251), .B2(n20707), .ZN(
        n20244) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20659), .ZN(n20243) );
  OAI211_X1 U23172 ( .C1(n20662), .C2(n20279), .A(n20244), .B(n20243), .ZN(
        P1_U3044) );
  AOI22_X1 U23173 ( .A1(n20714), .A2(n20252), .B1(n20251), .B2(n20713), .ZN(
        n20246) );
  AOI22_X1 U23174 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20715), .ZN(n20245) );
  OAI211_X1 U23175 ( .C1(n20718), .C2(n20279), .A(n20246), .B(n20245), .ZN(
        P1_U3045) );
  AOI22_X1 U23176 ( .A1(n20720), .A2(n20252), .B1(n20251), .B2(n20719), .ZN(
        n20248) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20721), .ZN(n20247) );
  OAI211_X1 U23178 ( .C1(n20724), .C2(n20279), .A(n20248), .B(n20247), .ZN(
        P1_U3046) );
  AOI22_X1 U23179 ( .A1(n20726), .A2(n20252), .B1(n20251), .B2(n20725), .ZN(
        n20250) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20727), .ZN(n20249) );
  OAI211_X1 U23181 ( .C1(n20732), .C2(n20279), .A(n20250), .B(n20249), .ZN(
        P1_U3047) );
  AOI22_X1 U23182 ( .A1(n20736), .A2(n20252), .B1(n20251), .B2(n20734), .ZN(
        n20256) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20671), .ZN(n20255) );
  OAI211_X1 U23184 ( .C1(n20676), .C2(n20279), .A(n20256), .B(n20255), .ZN(
        P1_U3048) );
  NAND2_X1 U23185 ( .A1(n20606), .A2(n20830), .ZN(n20642) );
  NOR2_X2 U23186 ( .A1(n20294), .A2(n20642), .ZN(n20316) );
  NAND2_X1 U23187 ( .A1(n20279), .A2(n20682), .ZN(n20257) );
  OAI21_X1 U23188 ( .B1(n20316), .B2(n20257), .A(n20557), .ZN(n20259) );
  NOR2_X1 U23189 ( .A1(n20258), .A2(n14182), .ZN(n20263) );
  NOR3_X1 U23190 ( .A1(n20490), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20296) );
  NAND2_X1 U23191 ( .A1(n20834), .A2(n20296), .ZN(n20278) );
  INV_X1 U23192 ( .A(n20278), .ZN(n20283) );
  AOI22_X1 U23193 ( .A1(n20316), .A2(n20610), .B1(n20686), .B2(n20283), .ZN(
        n20266) );
  INV_X1 U23194 ( .A(n20259), .ZN(n20264) );
  NOR2_X1 U23195 ( .A1(n10263), .A2(n20260), .ZN(n20378) );
  AOI211_X1 U23196 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20278), .A(n20378), 
        .B(n20261), .ZN(n20262) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20691), .ZN(n20265) );
  OAI211_X1 U23198 ( .C1(n20288), .C2(n20571), .A(n20266), .B(n20265), .ZN(
        P1_U3049) );
  INV_X1 U23199 ( .A(n20695), .ZN(n20574) );
  AOI22_X1 U23200 ( .A1(n20284), .A2(n20697), .B1(n20696), .B2(n20283), .ZN(
        n20268) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20285), .B1(
        n20316), .B2(n20614), .ZN(n20267) );
  OAI211_X1 U23202 ( .C1(n20288), .C2(n20574), .A(n20268), .B(n20267), .ZN(
        P1_U3050) );
  INV_X1 U23203 ( .A(n20701), .ZN(n20577) );
  AOI22_X1 U23204 ( .A1(n20316), .A2(n20618), .B1(n20702), .B2(n20283), .ZN(
        n20270) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20703), .ZN(n20269) );
  OAI211_X1 U23206 ( .C1(n20288), .C2(n20577), .A(n20270), .B(n20269), .ZN(
        P1_U3051) );
  INV_X1 U23207 ( .A(n20707), .ZN(n20580) );
  AOI22_X1 U23208 ( .A1(n20316), .A2(n20709), .B1(n20708), .B2(n20283), .ZN(
        n20272) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20659), .ZN(n20271) );
  OAI211_X1 U23210 ( .C1(n20288), .C2(n20580), .A(n20272), .B(n20271), .ZN(
        P1_U3052) );
  INV_X1 U23211 ( .A(n20713), .ZN(n20583) );
  AOI22_X1 U23212 ( .A1(n20284), .A2(n20715), .B1(n20714), .B2(n20283), .ZN(
        n20274) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20285), .B1(
        n20316), .B2(n20624), .ZN(n20273) );
  OAI211_X1 U23214 ( .C1(n20288), .C2(n20583), .A(n20274), .B(n20273), .ZN(
        P1_U3053) );
  INV_X1 U23215 ( .A(n20721), .ZN(n20631) );
  INV_X1 U23216 ( .A(n20720), .ZN(n20507) );
  OAI22_X1 U23217 ( .A1(n20279), .A2(n20631), .B1(n20507), .B2(n20278), .ZN(
        n20275) );
  INV_X1 U23218 ( .A(n20275), .ZN(n20277) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20285), .B1(
        n20316), .B2(n20628), .ZN(n20276) );
  OAI211_X1 U23220 ( .C1(n20288), .C2(n20586), .A(n20277), .B(n20276), .ZN(
        P1_U3054) );
  INV_X1 U23221 ( .A(n20725), .ZN(n20589) );
  INV_X1 U23222 ( .A(n20727), .ZN(n20635) );
  INV_X1 U23223 ( .A(n20726), .ZN(n20512) );
  OAI22_X1 U23224 ( .A1(n20279), .A2(n20635), .B1(n20512), .B2(n20278), .ZN(
        n20280) );
  INV_X1 U23225 ( .A(n20280), .ZN(n20282) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20285), .B1(
        n20316), .B2(n20632), .ZN(n20281) );
  OAI211_X1 U23227 ( .C1(n20288), .C2(n20589), .A(n20282), .B(n20281), .ZN(
        P1_U3055) );
  INV_X1 U23228 ( .A(n20734), .ZN(n20596) );
  AOI22_X1 U23229 ( .A1(n20316), .A2(n20737), .B1(n20736), .B2(n20283), .ZN(
        n20287) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20671), .ZN(n20286) );
  OAI211_X1 U23231 ( .C1(n20288), .C2(n20596), .A(n20287), .B(n20286), .ZN(
        P1_U3056) );
  INV_X1 U23232 ( .A(n20296), .ZN(n20292) );
  AND2_X1 U23233 ( .A1(n10570), .A2(n20289), .ZN(n20678) );
  NOR2_X1 U23234 ( .A1(n20524), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20315) );
  AOI21_X1 U23235 ( .B1(n20290), .B2(n20678), .A(n20315), .ZN(n20298) );
  INV_X1 U23236 ( .A(n20527), .ZN(n20291) );
  AOI21_X1 U23237 ( .B1(n20294), .B2(n20682), .A(n20291), .ZN(n20295) );
  OAI22_X1 U23238 ( .A1(n20260), .A2(n20292), .B1(n20298), .B2(n20295), .ZN(
        n20293) );
  NOR2_X2 U23239 ( .A1(n20294), .A2(n20533), .ZN(n20346) );
  AOI22_X1 U23240 ( .A1(n20346), .A2(n20610), .B1(n20686), .B2(n20315), .ZN(
        n20302) );
  INV_X1 U23241 ( .A(n20295), .ZN(n20299) );
  OAI21_X1 U23242 ( .B1(n20813), .B2(n20296), .A(n20689), .ZN(n20297) );
  AOI21_X1 U23243 ( .B1(n20299), .B2(n20298), .A(n20297), .ZN(n20300) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20691), .ZN(n20301) );
  OAI211_X1 U23245 ( .C1(n20320), .C2(n20571), .A(n20302), .B(n20301), .ZN(
        P1_U3057) );
  AOI22_X1 U23246 ( .A1(n20316), .A2(n20697), .B1(n20696), .B2(n20315), .ZN(
        n20304) );
  AOI22_X1 U23247 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20317), .B1(
        n20346), .B2(n20614), .ZN(n20303) );
  OAI211_X1 U23248 ( .C1(n20320), .C2(n20574), .A(n20304), .B(n20303), .ZN(
        P1_U3058) );
  AOI22_X1 U23249 ( .A1(n20316), .A2(n20703), .B1(n20702), .B2(n20315), .ZN(
        n20306) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20317), .B1(
        n20346), .B2(n20618), .ZN(n20305) );
  OAI211_X1 U23251 ( .C1(n20320), .C2(n20577), .A(n20306), .B(n20305), .ZN(
        P1_U3059) );
  AOI22_X1 U23252 ( .A1(n20346), .A2(n20709), .B1(n20708), .B2(n20315), .ZN(
        n20308) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20659), .ZN(n20307) );
  OAI211_X1 U23254 ( .C1(n20320), .C2(n20580), .A(n20308), .B(n20307), .ZN(
        P1_U3060) );
  AOI22_X1 U23255 ( .A1(n20316), .A2(n20715), .B1(n20714), .B2(n20315), .ZN(
        n20310) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20317), .B1(
        n20346), .B2(n20624), .ZN(n20309) );
  OAI211_X1 U23257 ( .C1(n20320), .C2(n20583), .A(n20310), .B(n20309), .ZN(
        P1_U3061) );
  AOI22_X1 U23258 ( .A1(n20316), .A2(n20721), .B1(n20720), .B2(n20315), .ZN(
        n20312) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20317), .B1(
        n20346), .B2(n20628), .ZN(n20311) );
  OAI211_X1 U23260 ( .C1(n20320), .C2(n20586), .A(n20312), .B(n20311), .ZN(
        P1_U3062) );
  AOI22_X1 U23261 ( .A1(n20316), .A2(n20727), .B1(n20726), .B2(n20315), .ZN(
        n20314) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20317), .B1(
        n20346), .B2(n20632), .ZN(n20313) );
  OAI211_X1 U23263 ( .C1(n20320), .C2(n20589), .A(n20314), .B(n20313), .ZN(
        P1_U3063) );
  AOI22_X1 U23264 ( .A1(n20346), .A2(n20737), .B1(n20736), .B2(n20315), .ZN(
        n20319) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20317), .B1(
        n20316), .B2(n20671), .ZN(n20318) );
  OAI211_X1 U23266 ( .C1(n20320), .C2(n20596), .A(n20319), .B(n20318), .ZN(
        P1_U3064) );
  NOR3_X1 U23267 ( .A1(n20562), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20353) );
  INV_X1 U23268 ( .A(n20353), .ZN(n20350) );
  NOR2_X1 U23269 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20350), .ZN(
        n20345) );
  INV_X1 U23270 ( .A(n20561), .ZN(n20644) );
  NOR2_X1 U23271 ( .A1(n13446), .A2(n20322), .ZN(n20403) );
  NAND3_X1 U23272 ( .A1(n20403), .A2(n20813), .A3(n14182), .ZN(n20323) );
  OAI21_X1 U23273 ( .B1(n20324), .B2(n20644), .A(n20323), .ZN(n20344) );
  AOI22_X1 U23274 ( .A1(n20686), .A2(n20345), .B1(n20685), .B2(n20344), .ZN(
        n20331) );
  INV_X1 U23275 ( .A(n20346), .ZN(n20325) );
  AOI21_X1 U23276 ( .B1(n20325), .B2(n20373), .A(n20814), .ZN(n20326) );
  AOI21_X1 U23277 ( .B1(n20403), .B2(n14182), .A(n20326), .ZN(n20327) );
  NOR2_X1 U23278 ( .A1(n20327), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20329) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20691), .ZN(n20330) );
  OAI211_X1 U23280 ( .C1(n20694), .C2(n20373), .A(n20331), .B(n20330), .ZN(
        P1_U3065) );
  AOI22_X1 U23281 ( .A1(n20696), .A2(n20345), .B1(n20695), .B2(n20344), .ZN(
        n20333) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20697), .ZN(n20332) );
  OAI211_X1 U23283 ( .C1(n20700), .C2(n20373), .A(n20333), .B(n20332), .ZN(
        P1_U3066) );
  AOI22_X1 U23284 ( .A1(n20702), .A2(n20345), .B1(n20701), .B2(n20344), .ZN(
        n20335) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20703), .ZN(n20334) );
  OAI211_X1 U23286 ( .C1(n20706), .C2(n20373), .A(n20335), .B(n20334), .ZN(
        P1_U3067) );
  AOI22_X1 U23287 ( .A1(n20708), .A2(n20345), .B1(n20707), .B2(n20344), .ZN(
        n20337) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20659), .ZN(n20336) );
  OAI211_X1 U23289 ( .C1(n20662), .C2(n20373), .A(n20337), .B(n20336), .ZN(
        P1_U3068) );
  AOI22_X1 U23290 ( .A1(n20714), .A2(n20345), .B1(n20713), .B2(n20344), .ZN(
        n20339) );
  AOI22_X1 U23291 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20715), .ZN(n20338) );
  OAI211_X1 U23292 ( .C1(n20718), .C2(n20373), .A(n20339), .B(n20338), .ZN(
        P1_U3069) );
  AOI22_X1 U23293 ( .A1(n20720), .A2(n20345), .B1(n20719), .B2(n20344), .ZN(
        n20341) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20721), .ZN(n20340) );
  OAI211_X1 U23295 ( .C1(n20724), .C2(n20373), .A(n20341), .B(n20340), .ZN(
        P1_U3070) );
  AOI22_X1 U23296 ( .A1(n20726), .A2(n20345), .B1(n20725), .B2(n20344), .ZN(
        n20343) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20727), .ZN(n20342) );
  OAI211_X1 U23298 ( .C1(n20732), .C2(n20373), .A(n20343), .B(n20342), .ZN(
        P1_U3071) );
  AOI22_X1 U23299 ( .A1(n20736), .A2(n20345), .B1(n20734), .B2(n20344), .ZN(
        n20349) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20671), .ZN(n20348) );
  OAI211_X1 U23301 ( .C1(n20676), .C2(n20373), .A(n20349), .B(n20348), .ZN(
        P1_U3072) );
  INV_X1 U23302 ( .A(n20691), .ZN(n20613) );
  NOR2_X1 U23303 ( .A1(n20834), .A2(n20350), .ZN(n20369) );
  AOI21_X1 U23304 ( .B1(n20403), .B2(n20461), .A(n20369), .ZN(n20351) );
  OAI22_X1 U23305 ( .A1(n20351), .A2(n20829), .B1(n20350), .B2(n20260), .ZN(
        n20368) );
  AOI22_X1 U23306 ( .A1(n20686), .A2(n20369), .B1(n20685), .B2(n20368), .ZN(
        n20355) );
  OAI211_X1 U23307 ( .C1(n20819), .C2(n20814), .A(n20813), .B(n20351), .ZN(
        n20352) );
  OAI211_X1 U23308 ( .C1(n20813), .C2(n20353), .A(n20689), .B(n20352), .ZN(
        n20370) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20370), .B1(
        n20397), .B2(n20610), .ZN(n20354) );
  OAI211_X1 U23310 ( .C1(n20613), .C2(n20373), .A(n20355), .B(n20354), .ZN(
        P1_U3073) );
  INV_X1 U23311 ( .A(n20697), .ZN(n20617) );
  AOI22_X1 U23312 ( .A1(n20696), .A2(n20369), .B1(n20695), .B2(n20368), .ZN(
        n20357) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20370), .B1(
        n20397), .B2(n20614), .ZN(n20356) );
  OAI211_X1 U23314 ( .C1(n20617), .C2(n20373), .A(n20357), .B(n20356), .ZN(
        P1_U3074) );
  INV_X1 U23315 ( .A(n20703), .ZN(n20621) );
  AOI22_X1 U23316 ( .A1(n20702), .A2(n20369), .B1(n20701), .B2(n20368), .ZN(
        n20359) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20370), .B1(
        n20397), .B2(n20618), .ZN(n20358) );
  OAI211_X1 U23318 ( .C1(n20621), .C2(n20373), .A(n20359), .B(n20358), .ZN(
        P1_U3075) );
  INV_X1 U23319 ( .A(n20659), .ZN(n20712) );
  AOI22_X1 U23320 ( .A1(n20708), .A2(n20369), .B1(n20707), .B2(n20368), .ZN(
        n20361) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20370), .B1(
        n20397), .B2(n20709), .ZN(n20360) );
  OAI211_X1 U23322 ( .C1(n20712), .C2(n20373), .A(n20361), .B(n20360), .ZN(
        P1_U3076) );
  INV_X1 U23323 ( .A(n20715), .ZN(n20627) );
  AOI22_X1 U23324 ( .A1(n20714), .A2(n20369), .B1(n20713), .B2(n20368), .ZN(
        n20363) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20370), .B1(
        n20397), .B2(n20624), .ZN(n20362) );
  OAI211_X1 U23326 ( .C1(n20627), .C2(n20373), .A(n20363), .B(n20362), .ZN(
        P1_U3077) );
  AOI22_X1 U23327 ( .A1(n20720), .A2(n20369), .B1(n20719), .B2(n20368), .ZN(
        n20365) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20370), .B1(
        n20397), .B2(n20628), .ZN(n20364) );
  OAI211_X1 U23329 ( .C1(n20631), .C2(n20373), .A(n20365), .B(n20364), .ZN(
        P1_U3078) );
  AOI22_X1 U23330 ( .A1(n20726), .A2(n20369), .B1(n20725), .B2(n20368), .ZN(
        n20367) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20370), .B1(
        n20397), .B2(n20632), .ZN(n20366) );
  OAI211_X1 U23332 ( .C1(n20635), .C2(n20373), .A(n20367), .B(n20366), .ZN(
        P1_U3079) );
  INV_X1 U23333 ( .A(n20671), .ZN(n20743) );
  AOI22_X1 U23334 ( .A1(n20736), .A2(n20369), .B1(n20734), .B2(n20368), .ZN(
        n20372) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20370), .B1(
        n20397), .B2(n20737), .ZN(n20371) );
  OAI211_X1 U23336 ( .C1(n20743), .C2(n20373), .A(n20372), .B(n20371), .ZN(
        P1_U3080) );
  INV_X1 U23337 ( .A(n20397), .ZN(n20374) );
  NAND2_X1 U23338 ( .A1(n20374), .A2(n20682), .ZN(n20375) );
  NOR2_X2 U23339 ( .A1(n20819), .A2(n20642), .ZN(n20427) );
  OAI21_X1 U23340 ( .B1(n20375), .B2(n20427), .A(n20557), .ZN(n20380) );
  AND2_X1 U23341 ( .A1(n20403), .A2(n20647), .ZN(n20377) );
  NOR2_X1 U23342 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20376), .ZN(
        n20396) );
  AOI22_X1 U23343 ( .A1(n20397), .A2(n20691), .B1(n20686), .B2(n20396), .ZN(
        n20383) );
  INV_X1 U23344 ( .A(n20377), .ZN(n20379) );
  AOI21_X1 U23345 ( .B1(n20380), .B2(n20379), .A(n20378), .ZN(n20381) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20398), .B1(
        n20427), .B2(n20610), .ZN(n20382) );
  OAI211_X1 U23347 ( .C1(n20401), .C2(n20571), .A(n20383), .B(n20382), .ZN(
        P1_U3081) );
  AOI22_X1 U23348 ( .A1(n20427), .A2(n20614), .B1(n20696), .B2(n20396), .ZN(
        n20385) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20398), .B1(
        n20397), .B2(n20697), .ZN(n20384) );
  OAI211_X1 U23350 ( .C1(n20401), .C2(n20574), .A(n20385), .B(n20384), .ZN(
        P1_U3082) );
  AOI22_X1 U23351 ( .A1(n20397), .A2(n20703), .B1(n20702), .B2(n20396), .ZN(
        n20387) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20398), .B1(
        n20427), .B2(n20618), .ZN(n20386) );
  OAI211_X1 U23353 ( .C1(n20401), .C2(n20577), .A(n20387), .B(n20386), .ZN(
        P1_U3083) );
  AOI22_X1 U23354 ( .A1(n20427), .A2(n20709), .B1(n20708), .B2(n20396), .ZN(
        n20389) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20398), .B1(
        n20397), .B2(n20659), .ZN(n20388) );
  OAI211_X1 U23356 ( .C1(n20401), .C2(n20580), .A(n20389), .B(n20388), .ZN(
        P1_U3084) );
  AOI22_X1 U23357 ( .A1(n20427), .A2(n20624), .B1(n20714), .B2(n20396), .ZN(
        n20391) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20398), .B1(
        n20397), .B2(n20715), .ZN(n20390) );
  OAI211_X1 U23359 ( .C1(n20401), .C2(n20583), .A(n20391), .B(n20390), .ZN(
        P1_U3085) );
  AOI22_X1 U23360 ( .A1(n20427), .A2(n20628), .B1(n20720), .B2(n20396), .ZN(
        n20393) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20398), .B1(
        n20397), .B2(n20721), .ZN(n20392) );
  OAI211_X1 U23362 ( .C1(n20401), .C2(n20586), .A(n20393), .B(n20392), .ZN(
        P1_U3086) );
  AOI22_X1 U23363 ( .A1(n20397), .A2(n20727), .B1(n20726), .B2(n20396), .ZN(
        n20395) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20398), .B1(
        n20427), .B2(n20632), .ZN(n20394) );
  OAI211_X1 U23365 ( .C1(n20401), .C2(n20589), .A(n20395), .B(n20394), .ZN(
        P1_U3087) );
  AOI22_X1 U23366 ( .A1(n20397), .A2(n20671), .B1(n20736), .B2(n20396), .ZN(
        n20400) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20398), .B1(
        n20427), .B2(n20737), .ZN(n20399) );
  OAI211_X1 U23368 ( .C1(n20401), .C2(n20596), .A(n20400), .B(n20399), .ZN(
        P1_U3088) );
  INV_X1 U23369 ( .A(n20402), .ZN(n20426) );
  AOI21_X1 U23370 ( .B1(n20403), .B2(n20678), .A(n20426), .ZN(n20407) );
  OR2_X1 U23371 ( .A1(n20407), .A2(n20829), .ZN(n20405) );
  NAND2_X1 U23372 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20410), .ZN(n20404) );
  NAND2_X1 U23373 ( .A1(n20405), .A2(n20404), .ZN(n20425) );
  AOI22_X1 U23374 ( .A1(n20686), .A2(n20426), .B1(n20685), .B2(n20425), .ZN(
        n20412) );
  INV_X1 U23375 ( .A(n20819), .ZN(n20406) );
  OAI21_X1 U23376 ( .B1(n20406), .B2(n20829), .A(n20527), .ZN(n20408) );
  NAND2_X1 U23377 ( .A1(n20408), .A2(n20407), .ZN(n20409) );
  OAI211_X1 U23378 ( .C1(n20410), .C2(n20813), .A(n20689), .B(n20409), .ZN(
        n20428) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20691), .ZN(n20411) );
  OAI211_X1 U23380 ( .C1(n20694), .C2(n20436), .A(n20412), .B(n20411), .ZN(
        P1_U3089) );
  AOI22_X1 U23381 ( .A1(n20696), .A2(n20426), .B1(n20695), .B2(n20425), .ZN(
        n20414) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20697), .ZN(n20413) );
  OAI211_X1 U23383 ( .C1(n20700), .C2(n20436), .A(n20414), .B(n20413), .ZN(
        P1_U3090) );
  AOI22_X1 U23384 ( .A1(n20702), .A2(n20426), .B1(n20701), .B2(n20425), .ZN(
        n20416) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20703), .ZN(n20415) );
  OAI211_X1 U23386 ( .C1(n20706), .C2(n20436), .A(n20416), .B(n20415), .ZN(
        P1_U3091) );
  AOI22_X1 U23387 ( .A1(n20708), .A2(n20426), .B1(n20707), .B2(n20425), .ZN(
        n20418) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20659), .ZN(n20417) );
  OAI211_X1 U23389 ( .C1(n20662), .C2(n20436), .A(n20418), .B(n20417), .ZN(
        P1_U3092) );
  AOI22_X1 U23390 ( .A1(n20714), .A2(n20426), .B1(n20713), .B2(n20425), .ZN(
        n20420) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20715), .ZN(n20419) );
  OAI211_X1 U23392 ( .C1(n20718), .C2(n20436), .A(n20420), .B(n20419), .ZN(
        P1_U3093) );
  AOI22_X1 U23393 ( .A1(n20720), .A2(n20426), .B1(n20719), .B2(n20425), .ZN(
        n20422) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20721), .ZN(n20421) );
  OAI211_X1 U23395 ( .C1(n20724), .C2(n20436), .A(n20422), .B(n20421), .ZN(
        P1_U3094) );
  AOI22_X1 U23396 ( .A1(n20726), .A2(n20426), .B1(n20725), .B2(n20425), .ZN(
        n20424) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20727), .ZN(n20423) );
  OAI211_X1 U23398 ( .C1(n20732), .C2(n20436), .A(n20424), .B(n20423), .ZN(
        P1_U3095) );
  AOI22_X1 U23399 ( .A1(n20736), .A2(n20426), .B1(n20734), .B2(n20425), .ZN(
        n20430) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20671), .ZN(n20429) );
  OAI211_X1 U23401 ( .C1(n20676), .C2(n20436), .A(n20430), .B(n20429), .ZN(
        P1_U3096) );
  INV_X1 U23402 ( .A(n20555), .ZN(n20432) );
  NOR3_X1 U23403 ( .A1(n20825), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20465) );
  INV_X1 U23404 ( .A(n20465), .ZN(n20462) );
  NOR2_X1 U23405 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20462), .ZN(
        n20456) );
  AND2_X1 U23406 ( .A1(n20817), .A2(n13446), .ZN(n20525) );
  AOI21_X1 U23407 ( .B1(n20525), .B2(n14182), .A(n20456), .ZN(n20438) );
  INV_X1 U23408 ( .A(n20487), .ZN(n20434) );
  NOR2_X1 U23409 ( .A1(n20434), .A2(n20433), .ZN(n20560) );
  INV_X1 U23410 ( .A(n20560), .ZN(n20564) );
  OAI22_X1 U23411 ( .A1(n20438), .A2(n20829), .B1(n20564), .B2(n20435), .ZN(
        n20455) );
  AOI22_X1 U23412 ( .A1(n20686), .A2(n20456), .B1(n20685), .B2(n20455), .ZN(
        n20442) );
  INV_X1 U23413 ( .A(n20485), .ZN(n20437) );
  OAI21_X1 U23414 ( .B1(n20437), .B2(n20457), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20439) );
  NAND2_X1 U23415 ( .A1(n20439), .A2(n20438), .ZN(n20440) );
  OAI211_X1 U23416 ( .C1(n20456), .C2(n20568), .A(n20492), .B(n20440), .ZN(
        n20458) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20691), .ZN(n20441) );
  OAI211_X1 U23418 ( .C1(n20694), .C2(n20485), .A(n20442), .B(n20441), .ZN(
        P1_U3097) );
  AOI22_X1 U23419 ( .A1(n20696), .A2(n20456), .B1(n20695), .B2(n20455), .ZN(
        n20444) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20697), .ZN(n20443) );
  OAI211_X1 U23421 ( .C1(n20700), .C2(n20485), .A(n20444), .B(n20443), .ZN(
        P1_U3098) );
  AOI22_X1 U23422 ( .A1(n20702), .A2(n20456), .B1(n20701), .B2(n20455), .ZN(
        n20446) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20703), .ZN(n20445) );
  OAI211_X1 U23424 ( .C1(n20706), .C2(n20485), .A(n20446), .B(n20445), .ZN(
        P1_U3099) );
  AOI22_X1 U23425 ( .A1(n20708), .A2(n20456), .B1(n20707), .B2(n20455), .ZN(
        n20448) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20659), .ZN(n20447) );
  OAI211_X1 U23427 ( .C1(n20662), .C2(n20485), .A(n20448), .B(n20447), .ZN(
        P1_U3100) );
  AOI22_X1 U23428 ( .A1(n20714), .A2(n20456), .B1(n20713), .B2(n20455), .ZN(
        n20450) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20715), .ZN(n20449) );
  OAI211_X1 U23430 ( .C1(n20718), .C2(n20485), .A(n20450), .B(n20449), .ZN(
        P1_U3101) );
  AOI22_X1 U23431 ( .A1(n20720), .A2(n20456), .B1(n20719), .B2(n20455), .ZN(
        n20452) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20721), .ZN(n20451) );
  OAI211_X1 U23433 ( .C1(n20724), .C2(n20485), .A(n20452), .B(n20451), .ZN(
        P1_U3102) );
  AOI22_X1 U23434 ( .A1(n20726), .A2(n20456), .B1(n20725), .B2(n20455), .ZN(
        n20454) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20727), .ZN(n20453) );
  OAI211_X1 U23436 ( .C1(n20732), .C2(n20485), .A(n20454), .B(n20453), .ZN(
        P1_U3103) );
  AOI22_X1 U23437 ( .A1(n20736), .A2(n20456), .B1(n20734), .B2(n20455), .ZN(
        n20460) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20671), .ZN(n20459) );
  OAI211_X1 U23439 ( .C1(n20676), .C2(n20485), .A(n20460), .B(n20459), .ZN(
        P1_U3104) );
  NOR2_X1 U23440 ( .A1(n20834), .A2(n20462), .ZN(n20481) );
  AOI21_X1 U23441 ( .B1(n20525), .B2(n20461), .A(n20481), .ZN(n20463) );
  OAI22_X1 U23442 ( .A1(n20463), .A2(n20829), .B1(n20462), .B2(n20260), .ZN(
        n20480) );
  AOI22_X1 U23443 ( .A1(n20686), .A2(n20481), .B1(n20685), .B2(n20480), .ZN(
        n20467) );
  OAI211_X1 U23444 ( .C1(n20534), .C2(n20814), .A(n20813), .B(n20463), .ZN(
        n20464) );
  OAI211_X1 U23445 ( .C1(n20813), .C2(n20465), .A(n20689), .B(n20464), .ZN(
        n20482) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20482), .B1(
        n20518), .B2(n20610), .ZN(n20466) );
  OAI211_X1 U23447 ( .C1(n20613), .C2(n20485), .A(n20467), .B(n20466), .ZN(
        P1_U3105) );
  AOI22_X1 U23448 ( .A1(n20696), .A2(n20481), .B1(n20695), .B2(n20480), .ZN(
        n20469) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20482), .B1(
        n20518), .B2(n20614), .ZN(n20468) );
  OAI211_X1 U23450 ( .C1(n20617), .C2(n20485), .A(n20469), .B(n20468), .ZN(
        P1_U3106) );
  AOI22_X1 U23451 ( .A1(n20702), .A2(n20481), .B1(n20701), .B2(n20480), .ZN(
        n20471) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20482), .B1(
        n20518), .B2(n20618), .ZN(n20470) );
  OAI211_X1 U23453 ( .C1(n20621), .C2(n20485), .A(n20471), .B(n20470), .ZN(
        P1_U3107) );
  AOI22_X1 U23454 ( .A1(n20708), .A2(n20481), .B1(n20707), .B2(n20480), .ZN(
        n20473) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20482), .B1(
        n20518), .B2(n20709), .ZN(n20472) );
  OAI211_X1 U23456 ( .C1(n20712), .C2(n20485), .A(n20473), .B(n20472), .ZN(
        P1_U3108) );
  AOI22_X1 U23457 ( .A1(n20714), .A2(n20481), .B1(n20713), .B2(n20480), .ZN(
        n20475) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20482), .B1(
        n20518), .B2(n20624), .ZN(n20474) );
  OAI211_X1 U23459 ( .C1(n20627), .C2(n20485), .A(n20475), .B(n20474), .ZN(
        P1_U3109) );
  AOI22_X1 U23460 ( .A1(n20720), .A2(n20481), .B1(n20719), .B2(n20480), .ZN(
        n20477) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20482), .B1(
        n20518), .B2(n20628), .ZN(n20476) );
  OAI211_X1 U23462 ( .C1(n20631), .C2(n20485), .A(n20477), .B(n20476), .ZN(
        P1_U3110) );
  AOI22_X1 U23463 ( .A1(n20726), .A2(n20481), .B1(n20725), .B2(n20480), .ZN(
        n20479) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20482), .B1(
        n20518), .B2(n20632), .ZN(n20478) );
  OAI211_X1 U23465 ( .C1(n20635), .C2(n20485), .A(n20479), .B(n20478), .ZN(
        P1_U3111) );
  AOI22_X1 U23466 ( .A1(n20736), .A2(n20481), .B1(n20734), .B2(n20480), .ZN(
        n20484) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20482), .B1(
        n20518), .B2(n20737), .ZN(n20483) );
  OAI211_X1 U23468 ( .C1(n20743), .C2(n20485), .A(n20484), .B(n20483), .ZN(
        P1_U3112) );
  NAND3_X1 U23469 ( .A1(n20554), .A2(n20513), .A3(n20813), .ZN(n20486) );
  NAND2_X1 U23470 ( .A1(n20486), .A2(n20557), .ZN(n20495) );
  AND2_X1 U23471 ( .A1(n20525), .A2(n20647), .ZN(n20491) );
  OR2_X1 U23472 ( .A1(n20487), .A2(n20825), .ZN(n20643) );
  INV_X1 U23473 ( .A(n20643), .ZN(n20488) );
  NOR3_X1 U23474 ( .A1(n20825), .A2(n20490), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20532) );
  INV_X1 U23475 ( .A(n20532), .ZN(n20526) );
  NOR2_X1 U23476 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20526), .ZN(
        n20517) );
  AOI22_X1 U23477 ( .A1(n20519), .A2(n20610), .B1(n20686), .B2(n20517), .ZN(
        n20498) );
  INV_X1 U23478 ( .A(n20491), .ZN(n20494) );
  NAND2_X1 U23479 ( .A1(n20643), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20650) );
  OAI211_X1 U23480 ( .C1(n20568), .C2(n20517), .A(n20650), .B(n20492), .ZN(
        n20493) );
  AOI21_X1 U23481 ( .B1(n20495), .B2(n20494), .A(n20493), .ZN(n20496) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20520), .B1(
        n20518), .B2(n20691), .ZN(n20497) );
  OAI211_X1 U23483 ( .C1(n20523), .C2(n20571), .A(n20498), .B(n20497), .ZN(
        P1_U3113) );
  AOI22_X1 U23484 ( .A1(n20519), .A2(n20614), .B1(n20696), .B2(n20517), .ZN(
        n20500) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20520), .B1(
        n20518), .B2(n20697), .ZN(n20499) );
  OAI211_X1 U23486 ( .C1(n20523), .C2(n20574), .A(n20500), .B(n20499), .ZN(
        P1_U3114) );
  AOI22_X1 U23487 ( .A1(n20519), .A2(n20618), .B1(n20702), .B2(n20517), .ZN(
        n20502) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20520), .B1(
        n20518), .B2(n20703), .ZN(n20501) );
  OAI211_X1 U23489 ( .C1(n20523), .C2(n20577), .A(n20502), .B(n20501), .ZN(
        P1_U3115) );
  AOI22_X1 U23490 ( .A1(n20519), .A2(n20709), .B1(n20708), .B2(n20517), .ZN(
        n20504) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20520), .B1(
        n20518), .B2(n20659), .ZN(n20503) );
  OAI211_X1 U23492 ( .C1(n20523), .C2(n20580), .A(n20504), .B(n20503), .ZN(
        P1_U3116) );
  AOI22_X1 U23493 ( .A1(n20519), .A2(n20624), .B1(n20714), .B2(n20517), .ZN(
        n20506) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20520), .B1(
        n20518), .B2(n20715), .ZN(n20505) );
  OAI211_X1 U23495 ( .C1(n20523), .C2(n20583), .A(n20506), .B(n20505), .ZN(
        P1_U3117) );
  INV_X1 U23496 ( .A(n20517), .ZN(n20511) );
  OAI22_X1 U23497 ( .A1(n20513), .A2(n20631), .B1(n20507), .B2(n20511), .ZN(
        n20508) );
  INV_X1 U23498 ( .A(n20508), .ZN(n20510) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20520), .B1(
        n20519), .B2(n20628), .ZN(n20509) );
  OAI211_X1 U23500 ( .C1(n20523), .C2(n20586), .A(n20510), .B(n20509), .ZN(
        P1_U3118) );
  OAI22_X1 U23501 ( .A1(n20513), .A2(n20635), .B1(n20512), .B2(n20511), .ZN(
        n20514) );
  INV_X1 U23502 ( .A(n20514), .ZN(n20516) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20520), .B1(
        n20519), .B2(n20632), .ZN(n20515) );
  OAI211_X1 U23504 ( .C1(n20523), .C2(n20589), .A(n20516), .B(n20515), .ZN(
        P1_U3119) );
  AOI22_X1 U23505 ( .A1(n20518), .A2(n20671), .B1(n20736), .B2(n20517), .ZN(
        n20522) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20520), .B1(
        n20519), .B2(n20737), .ZN(n20521) );
  OAI211_X1 U23507 ( .C1(n20523), .C2(n20596), .A(n20522), .B(n20521), .ZN(
        P1_U3120) );
  NOR2_X1 U23508 ( .A1(n20524), .A2(n20825), .ZN(n20550) );
  AOI21_X1 U23509 ( .B1(n20525), .B2(n20678), .A(n20550), .ZN(n20529) );
  OAI22_X1 U23510 ( .A1(n20529), .A2(n20829), .B1(n20526), .B2(n20260), .ZN(
        n20549) );
  AOI22_X1 U23511 ( .A1(n20686), .A2(n20550), .B1(n20685), .B2(n20549), .ZN(
        n20536) );
  OAI21_X1 U23512 ( .B1(n20528), .B2(n20829), .A(n20527), .ZN(n20530) );
  NAND2_X1 U23513 ( .A1(n20530), .A2(n20529), .ZN(n20531) );
  OAI211_X1 U23514 ( .C1(n20813), .C2(n20532), .A(n20689), .B(n20531), .ZN(
        n20551) );
  OR2_X1 U23515 ( .A1(n20534), .A2(n20533), .ZN(n20556) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20551), .B1(
        n20592), .B2(n20610), .ZN(n20535) );
  OAI211_X1 U23517 ( .C1(n20613), .C2(n20554), .A(n20536), .B(n20535), .ZN(
        P1_U3121) );
  AOI22_X1 U23518 ( .A1(n20696), .A2(n20550), .B1(n20695), .B2(n20549), .ZN(
        n20538) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20551), .B1(
        n20592), .B2(n20614), .ZN(n20537) );
  OAI211_X1 U23520 ( .C1(n20617), .C2(n20554), .A(n20538), .B(n20537), .ZN(
        P1_U3122) );
  AOI22_X1 U23521 ( .A1(n20702), .A2(n20550), .B1(n20701), .B2(n20549), .ZN(
        n20540) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20551), .B1(
        n20592), .B2(n20618), .ZN(n20539) );
  OAI211_X1 U23523 ( .C1(n20621), .C2(n20554), .A(n20540), .B(n20539), .ZN(
        P1_U3123) );
  AOI22_X1 U23524 ( .A1(n20708), .A2(n20550), .B1(n20707), .B2(n20549), .ZN(
        n20542) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20551), .B1(
        n20592), .B2(n20709), .ZN(n20541) );
  OAI211_X1 U23526 ( .C1(n20712), .C2(n20554), .A(n20542), .B(n20541), .ZN(
        P1_U3124) );
  AOI22_X1 U23527 ( .A1(n20714), .A2(n20550), .B1(n20713), .B2(n20549), .ZN(
        n20544) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20551), .B1(
        n20592), .B2(n20624), .ZN(n20543) );
  OAI211_X1 U23529 ( .C1(n20627), .C2(n20554), .A(n20544), .B(n20543), .ZN(
        P1_U3125) );
  AOI22_X1 U23530 ( .A1(n20720), .A2(n20550), .B1(n20719), .B2(n20549), .ZN(
        n20546) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20551), .B1(
        n20592), .B2(n20628), .ZN(n20545) );
  OAI211_X1 U23532 ( .C1(n20631), .C2(n20554), .A(n20546), .B(n20545), .ZN(
        P1_U3126) );
  AOI22_X1 U23533 ( .A1(n20726), .A2(n20550), .B1(n20725), .B2(n20549), .ZN(
        n20548) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20551), .B1(
        n20592), .B2(n20632), .ZN(n20547) );
  OAI211_X1 U23535 ( .C1(n20635), .C2(n20554), .A(n20548), .B(n20547), .ZN(
        P1_U3127) );
  AOI22_X1 U23536 ( .A1(n20736), .A2(n20550), .B1(n20734), .B2(n20549), .ZN(
        n20553) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20551), .B1(
        n20592), .B2(n20737), .ZN(n20552) );
  OAI211_X1 U23538 ( .C1(n20743), .C2(n20554), .A(n20553), .B(n20552), .ZN(
        P1_U3128) );
  NAND3_X1 U23539 ( .A1(n20556), .A2(n20813), .A3(n20641), .ZN(n20558) );
  NAND2_X1 U23540 ( .A1(n20558), .A2(n20557), .ZN(n20566) );
  OR2_X1 U23541 ( .A1(n13446), .A2(n20559), .ZN(n20598) );
  NOR2_X1 U23542 ( .A1(n20598), .A2(n20647), .ZN(n20563) );
  NOR3_X1 U23543 ( .A1(n20562), .A2(n20825), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20608) );
  INV_X1 U23544 ( .A(n20608), .ZN(n20601) );
  NOR2_X1 U23545 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20601), .ZN(
        n20590) );
  AOI22_X1 U23546 ( .A1(n20591), .A2(n20610), .B1(n20686), .B2(n20590), .ZN(
        n20570) );
  INV_X1 U23547 ( .A(n20563), .ZN(n20565) );
  AOI22_X1 U23548 ( .A1(n20566), .A2(n20565), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20564), .ZN(n20567) );
  OAI211_X1 U23549 ( .C1(n20590), .C2(n20568), .A(n20651), .B(n20567), .ZN(
        n20593) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20691), .ZN(n20569) );
  OAI211_X1 U23551 ( .C1(n20597), .C2(n20571), .A(n20570), .B(n20569), .ZN(
        P1_U3129) );
  AOI22_X1 U23552 ( .A1(n20591), .A2(n20614), .B1(n20590), .B2(n20696), .ZN(
        n20573) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20697), .ZN(n20572) );
  OAI211_X1 U23554 ( .C1(n20597), .C2(n20574), .A(n20573), .B(n20572), .ZN(
        P1_U3130) );
  AOI22_X1 U23555 ( .A1(n20591), .A2(n20618), .B1(n20590), .B2(n20702), .ZN(
        n20576) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20703), .ZN(n20575) );
  OAI211_X1 U23557 ( .C1(n20597), .C2(n20577), .A(n20576), .B(n20575), .ZN(
        P1_U3131) );
  AOI22_X1 U23558 ( .A1(n20591), .A2(n20709), .B1(n20590), .B2(n20708), .ZN(
        n20579) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20659), .ZN(n20578) );
  OAI211_X1 U23560 ( .C1(n20597), .C2(n20580), .A(n20579), .B(n20578), .ZN(
        P1_U3132) );
  AOI22_X1 U23561 ( .A1(n20591), .A2(n20624), .B1(n20590), .B2(n20714), .ZN(
        n20582) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20715), .ZN(n20581) );
  OAI211_X1 U23563 ( .C1(n20597), .C2(n20583), .A(n20582), .B(n20581), .ZN(
        P1_U3133) );
  AOI22_X1 U23564 ( .A1(n20591), .A2(n20628), .B1(n20590), .B2(n20720), .ZN(
        n20585) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20721), .ZN(n20584) );
  OAI211_X1 U23566 ( .C1(n20597), .C2(n20586), .A(n20585), .B(n20584), .ZN(
        P1_U3134) );
  AOI22_X1 U23567 ( .A1(n20591), .A2(n20632), .B1(n20590), .B2(n20726), .ZN(
        n20588) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20727), .ZN(n20587) );
  OAI211_X1 U23569 ( .C1(n20597), .C2(n20589), .A(n20588), .B(n20587), .ZN(
        P1_U3135) );
  AOI22_X1 U23570 ( .A1(n20591), .A2(n20737), .B1(n20590), .B2(n20736), .ZN(
        n20595) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20671), .ZN(n20594) );
  OAI211_X1 U23572 ( .C1(n20597), .C2(n20596), .A(n20595), .B(n20594), .ZN(
        P1_U3136) );
  NOR2_X1 U23573 ( .A1(n20834), .A2(n20601), .ZN(n20637) );
  INV_X1 U23574 ( .A(n20598), .ZN(n20648) );
  NAND2_X1 U23575 ( .A1(n20648), .A2(n20682), .ZN(n20680) );
  OR2_X1 U23576 ( .A1(n20680), .A2(n20599), .ZN(n20604) );
  INV_X1 U23577 ( .A(n20637), .ZN(n20600) );
  OAI22_X1 U23578 ( .A1(n20601), .A2(n20260), .B1(n20829), .B2(n20600), .ZN(
        n20602) );
  INV_X1 U23579 ( .A(n20602), .ZN(n20603) );
  NAND2_X1 U23580 ( .A1(n20604), .A2(n20603), .ZN(n20636) );
  AOI22_X1 U23581 ( .A1(n20686), .A2(n20637), .B1(n20685), .B2(n20636), .ZN(
        n20612) );
  OR3_X1 U23582 ( .A1(n20688), .A2(n20606), .A3(n20605), .ZN(n20821) );
  INV_X1 U23583 ( .A(n20821), .ZN(n20607) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20638), .B1(
        n20672), .B2(n20610), .ZN(n20611) );
  OAI211_X1 U23585 ( .C1(n20613), .C2(n20641), .A(n20612), .B(n20611), .ZN(
        P1_U3137) );
  AOI22_X1 U23586 ( .A1(n20696), .A2(n20637), .B1(n20695), .B2(n20636), .ZN(
        n20616) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20638), .B1(
        n20672), .B2(n20614), .ZN(n20615) );
  OAI211_X1 U23588 ( .C1(n20617), .C2(n20641), .A(n20616), .B(n20615), .ZN(
        P1_U3138) );
  AOI22_X1 U23589 ( .A1(n20702), .A2(n20637), .B1(n20701), .B2(n20636), .ZN(
        n20620) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20638), .B1(
        n20672), .B2(n20618), .ZN(n20619) );
  OAI211_X1 U23591 ( .C1(n20621), .C2(n20641), .A(n20620), .B(n20619), .ZN(
        P1_U3139) );
  AOI22_X1 U23592 ( .A1(n20708), .A2(n20637), .B1(n20707), .B2(n20636), .ZN(
        n20623) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20638), .B1(
        n20672), .B2(n20709), .ZN(n20622) );
  OAI211_X1 U23594 ( .C1(n20712), .C2(n20641), .A(n20623), .B(n20622), .ZN(
        P1_U3140) );
  AOI22_X1 U23595 ( .A1(n20714), .A2(n20637), .B1(n20713), .B2(n20636), .ZN(
        n20626) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20638), .B1(
        n20672), .B2(n20624), .ZN(n20625) );
  OAI211_X1 U23597 ( .C1(n20627), .C2(n20641), .A(n20626), .B(n20625), .ZN(
        P1_U3141) );
  AOI22_X1 U23598 ( .A1(n20720), .A2(n20637), .B1(n20719), .B2(n20636), .ZN(
        n20630) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20638), .B1(
        n20672), .B2(n20628), .ZN(n20629) );
  OAI211_X1 U23600 ( .C1(n20631), .C2(n20641), .A(n20630), .B(n20629), .ZN(
        P1_U3142) );
  AOI22_X1 U23601 ( .A1(n20726), .A2(n20637), .B1(n20725), .B2(n20636), .ZN(
        n20634) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20638), .B1(
        n20672), .B2(n20632), .ZN(n20633) );
  OAI211_X1 U23603 ( .C1(n20635), .C2(n20641), .A(n20634), .B(n20633), .ZN(
        P1_U3143) );
  AOI22_X1 U23604 ( .A1(n20736), .A2(n20637), .B1(n20734), .B2(n20636), .ZN(
        n20640) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20638), .B1(
        n20672), .B2(n20737), .ZN(n20639) );
  OAI211_X1 U23606 ( .C1(n20743), .C2(n20641), .A(n20640), .B(n20639), .ZN(
        P1_U3144) );
  NOR2_X1 U23607 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20687), .ZN(
        n20670) );
  OAI22_X1 U23608 ( .A1(n20680), .A2(n14182), .B1(n20644), .B2(n20643), .ZN(
        n20669) );
  AOI22_X1 U23609 ( .A1(n20686), .A2(n20670), .B1(n20685), .B2(n20669), .ZN(
        n20654) );
  AOI21_X1 U23610 ( .B1(n20742), .B2(n20645), .A(n20814), .ZN(n20646) );
  AOI21_X1 U23611 ( .B1(n20648), .B2(n20647), .A(n20646), .ZN(n20649) );
  NOR2_X1 U23612 ( .A1(n20649), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20652) );
  AOI22_X1 U23613 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20673), .B1(
        n20672), .B2(n20691), .ZN(n20653) );
  OAI211_X1 U23614 ( .C1(n20694), .C2(n20742), .A(n20654), .B(n20653), .ZN(
        P1_U3145) );
  AOI22_X1 U23615 ( .A1(n20696), .A2(n20670), .B1(n20695), .B2(n20669), .ZN(
        n20656) );
  AOI22_X1 U23616 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20673), .B1(
        n20672), .B2(n20697), .ZN(n20655) );
  OAI211_X1 U23617 ( .C1(n20700), .C2(n20742), .A(n20656), .B(n20655), .ZN(
        P1_U3146) );
  AOI22_X1 U23618 ( .A1(n20702), .A2(n20670), .B1(n20701), .B2(n20669), .ZN(
        n20658) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20673), .B1(
        n20672), .B2(n20703), .ZN(n20657) );
  OAI211_X1 U23620 ( .C1(n20706), .C2(n20742), .A(n20658), .B(n20657), .ZN(
        P1_U3147) );
  AOI22_X1 U23621 ( .A1(n20708), .A2(n20670), .B1(n20707), .B2(n20669), .ZN(
        n20661) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20673), .B1(
        n20672), .B2(n20659), .ZN(n20660) );
  OAI211_X1 U23623 ( .C1(n20662), .C2(n20742), .A(n20661), .B(n20660), .ZN(
        P1_U3148) );
  AOI22_X1 U23624 ( .A1(n20714), .A2(n20670), .B1(n20713), .B2(n20669), .ZN(
        n20664) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20673), .B1(
        n20672), .B2(n20715), .ZN(n20663) );
  OAI211_X1 U23626 ( .C1(n20718), .C2(n20742), .A(n20664), .B(n20663), .ZN(
        P1_U3149) );
  AOI22_X1 U23627 ( .A1(n20720), .A2(n20670), .B1(n20719), .B2(n20669), .ZN(
        n20666) );
  AOI22_X1 U23628 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20673), .B1(
        n20672), .B2(n20721), .ZN(n20665) );
  OAI211_X1 U23629 ( .C1(n20724), .C2(n20742), .A(n20666), .B(n20665), .ZN(
        P1_U3150) );
  AOI22_X1 U23630 ( .A1(n20726), .A2(n20670), .B1(n20725), .B2(n20669), .ZN(
        n20668) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20673), .B1(
        n20672), .B2(n20727), .ZN(n20667) );
  OAI211_X1 U23632 ( .C1(n20732), .C2(n20742), .A(n20668), .B(n20667), .ZN(
        P1_U3151) );
  AOI22_X1 U23633 ( .A1(n20736), .A2(n20670), .B1(n20734), .B2(n20669), .ZN(
        n20675) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20673), .B1(
        n20672), .B2(n20671), .ZN(n20674) );
  OAI211_X1 U23635 ( .C1(n20676), .C2(n20742), .A(n20675), .B(n20674), .ZN(
        P1_U3152) );
  INV_X1 U23636 ( .A(n20677), .ZN(n20735) );
  INV_X1 U23637 ( .A(n20678), .ZN(n20679) );
  OR2_X1 U23638 ( .A1(n20680), .A2(n20679), .ZN(n20684) );
  AOI22_X1 U23639 ( .A1(n20682), .A2(n20735), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20681), .ZN(n20683) );
  NAND2_X1 U23640 ( .A1(n20684), .A2(n20683), .ZN(n20733) );
  AOI22_X1 U23641 ( .A1(n20686), .A2(n20735), .B1(n20685), .B2(n20733), .ZN(
        n20693) );
  OAI21_X1 U23642 ( .B1(n20688), .B2(n20818), .A(n20687), .ZN(n20690) );
  NAND2_X1 U23643 ( .A1(n20690), .A2(n20689), .ZN(n20739) );
  INV_X1 U23644 ( .A(n20742), .ZN(n20728) );
  AOI22_X1 U23645 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20739), .B1(
        n20728), .B2(n20691), .ZN(n20692) );
  OAI211_X1 U23646 ( .C1(n20694), .C2(n20731), .A(n20693), .B(n20692), .ZN(
        P1_U3153) );
  AOI22_X1 U23647 ( .A1(n20696), .A2(n20735), .B1(n20695), .B2(n20733), .ZN(
        n20699) );
  AOI22_X1 U23648 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20739), .B1(
        n20728), .B2(n20697), .ZN(n20698) );
  OAI211_X1 U23649 ( .C1(n20700), .C2(n20731), .A(n20699), .B(n20698), .ZN(
        P1_U3154) );
  AOI22_X1 U23650 ( .A1(n20702), .A2(n20735), .B1(n20701), .B2(n20733), .ZN(
        n20705) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20739), .B1(
        n20728), .B2(n20703), .ZN(n20704) );
  OAI211_X1 U23652 ( .C1(n20706), .C2(n20731), .A(n20705), .B(n20704), .ZN(
        P1_U3155) );
  AOI22_X1 U23653 ( .A1(n20708), .A2(n20735), .B1(n20707), .B2(n20733), .ZN(
        n20711) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20739), .B1(
        n20738), .B2(n20709), .ZN(n20710) );
  OAI211_X1 U23655 ( .C1(n20712), .C2(n20742), .A(n20711), .B(n20710), .ZN(
        P1_U3156) );
  AOI22_X1 U23656 ( .A1(n20714), .A2(n20735), .B1(n20713), .B2(n20733), .ZN(
        n20717) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20739), .B1(
        n20728), .B2(n20715), .ZN(n20716) );
  OAI211_X1 U23658 ( .C1(n20718), .C2(n20731), .A(n20717), .B(n20716), .ZN(
        P1_U3157) );
  AOI22_X1 U23659 ( .A1(n20720), .A2(n20735), .B1(n20719), .B2(n20733), .ZN(
        n20723) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20739), .B1(
        n20728), .B2(n20721), .ZN(n20722) );
  OAI211_X1 U23661 ( .C1(n20724), .C2(n20731), .A(n20723), .B(n20722), .ZN(
        P1_U3158) );
  AOI22_X1 U23662 ( .A1(n20726), .A2(n20735), .B1(n20725), .B2(n20733), .ZN(
        n20730) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20739), .B1(
        n20728), .B2(n20727), .ZN(n20729) );
  OAI211_X1 U23664 ( .C1(n20732), .C2(n20731), .A(n20730), .B(n20729), .ZN(
        P1_U3159) );
  AOI22_X1 U23665 ( .A1(n20736), .A2(n20735), .B1(n20734), .B2(n20733), .ZN(
        n20741) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20739), .B1(
        n20738), .B2(n20737), .ZN(n20740) );
  OAI211_X1 U23667 ( .C1(n20743), .C2(n20742), .A(n20741), .B(n20740), .ZN(
        P1_U3160) );
  NOR2_X1 U23668 ( .A1(n9880), .A2(n11284), .ZN(n20746) );
  INV_X1 U23669 ( .A(n20744), .ZN(n20745) );
  OAI21_X1 U23670 ( .B1(n20746), .B2(n20260), .A(n20745), .ZN(P1_U3163) );
  AND2_X1 U23671 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20747), .ZN(
        P1_U3164) );
  AND2_X1 U23672 ( .A1(n20747), .A2(P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(
        P1_U3165) );
  AND2_X1 U23673 ( .A1(n20747), .A2(P1_DATAWIDTH_REG_29__SCAN_IN), .ZN(
        P1_U3166) );
  AND2_X1 U23674 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20747), .ZN(
        P1_U3167) );
  AND2_X1 U23675 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20747), .ZN(
        P1_U3168) );
  AND2_X1 U23676 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20747), .ZN(
        P1_U3169) );
  AND2_X1 U23677 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20747), .ZN(
        P1_U3170) );
  AND2_X1 U23678 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20747), .ZN(
        P1_U3171) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20747), .ZN(
        P1_U3172) );
  AND2_X1 U23680 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20747), .ZN(
        P1_U3173) );
  AND2_X1 U23681 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20747), .ZN(
        P1_U3174) );
  AND2_X1 U23682 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20747), .ZN(
        P1_U3175) );
  AND2_X1 U23683 ( .A1(n20747), .A2(P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(
        P1_U3176) );
  AND2_X1 U23684 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20747), .ZN(
        P1_U3177) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20747), .ZN(
        P1_U3178) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20747), .ZN(
        P1_U3179) );
  AND2_X1 U23687 ( .A1(n20747), .A2(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(
        P1_U3180) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20747), .ZN(
        P1_U3181) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20747), .ZN(
        P1_U3182) );
  AND2_X1 U23690 ( .A1(n20747), .A2(P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(
        P1_U3183) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20747), .ZN(
        P1_U3184) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20747), .ZN(
        P1_U3185) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20747), .ZN(P1_U3186) );
  AND2_X1 U23694 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20747), .ZN(P1_U3187) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20747), .ZN(P1_U3188) );
  AND2_X1 U23696 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20747), .ZN(P1_U3189) );
  AND2_X1 U23697 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20747), .ZN(P1_U3190) );
  AND2_X1 U23698 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20747), .ZN(P1_U3191) );
  AND2_X1 U23699 ( .A1(n20747), .A2(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(P1_U3192) );
  AND2_X1 U23700 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20747), .ZN(P1_U3193) );
  OAI21_X1 U23701 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20759), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20748) );
  AOI21_X1 U23702 ( .B1(HOLD), .B2(n20749), .A(n20748), .ZN(n20752) );
  AOI21_X1 U23703 ( .B1(n20756), .B2(n20762), .A(n20750), .ZN(n20751) );
  OAI21_X1 U23704 ( .B1(n20845), .B2(n20752), .A(n20751), .ZN(P1_U3194) );
  NOR2_X1 U23705 ( .A1(NA), .A2(n20848), .ZN(n20754) );
  OAI211_X1 U23706 ( .C1(n20754), .C2(n20753), .A(HOLD), .B(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20761) );
  NOR2_X1 U23707 ( .A1(NA), .A2(n20755), .ZN(n20758) );
  OAI222_X1 U23708 ( .A1(n20759), .A2(P1_STATE_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_2__SCAN_IN), .B2(n20758), .C1(n20757), .C2(n20756), .ZN(
        n20760) );
  OAI221_X1 U23709 ( .B1(n20761), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20761), .C2(n20762), .A(n20760), .ZN(P1_U3196) );
  OR2_X1 U23710 ( .A1(n20762), .A2(n20799), .ZN(n20786) );
  NAND2_X1 U23711 ( .A1(n20762), .A2(n20845), .ZN(n20784) );
  INV_X1 U23712 ( .A(n20784), .ZN(n20801) );
  AOI22_X1 U23713 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20799), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20801), .ZN(n20763) );
  OAI21_X1 U23714 ( .B1(n20836), .B2(n20786), .A(n20763), .ZN(P1_U3197) );
  INV_X1 U23715 ( .A(n20786), .ZN(n20802) );
  AOI22_X1 U23716 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20799), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20802), .ZN(n20764) );
  OAI21_X1 U23717 ( .B1(n20767), .B2(n20784), .A(n20764), .ZN(P1_U3198) );
  OAI222_X1 U23718 ( .A1(n20786), .A2(n20767), .B1(n20766), .B2(n20845), .C1(
        n20765), .C2(n20784), .ZN(P1_U3199) );
  AOI222_X1 U23719 ( .A1(n20801), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20802), .ZN(n20768) );
  INV_X1 U23720 ( .A(n20768), .ZN(P1_U3200) );
  AOI222_X1 U23721 ( .A1(n20802), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20801), .ZN(n20769) );
  INV_X1 U23722 ( .A(n20769), .ZN(P1_U3201) );
  AOI222_X1 U23723 ( .A1(n20802), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20801), .ZN(n20770) );
  INV_X1 U23724 ( .A(n20770), .ZN(P1_U3202) );
  AOI222_X1 U23725 ( .A1(n20802), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20801), .ZN(n20771) );
  INV_X1 U23726 ( .A(n20771), .ZN(P1_U3203) );
  AOI22_X1 U23727 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20799), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20801), .ZN(n20772) );
  OAI21_X1 U23728 ( .B1(n20773), .B2(n20786), .A(n20772), .ZN(P1_U3204) );
  AOI22_X1 U23729 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20799), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20802), .ZN(n20774) );
  OAI21_X1 U23730 ( .B1(n20775), .B2(n20784), .A(n20774), .ZN(P1_U3205) );
  AOI222_X1 U23731 ( .A1(n20801), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20802), .ZN(n20776) );
  INV_X1 U23732 ( .A(n20776), .ZN(P1_U3206) );
  AOI222_X1 U23733 ( .A1(n20802), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20801), .ZN(n20777) );
  INV_X1 U23734 ( .A(n20777), .ZN(P1_U3207) );
  AOI22_X1 U23735 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20799), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n20801), .ZN(n20778) );
  OAI21_X1 U23736 ( .B1(n20779), .B2(n20786), .A(n20778), .ZN(P1_U3208) );
  AOI22_X1 U23737 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20799), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n20802), .ZN(n20780) );
  OAI21_X1 U23738 ( .B1(n20781), .B2(n20784), .A(n20780), .ZN(P1_U3209) );
  AOI222_X1 U23739 ( .A1(n20801), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20802), .ZN(n20782) );
  INV_X1 U23740 ( .A(n20782), .ZN(P1_U3210) );
  AOI222_X1 U23741 ( .A1(n20802), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20801), .ZN(n20783) );
  INV_X1 U23742 ( .A(n20783), .ZN(P1_U3211) );
  INV_X1 U23743 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20947) );
  OAI222_X1 U23744 ( .A1(n20786), .A2(n20963), .B1(n20947), .B2(n20845), .C1(
        n20785), .C2(n20784), .ZN(P1_U3212) );
  AOI222_X1 U23745 ( .A1(n20802), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20801), .ZN(n20787) );
  INV_X1 U23746 ( .A(n20787), .ZN(P1_U3213) );
  AOI222_X1 U23747 ( .A1(n20802), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20801), .ZN(n20788) );
  INV_X1 U23748 ( .A(n20788), .ZN(P1_U3214) );
  AOI222_X1 U23749 ( .A1(n20801), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20802), .ZN(n20789) );
  INV_X1 U23750 ( .A(n20789), .ZN(P1_U3215) );
  AOI222_X1 U23751 ( .A1(n20802), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20801), .ZN(n20790) );
  INV_X1 U23752 ( .A(n20790), .ZN(P1_U3216) );
  AOI222_X1 U23753 ( .A1(n20802), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20801), .ZN(n20791) );
  INV_X1 U23754 ( .A(n20791), .ZN(P1_U3217) );
  AOI222_X1 U23755 ( .A1(n20802), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20801), .ZN(n20792) );
  INV_X1 U23756 ( .A(n20792), .ZN(P1_U3218) );
  AOI222_X1 U23757 ( .A1(n20801), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20802), .ZN(n20793) );
  INV_X1 U23758 ( .A(n20793), .ZN(P1_U3219) );
  AOI222_X1 U23759 ( .A1(n20802), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20801), .ZN(n20794) );
  INV_X1 U23760 ( .A(n20794), .ZN(P1_U3220) );
  AOI222_X1 U23761 ( .A1(n20802), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20801), .ZN(n20795) );
  INV_X1 U23762 ( .A(n20795), .ZN(P1_U3221) );
  AOI222_X1 U23763 ( .A1(n20802), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20801), .ZN(n20796) );
  INV_X1 U23764 ( .A(n20796), .ZN(P1_U3222) );
  AOI222_X1 U23765 ( .A1(n20802), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20801), .ZN(n20797) );
  INV_X1 U23766 ( .A(n20797), .ZN(P1_U3223) );
  AOI222_X1 U23767 ( .A1(n20802), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20801), .ZN(n20798) );
  INV_X1 U23768 ( .A(n20798), .ZN(P1_U3224) );
  AOI222_X1 U23769 ( .A1(n20801), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20802), .ZN(n20800) );
  INV_X1 U23770 ( .A(n20800), .ZN(P1_U3225) );
  AOI222_X1 U23771 ( .A1(n20802), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20799), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20801), .ZN(n20803) );
  INV_X1 U23772 ( .A(n20803), .ZN(P1_U3226) );
  OAI22_X1 U23773 ( .A1(n20799), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20845), .ZN(n20804) );
  INV_X1 U23774 ( .A(n20804), .ZN(P1_U3458) );
  OAI22_X1 U23775 ( .A1(n20799), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20845), .ZN(n20805) );
  INV_X1 U23776 ( .A(n20805), .ZN(P1_U3459) );
  OAI22_X1 U23777 ( .A1(n20799), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20845), .ZN(n20806) );
  INV_X1 U23778 ( .A(n20806), .ZN(P1_U3460) );
  OAI22_X1 U23779 ( .A1(n20799), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20845), .ZN(n20807) );
  INV_X1 U23780 ( .A(n20807), .ZN(P1_U3461) );
  OAI21_X1 U23781 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20811), .A(n20809), 
        .ZN(n20808) );
  INV_X1 U23782 ( .A(n20808), .ZN(P1_U3464) );
  OAI21_X1 U23783 ( .B1(n20811), .B2(n20810), .A(n20809), .ZN(P1_U3465) );
  INV_X1 U23784 ( .A(n20835), .ZN(n20826) );
  OAI211_X1 U23785 ( .C1(n20815), .C2(n20814), .A(n10607), .B(n20813), .ZN(
        n20823) );
  INV_X1 U23786 ( .A(n20828), .ZN(n20816) );
  NAND2_X1 U23787 ( .A1(n20817), .A2(n20816), .ZN(n20822) );
  OR2_X1 U23788 ( .A1(n20819), .A2(n20818), .ZN(n20820) );
  AND4_X1 U23789 ( .A1(n20823), .A2(n20822), .A3(n20821), .A4(n20820), .ZN(
        n20824) );
  AOI22_X1 U23790 ( .A1(n20826), .A2(n20825), .B1(n20824), .B2(n20835), .ZN(
        P1_U3475) );
  OAI22_X1 U23791 ( .A1(n20830), .A2(n20829), .B1(n20828), .B2(n20827), .ZN(
        n20831) );
  OAI21_X1 U23792 ( .B1(n20832), .B2(n20831), .A(n20835), .ZN(n20833) );
  OAI21_X1 U23793 ( .B1(n20835), .B2(n20834), .A(n20833), .ZN(P1_U3478) );
  AOI21_X1 U23794 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20837) );
  AOI22_X1 U23795 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20837), .B2(n20836), .ZN(n20840) );
  INV_X1 U23796 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20839) );
  AOI22_X1 U23797 ( .A1(n20843), .A2(n20840), .B1(n20839), .B2(n20838), .ZN(
        P1_U3481) );
  INV_X1 U23798 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20842) );
  OAI21_X1 U23799 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20843), .ZN(n20841) );
  OAI21_X1 U23800 ( .B1(n20843), .B2(n20842), .A(n20841), .ZN(P1_U3482) );
  AOI22_X1 U23801 ( .A1(n20845), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20844), 
        .B2(n20799), .ZN(P1_U3483) );
  AOI211_X1 U23802 ( .C1(n20849), .C2(n20848), .A(n20847), .B(n20846), .ZN(
        n20856) );
  OAI211_X1 U23803 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20851), .A(n20850), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20853) );
  AOI21_X1 U23804 ( .B1(n20853), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20852), 
        .ZN(n20855) );
  NAND2_X1 U23805 ( .A1(n20856), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20854) );
  OAI21_X1 U23806 ( .B1(n20856), .B2(n20855), .A(n20854), .ZN(P1_U3485) );
  MUX2_X1 U23807 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20799), .Z(P1_U3486) );
  INV_X1 U23808 ( .A(keyinput65), .ZN(n20858) );
  AOI22_X1 U23809 ( .A1(n20859), .A2(keyinput55), .B1(
        P3_DATAWIDTH_REG_1__SCAN_IN), .B2(n20858), .ZN(n20857) );
  OAI221_X1 U23810 ( .B1(n20859), .B2(keyinput55), .C1(n20858), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(n20857), .ZN(n20871) );
  AOI22_X1 U23811 ( .A1(n11837), .A2(keyinput59), .B1(keyinput50), .B2(n20861), 
        .ZN(n20860) );
  OAI221_X1 U23812 ( .B1(n11837), .B2(keyinput59), .C1(n20861), .C2(keyinput50), .A(n20860), .ZN(n20870) );
  INV_X1 U23813 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U23814 ( .A1(n20864), .A2(keyinput123), .B1(n20863), .B2(keyinput45), .ZN(n20862) );
  OAI221_X1 U23815 ( .B1(n20864), .B2(keyinput123), .C1(n20863), .C2(
        keyinput45), .A(n20862), .ZN(n20869) );
  INV_X1 U23816 ( .A(keyinput22), .ZN(n20865) );
  XOR2_X1 U23817 ( .A(P3_DATAWIDTH_REG_4__SCAN_IN), .B(n20865), .Z(n20867) );
  XNOR2_X1 U23818 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B(keyinput9), .ZN(
        n20866) );
  NAND2_X1 U23819 ( .A1(n20867), .A2(n20866), .ZN(n20868) );
  NOR4_X1 U23820 ( .A1(n20871), .A2(n20870), .A3(n20869), .A4(n20868), .ZN(
        n20922) );
  AOI22_X1 U23821 ( .A1(n20874), .A2(keyinput101), .B1(keyinput70), .B2(n20873), .ZN(n20872) );
  OAI221_X1 U23822 ( .B1(n20874), .B2(keyinput101), .C1(n20873), .C2(
        keyinput70), .A(n20872), .ZN(n20887) );
  INV_X1 U23823 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n20876) );
  AOI22_X1 U23824 ( .A1(n20877), .A2(keyinput99), .B1(keyinput127), .B2(n20876), .ZN(n20875) );
  OAI221_X1 U23825 ( .B1(n20877), .B2(keyinput99), .C1(n20876), .C2(
        keyinput127), .A(n20875), .ZN(n20886) );
  INV_X1 U23826 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n20880) );
  AOI22_X1 U23827 ( .A1(n20880), .A2(keyinput122), .B1(n20879), .B2(keyinput95), .ZN(n20878) );
  OAI221_X1 U23828 ( .B1(n20880), .B2(keyinput122), .C1(n20879), .C2(
        keyinput95), .A(n20878), .ZN(n20885) );
  INV_X1 U23829 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n20882) );
  AOI22_X1 U23830 ( .A1(n20883), .A2(keyinput84), .B1(n20882), .B2(keyinput114), .ZN(n20881) );
  OAI221_X1 U23831 ( .B1(n20883), .B2(keyinput84), .C1(n20882), .C2(
        keyinput114), .A(n20881), .ZN(n20884) );
  NOR4_X1 U23832 ( .A1(n20887), .A2(n20886), .A3(n20885), .A4(n20884), .ZN(
        n20921) );
  INV_X1 U23833 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U23834 ( .A1(n20890), .A2(keyinput30), .B1(n20889), .B2(keyinput87), 
        .ZN(n20888) );
  OAI221_X1 U23835 ( .B1(n20890), .B2(keyinput30), .C1(n20889), .C2(keyinput87), .A(n20888), .ZN(n20903) );
  INV_X1 U23836 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n20893) );
  INV_X1 U23837 ( .A(keyinput25), .ZN(n20892) );
  AOI22_X1 U23838 ( .A1(n20893), .A2(keyinput105), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n20892), .ZN(n20891) );
  OAI221_X1 U23839 ( .B1(n20893), .B2(keyinput105), .C1(n20892), .C2(
        P3_ADDRESS_REG_3__SCAN_IN), .A(n20891), .ZN(n20902) );
  INV_X1 U23840 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20896) );
  AOI22_X1 U23841 ( .A1(n20896), .A2(keyinput104), .B1(n20895), .B2(keyinput86), .ZN(n20894) );
  OAI221_X1 U23842 ( .B1(n20896), .B2(keyinput104), .C1(n20895), .C2(
        keyinput86), .A(n20894), .ZN(n20901) );
  INV_X1 U23843 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n20898) );
  AOI22_X1 U23844 ( .A1(n20899), .A2(keyinput125), .B1(keyinput11), .B2(n20898), .ZN(n20897) );
  OAI221_X1 U23845 ( .B1(n20899), .B2(keyinput125), .C1(n20898), .C2(
        keyinput11), .A(n20897), .ZN(n20900) );
  NOR4_X1 U23846 ( .A1(n20903), .A2(n20902), .A3(n20901), .A4(n20900), .ZN(
        n20920) );
  INV_X1 U23847 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20906) );
  INV_X1 U23848 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U23849 ( .A1(n20906), .A2(keyinput8), .B1(n20905), .B2(keyinput94), 
        .ZN(n20904) );
  OAI221_X1 U23850 ( .B1(n20906), .B2(keyinput8), .C1(n20905), .C2(keyinput94), 
        .A(n20904), .ZN(n20918) );
  AOI22_X1 U23851 ( .A1(n20909), .A2(keyinput0), .B1(n20908), .B2(keyinput14), 
        .ZN(n20907) );
  OAI221_X1 U23852 ( .B1(n20909), .B2(keyinput0), .C1(n20908), .C2(keyinput14), 
        .A(n20907), .ZN(n20917) );
  AOI22_X1 U23853 ( .A1(n20912), .A2(keyinput5), .B1(n20911), .B2(keyinput118), 
        .ZN(n20910) );
  OAI221_X1 U23854 ( .B1(n20912), .B2(keyinput5), .C1(n20911), .C2(keyinput118), .A(n20910), .ZN(n20916) );
  AOI22_X1 U23855 ( .A1(n20914), .A2(keyinput121), .B1(n12846), .B2(keyinput41), .ZN(n20913) );
  OAI221_X1 U23856 ( .B1(n20914), .B2(keyinput121), .C1(n12846), .C2(
        keyinput41), .A(n20913), .ZN(n20915) );
  NOR4_X1 U23857 ( .A1(n20918), .A2(n20917), .A3(n20916), .A4(n20915), .ZN(
        n20919) );
  NAND4_X1 U23858 ( .A1(n20922), .A2(n20921), .A3(n20920), .A4(n20919), .ZN(
        n21174) );
  INV_X1 U23859 ( .A(keyinput17), .ZN(n20924) );
  AOI22_X1 U23860 ( .A1(n20925), .A2(keyinput115), .B1(
        P3_ADDRESS_REG_23__SCAN_IN), .B2(n20924), .ZN(n20923) );
  OAI221_X1 U23861 ( .B1(n20925), .B2(keyinput115), .C1(n20924), .C2(
        P3_ADDRESS_REG_23__SCAN_IN), .A(n20923), .ZN(n20936) );
  INV_X1 U23862 ( .A(keyinput88), .ZN(n20927) );
  AOI22_X1 U23863 ( .A1(n20928), .A2(keyinput38), .B1(
        P3_DATAWIDTH_REG_7__SCAN_IN), .B2(n20927), .ZN(n20926) );
  OAI221_X1 U23864 ( .B1(n20928), .B2(keyinput38), .C1(n20927), .C2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A(n20926), .ZN(n20935) );
  INV_X1 U23865 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n20930) );
  AOI22_X1 U23866 ( .A1(n20930), .A2(keyinput26), .B1(n11465), .B2(keyinput80), 
        .ZN(n20929) );
  OAI221_X1 U23867 ( .B1(n20930), .B2(keyinput26), .C1(n11465), .C2(keyinput80), .A(n20929), .ZN(n20934) );
  AOI22_X1 U23868 ( .A1(n10101), .A2(keyinput77), .B1(n20932), .B2(keyinput56), 
        .ZN(n20931) );
  OAI221_X1 U23869 ( .B1(n10101), .B2(keyinput77), .C1(n20932), .C2(keyinput56), .A(n20931), .ZN(n20933) );
  NOR4_X1 U23870 ( .A1(n20936), .A2(n20935), .A3(n20934), .A4(n20933), .ZN(
        n20988) );
  INV_X1 U23871 ( .A(keyinput20), .ZN(n20938) );
  AOI22_X1 U23872 ( .A1(n20939), .A2(keyinput40), .B1(
        P2_DATAWIDTH_REG_25__SCAN_IN), .B2(n20938), .ZN(n20937) );
  OAI221_X1 U23873 ( .B1(n20939), .B2(keyinput40), .C1(n20938), .C2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A(n20937), .ZN(n20952) );
  AOI22_X1 U23874 ( .A1(n20942), .A2(keyinput24), .B1(keyinput93), .B2(n20941), 
        .ZN(n20940) );
  OAI221_X1 U23875 ( .B1(n20942), .B2(keyinput24), .C1(n20941), .C2(keyinput93), .A(n20940), .ZN(n20951) );
  INV_X1 U23876 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n20945) );
  AOI22_X1 U23877 ( .A1(n20945), .A2(keyinput66), .B1(n20944), .B2(keyinput52), 
        .ZN(n20943) );
  OAI221_X1 U23878 ( .B1(n20945), .B2(keyinput66), .C1(n20944), .C2(keyinput52), .A(n20943), .ZN(n20950) );
  AOI22_X1 U23879 ( .A1(n20948), .A2(keyinput43), .B1(keyinput67), .B2(n20947), 
        .ZN(n20946) );
  OAI221_X1 U23880 ( .B1(n20948), .B2(keyinput43), .C1(n20947), .C2(keyinput67), .A(n20946), .ZN(n20949) );
  NOR4_X1 U23881 ( .A1(n20952), .A2(n20951), .A3(n20950), .A4(n20949), .ZN(
        n20987) );
  AOI22_X1 U23882 ( .A1(n20955), .A2(keyinput90), .B1(keyinput3), .B2(n20954), 
        .ZN(n20953) );
  OAI221_X1 U23883 ( .B1(n20955), .B2(keyinput90), .C1(n20954), .C2(keyinput3), 
        .A(n20953), .ZN(n20968) );
  INV_X1 U23884 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n20958) );
  INV_X1 U23885 ( .A(keyinput57), .ZN(n20957) );
  AOI22_X1 U23886 ( .A1(n20958), .A2(keyinput119), .B1(
        P1_DATAWIDTH_REG_29__SCAN_IN), .B2(n20957), .ZN(n20956) );
  OAI221_X1 U23887 ( .B1(n20958), .B2(keyinput119), .C1(n20957), .C2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A(n20956), .ZN(n20967) );
  AOI22_X1 U23888 ( .A1(n20961), .A2(keyinput23), .B1(keyinput92), .B2(n20960), 
        .ZN(n20959) );
  OAI221_X1 U23889 ( .B1(n20961), .B2(keyinput23), .C1(n20960), .C2(keyinput92), .A(n20959), .ZN(n20966) );
  INV_X1 U23890 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n20964) );
  AOI22_X1 U23891 ( .A1(n20964), .A2(keyinput53), .B1(keyinput110), .B2(n20963), .ZN(n20962) );
  OAI221_X1 U23892 ( .B1(n20964), .B2(keyinput53), .C1(n20963), .C2(
        keyinput110), .A(n20962), .ZN(n20965) );
  NOR4_X1 U23893 ( .A1(n20968), .A2(n20967), .A3(n20966), .A4(n20965), .ZN(
        n20986) );
  AOI22_X1 U23894 ( .A1(n20971), .A2(keyinput72), .B1(n20970), .B2(keyinput36), 
        .ZN(n20969) );
  OAI221_X1 U23895 ( .B1(n20971), .B2(keyinput72), .C1(n20970), .C2(keyinput36), .A(n20969), .ZN(n20984) );
  INV_X1 U23896 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n20974) );
  AOI22_X1 U23897 ( .A1(n20974), .A2(keyinput27), .B1(n20973), .B2(keyinput46), 
        .ZN(n20972) );
  OAI221_X1 U23898 ( .B1(n20974), .B2(keyinput27), .C1(n20973), .C2(keyinput46), .A(n20972), .ZN(n20983) );
  INV_X1 U23899 ( .A(keyinput33), .ZN(n20976) );
  AOI22_X1 U23900 ( .A1(n20977), .A2(keyinput97), .B1(
        P1_DATAWIDTH_REG_19__SCAN_IN), .B2(n20976), .ZN(n20975) );
  OAI221_X1 U23901 ( .B1(n20977), .B2(keyinput97), .C1(n20976), .C2(
        P1_DATAWIDTH_REG_19__SCAN_IN), .A(n20975), .ZN(n20982) );
  INV_X1 U23902 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20980) );
  INV_X1 U23903 ( .A(keyinput10), .ZN(n20979) );
  AOI22_X1 U23904 ( .A1(n20980), .A2(keyinput82), .B1(P2_BE_N_REG_2__SCAN_IN), 
        .B2(n20979), .ZN(n20978) );
  OAI221_X1 U23905 ( .B1(n20980), .B2(keyinput82), .C1(n20979), .C2(
        P2_BE_N_REG_2__SCAN_IN), .A(n20978), .ZN(n20981) );
  NOR4_X1 U23906 ( .A1(n20984), .A2(n20983), .A3(n20982), .A4(n20981), .ZN(
        n20985) );
  NAND4_X1 U23907 ( .A1(n20988), .A2(n20987), .A3(n20986), .A4(n20985), .ZN(
        n21173) );
  INV_X1 U23908 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U23909 ( .A1(n11835), .A2(keyinput39), .B1(keyinput44), .B2(n20990), 
        .ZN(n20989) );
  OAI221_X1 U23910 ( .B1(n11835), .B2(keyinput39), .C1(n20990), .C2(keyinput44), .A(n20989), .ZN(n21002) );
  AOI22_X1 U23911 ( .A1(n20992), .A2(keyinput7), .B1(n10613), .B2(keyinput69), 
        .ZN(n20991) );
  OAI221_X1 U23912 ( .B1(n20992), .B2(keyinput7), .C1(n10613), .C2(keyinput69), 
        .A(n20991), .ZN(n21001) );
  INV_X1 U23913 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20994) );
  AOI22_X1 U23914 ( .A1(n20995), .A2(keyinput81), .B1(n20994), .B2(keyinput16), 
        .ZN(n20993) );
  OAI221_X1 U23915 ( .B1(n20995), .B2(keyinput81), .C1(n20994), .C2(keyinput16), .A(n20993), .ZN(n21000) );
  INV_X1 U23916 ( .A(keyinput58), .ZN(n20997) );
  AOI22_X1 U23917 ( .A1(n20998), .A2(keyinput71), .B1(P3_DATAO_REG_20__SCAN_IN), .B2(n20997), .ZN(n20996) );
  OAI221_X1 U23918 ( .B1(n20998), .B2(keyinput71), .C1(n20997), .C2(
        P3_DATAO_REG_20__SCAN_IN), .A(n20996), .ZN(n20999) );
  NOR4_X1 U23919 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21051) );
  INV_X1 U23920 ( .A(keyinput28), .ZN(n21004) );
  AOI22_X1 U23921 ( .A1(n21005), .A2(keyinput109), .B1(
        P2_DATAWIDTH_REG_17__SCAN_IN), .B2(n21004), .ZN(n21003) );
  OAI221_X1 U23922 ( .B1(n21005), .B2(keyinput109), .C1(n21004), .C2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A(n21003), .ZN(n21018) );
  AOI22_X1 U23923 ( .A1(n21008), .A2(keyinput32), .B1(n21007), .B2(keyinput37), 
        .ZN(n21006) );
  OAI221_X1 U23924 ( .B1(n21008), .B2(keyinput32), .C1(n21007), .C2(keyinput37), .A(n21006), .ZN(n21017) );
  AOI22_X1 U23925 ( .A1(n21011), .A2(keyinput31), .B1(n21010), .B2(keyinput124), .ZN(n21009) );
  OAI221_X1 U23926 ( .B1(n21011), .B2(keyinput31), .C1(n21010), .C2(
        keyinput124), .A(n21009), .ZN(n21016) );
  AOI22_X1 U23927 ( .A1(n21014), .A2(keyinput60), .B1(keyinput85), .B2(n21013), 
        .ZN(n21012) );
  OAI221_X1 U23928 ( .B1(n21014), .B2(keyinput60), .C1(n21013), .C2(keyinput85), .A(n21012), .ZN(n21015) );
  NOR4_X1 U23929 ( .A1(n21018), .A2(n21017), .A3(n21016), .A4(n21015), .ZN(
        n21050) );
  INV_X1 U23930 ( .A(keyinput126), .ZN(n21021) );
  INV_X1 U23931 ( .A(keyinput111), .ZN(n21020) );
  AOI22_X1 U23932 ( .A1(n21021), .A2(P1_DATAWIDTH_REG_12__SCAN_IN), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n21020), .ZN(n21019) );
  OAI221_X1 U23933 ( .B1(n21021), .B2(P1_DATAWIDTH_REG_12__SCAN_IN), .C1(
        n21020), .C2(P3_ADDRESS_REG_4__SCAN_IN), .A(n21019), .ZN(n21032) );
  INV_X1 U23934 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n21023) );
  AOI22_X1 U23935 ( .A1(n21023), .A2(keyinput98), .B1(keyinput1), .B2(n11105), 
        .ZN(n21022) );
  OAI221_X1 U23936 ( .B1(n21023), .B2(keyinput98), .C1(n11105), .C2(keyinput1), 
        .A(n21022), .ZN(n21031) );
  AOI22_X1 U23937 ( .A1(n21025), .A2(keyinput78), .B1(n11986), .B2(keyinput107), .ZN(n21024) );
  OAI221_X1 U23938 ( .B1(n21025), .B2(keyinput78), .C1(n11986), .C2(
        keyinput107), .A(n21024), .ZN(n21030) );
  INV_X1 U23939 ( .A(keyinput29), .ZN(n21026) );
  XOR2_X1 U23940 ( .A(P1_DATAWIDTH_REG_30__SCAN_IN), .B(n21026), .Z(n21028) );
  XNOR2_X1 U23941 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B(keyinput49), .ZN(
        n21027) );
  NAND2_X1 U23942 ( .A1(n21028), .A2(n21027), .ZN(n21029) );
  NOR4_X1 U23943 ( .A1(n21032), .A2(n21031), .A3(n21030), .A4(n21029), .ZN(
        n21049) );
  INV_X1 U23944 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n21035) );
  INV_X1 U23945 ( .A(keyinput12), .ZN(n21034) );
  AOI22_X1 U23946 ( .A1(n21035), .A2(keyinput47), .B1(
        P1_DATAWIDTH_REG_3__SCAN_IN), .B2(n21034), .ZN(n21033) );
  OAI221_X1 U23947 ( .B1(n21035), .B2(keyinput47), .C1(n21034), .C2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A(n21033), .ZN(n21047) );
  AOI22_X1 U23948 ( .A1(n21038), .A2(keyinput96), .B1(keyinput48), .B2(n21037), 
        .ZN(n21036) );
  OAI221_X1 U23949 ( .B1(n21038), .B2(keyinput96), .C1(n21037), .C2(keyinput48), .A(n21036), .ZN(n21046) );
  INV_X1 U23950 ( .A(keyinput102), .ZN(n21041) );
  INV_X1 U23951 ( .A(keyinput117), .ZN(n21040) );
  AOI22_X1 U23952 ( .A1(n21041), .A2(P3_DATAWIDTH_REG_26__SCAN_IN), .B1(
        P2_DATAWIDTH_REG_23__SCAN_IN), .B2(n21040), .ZN(n21039) );
  OAI221_X1 U23953 ( .B1(n21041), .B2(P3_DATAWIDTH_REG_26__SCAN_IN), .C1(
        n21040), .C2(P2_DATAWIDTH_REG_23__SCAN_IN), .A(n21039), .ZN(n21045) );
  XNOR2_X1 U23954 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B(keyinput120), .ZN(
        n21043) );
  XNOR2_X1 U23955 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B(keyinput100), .ZN(
        n21042) );
  NAND2_X1 U23956 ( .A1(n21043), .A2(n21042), .ZN(n21044) );
  NOR4_X1 U23957 ( .A1(n21047), .A2(n21046), .A3(n21045), .A4(n21044), .ZN(
        n21048) );
  NAND4_X1 U23958 ( .A1(n21051), .A2(n21050), .A3(n21049), .A4(n21048), .ZN(
        n21172) );
  NOR4_X1 U23959 ( .A1(keyinput105), .A2(keyinput121), .A3(keyinput125), .A4(
        keyinput8), .ZN(n21062) );
  NOR4_X1 U23960 ( .A1(keyinput61), .A2(keyinput65), .A3(keyinput89), .A4(
        keyinput101), .ZN(n21061) );
  INV_X1 U23961 ( .A(keyinput9), .ZN(n21052) );
  NOR4_X1 U23962 ( .A1(keyinput70), .A2(keyinput91), .A3(keyinput87), .A4(
        n21052), .ZN(n21053) );
  NAND3_X1 U23963 ( .A1(keyinput13), .A2(keyinput21), .A3(n21053), .ZN(n21059)
         );
  NOR4_X1 U23964 ( .A1(keyinput34), .A2(keyinput51), .A3(keyinput55), .A4(
        keyinput54), .ZN(n21057) );
  NOR4_X1 U23965 ( .A1(keyinput68), .A2(keyinput116), .A3(keyinput112), .A4(
        keyinput64), .ZN(n21056) );
  NOR4_X1 U23966 ( .A1(keyinput18), .A2(keyinput99), .A3(keyinput103), .A4(
        keyinput122), .ZN(n21055) );
  NOR4_X1 U23967 ( .A1(keyinput42), .A2(keyinput15), .A3(keyinput6), .A4(
        keyinput30), .ZN(n21054) );
  NAND4_X1 U23968 ( .A1(n21057), .A2(n21056), .A3(n21055), .A4(n21054), .ZN(
        n21058) );
  NOR4_X1 U23969 ( .A1(keyinput127), .A2(keyinput123), .A3(n21059), .A4(n21058), .ZN(n21060) );
  NAND3_X1 U23970 ( .A1(n21062), .A2(n21061), .A3(n21060), .ZN(n21170) );
  NOR4_X1 U23971 ( .A1(keyinput126), .A2(keyinput111), .A3(keyinput98), .A4(
        keyinput1), .ZN(n21063) );
  NAND3_X1 U23972 ( .A1(keyinput78), .A2(keyinput107), .A3(n21063), .ZN(n21076) );
  NOR2_X1 U23973 ( .A1(keyinput60), .A2(keyinput124), .ZN(n21064) );
  NAND3_X1 U23974 ( .A1(keyinput85), .A2(keyinput31), .A3(n21064), .ZN(n21065)
         );
  NOR3_X1 U23975 ( .A1(keyinput32), .A2(keyinput37), .A3(n21065), .ZN(n21074)
         );
  NOR3_X1 U23976 ( .A1(keyinput58), .A2(keyinput16), .A3(keyinput81), .ZN(
        n21066) );
  NAND2_X1 U23977 ( .A1(keyinput71), .A2(n21066), .ZN(n21072) );
  INV_X1 U23978 ( .A(keyinput7), .ZN(n21067) );
  NAND4_X1 U23979 ( .A1(keyinput69), .A2(keyinput39), .A3(keyinput44), .A4(
        n21067), .ZN(n21071) );
  NAND4_X1 U23980 ( .A1(keyinput96), .A2(keyinput48), .A3(keyinput12), .A4(
        keyinput47), .ZN(n21070) );
  NOR2_X1 U23981 ( .A1(keyinput102), .A2(keyinput100), .ZN(n21068) );
  NAND3_X1 U23982 ( .A1(keyinput117), .A2(keyinput120), .A3(n21068), .ZN(
        n21069) );
  NOR4_X1 U23983 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n21069), .ZN(
        n21073) );
  NAND4_X1 U23984 ( .A1(keyinput109), .A2(keyinput28), .A3(n21074), .A4(n21073), .ZN(n21075) );
  NOR4_X1 U23985 ( .A1(keyinput29), .A2(keyinput49), .A3(n21076), .A4(n21075), 
        .ZN(n21102) );
  NAND2_X1 U23986 ( .A1(keyinput26), .A2(keyinput115), .ZN(n21077) );
  NOR3_X1 U23987 ( .A1(keyinput17), .A2(keyinput80), .A3(n21077), .ZN(n21078)
         );
  NAND3_X1 U23988 ( .A1(keyinput77), .A2(keyinput56), .A3(n21078), .ZN(n21090)
         );
  NOR2_X1 U23989 ( .A1(keyinput119), .A2(keyinput23), .ZN(n21079) );
  NAND3_X1 U23990 ( .A1(keyinput57), .A2(keyinput92), .A3(n21079), .ZN(n21080)
         );
  NOR3_X1 U23991 ( .A1(keyinput90), .A2(keyinput3), .A3(n21080), .ZN(n21088)
         );
  NOR3_X1 U23992 ( .A1(keyinput66), .A2(keyinput52), .A3(keyinput67), .ZN(
        n21081) );
  NAND2_X1 U23993 ( .A1(keyinput43), .A2(n21081), .ZN(n21086) );
  NAND4_X1 U23994 ( .A1(keyinput24), .A2(keyinput93), .A3(keyinput20), .A4(
        keyinput40), .ZN(n21085) );
  NOR2_X1 U23995 ( .A1(keyinput10), .A2(keyinput97), .ZN(n21082) );
  NAND3_X1 U23996 ( .A1(keyinput82), .A2(keyinput33), .A3(n21082), .ZN(n21084)
         );
  NAND4_X1 U23997 ( .A1(keyinput27), .A2(keyinput46), .A3(keyinput72), .A4(
        keyinput36), .ZN(n21083) );
  NOR4_X1 U23998 ( .A1(n21086), .A2(n21085), .A3(n21084), .A4(n21083), .ZN(
        n21087) );
  NAND4_X1 U23999 ( .A1(keyinput53), .A2(keyinput110), .A3(n21088), .A4(n21087), .ZN(n21089) );
  NOR4_X1 U24000 ( .A1(keyinput88), .A2(keyinput38), .A3(n21090), .A4(n21089), 
        .ZN(n21101) );
  NAND4_X1 U24001 ( .A1(keyinput22), .A2(keyinput19), .A3(keyinput106), .A4(
        keyinput118), .ZN(n21094) );
  NAND4_X1 U24002 ( .A1(keyinput50), .A2(keyinput14), .A3(keyinput11), .A4(
        keyinput2), .ZN(n21093) );
  NAND4_X1 U24003 ( .A1(keyinput95), .A2(keyinput83), .A3(keyinput94), .A4(
        keyinput86), .ZN(n21092) );
  NAND4_X1 U24004 ( .A1(keyinput114), .A2(keyinput74), .A3(keyinput75), .A4(
        keyinput79), .ZN(n21091) );
  NOR4_X1 U24005 ( .A1(n21094), .A2(n21093), .A3(n21092), .A4(n21091), .ZN(
        n21100) );
  NAND4_X1 U24006 ( .A1(keyinput73), .A2(keyinput113), .A3(keyinput4), .A4(
        keyinput76), .ZN(n21098) );
  NAND4_X1 U24007 ( .A1(keyinput5), .A2(keyinput25), .A3(keyinput45), .A4(
        keyinput41), .ZN(n21097) );
  NAND4_X1 U24008 ( .A1(keyinput0), .A2(keyinput62), .A3(keyinput63), .A4(
        keyinput35), .ZN(n21096) );
  NAND4_X1 U24009 ( .A1(keyinput84), .A2(keyinput104), .A3(keyinput108), .A4(
        keyinput59), .ZN(n21095) );
  NOR4_X1 U24010 ( .A1(n21098), .A2(n21097), .A3(n21096), .A4(n21095), .ZN(
        n21099) );
  NAND4_X1 U24011 ( .A1(n21102), .A2(n21101), .A3(n21100), .A4(n21099), .ZN(
        n21169) );
  INV_X1 U24012 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n21104) );
  AOI22_X1 U24013 ( .A1(n10708), .A2(keyinput64), .B1(n21104), .B2(keyinput18), 
        .ZN(n21103) );
  OAI221_X1 U24014 ( .B1(n10708), .B2(keyinput64), .C1(n21104), .C2(keyinput18), .A(n21103), .ZN(n21117) );
  INV_X1 U24015 ( .A(keyinput34), .ZN(n21106) );
  AOI22_X1 U24016 ( .A1(n21107), .A2(keyinput6), .B1(
        P3_DATAWIDTH_REG_13__SCAN_IN), .B2(n21106), .ZN(n21105) );
  OAI221_X1 U24017 ( .B1(n21107), .B2(keyinput6), .C1(n21106), .C2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A(n21105), .ZN(n21116) );
  AOI22_X1 U24018 ( .A1(n21110), .A2(keyinput42), .B1(n21109), .B2(keyinput108), .ZN(n21108) );
  OAI221_X1 U24019 ( .B1(n21110), .B2(keyinput42), .C1(n21109), .C2(
        keyinput108), .A(n21108), .ZN(n21115) );
  AOI22_X1 U24020 ( .A1(n21113), .A2(keyinput68), .B1(n21112), .B2(keyinput113), .ZN(n21111) );
  OAI221_X1 U24021 ( .B1(n21113), .B2(keyinput68), .C1(n21112), .C2(
        keyinput113), .A(n21111), .ZN(n21114) );
  NOR4_X1 U24022 ( .A1(n21117), .A2(n21116), .A3(n21115), .A4(n21114), .ZN(
        n21168) );
  OAI22_X1 U24023 ( .A1(n21120), .A2(keyinput73), .B1(n21119), .B2(keyinput62), 
        .ZN(n21118) );
  AOI221_X1 U24024 ( .B1(n21120), .B2(keyinput73), .C1(keyinput62), .C2(n21119), .A(n21118), .ZN(n21133) );
  INV_X1 U24025 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21123) );
  INV_X1 U24026 ( .A(keyinput103), .ZN(n21122) );
  OAI22_X1 U24027 ( .A1(n21123), .A2(keyinput19), .B1(n21122), .B2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21121) );
  AOI221_X1 U24028 ( .B1(n21123), .B2(keyinput19), .C1(
        P1_DATAWIDTH_REG_15__SCAN_IN), .C2(n21122), .A(n21121), .ZN(n21132) );
  INV_X1 U24029 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n21126) );
  OAI22_X1 U24030 ( .A1(n21126), .A2(keyinput112), .B1(n21125), .B2(keyinput91), .ZN(n21124) );
  AOI221_X1 U24031 ( .B1(n21126), .B2(keyinput112), .C1(keyinput91), .C2(
        n21125), .A(n21124), .ZN(n21131) );
  INV_X1 U24032 ( .A(keyinput13), .ZN(n21128) );
  OAI22_X1 U24033 ( .A1(n21129), .A2(keyinput76), .B1(n21128), .B2(
        P3_DATAO_REG_28__SCAN_IN), .ZN(n21127) );
  AOI221_X1 U24034 ( .B1(n21129), .B2(keyinput76), .C1(
        P3_DATAO_REG_28__SCAN_IN), .C2(n21128), .A(n21127), .ZN(n21130) );
  NAND4_X1 U24035 ( .A1(n21133), .A2(n21132), .A3(n21131), .A4(n21130), .ZN(
        n21166) );
  INV_X1 U24036 ( .A(P3_LWORD_REG_9__SCAN_IN), .ZN(n21136) );
  AOI22_X1 U24037 ( .A1(n21136), .A2(keyinput75), .B1(n21135), .B2(keyinput83), 
        .ZN(n21134) );
  OAI221_X1 U24038 ( .B1(n21136), .B2(keyinput75), .C1(n21135), .C2(keyinput83), .A(n21134), .ZN(n21165) );
  INV_X1 U24039 ( .A(keyinput106), .ZN(n21138) );
  OAI22_X1 U24040 ( .A1(n21139), .A2(keyinput54), .B1(n21138), .B2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21137) );
  AOI221_X1 U24041 ( .B1(n21139), .B2(keyinput54), .C1(
        P2_DATAWIDTH_REG_12__SCAN_IN), .C2(n21138), .A(n21137), .ZN(n21147) );
  INV_X1 U24042 ( .A(P3_LWORD_REG_3__SCAN_IN), .ZN(n21142) );
  INV_X1 U24043 ( .A(keyinput35), .ZN(n21141) );
  OAI22_X1 U24044 ( .A1(n21142), .A2(keyinput2), .B1(n21141), .B2(
        P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21140) );
  AOI221_X1 U24045 ( .B1(n21142), .B2(keyinput2), .C1(
        P2_BYTEENABLE_REG_3__SCAN_IN), .C2(n21141), .A(n21140), .ZN(n21146) );
  OAI22_X1 U24046 ( .A1(n21144), .A2(keyinput89), .B1(n11288), .B2(keyinput63), 
        .ZN(n21143) );
  AOI221_X1 U24047 ( .B1(n21144), .B2(keyinput89), .C1(keyinput63), .C2(n11288), .A(n21143), .ZN(n21145) );
  NAND3_X1 U24048 ( .A1(n21147), .A2(n21146), .A3(n21145), .ZN(n21164) );
  INV_X1 U24049 ( .A(keyinput79), .ZN(n21149) );
  OAI22_X1 U24050 ( .A1(n12548), .A2(keyinput4), .B1(n21149), .B2(
        P3_ADDRESS_REG_0__SCAN_IN), .ZN(n21148) );
  AOI221_X1 U24051 ( .B1(n12548), .B2(keyinput4), .C1(
        P3_ADDRESS_REG_0__SCAN_IN), .C2(n21149), .A(n21148), .ZN(n21162) );
  INV_X1 U24052 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n21151) );
  OAI22_X1 U24053 ( .A1(n21152), .A2(keyinput15), .B1(n21151), .B2(keyinput74), 
        .ZN(n21150) );
  AOI221_X1 U24054 ( .B1(n21152), .B2(keyinput15), .C1(keyinput74), .C2(n21151), .A(n21150), .ZN(n21161) );
  OAI22_X1 U24055 ( .A1(n21155), .A2(keyinput116), .B1(n21154), .B2(keyinput51), .ZN(n21153) );
  AOI221_X1 U24056 ( .B1(n21155), .B2(keyinput116), .C1(keyinput51), .C2(
        n21154), .A(n21153), .ZN(n21160) );
  INV_X1 U24057 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n21157) );
  OAI22_X1 U24058 ( .A1(n21158), .A2(keyinput61), .B1(n21157), .B2(keyinput21), 
        .ZN(n21156) );
  AOI221_X1 U24059 ( .B1(n21158), .B2(keyinput61), .C1(keyinput21), .C2(n21157), .A(n21156), .ZN(n21159) );
  NAND4_X1 U24060 ( .A1(n21162), .A2(n21161), .A3(n21160), .A4(n21159), .ZN(
        n21163) );
  NOR4_X1 U24061 ( .A1(n21166), .A2(n21165), .A3(n21164), .A4(n21163), .ZN(
        n21167) );
  OAI211_X1 U24062 ( .C1(n21170), .C2(n21169), .A(n21168), .B(n21167), .ZN(
        n21171) );
  NOR4_X1 U24063 ( .A1(n21174), .A2(n21173), .A3(n21172), .A4(n21171), .ZN(
        n21176) );
  AOI22_X1 U24064 ( .A1(n16642), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(U215), .ZN(n21175) );
  XNOR2_X1 U24065 ( .A(n21176), .B(n21175), .ZN(U276) );
  INV_X1 U11197 ( .A(n14281), .ZN(n20207) );
  NAND2_X1 U11186 ( .A1(n10287), .A2(n10285), .ZN(n11195) );
  NAND2_X1 U11224 ( .A1(n14281), .A2(n20199), .ZN(n10435) );
  AND2_X2 U11244 ( .A1(n11538), .A2(n11795), .ZN(n12902) );
  CLKBUF_X1 U11246 ( .A(n10426), .Z(n12998) );
  CLKBUF_X1 U11252 ( .A(n11845), .Z(n13176) );
  NOR2_X1 U11253 ( .A1(n9780), .A2(n14011), .ZN(n12592) );
  CLKBUF_X2 U11260 ( .A(n17914), .Z(n9734) );
  INV_X1 U11262 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13370) );
  XNOR2_X1 U11539 ( .A(n12592), .B(n12591), .ZN(n14714) );
  NAND2_X4 U12240 ( .A1(n11789), .A2(n11772), .ZN(n21178) );
  INV_X1 U12431 ( .A(n15494), .ZN(n9735) );
  CLKBUF_X1 U12491 ( .A(n17544), .Z(n17584) );
  CLKBUF_X1 U12591 ( .A(n20093), .Z(n20849) );
endmodule

