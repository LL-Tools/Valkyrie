

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7362, n7363, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16567;

  OR2_X1 U7462 ( .A1(n15293), .A2(n9544), .ZN(n15284) );
  OAI21_X1 U7463 ( .B1(n12862), .B2(n7677), .A(n7674), .ZN(n14860) );
  INV_X1 U7464 ( .A(n14955), .ZN(n15003) );
  INV_X1 U7465 ( .A(n9746), .ZN(n9964) );
  BUF_X2 U7466 ( .A(n12021), .Z(n7370) );
  INV_X1 U7467 ( .A(n16360), .ZN(n12086) );
  BUF_X2 U7468 ( .A(n9107), .Z(n9530) );
  INV_X1 U7469 ( .A(n9386), .ZN(n9504) );
  AND2_X1 U7471 ( .A1(n7538), .A2(n9015), .ZN(n9050) );
  NAND2_X1 U7473 ( .A1(n7629), .A2(n7846), .ZN(n8591) );
  INV_X1 U7475 ( .A(n16567), .ZN(n7362) );
  NOR2_X1 U7476 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8658) );
  INV_X2 U7477 ( .A(n9530), .ZN(n9529) );
  NAND2_X1 U7478 ( .A1(n11308), .A2(n16130), .ZN(n13137) );
  NOR2_X1 U7479 ( .A1(n7515), .A2(n8821), .ZN(n8665) );
  INV_X1 U7480 ( .A(n9481), .ZN(n9512) );
  OAI21_X1 U7481 ( .B1(n9038), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9040) );
  INV_X1 U7482 ( .A(n13334), .ZN(n8565) );
  INV_X2 U7485 ( .A(n16261), .ZN(n14491) );
  INV_X2 U7486 ( .A(n15001), .ZN(n14925) );
  OR2_X1 U7487 ( .A1(n15484), .A2(n15365), .ZN(n15349) );
  OAI21_X1 U7488 ( .B1(n9196), .B2(n9030), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9041) );
  AND4_X1 U7489 ( .A1(n9735), .A2(n9734), .A3(n9733), .A4(n9732), .ZN(n12293)
         );
  INV_X2 U7490 ( .A(n8591), .ZN(n10976) );
  OAI21_X1 U7491 ( .B1(n14333), .B2(n14332), .A(n14390), .ZN(n14383) );
  NAND2_X1 U7492 ( .A1(n8859), .A2(n8858), .ZN(n14677) );
  AND4_X1 U7493 ( .A1(n9105), .A2(n9104), .A3(n9103), .A4(n9102), .ZN(n12048)
         );
  NAND2_X1 U7494 ( .A1(n9462), .A2(n9461), .ZN(n15274) );
  XNOR2_X1 U7495 ( .A(n9012), .B(n9008), .ZN(n9014) );
  NOR2_X1 U7496 ( .A1(n9082), .A2(n7710), .ZN(n11386) );
  XNOR2_X1 U7497 ( .A(n10046), .B(n10045), .ZN(n11774) );
  INV_X1 U7498 ( .A(n10259), .ZN(n13091) );
  INV_X1 U7499 ( .A(n15311), .ZN(n12559) );
  XNOR2_X1 U7500 ( .A(n15783), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15785) );
  NOR2_X2 U7502 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8346) );
  INV_X2 U7503 ( .A(n8674), .ZN(n8673) );
  OR2_X2 U7504 ( .A1(n10632), .A2(n10631), .ZN(n7448) );
  AND2_X1 U7506 ( .A1(n9044), .A2(n9045), .ZN(n8299) );
  OAI21_X2 U7507 ( .B1(n8733), .B2(n8732), .A(n8625), .ZN(n8726) );
  XNOR2_X2 U7508 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n15734) );
  AND2_X2 U7509 ( .A1(n13091), .A2(n10258), .ZN(n10296) );
  XNOR2_X1 U7510 ( .A(n9041), .B(P1_IR_REG_19__SCAN_IN), .ZN(n15311) );
  INV_X2 U7512 ( .A(n9781), .ZN(n10032) );
  OR2_X2 U7513 ( .A1(n14037), .A2(n14038), .ZN(n14039) );
  INV_X4 U7514 ( .A(n9122), .ZN(n9456) );
  AOI21_X2 U7515 ( .B1(n7540), .B2(n16488), .A(n7539), .ZN(n15434) );
  OAI22_X2 U7516 ( .A1(n12198), .A2(n12196), .B1(n12026), .B2(n12206), .ZN(
        n12216) );
  NAND3_X2 U7517 ( .A1(n13977), .A2(n14030), .A3(n13257), .ZN(n13125) );
  NOR2_X2 U7518 ( .A1(n13124), .A2(n13123), .ZN(n13257) );
  OR2_X2 U7519 ( .A1(n15550), .A2(n9608), .ZN(n11496) );
  OAI21_X2 U7520 ( .B1(n14103), .B2(n13299), .A(n13300), .ZN(n14099) );
  NAND2_X2 U7521 ( .A1(n10079), .A2(n13129), .ZN(n14103) );
  INV_X1 U7522 ( .A(n9059), .ZN(n9358) );
  XNOR2_X2 U7523 ( .A(n15748), .B(n8038), .ZN(n15750) );
  NAND2_X2 U7524 ( .A1(n7524), .A2(n15742), .ZN(n15748) );
  AOI21_X2 U7525 ( .B1(n16061), .B2(n13935), .A(n13934), .ZN(n13937) );
  INV_X4 U7526 ( .A(n9335), .ZN(n7366) );
  XNOR2_X2 U7527 ( .A(n15758), .B(n15759), .ZN(n15763) );
  XNOR2_X2 U7528 ( .A(n15757), .B(n8036), .ZN(n15759) );
  NAND2_X2 U7530 ( .A1(n9598), .A2(n15689), .ZN(n9059) );
  NAND2_X2 U7531 ( .A1(n7523), .A2(n15892), .ZN(n15783) );
  INV_X2 U7533 ( .A(n9011), .ZN(n9009) );
  OAI21_X2 U7534 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(n11864), .A(n9654), .ZN(
        n9867) );
  XNOR2_X2 U7535 ( .A(n8954), .B(P2_IR_REG_29__SCAN_IN), .ZN(n10258) );
  XNOR2_X2 U7536 ( .A(n15824), .B(n15823), .ZN(n15825) );
  NAND2_X2 U7537 ( .A1(n15818), .A2(n7532), .ZN(n15824) );
  NAND2_X1 U7538 ( .A1(n14023), .A2(n8245), .ZN(n14006) );
  OR2_X1 U7539 ( .A1(n14255), .A2(n14010), .ZN(n13246) );
  OAI22_X1 U7540 ( .A1(n8861), .A2(n8860), .B1(SI_17_), .B2(n8632), .ZN(n8633)
         );
  CLKBUF_X2 U7541 ( .A(n10129), .Z(n10191) );
  AND2_X1 U7542 ( .A1(n13157), .A2(n13158), .ZN(n13306) );
  INV_X2 U7543 ( .A(n10122), .ZN(n11308) );
  XNOR2_X1 U7544 ( .A(n13472), .B(n16333), .ZN(n13164) );
  INV_X2 U7545 ( .A(n12136), .ZN(n16179) );
  INV_X1 U7546 ( .A(n14471), .ZN(n11695) );
  INV_X4 U7547 ( .A(n11987), .ZN(n7367) );
  NAND2_X1 U7548 ( .A1(n9488), .A2(n12559), .ZN(n11580) );
  AND2_X1 U7549 ( .A1(n8950), .A2(n8949), .ZN(n12739) );
  XNOR2_X1 U7550 ( .A(n8943), .B(n8942), .ZN(n12877) );
  NAND2_X1 U7551 ( .A1(n10984), .A2(P1_U3086), .ZN(n15558) );
  INV_X2 U7552 ( .A(n10976), .ZN(n10983) );
  NAND2_X1 U7553 ( .A1(n8364), .A2(n7440), .ZN(n9614) );
  BUF_X1 U7554 ( .A(n9098), .Z(n7537) );
  NOR2_X1 U7555 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8997) );
  OAI21_X1 U7556 ( .B1(n14500), .B2(n14499), .A(n14498), .ZN(n14693) );
  NAND2_X1 U7557 ( .A1(n7849), .A2(n7847), .ZN(n14528) );
  OAI21_X1 U7558 ( .B1(n14934), .B2(n7683), .A(n7680), .ZN(n15028) );
  NAND2_X1 U7559 ( .A1(n14015), .A2(n14014), .ZN(n14017) );
  NAND3_X1 U7560 ( .A1(n7610), .A2(n7608), .A3(n14397), .ZN(n14409) );
  NAND2_X1 U7561 ( .A1(n8032), .A2(n15877), .ZN(n15880) );
  NAND2_X1 U7562 ( .A1(n9444), .A2(n9443), .ZN(n9544) );
  NAND2_X1 U7563 ( .A1(n13987), .A2(n13999), .ZN(n13250) );
  NAND2_X1 U7564 ( .A1(n14039), .A2(n9965), .ZN(n14025) );
  NAND2_X1 U7565 ( .A1(n9983), .A2(n9982), .ZN(n14260) );
  OAI21_X1 U7566 ( .B1(n10534), .B2(n7865), .A(n7864), .ZN(n12934) );
  NAND2_X1 U7567 ( .A1(n9943), .A2(n10183), .ZN(n14058) );
  NAND2_X1 U7568 ( .A1(n12579), .A2(n12578), .ZN(n12675) );
  AOI21_X1 U7569 ( .B1(n9979), .B2(n9670), .A(n9669), .ZN(n9994) );
  NAND2_X1 U7570 ( .A1(n8712), .A2(n8711), .ZN(n14645) );
  OAI21_X1 U7571 ( .B1(n9966), .B2(n14820), .A(n7401), .ZN(n9979) );
  OR2_X1 U7572 ( .A1(n12403), .A2(n8050), .ZN(n7624) );
  NAND2_X2 U7573 ( .A1(n8705), .A2(n8704), .ZN(n14742) );
  OR2_X1 U7574 ( .A1(n12337), .A2(n8923), .ZN(n8712) );
  NAND2_X1 U7575 ( .A1(n7514), .A2(n8708), .ZN(n12337) );
  INV_X1 U7576 ( .A(n8030), .ZN(n15832) );
  NAND2_X1 U7577 ( .A1(n7649), .A2(n8635), .ZN(n7514) );
  CLKBUF_X1 U7578 ( .A(n9934), .Z(n7531) );
  NAND2_X1 U7579 ( .A1(n7552), .A2(n8707), .ZN(n8708) );
  OR2_X1 U7580 ( .A1(n12801), .A2(n12802), .ZN(n7589) );
  NAND2_X1 U7581 ( .A1(n8634), .A2(n8706), .ZN(n7650) );
  NAND2_X1 U7582 ( .A1(n8633), .A2(n11374), .ZN(n8634) );
  OR2_X1 U7583 ( .A1(n8633), .A2(n11374), .ZN(n8635) );
  AND2_X1 U7584 ( .A1(n11890), .A2(n10525), .ZN(n12196) );
  NAND2_X1 U7585 ( .A1(n9660), .A2(n9659), .ZN(n9920) );
  NAND2_X1 U7586 ( .A1(n11519), .A2(n11520), .ZN(n11711) );
  NAND2_X1 U7587 ( .A1(n8849), .A2(n8848), .ZN(n12254) );
  NAND2_X1 U7588 ( .A1(n9199), .A2(n9198), .ZN(n16421) );
  NAND2_X1 U7589 ( .A1(n8833), .A2(n8832), .ZN(n12058) );
  AND2_X1 U7590 ( .A1(n10004), .A2(n10003), .ZN(n14010) );
  INV_X2 U7591 ( .A(n14169), .ZN(n14164) );
  NAND2_X1 U7592 ( .A1(n8761), .A2(n8073), .ZN(n8612) );
  NAND2_X1 U7593 ( .A1(n8786), .A2(n8785), .ZN(n12101) );
  NAND2_X1 U7594 ( .A1(n8759), .A2(n8758), .ZN(n8761) );
  NAND2_X2 U7595 ( .A1(n11745), .A2(n16117), .ZN(n14675) );
  NAND2_X1 U7596 ( .A1(n9100), .A2(n7694), .ZN(n11816) );
  NAND2_X1 U7597 ( .A1(n11570), .A2(n9549), .ZN(n11793) );
  OR2_X1 U7598 ( .A1(n9960), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U7599 ( .A1(n9093), .A2(n9092), .ZN(n14985) );
  NAND2_X1 U7600 ( .A1(n9085), .A2(n9084), .ZN(n11802) );
  OAI21_X2 U7601 ( .B1(n10986), .B2(n8923), .A(n8803), .ZN(n16270) );
  NAND2_X1 U7602 ( .A1(n11568), .A2(n11567), .ZN(n11788) );
  AND2_X1 U7603 ( .A1(n13153), .A2(n13154), .ZN(n13308) );
  OAI21_X1 U7604 ( .B1(n8796), .B2(n8798), .A(n8797), .ZN(n10986) );
  XNOR2_X1 U7605 ( .A(n15767), .B(n8035), .ZN(n15769) );
  AND2_X2 U7606 ( .A1(n11038), .A2(n15269), .ZN(n14955) );
  NAND2_X1 U7607 ( .A1(n8033), .A2(n15766), .ZN(n15767) );
  CLKBUF_X1 U7608 ( .A(n10571), .Z(n14473) );
  AND3_X2 U7609 ( .A1(n9680), .A2(n9679), .A3(n9678), .ZN(n10122) );
  AND3_X1 U7610 ( .A1(n9742), .A2(n9741), .A3(n9740), .ZN(n12333) );
  AND3_X1 U7611 ( .A1(n9713), .A2(n9712), .A3(n9711), .ZN(n12128) );
  AND3_X1 U7612 ( .A1(n9727), .A2(n9726), .A3(n9725), .ZN(n12141) );
  NAND3_X2 U7613 ( .A1(n8825), .A2(n7924), .A3(n8824), .ZN(n11752) );
  NAND2_X2 U7614 ( .A1(n9054), .A2(n9055), .ZN(n15143) );
  CLKBUF_X1 U7615 ( .A(n11983), .Z(n10036) );
  NAND2_X1 U7616 ( .A1(n11496), .A2(n11579), .ZN(n15000) );
  NAND4_X1 U7617 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n14469) );
  INV_X1 U7618 ( .A(n9507), .ZN(n9455) );
  OR2_X1 U7619 ( .A1(n9386), .A2(n9048), .ZN(n9055) );
  AND3_X1 U7620 ( .A1(n9053), .A2(n9052), .A3(n9051), .ZN(n9054) );
  INV_X2 U7621 ( .A(n10641), .ZN(n10577) );
  BUF_X2 U7622 ( .A(n9729), .Z(n11983) );
  NAND2_X2 U7623 ( .A1(n9013), .A2(n13090), .ZN(n9386) );
  CLKBUF_X3 U7624 ( .A(n9049), .Z(n9507) );
  XNOR2_X1 U7625 ( .A(n8449), .B(n8448), .ZN(n11452) );
  AND2_X1 U7626 ( .A1(n9622), .A2(n13356), .ZN(n9729) );
  AND2_X1 U7627 ( .A1(n14317), .A2(n13356), .ZN(n9746) );
  NAND2_X2 U7628 ( .A1(n8827), .A2(n10976), .ZN(n8864) );
  AND2_X1 U7629 ( .A1(n9622), .A2(n9621), .ZN(n9692) );
  XNOR2_X1 U7630 ( .A(n9603), .B(n9602), .ZN(n15550) );
  AND2_X1 U7631 ( .A1(n10054), .A2(n10976), .ZN(n9739) );
  BUF_X2 U7632 ( .A(n9014), .Z(n13090) );
  CLKBUF_X1 U7633 ( .A(n9488), .Z(n15559) );
  OAI21_X1 U7634 ( .B1(n9604), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9603) );
  XNOR2_X1 U7635 ( .A(n8702), .B(n8937), .ZN(n10842) );
  INV_X1 U7636 ( .A(n9481), .ZN(n7368) );
  NAND2_X1 U7637 ( .A1(n14796), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8953) );
  INV_X1 U7638 ( .A(n12877), .ZN(n10825) );
  CLKBUF_X1 U7639 ( .A(n9489), .Z(n11564) );
  NAND2_X1 U7640 ( .A1(n8458), .A2(n9614), .ZN(n13335) );
  OR2_X1 U7641 ( .A1(n8443), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U7642 ( .A1(n8701), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U7643 ( .A1(n9618), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U7644 ( .A1(n9619), .A2(n9618), .ZN(n14317) );
  MUX2_X1 U7645 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8456), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8458) );
  NAND2_X1 U7646 ( .A1(n8940), .A2(n8973), .ZN(n12987) );
  MUX2_X1 U7647 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8675), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n8676) );
  NAND2_X1 U7648 ( .A1(n9011), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U7649 ( .A1(n8677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8678) );
  OR2_X1 U7650 ( .A1(n9795), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9807) );
  OR2_X1 U7651 ( .A1(n15741), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n7524) );
  INV_X4 U7652 ( .A(n10976), .ZN(n10984) );
  XNOR2_X1 U7653 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(n15740), .ZN(n15741) );
  NOR2_X1 U7654 ( .A1(n7537), .A2(n7763), .ZN(n9190) );
  NAND2_X1 U7655 ( .A1(n7527), .A2(n7525), .ZN(n15740) );
  INV_X2 U7656 ( .A(n8699), .ZN(n7369) );
  NAND2_X1 U7657 ( .A1(n8584), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7846) );
  AND2_X1 U7658 ( .A1(n8345), .A2(n8183), .ZN(n8182) );
  AND2_X1 U7659 ( .A1(n8359), .A2(n8356), .ZN(n7522) );
  NAND4_X1 U7660 ( .A1(n8997), .A2(n8996), .A3(n8995), .A4(n9144), .ZN(n7763)
         );
  AND2_X1 U7661 ( .A1(n7888), .A2(n7887), .ZN(n7582) );
  AND2_X1 U7662 ( .A1(n8362), .A2(n8454), .ZN(n8244) );
  AND3_X1 U7663 ( .A1(n9001), .A2(n13878), .A3(n9000), .ZN(n9004) );
  INV_X1 U7664 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8406) );
  INV_X1 U7665 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8661) );
  INV_X1 U7666 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9599) );
  XNOR2_X1 U7667 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9683) );
  INV_X1 U7668 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9036) );
  INV_X1 U7669 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8942) );
  INV_X1 U7670 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9039) );
  INV_X1 U7671 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8772) );
  INV_X1 U7672 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8403) );
  NOR2_X1 U7673 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8944) );
  INV_X1 U7674 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8345) );
  INV_X1 U7675 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8843) );
  INV_X1 U7676 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n13875) );
  INV_X1 U7677 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8836) );
  INV_X1 U7678 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8945) );
  INV_X4 U7679 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7680 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8581) );
  INV_X1 U7681 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9629) );
  INV_X4 U7682 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7683 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8349) );
  NOR2_X1 U7684 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8348) );
  INV_X1 U7685 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8356) );
  INV_X1 U7686 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8378) );
  XNOR2_X1 U7687 ( .A(n7583), .B(P3_IR_REG_2__SCAN_IN), .ZN(n12021) );
  AND2_X1 U7688 ( .A1(n10011), .A2(n13664), .ZN(n13961) );
  NOR2_X2 U7689 ( .A1(n10012), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10011) );
  NOR2_X2 U7690 ( .A1(n11833), .A2(n11838), .ZN(n12069) );
  OAI21_X2 U7691 ( .B1(n9878), .B2(n8231), .A(n8229), .ZN(n14119) );
  NAND2_X2 U7692 ( .A1(n9628), .A2(n9627), .ZN(n13116) );
  OR2_X1 U7693 ( .A1(n13987), .A2(n13999), .ZN(n13249) );
  AND2_X2 U7694 ( .A1(n10020), .A2(n10019), .ZN(n13999) );
  NOR2_X2 U7695 ( .A1(n15349), .A2(n15334), .ZN(n15337) );
  OR2_X1 U7696 ( .A1(n14199), .A2(n14073), .ZN(n13237) );
  INV_X1 U7697 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U7698 ( .A1(n7855), .A2(n7856), .ZN(n7853) );
  AOI21_X1 U7699 ( .B1(n13430), .B2(n14073), .A(n10190), .ZN(n13412) );
  OAI21_X1 U7700 ( .B1(n14250), .B2(n16188), .A(n13117), .ZN(n8241) );
  INV_X1 U7701 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U7702 ( .A1(n10701), .A2(n7419), .ZN(n8172) );
  NAND2_X1 U7703 ( .A1(n7520), .A2(n7519), .ZN(n8170) );
  INV_X1 U7704 ( .A(n10733), .ZN(n8128) );
  AND2_X1 U7705 ( .A1(n14220), .A2(n14147), .ZN(n13133) );
  OR2_X1 U7706 ( .A1(n8197), .A2(n8195), .ZN(n8194) );
  INV_X1 U7707 ( .A(n13358), .ZN(n8195) );
  AND2_X1 U7708 ( .A1(n7411), .A2(n13358), .ZN(n8196) );
  OR2_X1 U7709 ( .A1(n13236), .A2(n13207), .ZN(n13265) );
  AND2_X1 U7710 ( .A1(n13184), .A2(n13192), .ZN(n13313) );
  NAND2_X1 U7711 ( .A1(n10122), .A2(n10121), .ZN(n13143) );
  INV_X1 U7712 ( .A(n9777), .ZN(n9721) );
  AND2_X1 U7713 ( .A1(n13338), .A2(n10118), .ZN(n13207) );
  INV_X1 U7714 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8360) );
  INV_X1 U7715 ( .A(n9645), .ZN(n7979) );
  INV_X1 U7716 ( .A(n10801), .ZN(n7952) );
  INV_X1 U7717 ( .A(n7960), .ZN(n7955) );
  NOR2_X1 U7718 ( .A1(n12037), .A2(n12254), .ZN(n7749) );
  NAND2_X1 U7719 ( .A1(n10547), .A2(n7850), .ZN(n7849) );
  AND2_X1 U7720 ( .A1(n12575), .A2(n12456), .ZN(n7703) );
  NOR2_X1 U7721 ( .A1(n11826), .A2(n8253), .ZN(n8252) );
  INV_X1 U7722 ( .A(n15422), .ZN(n13075) );
  NAND2_X1 U7723 ( .A1(n8909), .A2(n8908), .ZN(n8916) );
  OR2_X1 U7724 ( .A1(n8905), .A2(n8904), .ZN(n8909) );
  OAI21_X1 U7725 ( .B1(n8102), .B2(n8100), .A(n8098), .ZN(n8901) );
  INV_X1 U7726 ( .A(n8099), .ZN(n8098) );
  OAI21_X1 U7727 ( .B1(n8646), .B2(n8100), .A(n8880), .ZN(n8099) );
  INV_X1 U7728 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9005) );
  AOI21_X1 U7729 ( .B1(n8634), .B2(n7421), .A(n8076), .ZN(n7648) );
  NAND2_X1 U7730 ( .A1(n8077), .A2(n8643), .ZN(n8076) );
  AND2_X1 U7731 ( .A1(n8714), .A2(n8628), .ZN(n8067) );
  NAND2_X1 U7732 ( .A1(n7657), .A2(n7656), .ZN(n7655) );
  INV_X1 U7733 ( .A(n7658), .ZN(n7657) );
  AOI21_X1 U7734 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15806), .A(n15805), .ZN(
        n15812) );
  NOR2_X1 U7735 ( .A1(n15804), .A2(n15803), .ZN(n15805) );
  AOI21_X1 U7736 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n15822), .A(n15821), .ZN(
        n15827) );
  NOR2_X1 U7737 ( .A1(n15820), .A2(n15819), .ZN(n15821) );
  NAND2_X1 U7738 ( .A1(n13980), .A2(n13242), .ZN(n13294) );
  AOI21_X1 U7739 ( .B1(n8222), .B2(n8224), .A(n7424), .ZN(n8220) );
  NAND2_X1 U7740 ( .A1(n12412), .A2(n7422), .ZN(n7559) );
  INV_X1 U7741 ( .A(n13175), .ZN(n7560) );
  AND2_X1 U7742 ( .A1(n10054), .A2(n10984), .ZN(n9777) );
  INV_X1 U7743 ( .A(n9739), .ZN(n9781) );
  INV_X1 U7744 ( .A(n10054), .ZN(n9908) );
  INV_X1 U7745 ( .A(n9721), .ZN(n9995) );
  INV_X1 U7746 ( .A(n16180), .ZN(n14161) );
  NAND2_X1 U7747 ( .A1(n10226), .A2(n13207), .ZN(n14159) );
  INV_X2 U7748 ( .A(n9721), .ZN(n13279) );
  INV_X1 U7749 ( .A(n14156), .ZN(n16183) );
  INV_X1 U7750 ( .A(n12996), .ZN(n16441) );
  OR2_X1 U7751 ( .A1(n13338), .A2(n10118), .ZN(n16467) );
  NAND2_X2 U7752 ( .A1(n12984), .A2(n13335), .ZN(n10054) );
  OAI21_X1 U7753 ( .B1(n12633), .B2(n10086), .A(n12880), .ZN(n11024) );
  OAI21_X1 U7754 ( .B1(n10008), .B2(n10006), .A(n8041), .ZN(n10028) );
  NAND2_X1 U7755 ( .A1(n13087), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8041) );
  INV_X1 U7756 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8183) );
  NOR2_X1 U7757 ( .A1(n8351), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U7758 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n12561), .ZN(n9659) );
  XNOR2_X1 U7759 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9789) );
  INV_X1 U7760 ( .A(n8377), .ZN(n8425) );
  CLKBUF_X1 U7761 ( .A(n8376), .Z(n8377) );
  INV_X1 U7762 ( .A(n12400), .ZN(n12431) );
  NAND2_X1 U7763 ( .A1(n8053), .A2(n8055), .ZN(n8051) );
  INV_X1 U7764 ( .A(n12389), .ZN(n8055) );
  NOR2_X1 U7765 ( .A1(n10929), .A2(n8058), .ZN(n8057) );
  INV_X1 U7766 ( .A(n10922), .ZN(n8058) );
  NAND2_X1 U7767 ( .A1(n7617), .A2(n7416), .ZN(n10945) );
  INV_X1 U7768 ( .A(n10946), .ZN(n7616) );
  NAND2_X1 U7769 ( .A1(n7601), .A2(n7600), .ZN(n10953) );
  INV_X1 U7770 ( .A(n10954), .ZN(n7600) );
  INV_X1 U7771 ( .A(n10955), .ZN(n7601) );
  NAND3_X1 U7772 ( .A1(n10945), .A2(n10895), .A3(n12407), .ZN(n12403) );
  OR2_X1 U7773 ( .A1(n12030), .A2(n7621), .ZN(n7617) );
  INV_X1 U7774 ( .A(n12032), .ZN(n7621) );
  NOR2_X1 U7775 ( .A1(n10933), .A2(n15568), .ZN(n10940) );
  OR2_X1 U7776 ( .A1(n14695), .A2(n14369), .ZN(n10495) );
  OR2_X1 U7777 ( .A1(n14556), .A2(n14557), .ZN(n14554) );
  INV_X1 U7778 ( .A(n7862), .ZN(n7858) );
  NAND2_X1 U7779 ( .A1(n14625), .A2(n10539), .ZN(n14605) );
  NAND2_X1 U7780 ( .A1(n12661), .A2(n12666), .ZN(n10534) );
  NAND2_X1 U7781 ( .A1(n12665), .A2(n10398), .ZN(n7941) );
  AOI21_X1 U7782 ( .B1(n10316), .B2(n7382), .A(n7445), .ZN(n11457) );
  OAI21_X1 U7783 ( .B1(n12098), .B2(n7434), .A(n10521), .ZN(n11453) );
  INV_X1 U7784 ( .A(n16107), .ZN(n16256) );
  INV_X1 U7785 ( .A(n8864), .ZN(n8819) );
  AND2_X1 U7786 ( .A1(n12987), .A2(n12877), .ZN(n16105) );
  CLKBUF_X1 U7787 ( .A(n8819), .Z(n8934) );
  OR2_X1 U7788 ( .A1(n14813), .A2(n8971), .ZN(n8989) );
  NOR2_X1 U7789 ( .A1(n14835), .A2(n7679), .ZN(n7678) );
  INV_X1 U7790 ( .A(n12861), .ZN(n7679) );
  OR2_X1 U7791 ( .A1(n14921), .A2(n14920), .ZN(n14971) );
  AND4_X1 U7792 ( .A1(n9442), .A2(n9441), .A3(n9440), .A4(n9439), .ZN(n15056)
         );
  INV_X1 U7793 ( .A(n9014), .ZN(n7538) );
  NOR2_X1 U7794 ( .A1(n9015), .A2(n9014), .ZN(n9049) );
  NAND2_X1 U7795 ( .A1(n8266), .A2(n7439), .ZN(n15277) );
  INV_X1 U7796 ( .A(n8336), .ZN(n8265) );
  INV_X1 U7797 ( .A(n7646), .ZN(n15332) );
  INV_X1 U7798 ( .A(n7785), .ZN(n7784) );
  NAND2_X1 U7799 ( .A1(n7785), .A2(n7788), .ZN(n7783) );
  NAND2_X1 U7800 ( .A1(n15507), .A2(n13065), .ZN(n15377) );
  NAND2_X1 U7801 ( .A1(n11590), .A2(n11589), .ZN(n16248) );
  NAND2_X1 U7802 ( .A1(n9600), .A2(n8291), .ZN(n9011) );
  NOR2_X1 U7803 ( .A1(n8292), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n8291) );
  XNOR2_X1 U7804 ( .A(n8932), .B(n8931), .ZN(n14794) );
  INV_X1 U7805 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9001) );
  INV_X1 U7806 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U7807 ( .A1(n8797), .A2(n8072), .ZN(n8070) );
  AND2_X1 U7808 ( .A1(n8597), .A2(n8596), .ZN(n8072) );
  NAND2_X1 U7809 ( .A1(n8787), .A2(n8597), .ZN(n8071) );
  AOI21_X1 U7810 ( .B1(n15842), .B2(n15841), .A(P2_ADDR_REG_14__SCAN_IN), .ZN(
        n7965) );
  AND3_X1 U7811 ( .A1(n9954), .A2(n9953), .A3(n9952), .ZN(n14073) );
  INV_X1 U7812 ( .A(n12984), .ZN(n13334) );
  NAND2_X1 U7813 ( .A1(n13991), .A2(n7905), .ZN(n13106) );
  NAND2_X1 U7814 ( .A1(n13991), .A2(n13246), .ZN(n13104) );
  NAND2_X1 U7815 ( .A1(n13991), .A2(n13995), .ZN(n14257) );
  AOI21_X2 U7816 ( .B1(n14383), .B2(n14379), .A(n14381), .ZN(n14435) );
  NAND2_X1 U7817 ( .A1(n12862), .A2(n7678), .ZN(n8161) );
  NAND2_X1 U7818 ( .A1(n9372), .A2(n9371), .ZN(n15484) );
  NAND2_X1 U7819 ( .A1(n11067), .A2(n16104), .ZN(n16551) );
  NAND2_X1 U7820 ( .A1(n9612), .A2(n13013), .ZN(n8305) );
  AOI22_X1 U7821 ( .A1(n16225), .A2(n10577), .B1(n10747), .B2(n14472), .ZN(
        n10584) );
  NAND2_X1 U7822 ( .A1(n7437), .A2(n10627), .ZN(n8153) );
  NAND2_X1 U7823 ( .A1(n10636), .A2(n10638), .ZN(n8164) );
  INV_X1 U7824 ( .A(n9182), .ZN(n8297) );
  AOI21_X1 U7825 ( .B1(n7834), .B2(n7833), .A(n7830), .ZN(n13701) );
  NAND2_X1 U7826 ( .A1(n7832), .A2(n7831), .ZN(n7830) );
  AOI21_X1 U7827 ( .B1(SI_14_), .B2(keyinput_18), .A(n13694), .ZN(n7833) );
  OAI21_X1 U7828 ( .B1(n13688), .B2(n13689), .A(n7835), .ZN(n7834) );
  OAI21_X1 U7829 ( .B1(n13727), .B2(n13726), .A(n13725), .ZN(n13731) );
  OAI22_X1 U7830 ( .A1(n13734), .A2(keyinput_40), .B1(n13735), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n7812) );
  OAI21_X1 U7831 ( .B1(n7809), .B2(n7506), .A(n7807), .ZN(n13747) );
  NOR2_X1 U7832 ( .A1(n13746), .A2(n7808), .ZN(n7807) );
  INV_X1 U7833 ( .A(n10693), .ZN(n7519) );
  NOR2_X1 U7834 ( .A1(n10713), .A2(n7381), .ZN(n8159) );
  OR2_X1 U7835 ( .A1(n8322), .A2(n9363), .ZN(n8321) );
  INV_X1 U7836 ( .A(n9362), .ZN(n8322) );
  NAND2_X1 U7837 ( .A1(n10720), .A2(n7516), .ZN(n10727) );
  NAND2_X1 U7838 ( .A1(n7518), .A2(n7517), .ZN(n7516) );
  INV_X1 U7839 ( .A(n10718), .ZN(n7517) );
  OR2_X1 U7840 ( .A1(n9407), .A2(n9409), .ZN(n8326) );
  OR2_X1 U7841 ( .A1(n8014), .A2(n8013), .ZN(n8012) );
  NAND2_X1 U7842 ( .A1(n8015), .A2(n13127), .ZN(n8014) );
  INV_X1 U7843 ( .A(n13238), .ZN(n8015) );
  INV_X1 U7844 ( .A(n10743), .ZN(n8147) );
  AND2_X1 U7845 ( .A1(n13302), .A2(n13164), .ZN(n10068) );
  OR2_X1 U7846 ( .A1(n14202), .A2(n14089), .ZN(n10184) );
  INV_X1 U7847 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8657) );
  INV_X1 U7848 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8656) );
  NOR2_X1 U7849 ( .A1(n15247), .A2(n7723), .ZN(n7722) );
  NAND2_X1 U7850 ( .A1(n8101), .A2(n7502), .ZN(n8100) );
  INV_X1 U7851 ( .A(n8881), .ZN(n8101) );
  OAI21_X1 U7852 ( .B1(n8645), .B2(n8648), .A(n7391), .ZN(n8102) );
  NAND2_X1 U7853 ( .A1(n7637), .A2(n8608), .ZN(n7636) );
  INV_X1 U7854 ( .A(n8610), .ZN(n7637) );
  AND2_X1 U7855 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  NAND2_X1 U7856 ( .A1(n8582), .A2(n8581), .ZN(n7629) );
  INV_X1 U7857 ( .A(n10157), .ZN(n10129) );
  AND2_X1 U7858 ( .A1(n13207), .A2(n13289), .ZN(n7982) );
  NAND2_X1 U7859 ( .A1(n7995), .A2(n13266), .ZN(n7993) );
  NOR2_X1 U7860 ( .A1(n13207), .A2(n10237), .ZN(n7983) );
  NOR2_X1 U7861 ( .A1(n13287), .A2(n13290), .ZN(n7995) );
  NAND2_X1 U7862 ( .A1(n13288), .A2(n13326), .ZN(n7984) );
  INV_X1 U7863 ( .A(n7581), .ZN(n7908) );
  AND2_X1 U7864 ( .A1(n10175), .A2(n14122), .ZN(n13299) );
  INV_X1 U7865 ( .A(n13222), .ZN(n13300) );
  NAND2_X1 U7866 ( .A1(n8232), .A2(n14144), .ZN(n8230) );
  INV_X1 U7867 ( .A(n13131), .ZN(n13129) );
  AND2_X1 U7868 ( .A1(n14130), .A2(n9879), .ZN(n8232) );
  INV_X1 U7869 ( .A(n13194), .ZN(n7895) );
  OAI21_X1 U7870 ( .B1(n12918), .B2(n7895), .A(n13197), .ZN(n7894) );
  NAND2_X1 U7871 ( .A1(n9794), .A2(n8235), .ZN(n8234) );
  INV_X1 U7872 ( .A(n9782), .ZN(n8235) );
  OR2_X1 U7873 ( .A1(n13137), .A2(n9691), .ZN(n8226) );
  NAND2_X1 U7874 ( .A1(n14099), .A2(n14098), .ZN(n7900) );
  NAND2_X1 U7875 ( .A1(n9662), .A2(n9661), .ZN(n9934) );
  NAND2_X1 U7876 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n12771), .ZN(n9661) );
  INV_X1 U7877 ( .A(n8000), .ZN(n7999) );
  OAI21_X1 U7878 ( .B1(n9865), .B2(n8001), .A(n9880), .ZN(n8000) );
  INV_X1 U7879 ( .A(n9655), .ZN(n8001) );
  INV_X1 U7880 ( .A(n7978), .ZN(n7977) );
  OAI21_X1 U7881 ( .B1(n9801), .B2(n7979), .A(n9813), .ZN(n7978) );
  INV_X1 U7882 ( .A(n9631), .ZN(n8004) );
  AND3_X2 U7883 ( .A1(n10795), .A2(n11753), .A3(n10835), .ZN(n10641) );
  NOR2_X1 U7884 ( .A1(n7754), .A2(n10455), .ZN(n7753) );
  NOR2_X1 U7885 ( .A1(n12936), .A2(n14791), .ZN(n12935) );
  INV_X1 U7886 ( .A(n10535), .ZN(n7867) );
  AOI21_X1 U7887 ( .B1(n7940), .B2(n7938), .A(n7937), .ZN(n7936) );
  INV_X1 U7888 ( .A(n10398), .ZN(n7938) );
  INV_X1 U7889 ( .A(n12743), .ZN(n7937) );
  AND2_X1 U7890 ( .A1(n7413), .A2(n12627), .ZN(n7940) );
  INV_X1 U7891 ( .A(n12426), .ZN(n7954) );
  NOR2_X1 U7892 ( .A1(n12255), .A2(n7958), .ZN(n7957) );
  INV_X1 U7893 ( .A(n10367), .ZN(n7958) );
  NOR2_X1 U7894 ( .A1(n10368), .A2(n7961), .ZN(n7960) );
  INV_X1 U7895 ( .A(n10358), .ZN(n7961) );
  OR2_X1 U7896 ( .A1(n10361), .A2(n10360), .ZN(n10369) );
  XNOR2_X1 U7897 ( .A(n16225), .B(n14472), .ZN(n10807) );
  INV_X1 U7898 ( .A(n14584), .ZN(n8872) );
  AND2_X1 U7899 ( .A1(n8670), .A2(n8671), .ZN(n7521) );
  NOR2_X1 U7900 ( .A1(n11868), .A2(n8138), .ZN(n8137) );
  INV_X1 U7901 ( .A(n11709), .ZN(n8138) );
  AND2_X1 U7902 ( .A1(n7686), .A2(n14940), .ZN(n7684) );
  INV_X1 U7903 ( .A(n7688), .ZN(n7682) );
  NAND2_X1 U7904 ( .A1(n9412), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9411) );
  INV_X1 U7905 ( .A(n14904), .ZN(n8151) );
  INV_X1 U7906 ( .A(n14917), .ZN(n8152) );
  AND2_X1 U7907 ( .A1(n8149), .A2(n7662), .ZN(n7661) );
  NAND2_X1 U7908 ( .A1(n14992), .A2(n7663), .ZN(n7662) );
  INV_X1 U7909 ( .A(n14891), .ZN(n7663) );
  INV_X1 U7910 ( .A(n14992), .ZN(n7664) );
  INV_X1 U7911 ( .A(n7678), .ZN(n7676) );
  OR2_X1 U7912 ( .A1(n15274), .A2(n15428), .ZN(n7775) );
  AOI21_X1 U7913 ( .B1(n15262), .B2(n7714), .A(n7720), .ZN(n7719) );
  NOR2_X1 U7914 ( .A1(n7723), .A2(n7371), .ZN(n7714) );
  INV_X1 U7915 ( .A(n7719), .ZN(n7717) );
  INV_X1 U7916 ( .A(n7722), .ZN(n7721) );
  NAND2_X1 U7917 ( .A1(n8252), .A2(n8250), .ZN(n8249) );
  INV_X1 U7918 ( .A(n11585), .ZN(n8250) );
  OR2_X1 U7919 ( .A1(n7690), .A2(n12875), .ZN(n11579) );
  AND2_X1 U7920 ( .A1(n7691), .A2(n7469), .ZN(n12269) );
  INV_X1 U7921 ( .A(n12875), .ZN(n11588) );
  INV_X1 U7922 ( .A(n9596), .ZN(n9600) );
  NAND2_X1 U7923 ( .A1(n8293), .A2(n9028), .ZN(n8292) );
  INV_X1 U7924 ( .A(n9007), .ZN(n8293) );
  NOR2_X2 U7925 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7760) );
  XNOR2_X1 U7926 ( .A(n8901), .B(SI_26_), .ZN(n8886) );
  NOR2_X1 U7927 ( .A1(n8640), .A2(n8085), .ZN(n8084) );
  NOR2_X1 U7928 ( .A1(n8639), .A2(SI_20_), .ZN(n8640) );
  INV_X1 U7929 ( .A(n8638), .ZN(n8085) );
  INV_X1 U7930 ( .A(n8082), .ZN(n8081) );
  AOI21_X1 U7931 ( .B1(n8084), .B2(n8698), .A(n8083), .ZN(n8082) );
  NOR2_X1 U7932 ( .A1(n8692), .A2(n13668), .ZN(n8083) );
  NAND2_X1 U7933 ( .A1(n7403), .A2(n8618), .ZN(n8094) );
  NAND2_X1 U7934 ( .A1(n8614), .A2(SI_10_), .ZN(n8615) );
  NAND2_X1 U7935 ( .A1(n8749), .A2(n13506), .ZN(n8613) );
  NAND2_X1 U7936 ( .A1(n8612), .A2(n8611), .ZN(n8749) );
  NAND2_X1 U7937 ( .A1(n7632), .A2(n8608), .ZN(n8750) );
  NAND2_X1 U7938 ( .A1(n8612), .A2(n8610), .ZN(n7632) );
  NAND2_X1 U7939 ( .A1(n7841), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U7940 ( .A1(n7844), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7842) );
  INV_X1 U7941 ( .A(n7629), .ZN(n7844) );
  INV_X1 U7942 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15758) );
  INV_X1 U7943 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15772) );
  AOI22_X1 U7944 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15982), .B1(n15778), .B2(
        n15777), .ZN(n15779) );
  OR2_X1 U7945 ( .A1(n15982), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n15778) );
  INV_X1 U7946 ( .A(n8198), .ZN(n8197) );
  OAI22_X1 U7947 ( .A1(n13449), .A2(n8200), .B1(n13462), .B2(n10201), .ZN(
        n8198) );
  INV_X1 U7948 ( .A(n13389), .ZN(n8199) );
  NOR2_X1 U7949 ( .A1(n13001), .A2(n7574), .ZN(n7573) );
  INV_X1 U7950 ( .A(n10162), .ZN(n7574) );
  OR2_X1 U7951 ( .A1(n12925), .A2(n12924), .ZN(n7575) );
  INV_X1 U7952 ( .A(n7488), .ZN(n8204) );
  OAI21_X1 U7953 ( .B1(n10199), .B2(n11883), .A(n8214), .ZN(n11413) );
  NAND2_X1 U7954 ( .A1(n11884), .A2(n11883), .ZN(n8214) );
  NAND2_X1 U7955 ( .A1(n12222), .A2(n8215), .ZN(n12509) );
  NOR2_X1 U7956 ( .A1(n12512), .A2(n8216), .ZN(n8215) );
  INV_X1 U7957 ( .A(n10147), .ZN(n8216) );
  AND2_X1 U7958 ( .A1(n13201), .A2(n13200), .ZN(n13197) );
  NAND2_X1 U7959 ( .A1(n11846), .A2(n11845), .ZN(n8218) );
  AND2_X1 U7960 ( .A1(n13038), .A2(n8213), .ZN(n8212) );
  INV_X1 U7961 ( .A(n8342), .ZN(n8213) );
  AND4_X1 U7962 ( .A1(n9761), .A2(n9760), .A3(n9759), .A4(n9758), .ZN(n12294)
         );
  AND2_X1 U7963 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  OR2_X1 U7964 ( .A1(n15906), .A2(n7586), .ZN(n7585) );
  AND2_X1 U7965 ( .A1(n8413), .A2(n10965), .ZN(n7586) );
  OR2_X1 U7966 ( .A1(n15943), .A2(n8420), .ZN(n7591) );
  NAND2_X1 U7967 ( .A1(n7591), .A2(n7590), .ZN(n7917) );
  INV_X1 U7968 ( .A(n15966), .ZN(n7590) );
  AND2_X1 U7969 ( .A1(n7917), .A2(n7916), .ZN(n8421) );
  NAND2_X1 U7970 ( .A1(n10973), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U7971 ( .A1(n7599), .A2(n7598), .ZN(n7919) );
  INV_X1 U7972 ( .A(n16003), .ZN(n7598) );
  AOI21_X1 U7973 ( .B1(n8431), .B2(n8552), .A(n7922), .ZN(n7921) );
  INV_X1 U7974 ( .A(n8555), .ZN(n7922) );
  INV_X1 U7975 ( .A(n13898), .ZN(n7587) );
  NAND2_X1 U7976 ( .A1(n12803), .A2(n8482), .ZN(n13901) );
  XNOR2_X1 U7977 ( .A(n8483), .B(n13929), .ZN(n13924) );
  NAND2_X1 U7978 ( .A1(n13924), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13923) );
  NOR2_X1 U7979 ( .A1(n14014), .A2(n8246), .ZN(n8245) );
  INV_X1 U7980 ( .A(n9978), .ZN(n8246) );
  AND2_X1 U7981 ( .A1(n14023), .A2(n9978), .ZN(n14008) );
  NAND2_X1 U7982 ( .A1(n14141), .A2(n8232), .ZN(n14129) );
  NAND2_X1 U7983 ( .A1(n9841), .A2(n10161), .ZN(n13025) );
  OR2_X1 U7984 ( .A1(n13017), .A2(n9839), .ZN(n9841) );
  OAI21_X1 U7985 ( .B1(n12915), .B2(n10159), .A(n10160), .ZN(n13017) );
  AND2_X1 U7986 ( .A1(n13313), .A2(n13181), .ZN(n7558) );
  AND4_X1 U7987 ( .A1(n9774), .A2(n9773), .A3(n9772), .A4(n9771), .ZN(n12588)
         );
  NAND2_X1 U7988 ( .A1(n9768), .A2(n7405), .ZN(n12409) );
  AND2_X1 U7989 ( .A1(n13175), .A2(n13176), .ZN(n13173) );
  NAND2_X1 U7990 ( .A1(n12291), .A2(n13167), .ZN(n12442) );
  AND3_X1 U7991 ( .A1(n9702), .A2(n9701), .A3(n9700), .ZN(n11645) );
  OR2_X1 U7992 ( .A1(n9721), .A2(SI_2_), .ZN(n9702) );
  OR2_X1 U7993 ( .A1(n10054), .A2(n7889), .ZN(n9684) );
  NAND2_X1 U7994 ( .A1(n7900), .A2(n7897), .ZN(n14068) );
  AND2_X1 U7995 ( .A1(n10225), .A2(n13207), .ZN(n16180) );
  INV_X1 U7996 ( .A(n14159), .ZN(n16178) );
  OAI22_X1 U7997 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n14800), .B1(n13270), 
        .B2(n13269), .ZN(n13276) );
  AND3_X2 U7998 ( .A1(n8361), .A2(n8376), .A3(n7414), .ZN(n8364) );
  AND2_X1 U7999 ( .A1(n8244), .A2(n8460), .ZN(n8243) );
  AOI21_X1 U8000 ( .B1(n9672), .B2(n9993), .A(n9671), .ZN(n10008) );
  INV_X1 U8001 ( .A(n9994), .ZN(n9672) );
  INV_X1 U8002 ( .A(n8364), .ZN(n8370) );
  XNOR2_X1 U8003 ( .A(n9668), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n9966) );
  INV_X1 U8004 ( .A(n8028), .ZN(n8022) );
  INV_X1 U8005 ( .A(n8025), .ZN(n8024) );
  OAI21_X1 U8006 ( .B1(n8027), .B2(n9663), .A(n8026), .ZN(n8025) );
  NAND2_X1 U8007 ( .A1(n8029), .A2(n8028), .ZN(n8023) );
  INV_X1 U8008 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U8009 ( .A1(n9658), .A2(n9657), .ZN(n9907) );
  NAND2_X1 U8010 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n12336), .ZN(n9657) );
  NAND2_X1 U8011 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n12023), .ZN(n9655) );
  INV_X1 U8012 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9644) );
  INV_X1 U8013 ( .A(n7973), .ZN(n7972) );
  INV_X1 U8014 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9641) );
  INV_X1 U8015 ( .A(n8186), .ZN(n8180) );
  XNOR2_X1 U8016 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9775) );
  NAND2_X1 U8017 ( .A1(n9640), .A2(n9639), .ZN(n9776) );
  OAI21_X1 U8018 ( .B1(n9752), .B2(n9638), .A(n9637), .ZN(n9763) );
  AND2_X1 U8019 ( .A1(n11010), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9638) );
  XNOR2_X1 U8020 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9762) );
  XNOR2_X1 U8021 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9708) );
  NAND2_X1 U8022 ( .A1(n9683), .A2(n9682), .ZN(n9681) );
  NOR3_X1 U8023 ( .A1(n14818), .A2(n14813), .A3(n14815), .ZN(n10829) );
  AOI21_X1 U8024 ( .B1(n8054), .B2(n12389), .A(n7450), .ZN(n8053) );
  INV_X1 U8025 ( .A(n10898), .ZN(n8054) );
  INV_X1 U8026 ( .A(n14467), .ZN(n11505) );
  NAND2_X1 U8027 ( .A1(n8061), .A2(n8065), .ZN(n8060) );
  NOR2_X1 U8028 ( .A1(n14359), .A2(n10917), .ZN(n8065) );
  OR2_X1 U8029 ( .A1(n8063), .A2(n12909), .ZN(n8061) );
  NAND2_X1 U8030 ( .A1(n8059), .A2(n7612), .ZN(n7611) );
  INV_X1 U8031 ( .A(n7614), .ZN(n7612) );
  XNOR2_X1 U8032 ( .A(n14742), .B(n10854), .ZN(n14399) );
  AOI21_X1 U8033 ( .B1(n7620), .B2(n12032), .A(n7451), .ZN(n7619) );
  INV_X1 U8034 ( .A(n10887), .ZN(n7620) );
  AND2_X1 U8035 ( .A1(n8043), .A2(n10871), .ZN(n7628) );
  INV_X1 U8036 ( .A(n11654), .ZN(n8043) );
  AND2_X1 U8037 ( .A1(n7626), .A2(n7623), .ZN(n7622) );
  INV_X1 U8038 ( .A(n12898), .ZN(n7623) );
  AND2_X1 U8039 ( .A1(n10467), .A2(n10466), .ZN(n14439) );
  NAND2_X1 U8040 ( .A1(n10296), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10303) );
  NOR2_X1 U8041 ( .A1(n7875), .A2(n7874), .ZN(n7873) );
  INV_X1 U8042 ( .A(n10551), .ZN(n7875) );
  NOR2_X1 U8043 ( .A1(n7943), .A2(n14499), .ZN(n7942) );
  INV_X1 U8044 ( .A(n10484), .ZN(n7943) );
  NAND2_X1 U8045 ( .A1(n14528), .A2(n10550), .ZN(n14514) );
  NOR2_X1 U8046 ( .A1(n14573), .A2(n7751), .ZN(n14523) );
  NAND2_X1 U8047 ( .A1(n7753), .A2(n14521), .ZN(n7751) );
  OR2_X1 U8048 ( .A1(n10455), .A2(n14567), .ZN(n10456) );
  INV_X1 U8049 ( .A(n14558), .ZN(n14582) );
  NAND2_X1 U8050 ( .A1(n7458), .A2(n7952), .ZN(n7951) );
  AOI21_X1 U8051 ( .B1(n7857), .B2(n10540), .A(n7378), .ZN(n7855) );
  OR2_X1 U8052 ( .A1(n14739), .A2(n14629), .ZN(n7862) );
  INV_X1 U8053 ( .A(n14605), .ZN(n7861) );
  NAND2_X1 U8054 ( .A1(n14608), .A2(n14609), .ZN(n14607) );
  NAND2_X1 U8055 ( .A1(n14640), .A2(n7433), .ZN(n14625) );
  INV_X1 U8056 ( .A(n14623), .ZN(n10538) );
  XNOR2_X1 U8057 ( .A(n14742), .B(n14457), .ZN(n14623) );
  OAI21_X1 U8058 ( .B1(n12934), .B2(n12933), .A(n10536), .ZN(n14641) );
  XNOR2_X1 U8059 ( .A(n7745), .B(n14360), .ZN(n14650) );
  NAND2_X1 U8060 ( .A1(n14641), .A2(n14650), .ZN(n14640) );
  OR2_X1 U8061 ( .A1(n12795), .A2(n10412), .ZN(n12941) );
  NAND2_X1 U8062 ( .A1(n10534), .A2(n7868), .ZN(n12622) );
  NAND2_X1 U8063 ( .A1(n7941), .A2(n7940), .ZN(n12744) );
  NOR2_X1 U8064 ( .A1(n12902), .A2(n12663), .ZN(n12748) );
  NAND2_X1 U8065 ( .A1(n12493), .A2(n10391), .ZN(n12665) );
  NOR2_X1 U8066 ( .A1(n14677), .A2(n12504), .ZN(n7747) );
  NAND2_X1 U8067 ( .A1(n7959), .A2(n7957), .ZN(n12428) );
  NAND2_X1 U8068 ( .A1(n10359), .A2(n7960), .ZN(n7959) );
  NAND2_X1 U8069 ( .A1(n10350), .A2(n10349), .ZN(n12199) );
  OAI21_X1 U8070 ( .B1(n11453), .B2(n11456), .A(n10522), .ZN(n12082) );
  INV_X1 U8071 ( .A(n10844), .ZN(n11753) );
  INV_X1 U8072 ( .A(n14628), .ZN(n16108) );
  NAND2_X1 U8073 ( .A1(n10795), .A2(n10504), .ZN(n16107) );
  NAND2_X1 U8074 ( .A1(n13102), .A2(n14751), .ZN(n7926) );
  NOR2_X1 U8075 ( .A1(n7930), .A2(n10512), .ZN(n7928) );
  INV_X1 U8076 ( .A(n13100), .ZN(n7930) );
  NAND2_X1 U8077 ( .A1(n8870), .A2(n8869), .ZN(n14585) );
  OR2_X1 U8078 ( .A1(n11014), .A2(n8923), .ZN(n8767) );
  NAND2_X1 U8079 ( .A1(n8952), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8954) );
  INV_X1 U8080 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U8081 ( .A1(n8961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U8082 ( .A1(n8966), .A2(n8965), .ZN(n8964) );
  NAND2_X1 U8083 ( .A1(n7404), .A2(n8142), .ZN(n8973) );
  OAI21_X1 U8084 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(n8142), .A(n8143), .ZN(
        n8141) );
  NAND2_X1 U8085 ( .A1(n8142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U8086 ( .A1(n8699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8863) );
  INV_X1 U8087 ( .A(n8135), .ZN(n8134) );
  OAI21_X1 U8088 ( .B1(n11868), .B2(n8136), .A(n11867), .ZN(n8135) );
  NAND2_X1 U8089 ( .A1(n11710), .A2(n11709), .ZN(n8136) );
  NAND2_X1 U8090 ( .A1(n11711), .A2(n8137), .ZN(n8132) );
  NAND2_X1 U8091 ( .A1(n11471), .A2(n11470), .ZN(n11476) );
  AOI21_X1 U8092 ( .B1(n14963), .B2(n14960), .A(n14998), .ZN(n7672) );
  INV_X1 U8093 ( .A(n7672), .ZN(n7670) );
  NOR2_X1 U8094 ( .A1(n8117), .A2(n8113), .ZN(n8112) );
  INV_X1 U8095 ( .A(n12648), .ZN(n8113) );
  INV_X1 U8096 ( .A(n12652), .ZN(n8117) );
  INV_X1 U8097 ( .A(n12650), .ZN(n8116) );
  AND2_X1 U8098 ( .A1(n14971), .A2(n14922), .ZN(n15074) );
  NAND2_X1 U8099 ( .A1(n15028), .A2(n14949), .ZN(n15096) );
  NOR2_X1 U8100 ( .A1(n9263), .A2(n9262), .ZN(n9283) );
  AND4_X1 U8101 ( .A1(n9416), .A2(n9415), .A3(n9414), .A4(n9413), .ZN(n15057)
         );
  AND4_X1 U8102 ( .A1(n9218), .A2(n9217), .A3(n9216), .A4(n9215), .ZN(n12640)
         );
  AND4_X1 U8103 ( .A1(n9205), .A2(n9204), .A3(n9203), .A4(n9202), .ZN(n12343)
         );
  AND4_X1 U8104 ( .A1(n9127), .A2(n9126), .A3(n9125), .A4(n9124), .ZN(n11823)
         );
  OR2_X1 U8105 ( .A1(n15208), .A2(n15207), .ZN(n15209) );
  OR2_X1 U8106 ( .A1(n11671), .A2(n11672), .ZN(n11669) );
  INV_X2 U8107 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n13878) );
  OAI21_X1 U8108 ( .B1(n15247), .B2(n8289), .A(n13062), .ZN(n8287) );
  CLKBUF_X1 U8109 ( .A(n15258), .Z(n15259) );
  NAND2_X1 U8110 ( .A1(n13060), .A2(n15247), .ZN(n15260) );
  INV_X1 U8111 ( .A(n15258), .ZN(n13060) );
  AND2_X1 U8112 ( .A1(n7793), .A2(n13055), .ZN(n7534) );
  NAND2_X1 U8113 ( .A1(n7643), .A2(n13055), .ZN(n7641) );
  INV_X1 U8114 ( .A(n7791), .ZN(n7643) );
  OR2_X1 U8115 ( .A1(n9544), .A2(n15056), .ZN(n9545) );
  NAND2_X1 U8116 ( .A1(n9418), .A2(n9417), .ZN(n14928) );
  NAND2_X1 U8117 ( .A1(n7708), .A2(n7400), .ZN(n7707) );
  INV_X1 U8118 ( .A(n8262), .ZN(n7708) );
  NAND2_X1 U8119 ( .A1(n9381), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9400) );
  NOR2_X1 U8120 ( .A1(n15318), .A2(n8263), .ZN(n8262) );
  INV_X1 U8121 ( .A(n13071), .ZN(n8263) );
  NAND2_X1 U8122 ( .A1(n9391), .A2(n9390), .ZN(n15334) );
  OR2_X1 U8123 ( .A1(n15484), .A2(n13068), .ZN(n13069) );
  NAND2_X1 U8124 ( .A1(n15331), .A2(n15330), .ZN(n15329) );
  OR2_X1 U8125 ( .A1(n7789), .A2(n7786), .ZN(n7785) );
  INV_X1 U8126 ( .A(n13044), .ZN(n7786) );
  XNOR2_X1 U8127 ( .A(n15500), .B(n15128), .ZN(n15378) );
  INV_X1 U8128 ( .A(n16550), .ZN(n7769) );
  NAND2_X1 U8129 ( .A1(n9328), .A2(n9327), .ZN(n15508) );
  AND2_X1 U8130 ( .A1(n12959), .A2(n7412), .ZN(n7789) );
  NOR2_X1 U8131 ( .A1(n15397), .A2(n8261), .ZN(n8260) );
  INV_X1 U8132 ( .A(n12954), .ZN(n8261) );
  NAND2_X1 U8133 ( .A1(n12952), .A2(n12951), .ZN(n15395) );
  NAND2_X1 U8134 ( .A1(n12717), .A2(n12716), .ZN(n12952) );
  NAND2_X1 U8135 ( .A1(n12675), .A2(n12674), .ZN(n8285) );
  AND2_X1 U8136 ( .A1(n7700), .A2(n12687), .ZN(n7699) );
  OR2_X1 U8137 ( .A1(n7703), .A2(n7702), .ZN(n7700) );
  INV_X1 U8138 ( .A(n12687), .ZN(n12674) );
  NAND2_X1 U8139 ( .A1(n12457), .A2(n7703), .ZN(n12564) );
  NAND2_X1 U8140 ( .A1(n9220), .A2(n9219), .ZN(n12642) );
  NAND2_X1 U8141 ( .A1(n12269), .A2(n12268), .ZN(n12345) );
  NOR2_X1 U8142 ( .A1(n9184), .A2(n9183), .ZN(n9200) );
  NAND2_X1 U8143 ( .A1(n11824), .A2(n11823), .ZN(n8279) );
  NAND2_X1 U8144 ( .A1(n11578), .A2(n11577), .ZN(n11822) );
  NAND2_X1 U8145 ( .A1(n11808), .A2(n11585), .ZN(n8254) );
  AND2_X1 U8146 ( .A1(n11063), .A2(n9598), .ZN(n15099) );
  AND2_X1 U8147 ( .A1(n15560), .A2(n9059), .ZN(n15470) );
  AND2_X1 U8148 ( .A1(n11564), .A2(n12875), .ZN(n16086) );
  NAND2_X1 U8149 ( .A1(n8919), .A2(n8918), .ZN(n8929) );
  XNOR2_X1 U8150 ( .A(n8916), .B(n8915), .ZN(n13088) );
  NOR2_X1 U8151 ( .A1(n7537), .A2(n7763), .ZN(n7713) );
  INV_X1 U8152 ( .A(n8292), .ZN(n7712) );
  INV_X1 U8153 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9028) );
  AND3_X1 U8154 ( .A1(n7760), .A2(n8997), .A3(n9144), .ZN(n7758) );
  NOR2_X1 U8155 ( .A1(n9007), .A2(n7759), .ZN(n7756) );
  XNOR2_X1 U8156 ( .A(n8655), .B(n8654), .ZN(n14814) );
  NAND2_X1 U8157 ( .A1(n8075), .A2(n8644), .ZN(n8646) );
  AND3_X1 U8158 ( .A1(n9031), .A2(n7467), .A3(n9190), .ZN(n9032) );
  NAND2_X1 U8159 ( .A1(n9032), .A2(n13875), .ZN(n9038) );
  XNOR2_X1 U8160 ( .A(n8697), .B(n8698), .ZN(n12557) );
  NAND2_X1 U8161 ( .A1(n8068), .A2(n8628), .ZN(n8715) );
  INV_X1 U8162 ( .A(n8777), .ZN(n8069) );
  OAI21_X1 U8163 ( .B1(n15894), .B2(n15893), .A(P2_ADDR_REG_6__SCAN_IN), .ZN(
        n7523) );
  OAI21_X1 U8164 ( .B1(n15816), .B2(n15817), .A(P2_ADDR_REG_11__SCAN_IN), .ZN(
        n7532) );
  OAI21_X1 U8165 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15829), .A(n15828), .ZN(
        n15838) );
  AND2_X1 U8166 ( .A1(n7575), .A2(n7573), .ZN(n12999) );
  NAND2_X1 U8167 ( .A1(n9959), .A2(n9958), .ZN(n13367) );
  AND4_X1 U8168 ( .A1(n9788), .A2(n9787), .A3(n9786), .A4(n9785), .ZN(n12602)
         );
  NAND2_X1 U8169 ( .A1(n12601), .A2(n12600), .ZN(n12599) );
  INV_X1 U8170 ( .A(n8187), .ZN(n10204) );
  OAI21_X1 U8171 ( .B1(n13412), .B2(n8189), .A(n7444), .ZN(n8187) );
  AND4_X1 U8172 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), .ZN(n12780)
         );
  NAND2_X1 U8173 ( .A1(n13037), .A2(n10167), .ZN(n13396) );
  XNOR2_X1 U8174 ( .A(n10189), .B(n10187), .ZN(n13430) );
  NAND2_X1 U8175 ( .A1(n10211), .A2(n11923), .ZN(n13447) );
  AND4_X1 U8176 ( .A1(n9851), .A2(n9850), .A3(n9849), .A4(n9848), .ZN(n14160)
         );
  AND2_X1 U8177 ( .A1(n10209), .A2(n10208), .ZN(n13437) );
  NAND2_X1 U8178 ( .A1(n13331), .A2(n13332), .ZN(n7878) );
  XNOR2_X1 U8179 ( .A(n7880), .B(n11452), .ZN(n7879) );
  NOR2_X1 U8180 ( .A1(n13298), .A2(n13297), .ZN(n7880) );
  OR2_X1 U8181 ( .A1(n14306), .A2(n8463), .ZN(n13337) );
  OR2_X1 U8182 ( .A1(n13266), .A2(n13290), .ZN(n13336) );
  NAND2_X1 U8183 ( .A1(n9976), .A2(n9975), .ZN(n14042) );
  INV_X1 U8184 ( .A(n12602), .ZN(n13468) );
  NOR2_X1 U8185 ( .A1(n15944), .A2(n15945), .ZN(n15943) );
  NAND2_X1 U8186 ( .A1(n16036), .A2(n8477), .ZN(n12540) );
  OR2_X1 U8187 ( .A1(n16063), .A2(n16064), .ZN(n16061) );
  XNOR2_X1 U8188 ( .A(n7732), .B(n8573), .ZN(n7731) );
  NAND2_X1 U8189 ( .A1(n13948), .A2(n7733), .ZN(n7732) );
  NAND2_X1 U8190 ( .A1(n13943), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U8191 ( .A1(n8578), .A2(n7730), .ZN(n7729) );
  INV_X1 U8192 ( .A(n8494), .ZN(n7730) );
  AND2_X1 U8193 ( .A1(n8488), .A2(n8565), .ZN(n16079) );
  NOR2_X1 U8194 ( .A1(n16082), .A2(n7912), .ZN(n7910) );
  AND2_X1 U8195 ( .A1(n7914), .A2(n8575), .ZN(n7912) );
  NAND2_X1 U8196 ( .A1(n9947), .A2(n9946), .ZN(n14199) );
  NAND2_X1 U8197 ( .A1(n9885), .A2(n9884), .ZN(n14220) );
  AND3_X1 U8198 ( .A1(n9817), .A2(n9816), .A3(n9815), .ZN(n12996) );
  AND3_X1 U8199 ( .A1(n9793), .A2(n9792), .A3(n9791), .ZN(n16381) );
  INV_X1 U8200 ( .A(n14166), .ZN(n14097) );
  INV_X1 U8201 ( .A(n10022), .ZN(n14247) );
  NAND2_X1 U8202 ( .A1(n8242), .A2(n8240), .ZN(n14248) );
  NAND2_X1 U8203 ( .A1(n13115), .A2(n16183), .ZN(n8242) );
  INV_X1 U8204 ( .A(n8241), .ZN(n8240) );
  OR2_X1 U8205 ( .A1(n16447), .A2(n14254), .ZN(n7565) );
  AND2_X1 U8206 ( .A1(n7567), .A2(n7566), .ZN(n14253) );
  AOI21_X1 U8207 ( .B1(n14001), .B2(n16183), .A(n14000), .ZN(n7566) );
  NAND2_X1 U8208 ( .A1(n7568), .A2(n16475), .ZN(n7567) );
  AND2_X1 U8209 ( .A1(n10091), .A2(n10090), .ZN(n14305) );
  AND2_X1 U8210 ( .A1(n10089), .A2(n10088), .ZN(n14307) );
  NAND2_X1 U8211 ( .A1(n8464), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14306) );
  AND2_X1 U8212 ( .A1(n8244), .A2(n7577), .ZN(n7576) );
  NAND2_X1 U8213 ( .A1(n8893), .A2(n8892), .ZN(n14700) );
  NAND2_X1 U8214 ( .A1(n12403), .A2(n8053), .ZN(n7625) );
  NAND2_X1 U8215 ( .A1(n8687), .A2(n8686), .ZN(n14721) );
  NAND2_X1 U8216 ( .A1(n11771), .A2(n10862), .ZN(n10955) );
  NAND2_X1 U8217 ( .A1(n11629), .A2(n8042), .ZN(n11632) );
  AND2_X1 U8218 ( .A1(n11641), .A2(n10876), .ZN(n8042) );
  NAND2_X1 U8219 ( .A1(n11144), .A2(n11145), .ZN(n11764) );
  NAND2_X1 U8220 ( .A1(n14409), .A2(n10922), .ZN(n10928) );
  INV_X1 U8221 ( .A(n14463), .ZN(n12432) );
  NAND2_X1 U8222 ( .A1(n11679), .A2(n10884), .ZN(n12030) );
  NAND2_X1 U8223 ( .A1(n8052), .A2(n12389), .ZN(n12395) );
  NAND2_X1 U8224 ( .A1(n12403), .A2(n10898), .ZN(n8052) );
  NAND2_X1 U8225 ( .A1(n10931), .A2(n16117), .ZN(n14432) );
  XNOR2_X1 U8226 ( .A(n10553), .B(n10552), .ZN(n13102) );
  OAI21_X1 U8227 ( .B1(n14514), .B2(n7872), .A(n7871), .ZN(n10553) );
  AOI21_X1 U8228 ( .B1(n7873), .B2(n14503), .A(n7446), .ZN(n7871) );
  INV_X1 U8229 ( .A(n7873), .ZN(n7872) );
  INV_X1 U8230 ( .A(n16228), .ZN(n16403) );
  OR2_X1 U8231 ( .A1(n10932), .A2(n15568), .ZN(n16117) );
  NAND2_X1 U8232 ( .A1(n8936), .A2(n8935), .ZN(n14687) );
  INV_X1 U8233 ( .A(n14687), .ZN(n8991) );
  NAND2_X1 U8234 ( .A1(n8738), .A2(n8737), .ZN(n14666) );
  OAI21_X1 U8235 ( .B1(n8989), .B2(P2_D_REG_0__SCAN_IN), .A(n8988), .ZN(n15570) );
  NAND2_X1 U8236 ( .A1(n8087), .A2(n9029), .ZN(n15436) );
  NAND2_X1 U8237 ( .A1(n13086), .A2(n9512), .ZN(n8087) );
  NAND2_X1 U8238 ( .A1(n9274), .A2(n9273), .ZN(n16523) );
  AND2_X1 U8239 ( .A1(n14851), .A2(n14841), .ZN(n8160) );
  NAND2_X1 U8240 ( .A1(n8161), .A2(n14841), .ZN(n16518) );
  NAND2_X1 U8241 ( .A1(n9232), .A2(n9231), .ZN(n16482) );
  INV_X1 U8242 ( .A(n15102), .ZN(n16548) );
  INV_X1 U8243 ( .A(n15115), .ZN(n16546) );
  AND2_X1 U8244 ( .A1(n9518), .A2(n8305), .ZN(n8303) );
  AND2_X1 U8245 ( .A1(n9591), .A2(n9590), .ZN(n9595) );
  AND2_X1 U8246 ( .A1(n8307), .A2(n8305), .ZN(n8302) );
  AND2_X1 U8247 ( .A1(n9593), .A2(n9592), .ZN(n8307) );
  INV_X1 U8248 ( .A(n15057), .ZN(n15123) );
  INV_X1 U8249 ( .A(n12343), .ZN(n15136) );
  NAND2_X1 U8250 ( .A1(n13348), .A2(n15011), .ZN(n7539) );
  NAND2_X1 U8251 ( .A1(n13343), .A2(n16248), .ZN(n13348) );
  INV_X1 U8252 ( .A(n15470), .ZN(n15326) );
  AND2_X1 U8253 ( .A1(n15486), .A2(n13052), .ZN(n8294) );
  NAND2_X1 U8254 ( .A1(n11066), .A2(n15501), .ZN(n16104) );
  NAND2_X1 U8255 ( .A1(n7653), .A2(n7425), .ZN(n8247) );
  OR2_X1 U8256 ( .A1(n15426), .A2(n16243), .ZN(n7653) );
  NAND2_X1 U8257 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n7781) );
  OAI21_X1 U8258 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(n9010), .A(n7779), .ZN(
        n7778) );
  INV_X1 U8259 ( .A(n15768), .ZN(n8035) );
  INV_X1 U8260 ( .A(n15808), .ZN(n8017) );
  INV_X1 U8261 ( .A(n15852), .ZN(n7963) );
  NAND2_X1 U8262 ( .A1(n10608), .A2(n10607), .ZN(n8176) );
  AOI22_X1 U8263 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n13670) );
  NAND2_X1 U8264 ( .A1(n8310), .A2(n8309), .ZN(n9164) );
  NAND2_X1 U8265 ( .A1(n9149), .A2(n9151), .ZN(n8309) );
  OR2_X1 U8266 ( .A1(n9151), .A2(n9149), .ZN(n8311) );
  XNOR2_X1 U8267 ( .A(SI_23_), .B(keyinput_9), .ZN(n7825) );
  NAND2_X1 U8268 ( .A1(n13677), .A2(keyinput_6), .ZN(n7828) );
  NAND2_X1 U8269 ( .A1(n13678), .A2(SI_26_), .ZN(n7827) );
  INV_X1 U8270 ( .A(n10638), .ZN(n8168) );
  OAI21_X1 U8271 ( .B1(n7829), .B2(n7826), .A(n7824), .ZN(n13686) );
  NAND2_X1 U8272 ( .A1(n7828), .A2(n7827), .ZN(n7826) );
  NOR2_X1 U8273 ( .A1(n13682), .A2(n7825), .ZN(n7824) );
  AOI21_X1 U8274 ( .B1(keyinput_5), .B2(SI_27_), .A(n13676), .ZN(n7829) );
  NOR2_X1 U8275 ( .A1(n8297), .A2(n9180), .ZN(n8296) );
  INV_X1 U8276 ( .A(n9180), .ZN(n8295) );
  XNOR2_X1 U8277 ( .A(n13690), .B(n7836), .ZN(n7835) );
  INV_X1 U8278 ( .A(keyinput_15), .ZN(n7836) );
  NAND2_X1 U8279 ( .A1(n13695), .A2(keyinput_19), .ZN(n7832) );
  NAND2_X1 U8280 ( .A1(n13696), .A2(SI_13_), .ZN(n7831) );
  OR2_X1 U8281 ( .A1(n8329), .A2(n13710), .ZN(n7806) );
  AND2_X1 U8282 ( .A1(n13709), .A2(n7805), .ZN(n7804) );
  NAND2_X1 U8283 ( .A1(n13711), .A2(keyinput_25), .ZN(n7805) );
  INV_X1 U8284 ( .A(n13716), .ZN(n7801) );
  AND2_X1 U8285 ( .A1(n7799), .A2(n13712), .ZN(n7798) );
  NAND2_X1 U8286 ( .A1(n7800), .A2(n10969), .ZN(n7799) );
  INV_X1 U8287 ( .A(keyinput_30), .ZN(n7800) );
  INV_X1 U8288 ( .A(n10661), .ZN(n8163) );
  NAND2_X1 U8289 ( .A1(n9240), .A2(n8317), .ZN(n8316) );
  AOI21_X1 U8290 ( .B1(n7803), .B2(n7802), .A(n7797), .ZN(n13727) );
  INV_X1 U8291 ( .A(n13713), .ZN(n7802) );
  NAND2_X1 U8292 ( .A1(n7801), .A2(n7798), .ZN(n7797) );
  NAND2_X1 U8293 ( .A1(n7806), .A2(n7804), .ZN(n7803) );
  NAND2_X1 U8294 ( .A1(n10679), .A2(n7418), .ZN(n8175) );
  XNOR2_X1 U8295 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n7808) );
  AOI21_X1 U8296 ( .B1(n13733), .B2(n7811), .A(n7810), .ZN(n7809) );
  INV_X1 U8297 ( .A(n7812), .ZN(n7811) );
  INV_X1 U8298 ( .A(n13743), .ZN(n7810) );
  NAND2_X1 U8299 ( .A1(n8324), .A2(n9300), .ZN(n8323) );
  NAND2_X1 U8300 ( .A1(n13754), .A2(n13753), .ZN(n13759) );
  NOR2_X1 U8301 ( .A1(n10701), .A2(n7419), .ZN(n8173) );
  NAND2_X1 U8302 ( .A1(n9329), .A2(n9331), .ZN(n8308) );
  OAI21_X1 U8303 ( .B1(n13803), .B2(n13802), .A(n13801), .ZN(n13808) );
  AOI21_X1 U8304 ( .B1(n13794), .B2(n13793), .A(n13792), .ZN(n13803) );
  NAND2_X1 U8305 ( .A1(n10713), .A2(n7381), .ZN(n8155) );
  NAND2_X1 U8306 ( .A1(n7823), .A2(n7822), .ZN(n7821) );
  INV_X1 U8307 ( .A(n13819), .ZN(n7822) );
  NAND2_X1 U8308 ( .A1(n13820), .A2(n13821), .ZN(n7823) );
  AND2_X1 U8309 ( .A1(n7820), .A2(n7819), .ZN(n7818) );
  NAND2_X1 U8310 ( .A1(n13823), .A2(P3_DATAO_REG_8__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U8311 ( .A1(n13822), .A2(keyinput_88), .ZN(n7820) );
  NAND2_X1 U8312 ( .A1(n13827), .A2(n13826), .ZN(n7815) );
  NAND2_X1 U8313 ( .A1(keyinput_90), .A2(P3_DATAO_REG_6__SCAN_IN), .ZN(n7814)
         );
  AOI21_X1 U8314 ( .B1(n7817), .B2(n7816), .A(n7813), .ZN(n13835) );
  AOI22_X1 U8315 ( .A1(n13825), .A2(n13824), .B1(keyinput_89), .B2(
        P3_DATAO_REG_7__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U8316 ( .A1(n7815), .A2(n7814), .ZN(n7813) );
  NAND2_X1 U8317 ( .A1(n7821), .A2(n7818), .ZN(n7817) );
  INV_X1 U8318 ( .A(n10734), .ZN(n8127) );
  NAND2_X1 U8319 ( .A1(n10730), .A2(n8125), .ZN(n8123) );
  AND2_X1 U8320 ( .A1(n10734), .A2(n10729), .ZN(n8125) );
  AND2_X1 U8321 ( .A1(n10734), .A2(n10725), .ZN(n8126) );
  OR2_X1 U8322 ( .A1(n8328), .A2(n9408), .ZN(n8327) );
  INV_X1 U8323 ( .A(n9407), .ZN(n8328) );
  NAND2_X1 U8324 ( .A1(n9435), .A2(n8320), .ZN(n8319) );
  NOR2_X1 U8325 ( .A1(n13125), .A2(n8011), .ZN(n8010) );
  AND2_X1 U8326 ( .A1(n13234), .A2(n8012), .ZN(n8011) );
  OAI21_X1 U8327 ( .B1(n13262), .B2(n13266), .A(n13261), .ZN(n13263) );
  AND2_X1 U8328 ( .A1(n14287), .A2(n13442), .ZN(n13222) );
  AND2_X1 U8329 ( .A1(n13436), .A2(n14108), .ZN(n13131) );
  INV_X1 U8330 ( .A(n9957), .ZN(n8020) );
  INV_X1 U8331 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U8332 ( .A1(n10742), .A2(n8147), .ZN(n8146) );
  OAI22_X1 U8333 ( .A1(n14768), .A2(n10759), .B1(n14439), .B2(n10789), .ZN(
        n10745) );
  NOR2_X1 U8334 ( .A1(n14742), .A2(n7745), .ZN(n7744) );
  INV_X1 U8335 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8105) );
  INV_X1 U8336 ( .A(n7725), .ZN(n7723) );
  NAND2_X1 U8337 ( .A1(n15274), .A2(n14965), .ZN(n7727) );
  NAND2_X1 U8338 ( .A1(n15337), .A2(n15326), .ZN(n15307) );
  NAND2_X1 U8339 ( .A1(n8079), .A2(n8081), .ZN(n8077) );
  INV_X1 U8340 ( .A(SI_15_), .ZN(n13692) );
  NAND2_X1 U8341 ( .A1(n8037), .A2(n15751), .ZN(n15757) );
  AND2_X1 U8342 ( .A1(n10167), .A2(n7573), .ZN(n7572) );
  NAND2_X1 U8343 ( .A1(n8009), .A2(n8008), .ZN(n13328) );
  NOR2_X1 U8344 ( .A1(n13125), .A2(n8013), .ZN(n8008) );
  NAND2_X1 U8345 ( .A1(n12001), .A2(n8412), .ZN(n8413) );
  OR2_X1 U8346 ( .A1(n15936), .A2(n7736), .ZN(n8472) );
  NOR2_X1 U8347 ( .A1(n8512), .A2(n16282), .ZN(n7736) );
  OR2_X1 U8348 ( .A1(n15962), .A2(n7738), .ZN(n8474) );
  NOR2_X1 U8349 ( .A1(n15978), .A2(n16334), .ZN(n7738) );
  NAND2_X1 U8350 ( .A1(n12538), .A2(n8478), .ZN(n8479) );
  NAND2_X1 U8351 ( .A1(n12520), .A2(n8554), .ZN(n8481) );
  INV_X1 U8352 ( .A(n13133), .ZN(n10077) );
  INV_X1 U8353 ( .A(n8223), .ZN(n8222) );
  OAI21_X1 U8354 ( .B1(n9852), .B2(n8224), .A(n14154), .ZN(n8223) );
  INV_X1 U8355 ( .A(n9853), .ZN(n8224) );
  NAND2_X1 U8356 ( .A1(n12281), .A2(n7415), .ZN(n12440) );
  NAND2_X1 U8357 ( .A1(n10068), .A2(n7562), .ZN(n12280) );
  INV_X1 U8358 ( .A(n13157), .ZN(n7562) );
  NAND2_X1 U8359 ( .A1(n13164), .A2(n7561), .ZN(n12282) );
  INV_X1 U8360 ( .A(n13162), .ZN(n7561) );
  NAND2_X1 U8361 ( .A1(n14006), .A2(n10021), .ZN(n13969) );
  AND2_X1 U8362 ( .A1(n13246), .A2(n13245), .ZN(n13997) );
  OR2_X1 U8363 ( .A1(n11024), .A2(n10102), .ZN(n10108) );
  NAND2_X1 U8364 ( .A1(n9667), .A2(n9666), .ZN(n9668) );
  NAND2_X1 U8365 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n9665), .ZN(n9666) );
  NAND2_X1 U8366 ( .A1(n8021), .A2(n8019), .ZN(n9667) );
  AOI21_X1 U8367 ( .B1(n7501), .B2(n8023), .A(n8020), .ZN(n8019) );
  NAND2_X1 U8368 ( .A1(n9664), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8028) );
  INV_X1 U8369 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9664) );
  OAI21_X1 U8370 ( .B1(n9775), .B2(n7393), .A(n9789), .ZN(n7973) );
  NOR2_X1 U8371 ( .A1(n7393), .A2(n7970), .ZN(n7969) );
  INV_X1 U8372 ( .A(n9639), .ZN(n7970) );
  INV_X1 U8373 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7887) );
  INV_X1 U8374 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7888) );
  INV_X1 U8375 ( .A(n10751), .ZN(n10752) );
  OAI22_X1 U8376 ( .A1(n10768), .A2(n10770), .B1(n10763), .B2(n10764), .ZN(
        n10751) );
  NAND2_X1 U8377 ( .A1(n12935), .A2(n7744), .ZN(n7746) );
  NAND2_X1 U8378 ( .A1(n14782), .A2(n7741), .ZN(n14598) );
  AND2_X1 U8379 ( .A1(n12935), .A2(n7742), .ZN(n7741) );
  AND2_X1 U8380 ( .A1(n7743), .A2(n7744), .ZN(n7742) );
  OAI22_X1 U8381 ( .A1(n11757), .A2(n11756), .B1(n14473), .B2(n11752), .ZN(
        n16212) );
  NAND2_X1 U8382 ( .A1(n8676), .A2(n8952), .ZN(n8957) );
  INV_X1 U8383 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8939) );
  INV_X1 U8384 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8937) );
  AND2_X1 U8385 ( .A1(n8663), .A2(n8662), .ZN(n8719) );
  CLKBUF_X1 U8386 ( .A(n8716), .Z(n8717) );
  OR2_X1 U8387 ( .A1(n8830), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U8388 ( .A1(n8108), .A2(n8106), .ZN(n8107) );
  NAND2_X1 U8389 ( .A1(n8312), .A2(n8313), .ZN(n9467) );
  NAND2_X1 U8390 ( .A1(n8314), .A2(n9463), .ZN(n8313) );
  NAND2_X1 U8391 ( .A1(n7726), .A2(n7727), .ZN(n7725) );
  NOR2_X1 U8392 ( .A1(n14928), .A2(n15307), .ZN(n7768) );
  NOR2_X1 U8393 ( .A1(n16529), .A2(n7771), .ZN(n7770) );
  INV_X1 U8394 ( .A(n7772), .ZN(n7771) );
  NOR2_X1 U8395 ( .A1(n16493), .A2(n16523), .ZN(n7772) );
  INV_X1 U8396 ( .A(n12563), .ZN(n7702) );
  NAND2_X1 U8397 ( .A1(n8281), .A2(n8279), .ZN(n8276) );
  INV_X1 U8398 ( .A(n8279), .ZN(n8278) );
  AND2_X1 U8399 ( .A1(n16288), .A2(n12044), .ZN(n11594) );
  NAND2_X1 U8400 ( .A1(n12676), .A2(n7770), .ZN(n15406) );
  AND2_X1 U8401 ( .A1(n16086), .A2(n12770), .ZN(n11068) );
  INV_X1 U8402 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8998) );
  INV_X1 U8403 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8995) );
  INV_X1 U8404 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U8405 ( .A1(n8097), .A2(n7502), .ZN(n8882) );
  NAND2_X1 U8406 ( .A1(n8102), .A2(n8646), .ZN(n8097) );
  XNOR2_X1 U8407 ( .A(n8882), .B(SI_24_), .ZN(n8681) );
  XNOR2_X1 U8408 ( .A(n9040), .B(n9039), .ZN(n9489) );
  NOR2_X1 U8409 ( .A1(n8828), .A2(n8074), .ZN(n8073) );
  INV_X1 U8410 ( .A(n8605), .ZN(n8074) );
  AND2_X1 U8411 ( .A1(n8093), .A2(n7634), .ZN(n7633) );
  AND2_X1 U8412 ( .A1(n8096), .A2(n7465), .ZN(n8093) );
  OAI21_X1 U8413 ( .B1(n8611), .B2(SI_9_), .A(n7636), .ZN(n7635) );
  NAND2_X1 U8414 ( .A1(n7633), .A2(n7638), .ZN(n7631) );
  NOR2_X1 U8415 ( .A1(n8608), .A2(n13506), .ZN(n7638) );
  OAI21_X1 U8416 ( .B1(n10983), .B2(n7529), .A(n7528), .ZN(n8594) );
  NAND2_X1 U8417 ( .A1(n10983), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U8418 ( .A1(n7760), .A2(n8998), .ZN(n9098) );
  OAI21_X1 U8419 ( .B1(n10983), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n7513), .ZN(
        n8804) );
  NAND2_X1 U8420 ( .A1(n10983), .A2(n10989), .ZN(n7513) );
  NAND2_X1 U8421 ( .A1(n7838), .A2(SI_1_), .ZN(n8588) );
  NAND2_X1 U8422 ( .A1(n15782), .A2(n15781), .ZN(n15793) );
  OR2_X1 U8423 ( .A1(n15780), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n15781) );
  INV_X1 U8424 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15806) );
  OR2_X1 U8425 ( .A1(n15864), .A2(n15863), .ZN(n15870) );
  NOR2_X1 U8426 ( .A1(n9911), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U8427 ( .A1(n8194), .A2(n7430), .ZN(n8193) );
  NAND2_X1 U8428 ( .A1(n8196), .A2(n8201), .ZN(n8189) );
  AND2_X1 U8429 ( .A1(n8208), .A2(n7571), .ZN(n7570) );
  NAND2_X1 U8430 ( .A1(n7572), .A2(n12924), .ZN(n7571) );
  AND2_X1 U8431 ( .A1(n8209), .A2(n13395), .ZN(n8208) );
  OR2_X1 U8432 ( .A1(n8212), .A2(n8210), .ZN(n8209) );
  INV_X1 U8433 ( .A(n11731), .ZN(n10133) );
  NAND2_X1 U8434 ( .A1(n7555), .A2(n13378), .ZN(n10189) );
  NOR2_X1 U8435 ( .A1(n13380), .A2(n7557), .ZN(n7556) );
  INV_X1 U8436 ( .A(n10181), .ZN(n7557) );
  NAND2_X1 U8437 ( .A1(n8207), .A2(n7488), .ZN(n8206) );
  INV_X1 U8438 ( .A(n13405), .ZN(n8207) );
  NAND2_X1 U8439 ( .A1(n9886), .A2(n13748), .ZN(n9899) );
  NAND2_X1 U8440 ( .A1(n7994), .A2(n7991), .ZN(n7990) );
  INV_X1 U8441 ( .A(n13267), .ZN(n7994) );
  NAND2_X1 U8442 ( .A1(n7984), .A2(n7982), .ZN(n7992) );
  NAND2_X1 U8443 ( .A1(n7986), .A2(n13267), .ZN(n7985) );
  NAND2_X1 U8444 ( .A1(n7988), .A2(n7987), .ZN(n7986) );
  NAND2_X1 U8445 ( .A1(n7995), .A2(n13207), .ZN(n7988) );
  AND2_X1 U8446 ( .A1(n7981), .A2(n7980), .ZN(n7989) );
  NAND2_X1 U8447 ( .A1(n7995), .A2(n13326), .ZN(n7981) );
  NAND2_X1 U8448 ( .A1(n7884), .A2(n7883), .ZN(n11777) );
  NAND2_X1 U8449 ( .A1(n7889), .A2(n7885), .ZN(n7884) );
  XNOR2_X1 U8450 ( .A(n8413), .B(n15917), .ZN(n15905) );
  NOR2_X1 U8451 ( .A1(n15938), .A2(n15937), .ZN(n15936) );
  XNOR2_X1 U8452 ( .A(n8472), .B(n7735), .ZN(n15957) );
  NOR2_X1 U8453 ( .A1(n15923), .A2(n8340), .ZN(n8419) );
  NOR2_X1 U8454 ( .A1(n15964), .A2(n15963), .ZN(n15962) );
  XNOR2_X1 U8455 ( .A(n8474), .B(n7737), .ZN(n15997) );
  OR2_X1 U8456 ( .A1(n15983), .A2(n8422), .ZN(n7599) );
  AND2_X1 U8457 ( .A1(n7919), .A2(n7918), .ZN(n8423) );
  NAND2_X1 U8458 ( .A1(n16011), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7918) );
  NOR2_X1 U8459 ( .A1(n16022), .A2(n8424), .ZN(n12543) );
  OAI21_X1 U8460 ( .B1(n16022), .B2(n7593), .A(n7592), .ZN(n8430) );
  NAND2_X1 U8461 ( .A1(n12542), .A2(n8429), .ZN(n7592) );
  OR2_X1 U8462 ( .A1(n8424), .A2(n7594), .ZN(n7593) );
  INV_X1 U8463 ( .A(n8429), .ZN(n7594) );
  XNOR2_X1 U8464 ( .A(n8479), .B(n8550), .ZN(n12234) );
  XNOR2_X1 U8465 ( .A(n8481), .B(n7734), .ZN(n12804) );
  NAND2_X1 U8466 ( .A1(n12804), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12803) );
  OR2_X1 U8467 ( .A1(n12806), .A2(n12807), .ZN(n13905) );
  NAND2_X1 U8468 ( .A1(n7589), .A2(n7431), .ZN(n7588) );
  AND2_X1 U8469 ( .A1(n13896), .A2(n8438), .ZN(n8439) );
  NAND2_X1 U8470 ( .A1(n13923), .A2(n8485), .ZN(n16045) );
  INV_X1 U8471 ( .A(n8483), .ZN(n8484) );
  OR2_X1 U8472 ( .A1(n16070), .A2(n16071), .ZN(n16067) );
  NAND2_X1 U8473 ( .A1(n7915), .A2(n8447), .ZN(n7914) );
  AOI21_X1 U8474 ( .B1(n7905), .B2(n7904), .A(n7903), .ZN(n7902) );
  INV_X1 U8475 ( .A(n13250), .ZN(n7903) );
  INV_X1 U8476 ( .A(n10083), .ZN(n7904) );
  OR2_X1 U8477 ( .A1(n9998), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U8478 ( .A1(n14029), .A2(n13253), .ZN(n14015) );
  AND2_X1 U8479 ( .A1(n13256), .A2(n13253), .ZN(n14030) );
  NAND2_X1 U8480 ( .A1(n8339), .A2(n14030), .ZN(n14029) );
  OR2_X1 U8481 ( .A1(n9948), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9960) );
  AND2_X1 U8482 ( .A1(n9923), .A2(n13556), .ZN(n9937) );
  INV_X1 U8483 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n13740) );
  AND4_X1 U8484 ( .A1(n9942), .A2(n9941), .A3(n9940), .A4(n9939), .ZN(n14089)
         );
  AND4_X1 U8485 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(n14109)
         );
  INV_X1 U8486 ( .A(n8232), .ZN(n8231) );
  AND2_X1 U8487 ( .A1(n9905), .A2(n8230), .ZN(n8229) );
  AND2_X1 U8488 ( .A1(n13132), .A2(n13129), .ZN(n14116) );
  NAND2_X1 U8489 ( .A1(n9878), .A2(n9877), .ZN(n14141) );
  OR2_X1 U8490 ( .A1(n9846), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U8491 ( .A1(n9859), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9871) );
  AOI21_X1 U8492 ( .B1(n7893), .B2(n7895), .A(n7892), .ZN(n7891) );
  INV_X1 U8493 ( .A(n7894), .ZN(n7893) );
  OR2_X1 U8494 ( .A1(n9807), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U8495 ( .A1(n9818), .A2(n10155), .ZN(n12915) );
  AND2_X1 U8496 ( .A1(n13190), .A2(n13188), .ZN(n13312) );
  AOI21_X1 U8497 ( .B1(n9768), .B2(n8236), .A(n8233), .ZN(n12760) );
  NAND2_X1 U8498 ( .A1(n8234), .A2(n7432), .ZN(n8233) );
  AND2_X1 U8499 ( .A1(n7405), .A2(n9794), .ZN(n8236) );
  NAND2_X1 U8500 ( .A1(n9783), .A2(n13551), .ZN(n9795) );
  INV_X1 U8501 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n13551) );
  AND4_X1 U8502 ( .A1(n9800), .A2(n9799), .A3(n9798), .A4(n9797), .ZN(n12696)
         );
  NAND2_X1 U8503 ( .A1(n12409), .A2(n9782), .ZN(n12587) );
  INV_X1 U8504 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n13737) );
  NOR2_X1 U8505 ( .A1(n9756), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9769) );
  OR2_X1 U8506 ( .A1(n9744), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9756) );
  NAND2_X1 U8507 ( .A1(n8225), .A2(n9728), .ZN(n12323) );
  NOR2_X1 U8508 ( .A1(n13308), .A2(n12122), .ZN(n9714) );
  NAND2_X1 U8509 ( .A1(n7901), .A2(n10065), .ZN(n16174) );
  INV_X1 U8510 ( .A(n16177), .ZN(n10066) );
  INV_X1 U8511 ( .A(n14257), .ZN(n7568) );
  NAND2_X1 U8512 ( .A1(n7897), .A2(n9929), .ZN(n7896) );
  NAND2_X1 U8513 ( .A1(n7900), .A2(n10080), .ZN(n14066) );
  AND2_X1 U8514 ( .A1(n9910), .A2(n9909), .ZN(n10175) );
  NAND2_X1 U8515 ( .A1(n12917), .A2(n13194), .ZN(n13016) );
  NAND2_X1 U8516 ( .A1(n12919), .A2(n12918), .ZN(n12917) );
  AND3_X1 U8517 ( .A1(n9805), .A2(n9804), .A3(n9803), .ZN(n16411) );
  INV_X1 U8518 ( .A(n12128), .ZN(n16234) );
  INV_X1 U8519 ( .A(n8228), .ZN(n13307) );
  NOR2_X1 U8520 ( .A1(n10234), .A2(n10236), .ZN(n10224) );
  INV_X1 U8521 ( .A(n16467), .ZN(n16410) );
  AND2_X1 U8522 ( .A1(n10030), .A2(n10029), .ZN(n13270) );
  INV_X1 U8523 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8454) );
  INV_X1 U8524 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7577) );
  AND2_X1 U8525 ( .A1(n15553), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9669) );
  XNOR2_X1 U8526 ( .A(n8354), .B(n8353), .ZN(n8464) );
  OAI21_X1 U8527 ( .B1(n8450), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U8528 ( .A1(n8352), .A2(n8356), .ZN(n8450) );
  INV_X1 U8529 ( .A(n8452), .ZN(n8352) );
  AOI21_X1 U8530 ( .B1(n7999), .B2(n8001), .A(n7509), .ZN(n7997) );
  NAND2_X1 U8531 ( .A1(n9653), .A2(n9652), .ZN(n9856) );
  NAND2_X1 U8532 ( .A1(n7975), .A2(n7974), .ZN(n9826) );
  AOI21_X1 U8533 ( .B1(n7977), .B2(n7979), .A(n7497), .ZN(n7974) );
  NOR2_X1 U8534 ( .A1(n8387), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8382) );
  NOR2_X1 U8535 ( .A1(n8185), .A2(n8184), .ZN(n8393) );
  OR2_X1 U8536 ( .A1(n8417), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8399) );
  XNOR2_X1 U8537 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9736) );
  AOI21_X1 U8538 ( .B1(n8004), .B2(n9708), .A(n7453), .ZN(n8003) );
  XNOR2_X1 U8539 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9722) );
  AND2_X1 U8540 ( .A1(n9629), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9682) );
  OR2_X1 U8541 ( .A1(n14436), .A2(n14338), .ZN(n8046) );
  INV_X1 U8542 ( .A(n10853), .ZN(n10854) );
  OR2_X1 U8543 ( .A1(n10408), .A2(n12791), .ZN(n10415) );
  NAND2_X1 U8544 ( .A1(n10252), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10422) );
  INV_X1 U8545 ( .A(n10415), .ZN(n10252) );
  NOR2_X1 U8546 ( .A1(n8063), .A2(n7615), .ZN(n7614) );
  INV_X1 U8547 ( .A(n10911), .ZN(n7615) );
  XNOR2_X1 U8548 ( .A(n14645), .B(n10853), .ZN(n14358) );
  AOI21_X1 U8549 ( .B1(n8049), .B2(n7627), .A(n7452), .ZN(n7626) );
  INV_X1 U8550 ( .A(n8053), .ZN(n7627) );
  NAND2_X1 U8551 ( .A1(n10783), .A2(n10784), .ZN(n10785) );
  AND2_X1 U8552 ( .A1(n10493), .A2(n10492), .ZN(n14369) );
  NAND2_X1 U8553 ( .A1(n8912), .A2(n10761), .ZN(n14480) );
  INV_X1 U8554 ( .A(n10817), .ZN(n10552) );
  INV_X1 U8555 ( .A(n14490), .ZN(n8912) );
  AND2_X1 U8556 ( .A1(n8903), .A2(n8902), .ZN(n14493) );
  NOR2_X1 U8557 ( .A1(n7750), .A2(n14573), .ZN(n14507) );
  AND2_X1 U8558 ( .A1(n10487), .A2(n10471), .ZN(n14524) );
  AOI21_X1 U8559 ( .B1(n14557), .B2(n10457), .A(n7376), .ZN(n7946) );
  NOR2_X1 U8560 ( .A1(n14573), .A2(n10455), .ZN(n14549) );
  INV_X1 U8561 ( .A(n7855), .ZN(n7854) );
  NAND2_X1 U8562 ( .A1(n8871), .A2(n14777), .ZN(n14584) );
  AOI21_X1 U8563 ( .B1(n14608), .B2(n7950), .A(n7948), .ZN(n14566) );
  OAI21_X1 U8564 ( .B1(n7951), .B2(n7949), .A(n7442), .ZN(n7948) );
  AND2_X1 U8565 ( .A1(n7406), .A2(n14583), .ZN(n7950) );
  XNOR2_X1 U8566 ( .A(n14721), .B(n14582), .ZN(n14569) );
  OR2_X1 U8567 ( .A1(n10435), .A2(n10938), .ZN(n10437) );
  INV_X1 U8568 ( .A(n14598), .ZN(n8871) );
  OR2_X1 U8569 ( .A1(n7746), .A2(n14739), .ZN(n14612) );
  AOI21_X1 U8570 ( .B1(n14651), .B2(n10431), .A(n8333), .ZN(n14621) );
  INV_X1 U8571 ( .A(n14788), .ZN(n7745) );
  NAND2_X1 U8572 ( .A1(n12935), .A2(n14788), .ZN(n14642) );
  INV_X1 U8573 ( .A(n7866), .ZN(n7865) );
  AOI21_X1 U8574 ( .B1(n7866), .B2(n7869), .A(n7375), .ZN(n7864) );
  NOR2_X1 U8575 ( .A1(n12742), .A2(n7867), .ZN(n7866) );
  NAND2_X1 U8576 ( .A1(n7935), .A2(n7933), .ZN(n12943) );
  AOI21_X1 U8577 ( .B1(n7936), .B2(n7939), .A(n7934), .ZN(n7933) );
  INV_X1 U8578 ( .A(n7940), .ZN(n7939) );
  OR2_X1 U8579 ( .A1(n14666), .A2(n12662), .ZN(n12663) );
  NAND2_X1 U8580 ( .A1(n10249), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10383) );
  INV_X1 U8581 ( .A(n7957), .ZN(n7956) );
  AOI21_X1 U8582 ( .B1(n7957), .B2(n7955), .A(n7954), .ZN(n7953) );
  NAND2_X1 U8583 ( .A1(n7749), .A2(n12213), .ZN(n12423) );
  AND3_X1 U8584 ( .A1(n7749), .A2(n12213), .A3(n7748), .ZN(n12503) );
  NAND2_X1 U8585 ( .A1(n12213), .A2(n16434), .ZN(n12250) );
  OR2_X1 U8586 ( .A1(n10343), .A2(n11509), .ZN(n10352) );
  OR2_X1 U8587 ( .A1(n12083), .A2(n12058), .ZN(n12197) );
  NOR2_X1 U8588 ( .A1(n16400), .A2(n12197), .ZN(n12213) );
  NAND2_X1 U8589 ( .A1(n12084), .A2(n16360), .ZN(n12083) );
  NOR2_X1 U8590 ( .A1(n12099), .A2(n11906), .ZN(n12084) );
  NAND2_X1 U8591 ( .A1(n10316), .A2(n10315), .ZN(n12104) );
  NAND2_X1 U8592 ( .A1(n7510), .A2(n16323), .ZN(n12099) );
  OAI21_X1 U8593 ( .B1(n16253), .B2(n16254), .A(n10307), .ZN(n11857) );
  NOR2_X1 U8594 ( .A1(n16260), .A2(n16270), .ZN(n16264) );
  XNOR2_X1 U8595 ( .A(n16270), .B(n11695), .ZN(n16254) );
  NAND2_X1 U8596 ( .A1(n16213), .A2(n16214), .ZN(n16260) );
  NOR2_X1 U8597 ( .A1(n11752), .A2(n16106), .ZN(n16213) );
  INV_X1 U8598 ( .A(n10988), .ZN(n7925) );
  INV_X1 U8599 ( .A(n14493), .ZN(n14695) );
  NOR2_X1 U8600 ( .A1(n14529), .A2(n7848), .ZN(n7847) );
  INV_X1 U8601 ( .A(n10548), .ZN(n7848) );
  NAND2_X1 U8602 ( .A1(n7849), .A2(n10548), .ZN(n14530) );
  AND3_X1 U8603 ( .A1(n15564), .A2(n11739), .A3(n8987), .ZN(n10556) );
  XNOR2_X1 U8604 ( .A(n8975), .B(n8974), .ZN(n10935) );
  INV_X1 U8605 ( .A(n8957), .ZN(n11102) );
  NAND2_X1 U8606 ( .A1(n8960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8968) );
  OR2_X1 U8607 ( .A1(n8973), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8960) );
  INV_X1 U8608 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8967) );
  INV_X1 U8609 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8938) );
  OR2_X1 U8610 ( .A1(n8791), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8782) );
  AND2_X1 U8611 ( .A1(n8799), .A2(n8661), .ZN(n8801) );
  NAND2_X1 U8612 ( .A1(n8660), .A2(n8659), .ZN(n8821) );
  INV_X1 U8613 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8660) );
  INV_X1 U8614 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8659) );
  INV_X1 U8615 ( .A(n11874), .ZN(n8131) );
  OR2_X1 U8616 ( .A1(n9247), .A2(n9246), .ZN(n9263) );
  AND2_X1 U8617 ( .A1(n9200), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9213) );
  OAI21_X1 U8618 ( .B1(n7399), .B2(n8130), .A(n7660), .ZN(n12169) );
  INV_X1 U8619 ( .A(n12167), .ZN(n8130) );
  NAND2_X1 U8620 ( .A1(n8129), .A2(n11711), .ZN(n7660) );
  AND2_X1 U8621 ( .A1(n8137), .A2(n12167), .ZN(n8129) );
  NAND2_X1 U8622 ( .A1(n12169), .A2(n12170), .ZN(n12362) );
  INV_X1 U8623 ( .A(n7684), .ZN(n7683) );
  AND2_X1 U8624 ( .A1(n7681), .A2(n15027), .ZN(n7680) );
  NAND2_X1 U8625 ( .A1(n7684), .A2(n7682), .ZN(n7681) );
  NAND2_X1 U8626 ( .A1(n15052), .A2(n7687), .ZN(n7686) );
  AND2_X1 U8627 ( .A1(n15052), .A2(n14972), .ZN(n7688) );
  INV_X1 U8628 ( .A(n8107), .ZN(n11082) );
  NAND2_X1 U8629 ( .A1(n11036), .A2(n8110), .ZN(n11041) );
  NAND2_X1 U8630 ( .A1(n14955), .A2(n11565), .ZN(n8110) );
  NAND2_X1 U8631 ( .A1(n15085), .A2(n14891), .ZN(n14991) );
  NAND2_X1 U8632 ( .A1(n7665), .A2(n7398), .ZN(n14970) );
  OAI21_X1 U8633 ( .B1(n15085), .B2(n7664), .A(n7661), .ZN(n7665) );
  INV_X1 U8634 ( .A(n9437), .ZN(n9454) );
  INV_X1 U8635 ( .A(n8160), .ZN(n7677) );
  AOI21_X1 U8636 ( .B1(n8160), .B2(n7676), .A(n7675), .ZN(n7674) );
  INV_X1 U8637 ( .A(n14852), .ZN(n7675) );
  INV_X1 U8638 ( .A(n9465), .ZN(n7550) );
  AND4_X1 U8639 ( .A1(n9432), .A2(n9431), .A3(n9430), .A4(n9429), .ZN(n14833)
         );
  OR2_X1 U8640 ( .A1(n9386), .A2(n9043), .ZN(n9044) );
  NOR2_X1 U8641 ( .A1(n7428), .A2(n7373), .ZN(n8298) );
  NAND2_X1 U8642 ( .A1(n15187), .A2(n15186), .ZN(n15185) );
  AND2_X1 U8643 ( .A1(n15209), .A2(n11360), .ZN(n11363) );
  NAND2_X1 U8644 ( .A1(n11363), .A2(n11362), .ZN(n15717) );
  NAND2_X1 U8645 ( .A1(n11669), .A2(n11611), .ZN(n12304) );
  AOI21_X1 U8646 ( .B1(n12609), .B2(P1_REG1_REG_16__SCAN_IN), .A(n12608), .ZN(
        n12611) );
  XNOR2_X1 U8647 ( .A(n15217), .B(n7542), .ZN(n12972) );
  NOR2_X1 U8648 ( .A1(n12969), .A2(n7543), .ZN(n15217) );
  AND2_X1 U8649 ( .A1(n12970), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7543) );
  NAND2_X1 U8650 ( .A1(n9472), .A2(n9471), .ZN(n9583) );
  NAND2_X1 U8651 ( .A1(n9483), .A2(n9482), .ZN(n15241) );
  NOR2_X1 U8652 ( .A1(n15284), .A2(n7773), .ZN(n15242) );
  NAND2_X1 U8653 ( .A1(n15257), .A2(n7774), .ZN(n7773) );
  NOR2_X1 U8654 ( .A1(n7775), .A2(n13075), .ZN(n7774) );
  AOI21_X1 U8655 ( .B1(n15247), .B2(n7392), .A(n8258), .ZN(n8257) );
  OAI22_X1 U8656 ( .A1(n7717), .A2(n7716), .B1(n7719), .B2(n13344), .ZN(n7715)
         );
  NAND2_X1 U8657 ( .A1(n7724), .A2(n7725), .ZN(n15248) );
  NAND2_X1 U8658 ( .A1(n15277), .A2(n7371), .ZN(n7724) );
  NOR2_X1 U8659 ( .A1(n7380), .A2(n7640), .ZN(n7639) );
  INV_X1 U8660 ( .A(n13057), .ZN(n7640) );
  INV_X1 U8661 ( .A(n8266), .ZN(n15301) );
  NAND2_X1 U8662 ( .A1(n7768), .A2(n15299), .ZN(n15293) );
  INV_X1 U8663 ( .A(n7768), .ZN(n15308) );
  AOI21_X1 U8664 ( .B1(n7793), .B2(n7792), .A(n7454), .ZN(n7791) );
  INV_X1 U8665 ( .A(n7397), .ZN(n7792) );
  NAND2_X1 U8666 ( .A1(n7646), .A2(n7793), .ZN(n7645) );
  INV_X1 U8667 ( .A(n9400), .ZN(n9017) );
  OAI21_X1 U8668 ( .B1(n8269), .B2(n8343), .A(n8267), .ZN(n15346) );
  NAND2_X1 U8669 ( .A1(n15377), .A2(n8268), .ZN(n8267) );
  AND2_X1 U8670 ( .A1(n8271), .A2(n15378), .ZN(n8268) );
  NOR2_X1 U8671 ( .A1(n13067), .A2(n8270), .ZN(n8269) );
  INV_X1 U8672 ( .A(n13066), .ZN(n8270) );
  NOR2_X1 U8673 ( .A1(n9319), .A2(n9318), .ZN(n9351) );
  NAND2_X1 U8674 ( .A1(n15377), .A2(n15378), .ZN(n15376) );
  OR2_X1 U8675 ( .A1(n15404), .A2(n15508), .ZN(n15384) );
  OR2_X1 U8676 ( .A1(n9303), .A2(n9302), .ZN(n9319) );
  NAND2_X1 U8677 ( .A1(n12676), .A2(n12677), .ZN(n12678) );
  NAND2_X1 U8678 ( .A1(n9213), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9234) );
  OR2_X1 U8679 ( .A1(n9234), .A2(n9233), .ZN(n9247) );
  NOR2_X1 U8680 ( .A1(n12350), .A2(n12642), .ZN(n12461) );
  OR2_X1 U8681 ( .A1(n9170), .A2(n12174), .ZN(n9184) );
  INV_X1 U8682 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U8683 ( .A1(n7765), .A2(n7764), .ZN(n12273) );
  INV_X1 U8684 ( .A(n12183), .ZN(n7764) );
  NAND2_X1 U8685 ( .A1(n12184), .A2(n16374), .ZN(n12183) );
  AND2_X1 U8686 ( .A1(n12069), .A2(n16351), .ZN(n12184) );
  INV_X1 U8687 ( .A(n8252), .ZN(n8251) );
  AND2_X1 U8688 ( .A1(n8249), .A2(n11825), .ZN(n8248) );
  AND2_X1 U8689 ( .A1(n11063), .A2(n11285), .ZN(n15100) );
  NOR2_X1 U8690 ( .A1(n12045), .A2(n14985), .ZN(n12044) );
  OAI21_X1 U8691 ( .B1(n16139), .B2(n16143), .A(n8272), .ZN(n11794) );
  NAND3_X1 U8692 ( .A1(n9047), .A2(n8299), .A3(n8298), .ZN(n16143) );
  NAND2_X1 U8693 ( .A1(n9342), .A2(n9341), .ZN(n15500) );
  OR2_X1 U8694 ( .A1(n12337), .A2(n9481), .ZN(n9342) );
  NAND2_X1 U8695 ( .A1(n11798), .A2(n11060), .ZN(n16528) );
  INV_X1 U8696 ( .A(n16528), .ZN(n16448) );
  NAND2_X1 U8697 ( .A1(n9596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9597) );
  AND2_X1 U8698 ( .A1(n9008), .A2(n9010), .ZN(n7777) );
  NAND2_X1 U8699 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n7780), .ZN(n7779) );
  NAND2_X1 U8700 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n7780) );
  AOI21_X1 U8701 ( .B1(n8916), .B2(n8915), .A(n8914), .ZN(n8919) );
  OAI21_X1 U8702 ( .B1(n8901), .B2(n8900), .A(n8899), .ZN(n8905) );
  XNOR2_X1 U8703 ( .A(n8891), .B(n8890), .ZN(n13086) );
  NAND2_X1 U8704 ( .A1(n8889), .A2(n8888), .ZN(n8891) );
  INV_X1 U8705 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9602) );
  XNOR2_X1 U8706 ( .A(n9607), .B(P1_IR_REG_24__SCAN_IN), .ZN(n11056) );
  XNOR2_X1 U8707 ( .A(n8681), .B(n8875), .ZN(n14817) );
  INV_X1 U8708 ( .A(n9489), .ZN(n9488) );
  XNOR2_X1 U8709 ( .A(n8688), .B(n8689), .ZN(n12874) );
  NAND2_X1 U8710 ( .A1(n8634), .A2(n8635), .ZN(n7552) );
  INV_X1 U8711 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n13871) );
  AND2_X1 U8712 ( .A1(n8089), .A2(n8094), .ZN(n8851) );
  AND2_X1 U8713 ( .A1(n8096), .A2(n8618), .ZN(n8090) );
  NAND2_X1 U8714 ( .A1(n8088), .A2(n8615), .ZN(n8842) );
  OR2_X1 U8715 ( .A1(n9152), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U8716 ( .A1(n8761), .A2(n8605), .ZN(n8829) );
  OAI21_X1 U8717 ( .B1(n8591), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n7530), .ZN(
        n8586) );
  NAND2_X1 U8718 ( .A1(n8591), .A2(n9629), .ZN(n7530) );
  AND2_X1 U8719 ( .A1(n7962), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15735) );
  INV_X1 U8720 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7962) );
  INV_X1 U8721 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15730) );
  XNOR2_X1 U8722 ( .A(n15734), .B(n15735), .ZN(n15736) );
  OAI22_X1 U8723 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n15775), .B1(n15774), .B2(
        n15773), .ZN(n15777) );
  NOR2_X1 U8724 ( .A1(n15786), .A2(n15787), .ZN(n15788) );
  AOI21_X1 U8725 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15796), .A(n15795), .ZN(
        n15804) );
  NOR2_X1 U8726 ( .A1(n15794), .A2(n15793), .ZN(n15795) );
  OAI21_X1 U8727 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n15814), .A(n15813), .ZN(
        n15819) );
  AOI22_X1 U8728 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n15839), .B1(n15838), 
        .B2(n15837), .ZN(n15846) );
  NAND2_X1 U8729 ( .A1(n7575), .A2(n10162), .ZN(n13000) );
  AND2_X1 U8730 ( .A1(n12509), .A2(n10149), .ZN(n12601) );
  NAND2_X1 U8731 ( .A1(n11661), .A2(n11660), .ZN(n11659) );
  NAND2_X1 U8732 ( .A1(n8202), .A2(n8203), .ZN(n13372) );
  AOI21_X1 U8733 ( .B1(n8205), .B2(n8204), .A(n7492), .ZN(n8203) );
  NAND2_X1 U8734 ( .A1(n12224), .A2(n12223), .ZN(n12222) );
  NAND2_X1 U8735 ( .A1(n10182), .A2(n10181), .ZN(n13382) );
  NAND2_X1 U8736 ( .A1(n12693), .A2(n10156), .ZN(n12776) );
  NAND2_X1 U8737 ( .A1(n11659), .A2(n10132), .ZN(n11730) );
  NAND2_X1 U8738 ( .A1(n12222), .A2(n10147), .ZN(n12511) );
  AND4_X1 U8739 ( .A1(n9916), .A2(n9915), .A3(n9914), .A4(n9913), .ZN(n14122)
         );
  OAI21_X1 U8740 ( .B1(n12776), .B2(n12773), .A(n12772), .ZN(n12925) );
  AND4_X1 U8741 ( .A1(n9824), .A2(n9823), .A3(n9822), .A4(n9821), .ZN(n12928)
         );
  OR2_X1 U8742 ( .A1(n10227), .A2(n10225), .ZN(n13451) );
  NAND2_X1 U8743 ( .A1(n11412), .A2(n10125), .ZN(n11643) );
  AND4_X1 U8744 ( .A1(n9891), .A2(n9890), .A3(n9889), .A4(n9888), .ZN(n14147)
         );
  AND2_X1 U8745 ( .A1(n8206), .A2(n7409), .ZN(n13440) );
  NAND2_X1 U8746 ( .A1(n8206), .A2(n8205), .ZN(n13438) );
  AND2_X1 U8747 ( .A1(n10139), .A2(n10138), .ZN(n8217) );
  NAND2_X1 U8748 ( .A1(n8218), .A2(n10138), .ZN(n11993) );
  INV_X1 U8749 ( .A(n8190), .ZN(n13448) );
  NAND2_X1 U8750 ( .A1(n13389), .A2(n8201), .ZN(n8192) );
  NOR2_X1 U8751 ( .A1(n7374), .A2(n10198), .ZN(n8191) );
  NAND2_X1 U8752 ( .A1(n8211), .A2(n8212), .ZN(n13037) );
  NOR2_X1 U8753 ( .A1(n12999), .A2(n8342), .ZN(n13039) );
  NAND2_X1 U8754 ( .A1(n11411), .A2(n13341), .ZN(n13454) );
  AND2_X1 U8755 ( .A1(n11990), .A2(n10041), .ZN(n13974) );
  INV_X1 U8756 ( .A(n13999), .ZN(n13461) );
  INV_X1 U8757 ( .A(n14010), .ZN(n13462) );
  OAI211_X1 U8758 ( .C1(n9964), .C2(n14267), .A(n9963), .B(n9962), .ZN(n14056)
         );
  INV_X1 U8759 ( .A(n14073), .ZN(n14041) );
  INV_X1 U8760 ( .A(n14089), .ZN(n14055) );
  INV_X1 U8761 ( .A(n14109), .ZN(n13464) );
  INV_X1 U8762 ( .A(n14122), .ZN(n13442) );
  INV_X1 U8763 ( .A(n14146), .ZN(n13027) );
  OR2_X1 U8764 ( .A1(n14306), .A2(n10217), .ZN(n13471) );
  NAND2_X1 U8765 ( .A1(n7370), .A2(n16202), .ZN(n8407) );
  AND2_X1 U8766 ( .A1(n15905), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n15906) );
  AND2_X1 U8767 ( .A1(n7585), .A2(n7584), .ZN(n15923) );
  INV_X1 U8768 ( .A(n15924), .ZN(n7584) );
  INV_X1 U8769 ( .A(n7585), .ZN(n15925) );
  XNOR2_X1 U8770 ( .A(n8419), .B(n7735), .ZN(n15944) );
  INV_X1 U8771 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15982) );
  INV_X1 U8772 ( .A(n7591), .ZN(n15967) );
  INV_X1 U8773 ( .A(n7917), .ZN(n15965) );
  XNOR2_X1 U8774 ( .A(n8421), .B(n7737), .ZN(n15984) );
  NOR2_X1 U8775 ( .A1(n15984), .A2(n15985), .ZN(n15983) );
  INV_X1 U8776 ( .A(n7919), .ZN(n16002) );
  INV_X1 U8777 ( .A(n7599), .ZN(n16004) );
  NOR2_X1 U8778 ( .A1(n16024), .A2(n16023), .ZN(n16022) );
  XNOR2_X1 U8779 ( .A(n8423), .B(n8537), .ZN(n16023) );
  NAND2_X1 U8780 ( .A1(n12540), .A2(n12539), .ZN(n12538) );
  XNOR2_X1 U8781 ( .A(n8430), .B(n8550), .ZN(n12230) );
  NOR2_X1 U8782 ( .A1(n12229), .A2(n8431), .ZN(n12519) );
  NOR2_X1 U8783 ( .A1(n12519), .A2(n12518), .ZN(n12517) );
  INV_X1 U8784 ( .A(n7588), .ZN(n13899) );
  XNOR2_X1 U8785 ( .A(n8439), .B(n11075), .ZN(n13918) );
  NOR2_X1 U8786 ( .A1(n13918), .A2(n13919), .ZN(n13917) );
  OAI21_X1 U8787 ( .B1(n13918), .B2(n7596), .A(n7595), .ZN(n16056) );
  NAND2_X1 U8788 ( .A1(n7597), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U8789 ( .A1(n8440), .A2(n7597), .ZN(n7595) );
  INV_X1 U8790 ( .A(n16055), .ZN(n7597) );
  NAND2_X1 U8791 ( .A1(n7511), .A2(n7914), .ZN(n7913) );
  AND2_X1 U8792 ( .A1(n14013), .A2(n14012), .ZN(n14187) );
  NAND2_X1 U8793 ( .A1(n9936), .A2(n9935), .ZN(n14202) );
  NAND2_X1 U8794 ( .A1(n9922), .A2(n9921), .ZN(n14205) );
  NAND2_X1 U8795 ( .A1(n8221), .A2(n9853), .ZN(n14155) );
  NAND2_X1 U8796 ( .A1(n13025), .A2(n9852), .ZN(n8221) );
  NAND2_X1 U8797 ( .A1(n9845), .A2(n9844), .ZN(n14236) );
  INV_X1 U8798 ( .A(n12782), .ZN(n16468) );
  NAND2_X1 U8799 ( .A1(n7559), .A2(n13181), .ZN(n12757) );
  NAND2_X1 U8800 ( .A1(n12412), .A2(n13175), .ZN(n12586) );
  AND2_X1 U8801 ( .A1(n9768), .A2(n9767), .ZN(n12410) );
  AND3_X1 U8802 ( .A1(n9766), .A2(n9765), .A3(n9764), .ZN(n12449) );
  NAND2_X1 U8803 ( .A1(n11922), .A2(n16129), .ZN(n14166) );
  AOI21_X1 U8804 ( .B1(n14308), .B2(n10032), .A(n7507), .ZN(n14173) );
  INV_X1 U8805 ( .A(n16556), .ZN(n14176) );
  INV_X1 U8806 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8238) );
  INV_X1 U8807 ( .A(n16473), .ZN(n16470) );
  INV_X1 U8808 ( .A(n14173), .ZN(n16559) );
  AND2_X1 U8809 ( .A1(n9968), .A2(n9967), .ZN(n14265) );
  INV_X1 U8810 ( .A(n13367), .ZN(n14269) );
  INV_X1 U8811 ( .A(n10175), .ZN(n14287) );
  INV_X1 U8812 ( .A(n10028), .ZN(n10026) );
  XNOR2_X1 U8813 ( .A(n8363), .B(P3_IR_REG_26__SCAN_IN), .ZN(n12880) );
  INV_X1 U8814 ( .A(SI_25_), .ZN(n13680) );
  AND2_X1 U8815 ( .A1(n8367), .A2(n8366), .ZN(n12633) );
  NAND2_X1 U8816 ( .A1(n8370), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8365) );
  INV_X1 U8817 ( .A(SI_24_), .ZN(n13681) );
  NAND2_X1 U8818 ( .A1(n8371), .A2(n8370), .ZN(n12537) );
  NAND2_X1 U8819 ( .A1(n8374), .A2(n8361), .ZN(n8368) );
  INV_X1 U8820 ( .A(SI_23_), .ZN(n12149) );
  NAND2_X1 U8821 ( .A1(n8018), .A2(n7501), .ZN(n9956) );
  OR2_X1 U8822 ( .A1(n7531), .A2(n8023), .ZN(n8018) );
  AOI21_X1 U8823 ( .B1(n7531), .B2(n9663), .A(n8027), .ZN(n9945) );
  XNOR2_X1 U8824 ( .A(n8453), .B(n8356), .ZN(n11932) );
  INV_X1 U8825 ( .A(SI_20_), .ZN(n13668) );
  INV_X1 U8826 ( .A(SI_18_), .ZN(n11374) );
  NAND2_X1 U8827 ( .A1(n7998), .A2(n9655), .ZN(n9882) );
  NAND2_X1 U8828 ( .A1(n9867), .A2(n9865), .ZN(n7998) );
  INV_X1 U8829 ( .A(SI_12_), .ZN(n13699) );
  NAND2_X1 U8830 ( .A1(n7976), .A2(n9645), .ZN(n9814) );
  NAND2_X1 U8831 ( .A1(n9802), .A2(n9801), .ZN(n7976) );
  INV_X1 U8832 ( .A(n7971), .ZN(n9790) );
  AOI21_X1 U8833 ( .B1(n9776), .B2(n9775), .A(n7393), .ZN(n7971) );
  NAND2_X1 U8834 ( .A1(n7496), .A2(n8180), .ZN(n8390) );
  INV_X1 U8835 ( .A(SI_8_), .ZN(n13705) );
  INV_X1 U8836 ( .A(n9778), .ZN(n16011) );
  NAND2_X1 U8837 ( .A1(n8005), .A2(n9631), .ZN(n9710) );
  NAND2_X1 U8838 ( .A1(n14435), .A2(n7402), .ZN(n7603) );
  OAI21_X1 U8839 ( .B1(n14368), .B2(n7443), .A(n7605), .ZN(n7604) );
  NAND2_X1 U8840 ( .A1(n14368), .A2(n14339), .ZN(n7605) );
  NAND2_X1 U8841 ( .A1(n7607), .A2(n14339), .ZN(n7606) );
  INV_X1 U8842 ( .A(n14368), .ZN(n7607) );
  OAI21_X1 U8843 ( .B1(n14435), .B2(n8047), .A(n8044), .ZN(n8048) );
  OR2_X1 U8844 ( .A1(n14368), .A2(n14338), .ZN(n8047) );
  INV_X1 U8845 ( .A(n8045), .ZN(n8044) );
  OAI22_X1 U8846 ( .A1(n14368), .A2(n8046), .B1(n14366), .B2(n14367), .ZN(
        n8045) );
  NAND2_X1 U8847 ( .A1(n8724), .A2(n8723), .ZN(n12795) );
  NAND2_X1 U8848 ( .A1(n10867), .A2(n11422), .ZN(n11429) );
  NAND2_X1 U8849 ( .A1(n10912), .A2(n12909), .ZN(n12914) );
  NAND2_X1 U8850 ( .A1(n12789), .A2(n10911), .ZN(n10912) );
  NAND2_X1 U8851 ( .A1(n10953), .A2(n8056), .ZN(n11704) );
  AND2_X1 U8852 ( .A1(n11699), .A2(n10863), .ZN(n8056) );
  NAND2_X1 U8853 ( .A1(n11632), .A2(n10879), .ZN(n10880) );
  OR2_X1 U8854 ( .A1(n14427), .A2(n16261), .ZN(n14398) );
  NAND2_X1 U8855 ( .A1(n7611), .A2(n7609), .ZN(n7608) );
  AND2_X1 U8856 ( .A1(n8060), .A2(n7417), .ZN(n7609) );
  NAND2_X1 U8857 ( .A1(n8059), .A2(n7613), .ZN(n14401) );
  NAND2_X1 U8858 ( .A1(n12789), .A2(n7614), .ZN(n7613) );
  OR2_X1 U8859 ( .A1(n11400), .A2(n8923), .ZN(n8748) );
  XNOR2_X1 U8860 ( .A(n14325), .B(n14326), .ZN(n14412) );
  NAND2_X1 U8861 ( .A1(n7617), .A2(n7619), .ZN(n10947) );
  NAND2_X1 U8862 ( .A1(n7602), .A2(n11765), .ZN(n11771) );
  NAND2_X1 U8863 ( .A1(n11764), .A2(n10858), .ZN(n7602) );
  NAND2_X1 U8864 ( .A1(n12914), .A2(n10916), .ZN(n14429) );
  NAND2_X1 U8865 ( .A1(n11429), .A2(n10871), .ZN(n11655) );
  NAND2_X1 U8866 ( .A1(n14435), .A2(n14436), .ZN(n14434) );
  AND2_X1 U8867 ( .A1(n10940), .A2(n10926), .ZN(n14437) );
  NAND2_X1 U8868 ( .A1(n7624), .A2(n7626), .ZN(n12899) );
  NAND2_X1 U8869 ( .A1(n11143), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14442) );
  NOR3_X1 U8870 ( .A1(n10826), .A2(n10825), .A3(n13010), .ZN(n10827) );
  NOR4_X1 U8871 ( .A1(n10821), .A2(n14538), .A3(n14513), .A4(n10820), .ZN(
        n10823) );
  INV_X1 U8872 ( .A(n12739), .ZN(n10930) );
  NAND4_X1 U8873 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n14471) );
  NAND2_X1 U8874 ( .A1(n10302), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n10299) );
  NAND4_X2 U8875 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n14475) );
  NAND2_X1 U8876 ( .A1(n10506), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10288) );
  INV_X1 U8877 ( .A(n12843), .ZN(n12849) );
  NAND2_X1 U8878 ( .A1(n14512), .A2(n7873), .ZN(n14498) );
  AND2_X1 U8879 ( .A1(n14512), .A2(n10551), .ZN(n14500) );
  NAND2_X1 U8880 ( .A1(n7944), .A2(n10484), .ZN(n14486) );
  INV_X1 U8881 ( .A(n14700), .ZN(n14511) );
  OR3_X1 U8882 ( .A1(n14523), .A2(n14522), .A3(n14491), .ZN(n14707) );
  NAND2_X1 U8883 ( .A1(n14554), .A2(n10457), .ZN(n14535) );
  NAND2_X1 U8884 ( .A1(n7947), .A2(n7951), .ZN(n14579) );
  NAND2_X1 U8885 ( .A1(n14608), .A2(n7406), .ZN(n7947) );
  NAND2_X1 U8886 ( .A1(n14605), .A2(n7857), .ZN(n7852) );
  AND2_X1 U8887 ( .A1(n14607), .A2(n10434), .ZN(n14594) );
  NAND2_X1 U8888 ( .A1(n7859), .A2(n7862), .ZN(n14592) );
  NAND2_X1 U8889 ( .A1(n7861), .A2(n7860), .ZN(n7859) );
  NAND2_X1 U8890 ( .A1(n14640), .A2(n10537), .ZN(n14622) );
  NAND2_X1 U8891 ( .A1(n12622), .A2(n10535), .ZN(n12741) );
  AND2_X1 U8892 ( .A1(n7941), .A2(n7413), .ZN(n12628) );
  NAND2_X1 U8893 ( .A1(n7959), .A2(n10367), .ZN(n12244) );
  NAND2_X1 U8894 ( .A1(n10359), .A2(n10358), .ZN(n12210) );
  NAND2_X1 U8895 ( .A1(n12081), .A2(n10523), .ZN(n11892) );
  NAND2_X1 U8896 ( .A1(n11746), .A2(n12843), .ZN(n16228) );
  AND2_X1 U8897 ( .A1(n14675), .A2(n11743), .ZN(n16399) );
  AND2_X1 U8898 ( .A1(n14675), .A2(n11755), .ZN(n14678) );
  NAND2_X1 U8899 ( .A1(n8925), .A2(n8924), .ZN(n14691) );
  NAND2_X1 U8900 ( .A1(n7377), .A2(n7536), .ZN(n7863) );
  AND2_X1 U8901 ( .A1(n7926), .A2(n7928), .ZN(n7536) );
  AND2_X1 U8902 ( .A1(n7928), .A2(n16516), .ZN(n7927) );
  INV_X1 U8903 ( .A(n14585), .ZN(n14777) );
  INV_X1 U8904 ( .A(n14645), .ZN(n14788) );
  NAND2_X1 U8905 ( .A1(n8867), .A2(n8866), .ZN(n14791) );
  NAND2_X1 U8906 ( .A1(n8731), .A2(n8730), .ZN(n12902) );
  AND2_X1 U8907 ( .A1(n10935), .A2(n8976), .ZN(n15571) );
  AND2_X1 U8908 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10934), .ZN(n8976) );
  NOR2_X1 U8909 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n8066) );
  INV_X1 U8910 ( .A(n10258), .ZN(n14802) );
  NAND2_X1 U8911 ( .A1(n8964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8963) );
  OAI21_X1 U8912 ( .B1(n8966), .B2(n8965), .A(n8964), .ZN(n14815) );
  XNOR2_X1 U8913 ( .A(n8968), .B(n8967), .ZN(n14818) );
  NAND2_X1 U8914 ( .A1(n8139), .A2(n8140), .ZN(n8940) );
  INV_X1 U8915 ( .A(n8141), .ZN(n8140) );
  NAND2_X1 U8916 ( .A1(n7369), .A2(n7384), .ZN(n8139) );
  CLKBUF_X1 U8917 ( .A(n10842), .Z(n12843) );
  INV_X1 U8918 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11864) );
  INV_X1 U8919 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n11010) );
  INV_X1 U8920 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n11002) );
  INV_X1 U8921 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10989) );
  NAND2_X1 U8922 ( .A1(n8132), .A2(n8134), .ZN(n11875) );
  NAND2_X1 U8923 ( .A1(n8132), .A2(n7399), .ZN(n12168) );
  NAND2_X1 U8924 ( .A1(n14962), .A2(n14963), .ZN(n14999) );
  INV_X1 U8925 ( .A(n14981), .ZN(n7659) );
  NAND2_X1 U8926 ( .A1(n11476), .A2(n11475), .ZN(n14982) );
  NOR2_X1 U8927 ( .A1(n7670), .A2(n15009), .ZN(n7667) );
  OAI22_X1 U8928 ( .A1(n7670), .A2(n7669), .B1(n15009), .B2(n7672), .ZN(n7668)
         );
  NOR2_X1 U8929 ( .A1(n15009), .A2(n14963), .ZN(n7669) );
  INV_X1 U8930 ( .A(n15009), .ZN(n7671) );
  AND2_X1 U8931 ( .A1(n13078), .A2(n9506), .ZN(n15013) );
  NAND2_X1 U8932 ( .A1(n8111), .A2(n8114), .ZN(n12860) );
  AOI21_X1 U8933 ( .B1(n12652), .B2(n8116), .A(n8115), .ZN(n8114) );
  INV_X1 U8934 ( .A(n12720), .ZN(n8115) );
  NAND2_X1 U8935 ( .A1(n7685), .A2(n7686), .ZN(n15053) );
  NAND2_X1 U8936 ( .A1(n14934), .A2(n7688), .ZN(n7685) );
  NAND2_X1 U8937 ( .A1(n14934), .A2(n14972), .ZN(n15054) );
  NAND2_X1 U8938 ( .A1(n15065), .A2(n14904), .ZN(n15062) );
  NAND2_X1 U8939 ( .A1(n14991), .A2(n14992), .ZN(n15065) );
  NAND2_X1 U8940 ( .A1(n12862), .A2(n12861), .ZN(n14836) );
  NAND2_X1 U8941 ( .A1(n12651), .A2(n12652), .ZN(n12721) );
  NAND2_X1 U8942 ( .A1(n8118), .A2(n12650), .ZN(n12651) );
  NAND2_X1 U8943 ( .A1(n12649), .A2(n12648), .ZN(n8118) );
  XNOR2_X1 U8944 ( .A(n11474), .B(n11472), .ZN(n11470) );
  NAND2_X1 U8945 ( .A1(n11167), .A2(n11166), .ZN(n11471) );
  NAND2_X1 U8946 ( .A1(n8133), .A2(n11709), .ZN(n11869) );
  OR2_X1 U8947 ( .A1(n11711), .A2(n11710), .ZN(n8133) );
  INV_X1 U8948 ( .A(n16555), .ZN(n15104) );
  INV_X1 U8949 ( .A(n14833), .ZN(n15122) );
  INV_X1 U8950 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n11134) );
  AND4_X1 U8951 ( .A1(n9189), .A2(n9188), .A3(n9187), .A4(n9186), .ZN(n12365)
         );
  INV_X1 U8952 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n11016) );
  NAND4_X2 U8953 ( .A1(n9097), .A2(n9096), .A3(n9095), .A4(n9094), .ZN(n15141)
         );
  OR2_X1 U8954 ( .A1(n11496), .A2(n10841), .ZN(n15142) );
  OR2_X1 U8955 ( .A1(n11446), .A2(n11447), .ZN(n11444) );
  XNOR2_X1 U8956 ( .A(n7541), .B(n15705), .ZN(n15701) );
  INV_X1 U8957 ( .A(n12306), .ZN(n7541) );
  NAND2_X1 U8958 ( .A1(n15701), .A2(n16538), .ZN(n15700) );
  INV_X1 U8959 ( .A(n9583), .ZN(n15415) );
  INV_X1 U8960 ( .A(n15241), .ZN(n15418) );
  XNOR2_X1 U8961 ( .A(n8259), .B(n13074), .ZN(n15419) );
  OAI21_X1 U8962 ( .B1(n15248), .B2(n8256), .A(n8255), .ZN(n8259) );
  AOI21_X1 U8963 ( .B1(n8257), .B2(n7720), .A(n7438), .ZN(n8255) );
  INV_X1 U8964 ( .A(n8257), .ZN(n8256) );
  INV_X1 U8965 ( .A(n13074), .ZN(n13063) );
  NAND2_X1 U8966 ( .A1(n8288), .A2(n8286), .ZN(n13064) );
  INV_X1 U8967 ( .A(n8287), .ZN(n8286) );
  AOI21_X1 U8968 ( .B1(n13088), .B2(n9512), .A(n9493), .ZN(n15422) );
  AND2_X1 U8969 ( .A1(n7396), .A2(n13349), .ZN(n15429) );
  NAND2_X1 U8970 ( .A1(n15260), .A2(n8290), .ZN(n13347) );
  NAND2_X1 U8971 ( .A1(n15277), .A2(n13072), .ZN(n15267) );
  NAND2_X1 U8972 ( .A1(n14814), .A2(n9512), .ZN(n9444) );
  INV_X1 U8973 ( .A(n14928), .ZN(n15464) );
  NAND2_X1 U8974 ( .A1(n7706), .A2(n7707), .ZN(n15306) );
  NAND2_X1 U8975 ( .A1(n15332), .A2(n7397), .ZN(n7794) );
  NAND2_X1 U8976 ( .A1(n15329), .A2(n13071), .ZN(n15317) );
  INV_X1 U8977 ( .A(n15359), .ZN(n13050) );
  NAND2_X1 U8978 ( .A1(n9361), .A2(n9360), .ZN(n15370) );
  INV_X1 U8979 ( .A(n15500), .ZN(n15391) );
  NAND2_X1 U8980 ( .A1(n7782), .A2(n7785), .ZN(n15382) );
  NAND2_X1 U8981 ( .A1(n15395), .A2(n7787), .ZN(n7782) );
  NOR2_X1 U8982 ( .A1(n12959), .A2(n7693), .ZN(n7692) );
  INV_X1 U8983 ( .A(n12958), .ZN(n7693) );
  NAND2_X1 U8984 ( .A1(n15398), .A2(n12958), .ZN(n12960) );
  NAND2_X1 U8985 ( .A1(n7790), .A2(n7789), .ZN(n13045) );
  AND2_X1 U8986 ( .A1(n7790), .A2(n7412), .ZN(n12953) );
  NAND2_X1 U8987 ( .A1(n15395), .A2(n15397), .ZN(n7790) );
  NAND2_X1 U8988 ( .A1(n9309), .A2(n9308), .ZN(n16550) );
  NOR2_X1 U8989 ( .A1(n12582), .A2(n8283), .ZN(n8284) );
  INV_X1 U8990 ( .A(n12581), .ZN(n8283) );
  NAND2_X1 U8991 ( .A1(n8285), .A2(n12581), .ZN(n12583) );
  OR2_X1 U8992 ( .A1(n16153), .A2(n16532), .ZN(n15345) );
  NAND2_X1 U8993 ( .A1(n12564), .A2(n12563), .ZN(n12688) );
  AND2_X1 U8994 ( .A1(n12457), .A2(n12456), .ZN(n12458) );
  NAND2_X1 U8995 ( .A1(n12345), .A2(n12344), .ZN(n12348) );
  NAND2_X1 U8996 ( .A1(n8277), .A2(n8279), .ZN(n11968) );
  NAND2_X1 U8997 ( .A1(n11822), .A2(n8280), .ZN(n8277) );
  NAND2_X1 U8998 ( .A1(n8254), .A2(n11586), .ZN(n11827) );
  AOI21_X1 U8999 ( .B1(n7365), .B2(n15172), .A(n7695), .ZN(n7694) );
  NOR2_X1 U9000 ( .A1(n9513), .A2(n7696), .ZN(n7695) );
  INV_X1 U9001 ( .A(n15345), .ZN(n15374) );
  INV_X1 U9002 ( .A(n16156), .ZN(n16313) );
  OR2_X1 U9003 ( .A1(n16153), .A2(n16093), .ZN(n13351) );
  XNOR2_X1 U9004 ( .A(n8905), .B(n8904), .ZN(n14804) );
  NAND2_X1 U9005 ( .A1(n9025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9027) );
  INV_X1 U9006 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13087) );
  NAND2_X1 U9007 ( .A1(n7755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8273) );
  AND2_X1 U9008 ( .A1(n7758), .A2(n9004), .ZN(n7757) );
  NAND2_X1 U9009 ( .A1(n8103), .A2(n8646), .ZN(n8685) );
  XNOR2_X1 U9010 ( .A(n9406), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15560) );
  INV_X1 U9011 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12876) );
  XNOR2_X1 U9012 ( .A(n9037), .B(n9036), .ZN(n12875) );
  INV_X1 U9013 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n11132) );
  INV_X1 U9014 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n11013) );
  INV_X1 U9015 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U9016 ( .A1(n8070), .A2(n8071), .ZN(n8778) );
  XNOR2_X1 U9017 ( .A(n15736), .B(n7533), .ZN(n15897) );
  INV_X1 U9018 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7533) );
  INV_X1 U9019 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8034) );
  NAND2_X1 U9020 ( .A1(n15770), .A2(n15771), .ZN(n15894) );
  NAND2_X1 U9021 ( .A1(n15894), .A2(n15893), .ZN(n15892) );
  AND2_X1 U9022 ( .A1(n15788), .A2(n15789), .ZN(n15791) );
  NAND2_X1 U9023 ( .A1(n15810), .A2(n8016), .ZN(n15816) );
  AND2_X1 U9024 ( .A1(n7967), .A2(n7966), .ZN(n15842) );
  INV_X1 U9025 ( .A(n7964), .ZN(n15851) );
  OAI21_X1 U9026 ( .B1(n15869), .B2(n15868), .A(n15867), .ZN(n15875) );
  XNOR2_X1 U9027 ( .A(n15880), .B(n8031), .ZN(n15878) );
  INV_X1 U9028 ( .A(n15879), .ZN(n8031) );
  OAI21_X1 U9029 ( .B1(n14247), .B2(n13447), .A(n10230), .ZN(n10231) );
  AOI21_X1 U9030 ( .B1(n7879), .B2(n13333), .A(n7877), .ZN(n13342) );
  NAND2_X1 U9031 ( .A1(n16054), .A2(n7913), .ZN(n7911) );
  AOI21_X1 U9032 ( .B1(n7731), .B2(n16079), .A(n7729), .ZN(n8330) );
  NAND2_X1 U9033 ( .A1(n8239), .A2(n7423), .ZN(P3_U3486) );
  NAND2_X1 U9034 ( .A1(n14248), .A2(n16473), .ZN(n8239) );
  NOR2_X1 U9035 ( .A1(n16473), .A2(n8238), .ZN(n8237) );
  NOR2_X1 U9036 ( .A1(n10115), .A2(n10114), .ZN(n10116) );
  OAI21_X1 U9037 ( .B1(n14253), .B2(n16562), .A(n7563), .ZN(P3_U3453) );
  INV_X1 U9038 ( .A(n7564), .ZN(n7563) );
  OAI21_X1 U9039 ( .B1(n14257), .B2(n14303), .A(n7494), .ZN(n7564) );
  NAND2_X1 U9040 ( .A1(n7625), .A2(n8049), .ZN(n12384) );
  NAND2_X1 U9041 ( .A1(n7618), .A2(n12032), .ZN(n12039) );
  NAND2_X1 U9042 ( .A1(n12030), .A2(n10887), .ZN(n7618) );
  NAND2_X1 U9043 ( .A1(n7740), .A2(n7739), .ZN(P2_U3530) );
  AOI21_X1 U9044 ( .B1(n14687), .B2(n14757), .A(n7508), .ZN(n7739) );
  NAND2_X1 U9045 ( .A1(n14685), .A2(n16512), .ZN(n7740) );
  OAI21_X1 U9046 ( .B1(n8991), .B2(n14787), .A(n8990), .ZN(n8992) );
  NAND2_X1 U9047 ( .A1(n8161), .A2(n8160), .ZN(n16520) );
  INV_X1 U9048 ( .A(n8305), .ZN(n8304) );
  AND2_X1 U9049 ( .A1(n9595), .A2(n9612), .ZN(n8306) );
  NAND2_X1 U9050 ( .A1(n7652), .A2(n7503), .ZN(P1_U3557) );
  NAND2_X1 U9051 ( .A1(n8247), .A2(n16539), .ZN(n7652) );
  INV_X1 U9052 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U9053 ( .A1(n7698), .A2(n7504), .ZN(P1_U3556) );
  NAND2_X1 U9054 ( .A1(n15527), .A2(n16539), .ZN(n7698) );
  INV_X1 U9055 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U9056 ( .A1(n7767), .A2(n7505), .ZN(P1_U3525) );
  NAND2_X1 U9057 ( .A1(n8247), .A2(n16543), .ZN(n7767) );
  INV_X1 U9058 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U9059 ( .A1(n9009), .A2(n9008), .ZN(n15543) );
  OAI21_X1 U9060 ( .B1(n13122), .B2(n15556), .A(n7512), .ZN(P1_U3325) );
  OR2_X1 U9061 ( .A1(n15558), .A2(n13268), .ZN(n8275) );
  INV_X2 U9062 ( .A(n10351), .ZN(n10507) );
  INV_X1 U9063 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15542) );
  AND2_X1 U9064 ( .A1(n7727), .A2(n13072), .ZN(n7371) );
  NAND2_X1 U9065 ( .A1(n8683), .A2(n8682), .ZN(n10455) );
  NAND2_X1 U9066 ( .A1(n7658), .A2(SI_4_), .ZN(n8597) );
  XNOR2_X1 U9067 ( .A(n14700), .B(n14440), .ZN(n14513) );
  AND3_X1 U9068 ( .A1(n9003), .A2(n9291), .A3(n9002), .ZN(n7372) );
  AND2_X1 U9069 ( .A1(n9049), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7373) );
  INV_X1 U9070 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9010) );
  XNOR2_X1 U9071 ( .A(n14585), .B(n14455), .ZN(n14583) );
  INV_X1 U9072 ( .A(n14583), .ZN(n7949) );
  INV_X1 U9073 ( .A(n8834), .ZN(n8096) );
  AND2_X1 U9074 ( .A1(n13389), .A2(n8188), .ZN(n7374) );
  AND2_X1 U9075 ( .A1(n12795), .A2(n14459), .ZN(n7375) );
  AND2_X1 U9076 ( .A1(n14768), .A2(n14559), .ZN(n7376) );
  AND2_X1 U9077 ( .A1(n7929), .A2(n16512), .ZN(n7377) );
  AND2_X1 U9078 ( .A1(n14732), .A2(n14456), .ZN(n7378) );
  AND2_X1 U9079 ( .A1(n8335), .A2(n8942), .ZN(n7379) );
  INV_X1 U9080 ( .A(n7392), .ZN(n7720) );
  INV_X1 U9081 ( .A(n10302), .ZN(n10351) );
  AND2_X1 U9082 ( .A1(n13072), .A2(n9545), .ZN(n7380) );
  INV_X1 U9083 ( .A(n14677), .ZN(n7748) );
  AND2_X1 U9084 ( .A1(n10710), .A2(n10709), .ZN(n7381) );
  AND2_X1 U9085 ( .A1(n7455), .A2(n10315), .ZN(n7382) );
  AND2_X1 U9086 ( .A1(n11034), .A2(n11496), .ZN(n11037) );
  OR2_X1 U9087 ( .A1(n10656), .A2(n10655), .ZN(n7383) );
  AND2_X1 U9088 ( .A1(n7379), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n7384) );
  OAI21_X1 U9089 ( .B1(n8635), .B2(n8080), .A(n7648), .ZN(n7647) );
  OR2_X1 U9090 ( .A1(n10739), .A2(n10738), .ZN(n7385) );
  INV_X1 U9091 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8672) );
  AND2_X1 U9092 ( .A1(n7896), .A2(n10081), .ZN(n7386) );
  INV_X1 U9093 ( .A(n9565), .ZN(n8086) );
  XNOR2_X1 U9094 ( .A(n15457), .B(n14833), .ZN(n13055) );
  AND2_X1 U9095 ( .A1(n7794), .A2(n7796), .ZN(n7387) );
  OAI21_X1 U9096 ( .B1(n13325), .B2(n13955), .A(n13296), .ZN(n13287) );
  AND2_X1 U9097 ( .A1(n8196), .A2(n8188), .ZN(n7388) );
  AND2_X1 U9098 ( .A1(n15376), .A2(n13066), .ZN(n7389) );
  NOR2_X1 U9099 ( .A1(n12543), .A2(n12542), .ZN(n7390) );
  OR2_X1 U9100 ( .A1(n8104), .A2(n8648), .ZN(n7391) );
  INV_X2 U9101 ( .A(n13207), .ZN(n13266) );
  INV_X1 U9102 ( .A(n11932), .ZN(n10118) );
  INV_X1 U9103 ( .A(n15952), .ZN(n7735) );
  INV_X1 U9104 ( .A(n15305), .ZN(n7705) );
  OR2_X1 U9105 ( .A1(n15257), .A2(n8086), .ZN(n7392) );
  AND2_X1 U9106 ( .A1(n9641), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7393) );
  AND2_X1 U9107 ( .A1(n7964), .A2(n7963), .ZN(n7394) );
  NAND2_X1 U9108 ( .A1(n7650), .A2(n8635), .ZN(n8697) );
  INV_X1 U9109 ( .A(n8078), .ZN(n8688) );
  AND2_X1 U9110 ( .A1(n15062), .A2(n14917), .ZN(n7395) );
  INV_X1 U9111 ( .A(n12339), .ZN(n12268) );
  OR3_X1 U9112 ( .A1(n15284), .A2(n7775), .A3(n15436), .ZN(n7396) );
  XNOR2_X1 U9113 ( .A(n15428), .B(n15119), .ZN(n13344) );
  INV_X1 U9114 ( .A(n13344), .ZN(n8258) );
  INV_X1 U9115 ( .A(n10296), .ZN(n10407) );
  INV_X1 U9116 ( .A(n9050), .ZN(n9335) );
  AND2_X1 U9117 ( .A1(n13054), .A2(n13053), .ZN(n7397) );
  AND2_X1 U9118 ( .A1(n8148), .A2(n15074), .ZN(n7398) );
  AND2_X1 U9119 ( .A1(n8134), .A2(n8131), .ZN(n7399) );
  INV_X1 U9120 ( .A(n9098), .ZN(n7710) );
  NAND2_X1 U9121 ( .A1(n15470), .A2(n14919), .ZN(n7400) );
  INV_X1 U9122 ( .A(n16142), .ZN(n9047) );
  NAND2_X1 U9123 ( .A1(n14017), .A2(n10083), .ZN(n13991) );
  OR2_X1 U9124 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n9668), .ZN(n7401) );
  INV_X1 U9125 ( .A(n13073), .ZN(n7726) );
  AND2_X1 U9126 ( .A1(n14368), .A2(n14436), .ZN(n7402) );
  OR2_X1 U9127 ( .A1(n8841), .A2(n8095), .ZN(n7403) );
  AND2_X1 U9128 ( .A1(n7369), .A2(n7379), .ZN(n7404) );
  XNOR2_X1 U9129 ( .A(n15436), .B(n8086), .ZN(n15262) );
  INV_X1 U9130 ( .A(n15262), .ZN(n15247) );
  NAND2_X1 U9131 ( .A1(n14053), .A2(n13237), .ZN(n14036) );
  NAND4_X1 U9132 ( .A1(n9689), .A2(n9688), .A3(n9687), .A4(n9686), .ZN(n13893)
         );
  AND2_X1 U9133 ( .A1(n13304), .A2(n9767), .ZN(n7405) );
  NOR2_X1 U9134 ( .A1(n7795), .A2(n7705), .ZN(n7793) );
  AND2_X1 U9135 ( .A1(n7952), .A2(n14609), .ZN(n7406) );
  OR2_X1 U9136 ( .A1(n8619), .A2(SI_12_), .ZN(n7407) );
  NAND2_X1 U9137 ( .A1(n8696), .A2(n8695), .ZN(n14739) );
  NAND2_X1 U9138 ( .A1(n8885), .A2(n8884), .ZN(n14705) );
  INV_X1 U9139 ( .A(n14963), .ZN(n7673) );
  AND2_X1 U9140 ( .A1(n7852), .A2(n7855), .ZN(n7408) );
  XNOR2_X1 U9141 ( .A(n13064), .B(n13063), .ZN(n15426) );
  AND2_X1 U9142 ( .A1(n7929), .A2(n7931), .ZN(n13094) );
  NAND2_X1 U9143 ( .A1(n8873), .A2(n8872), .ZN(n14573) );
  INV_X1 U9144 ( .A(n14573), .ZN(n7752) );
  NAND2_X1 U9145 ( .A1(n8840), .A2(n8839), .ZN(n12037) );
  NAND2_X1 U9146 ( .A1(n10172), .A2(n14147), .ZN(n7409) );
  AND2_X1 U9147 ( .A1(n7752), .A2(n7753), .ZN(n7410) );
  NOR2_X1 U9148 ( .A1(n13449), .A2(n8199), .ZN(n7411) );
  INV_X1 U9149 ( .A(n9241), .ZN(n8317) );
  OR2_X1 U9150 ( .A1(n16550), .A2(n15130), .ZN(n7412) );
  INV_X1 U9151 ( .A(n9436), .ZN(n8320) );
  NAND2_X1 U9152 ( .A1(n9245), .A2(n9244), .ZN(n16493) );
  NAND2_X1 U9153 ( .A1(n14666), .A2(n10678), .ZN(n7413) );
  XNOR2_X1 U9154 ( .A(n14705), .B(n14453), .ZN(n14529) );
  NAND2_X1 U9155 ( .A1(n9434), .A2(n9433), .ZN(n15457) );
  AND2_X1 U9156 ( .A1(n8338), .A2(n7577), .ZN(n7414) );
  AND3_X1 U9157 ( .A1(n12280), .A2(n10069), .A3(n12282), .ZN(n7415) );
  AND2_X1 U9158 ( .A1(n7619), .A2(n7616), .ZN(n7416) );
  NAND2_X1 U9159 ( .A1(n14399), .A2(n10918), .ZN(n7417) );
  AND2_X1 U9160 ( .A1(n10676), .A2(n10675), .ZN(n7418) );
  AND2_X1 U9161 ( .A1(n10698), .A2(n10697), .ZN(n7419) );
  NAND2_X1 U9162 ( .A1(n9299), .A2(n9298), .ZN(n16529) );
  AND3_X1 U9163 ( .A1(n7990), .A2(n7989), .A3(n7985), .ZN(n7420) );
  AND2_X1 U9164 ( .A1(n8079), .A2(n8706), .ZN(n7421) );
  NOR2_X1 U9165 ( .A1(n10070), .A2(n7560), .ZN(n7422) );
  NOR2_X1 U9166 ( .A1(n13118), .A2(n8237), .ZN(n7423) );
  AND2_X1 U9167 ( .A1(n14229), .A2(n13027), .ZN(n7424) );
  NAND2_X1 U9168 ( .A1(n8748), .A2(n8747), .ZN(n12504) );
  AND2_X1 U9169 ( .A1(n15427), .A2(n15425), .ZN(n7425) );
  AND2_X1 U9170 ( .A1(n13056), .A2(n13055), .ZN(n7426) );
  AND2_X1 U9171 ( .A1(n8680), .A2(n8679), .ZN(n14768) );
  INV_X1 U9172 ( .A(n14768), .ZN(n7754) );
  INV_X1 U9173 ( .A(n10540), .ZN(n7860) );
  XOR2_X1 U9174 ( .A(n8577), .B(n8576), .Z(n7427) );
  INV_X1 U9175 ( .A(n9464), .ZN(n8314) );
  INV_X1 U9176 ( .A(n15428), .ZN(n15006) );
  NAND2_X1 U9177 ( .A1(n9515), .A2(n9514), .ZN(n15428) );
  AND2_X1 U9178 ( .A1(n9050), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7428) );
  INV_X1 U9179 ( .A(n7869), .ZN(n7868) );
  NAND2_X1 U9180 ( .A1(n7870), .A2(n10533), .ZN(n7869) );
  INV_X1 U9181 ( .A(n9301), .ZN(n8324) );
  AND2_X1 U9182 ( .A1(n7707), .A2(n7705), .ZN(n7429) );
  NAND2_X1 U9183 ( .A1(n10202), .A2(n13999), .ZN(n7430) );
  NAND2_X1 U9184 ( .A1(n11019), .A2(n8433), .ZN(n7431) );
  NAND2_X1 U9185 ( .A1(n12602), .A2(n10071), .ZN(n7432) );
  AND2_X1 U9186 ( .A1(n10538), .A2(n10537), .ZN(n7433) );
  NOR2_X1 U9187 ( .A1(n12101), .A2(n14469), .ZN(n7434) );
  NOR2_X1 U9188 ( .A1(n13917), .A2(n8440), .ZN(n7435) );
  AND2_X1 U9189 ( .A1(n7631), .A2(n8091), .ZN(n7436) );
  AND2_X1 U9190 ( .A1(n10625), .A2(n10624), .ZN(n7437) );
  AND2_X1 U9191 ( .A1(n15428), .A2(n15004), .ZN(n7438) );
  AND2_X1 U9192 ( .A1(n7380), .A2(n8265), .ZN(n7439) );
  AND2_X1 U9193 ( .A1(n8243), .A2(n7907), .ZN(n7440) );
  AND2_X1 U9194 ( .A1(n15329), .A2(n8262), .ZN(n7441) );
  OR2_X1 U9195 ( .A1(n14585), .A2(n14597), .ZN(n7442) );
  NOR2_X1 U9196 ( .A1(n14436), .A2(n14338), .ZN(n7443) );
  INV_X1 U9197 ( .A(n7788), .ZN(n7787) );
  NAND2_X1 U9198 ( .A1(n15397), .A2(n13044), .ZN(n7788) );
  NOR2_X1 U9199 ( .A1(n8193), .A2(n7388), .ZN(n7444) );
  NAND2_X1 U9200 ( .A1(n10495), .A2(n10494), .ZN(n14499) );
  INV_X1 U9201 ( .A(n14499), .ZN(n7874) );
  INV_X1 U9202 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9008) );
  AND2_X1 U9203 ( .A1(n16323), .A2(n14469), .ZN(n7445) );
  INV_X1 U9204 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8142) );
  AND2_X1 U9205 ( .A1(n14493), .A2(n14369), .ZN(n7446) );
  AND4_X1 U9206 ( .A1(n7522), .A2(n8355), .A3(n8357), .A4(n8358), .ZN(n7447)
         );
  INV_X1 U9207 ( .A(n9691), .ZN(n8227) );
  NAND2_X1 U9208 ( .A1(n8588), .A2(n7845), .ZN(n8815) );
  NAND2_X1 U9209 ( .A1(n15333), .A2(n13052), .ZN(n7449) );
  INV_X1 U9210 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7689) );
  AND2_X1 U9211 ( .A1(n12379), .A2(n10900), .ZN(n7450) );
  AND2_X1 U9212 ( .A1(n10890), .A2(n10889), .ZN(n7451) );
  AND2_X1 U9213 ( .A1(n10903), .A2(n10902), .ZN(n7452) );
  INV_X1 U9214 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9026) );
  INV_X1 U9215 ( .A(n7898), .ZN(n7897) );
  NAND2_X1 U9216 ( .A1(n7899), .A2(n10080), .ZN(n7898) );
  AND2_X1 U9217 ( .A1(n9632), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7453) );
  NOR2_X1 U9218 ( .A1(n14928), .A2(n15123), .ZN(n7454) );
  INV_X1 U9219 ( .A(n9030), .ZN(n9031) );
  NAND2_X1 U9220 ( .A1(n7372), .A2(n9004), .ZN(n9030) );
  NAND2_X1 U9221 ( .A1(n9038), .A2(n9035), .ZN(n12770) );
  INV_X1 U9222 ( .A(n12770), .ZN(n7690) );
  NAND2_X1 U9223 ( .A1(n12101), .A2(n10324), .ZN(n7455) );
  AND2_X1 U9224 ( .A1(n7400), .A2(n15330), .ZN(n7456) );
  INV_X1 U9225 ( .A(n8281), .ZN(n8280) );
  NOR2_X1 U9226 ( .A1(n11824), .A2(n11823), .ZN(n8281) );
  AND2_X1 U9227 ( .A1(n9697), .A2(n9708), .ZN(n7457) );
  NAND2_X1 U9228 ( .A1(n8597), .A2(n7655), .ZN(n8787) );
  NAND2_X1 U9229 ( .A1(n10443), .A2(n10434), .ZN(n7458) );
  OR2_X1 U9230 ( .A1(n15824), .A2(n15823), .ZN(n7459) );
  NAND2_X1 U9231 ( .A1(n10456), .A2(n10457), .ZN(n14557) );
  AND2_X1 U9232 ( .A1(n15332), .A2(n13053), .ZN(n7460) );
  OR2_X1 U9233 ( .A1(n7721), .A2(n8258), .ZN(n7461) );
  OR2_X1 U9234 ( .A1(n15464), .A2(n15123), .ZN(n7462) );
  OR2_X1 U9235 ( .A1(n10661), .A2(n10663), .ZN(n7463) );
  OR2_X1 U9236 ( .A1(n10679), .A2(n7418), .ZN(n7464) );
  AND2_X1 U9237 ( .A1(n8618), .A2(n7407), .ZN(n7465) );
  AND2_X1 U9238 ( .A1(n7770), .A2(n7769), .ZN(n7466) );
  AND2_X1 U9239 ( .A1(n8999), .A2(n7689), .ZN(n7467) );
  AND2_X1 U9240 ( .A1(n10960), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9241 ( .A1(n16388), .A2(n12365), .ZN(n7469) );
  INV_X1 U9242 ( .A(n10167), .ZN(n8210) );
  AND2_X1 U9243 ( .A1(n7710), .A2(n9004), .ZN(n7470) );
  AND2_X1 U9244 ( .A1(n9743), .A2(n9728), .ZN(n7471) );
  OR2_X1 U9245 ( .A1(n8324), .A2(n9300), .ZN(n7472) );
  OR2_X1 U9246 ( .A1(n8314), .A2(n9463), .ZN(n7473) );
  OR2_X1 U9247 ( .A1(n9331), .A2(n9329), .ZN(n7474) );
  OR2_X1 U9248 ( .A1(n9364), .A2(n9362), .ZN(n7475) );
  OR2_X1 U9249 ( .A1(n8317), .A2(n9240), .ZN(n7476) );
  AND2_X1 U9250 ( .A1(n7949), .A2(n7853), .ZN(n7477) );
  OR2_X1 U9251 ( .A1(n8163), .A2(n10662), .ZN(n7478) );
  AND2_X1 U9252 ( .A1(n7783), .A2(n15383), .ZN(n7479) );
  AND2_X1 U9253 ( .A1(n10524), .A2(n10523), .ZN(n7480) );
  OR2_X1 U9254 ( .A1(n8320), .A2(n9435), .ZN(n7481) );
  AND2_X1 U9255 ( .A1(n10133), .A2(n10132), .ZN(n7482) );
  INV_X1 U9256 ( .A(n8050), .ZN(n8049) );
  NAND2_X1 U9257 ( .A1(n8051), .A2(n12378), .ZN(n8050) );
  INV_X1 U9258 ( .A(n8290), .ZN(n8289) );
  AND2_X1 U9259 ( .A1(n13061), .A2(n8258), .ZN(n8290) );
  AND2_X1 U9260 ( .A1(n13439), .A2(n7409), .ZN(n8205) );
  OR2_X1 U9261 ( .A1(n10742), .A2(n8147), .ZN(n7483) );
  INV_X1 U9262 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8460) );
  OR2_X1 U9263 ( .A1(n10112), .A2(n13974), .ZN(n13295) );
  INV_X1 U9264 ( .A(n7906), .ZN(n7905) );
  NAND2_X1 U9265 ( .A1(n13111), .A2(n13246), .ZN(n7906) );
  OR2_X1 U9266 ( .A1(n7673), .A2(n7671), .ZN(n7484) );
  OR2_X1 U9267 ( .A1(n14252), .A2(n14251), .ZN(P3_U3454) );
  OR2_X1 U9268 ( .A1(n13990), .A2(n13989), .ZN(P3_U3206) );
  INV_X2 U9269 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U9270 ( .A(SI_4_), .ZN(n7656) );
  INV_X1 U9271 ( .A(n15992), .ZN(n7737) );
  INV_X1 U9272 ( .A(n11784), .ZN(n7889) );
  INV_X1 U9273 ( .A(n14038), .ZN(n8013) );
  INV_X1 U9274 ( .A(SI_1_), .ZN(n7839) );
  INV_X1 U9275 ( .A(n10195), .ZN(n8188) );
  NAND2_X1 U9276 ( .A1(n8691), .A2(n8690), .ZN(n14732) );
  INV_X1 U9277 ( .A(n14732), .ZN(n7743) );
  NAND2_X1 U9278 ( .A1(n8285), .A2(n8284), .ZN(n12714) );
  AND2_X1 U9279 ( .A1(n12676), .A2(n7772), .ZN(n7487) );
  XNOR2_X1 U9280 ( .A(n8886), .B(n8883), .ZN(n14811) );
  NAND2_X1 U9281 ( .A1(n13403), .A2(n13397), .ZN(n7488) );
  INV_X1 U9282 ( .A(n14069), .ZN(n7899) );
  NAND2_X1 U9283 ( .A1(n8700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8709) );
  INV_X1 U9284 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n7881) );
  INV_X1 U9285 ( .A(n15073), .ZN(n8150) );
  INV_X1 U9286 ( .A(n15051), .ZN(n7687) );
  AND2_X1 U9287 ( .A1(n12914), .A2(n8062), .ZN(n7489) );
  AND2_X1 U9288 ( .A1(n8911), .A2(n8910), .ZN(n10761) );
  INV_X1 U9289 ( .A(n10761), .ZN(n13098) );
  INV_X1 U9290 ( .A(n7857), .ZN(n7856) );
  NOR2_X1 U9291 ( .A1(n10541), .A2(n7858), .ZN(n7857) );
  AND2_X1 U9292 ( .A1(n10534), .A2(n10533), .ZN(n7490) );
  INV_X1 U9293 ( .A(n10512), .ZN(n7931) );
  NAND2_X1 U9294 ( .A1(n8269), .A2(n15376), .ZN(n7491) );
  INV_X1 U9295 ( .A(n7796), .ZN(n7795) );
  NAND2_X1 U9296 ( .A1(n15470), .A2(n15124), .ZN(n7796) );
  INV_X1 U9297 ( .A(n10196), .ZN(n8201) );
  INV_X1 U9298 ( .A(n8080), .ZN(n8079) );
  OAI21_X1 U9299 ( .B1(n8081), .B2(n8084), .A(n8641), .ZN(n8080) );
  AND2_X1 U9300 ( .A1(n10174), .A2(n14132), .ZN(n7492) );
  OR2_X1 U9301 ( .A1(n14247), .A2(n14227), .ZN(n7493) );
  INV_X1 U9302 ( .A(SI_9_), .ZN(n13506) );
  AND2_X1 U9303 ( .A1(n14256), .A2(n7565), .ZN(n7494) );
  INV_X1 U9304 ( .A(n10198), .ZN(n8200) );
  AND2_X1 U9305 ( .A1(n10197), .A2(n14027), .ZN(n10198) );
  OR2_X1 U9306 ( .A1(n14247), .A2(n14296), .ZN(n7495) );
  NOR2_X1 U9307 ( .A1(n8185), .A2(n7882), .ZN(n7496) );
  AND2_X1 U9308 ( .A1(n9646), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7497) );
  INV_X1 U9309 ( .A(n8868), .ZN(n8104) );
  OR2_X1 U9310 ( .A1(n14238), .A2(n13026), .ZN(n13201) );
  INV_X1 U9311 ( .A(n13201), .ZN(n7892) );
  AND2_X1 U9312 ( .A1(n12955), .A2(n12954), .ZN(n7498) );
  AND2_X1 U9313 ( .A1(n14376), .A2(n14377), .ZN(n7499) );
  INV_X1 U9314 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n7886) );
  AND2_X1 U9315 ( .A1(n14141), .A2(n9879), .ZN(n7500) );
  INV_X1 U9316 ( .A(n15000), .ZN(n11038) );
  INV_X1 U9317 ( .A(n16447), .ZN(n16562) );
  INV_X1 U9318 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n13555) );
  INV_X1 U9319 ( .A(n12627), .ZN(n7870) );
  OR2_X1 U9320 ( .A1(n8024), .A2(n8022), .ZN(n7501) );
  INV_X1 U9321 ( .A(n11019), .ZN(n7734) );
  NAND2_X1 U9322 ( .A1(n8647), .A2(SI_23_), .ZN(n7502) );
  OR2_X1 U9323 ( .A1(n16539), .A2(n7651), .ZN(n7503) );
  OR2_X1 U9324 ( .A1(n16539), .A2(n7697), .ZN(n7504) );
  OR2_X1 U9325 ( .A1(n16543), .A2(n7766), .ZN(n7505) );
  INV_X1 U9326 ( .A(n16388), .ZN(n7765) );
  NAND2_X1 U9327 ( .A1(n11963), .A2(n11962), .ZN(n12267) );
  OR2_X1 U9328 ( .A1(n13742), .A2(n13741), .ZN(n7506) );
  AND2_X1 U9329 ( .A1(n12941), .A2(n10413), .ZN(n12742) );
  INV_X1 U9330 ( .A(n12742), .ZN(n7934) );
  AND2_X1 U9331 ( .A1(n13279), .A2(SI_31_), .ZN(n7507) );
  AND2_X1 U9332 ( .A1(n14686), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7508) );
  AND2_X1 U9333 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n9656), .ZN(n7509) );
  INV_X1 U9334 ( .A(n8029), .ZN(n8027) );
  NAND2_X1 U9335 ( .A1(n12876), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8029) );
  INV_X1 U9336 ( .A(n15222), .ZN(n7542) );
  AND2_X1 U9337 ( .A1(n16298), .A2(n16264), .ZN(n7510) );
  INV_X1 U9338 ( .A(n9944), .ZN(n8026) );
  AND2_X1 U9339 ( .A1(n11774), .A2(n13330), .ZN(n13289) );
  OR2_X1 U9340 ( .A1(n7915), .A2(n8447), .ZN(n7511) );
  INV_X1 U9341 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8038) );
  INV_X1 U9342 ( .A(n11452), .ZN(n13330) );
  INV_X1 U9343 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n8036) );
  AND2_X1 U9344 ( .A1(n8275), .A2(n8274), .ZN(n7512) );
  INV_X1 U9345 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15886) );
  INV_X1 U9346 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7529) );
  INV_X1 U9347 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7696) );
  INV_X1 U9348 ( .A(n13234), .ZN(n7876) );
  AND2_X1 U9349 ( .A1(n11496), .A2(n10996), .ZN(n11555) );
  NAND2_X1 U9350 ( .A1(n8064), .A2(n10916), .ZN(n8063) );
  INV_X1 U9351 ( .A(n8615), .ZN(n8095) );
  NAND2_X1 U9352 ( .A1(n8094), .A2(n8850), .ZN(n8092) );
  NAND2_X1 U9353 ( .A1(n8092), .A2(n7407), .ZN(n8091) );
  OAI22_X1 U9354 ( .A1(n14412), .A2(n14410), .B1(n14326), .B2(n14325), .ZN(
        n14329) );
  AOI21_X1 U9355 ( .B1(n14348), .B2(n14347), .A(n14330), .ZN(n14392) );
  OAI21_X1 U9356 ( .B1(n14378), .B2(n14408), .A(n7499), .ZN(P2_U3192) );
  NAND2_X1 U9357 ( .A1(n8771), .A2(n8602), .ZN(n8759) );
  INV_X1 U9358 ( .A(n8060), .ZN(n8059) );
  NAND2_X1 U9359 ( .A1(n8814), .A2(n8588), .ZN(n8590) );
  NAND2_X1 U9360 ( .A1(n10848), .A2(n10847), .ZN(n14428) );
  NAND2_X1 U9361 ( .A1(n14409), .A2(n8057), .ZN(n14324) );
  NAND3_X1 U9362 ( .A1(n8105), .A2(n8661), .A3(n8809), .ZN(n7515) );
  INV_X1 U9363 ( .A(n10719), .ZN(n7518) );
  NAND2_X1 U9364 ( .A1(n10695), .A2(n10694), .ZN(n7520) );
  NAND2_X1 U9365 ( .A1(n7369), .A2(n7521), .ZN(n8674) );
  NAND2_X1 U9366 ( .A1(n12342), .A2(n12341), .ZN(n12453) );
  NAND2_X1 U9367 ( .A1(n11975), .A2(n11974), .ZN(n12263) );
  NAND2_X1 U9368 ( .A1(n12325), .A2(n9755), .ZN(n12291) );
  NAND2_X1 U9369 ( .A1(n11571), .A2(n11570), .ZN(n12040) );
  NAND2_X1 U9370 ( .A1(n14181), .A2(n7493), .ZN(P3_U3487) );
  NAND2_X1 U9371 ( .A1(n14246), .A2(n7495), .ZN(P3_U3455) );
  NAND2_X1 U9372 ( .A1(n7646), .A2(n7534), .ZN(n7642) );
  NAND2_X1 U9373 ( .A1(n12134), .A2(n12133), .ZN(n8225) );
  INV_X1 U9374 ( .A(n15431), .ZN(n7540) );
  NAND2_X1 U9375 ( .A1(n7654), .A2(n13059), .ZN(n15258) );
  INV_X1 U9376 ( .A(n15486), .ZN(n7535) );
  NAND2_X1 U9377 ( .A1(n15434), .A2(n15433), .ZN(n15527) );
  OAI211_X1 U9378 ( .C1(n11822), .C2(n8278), .A(n11967), .B(n8276), .ZN(n8282)
         );
  AOI21_X1 U9379 ( .B1(n13116), .B2(n10022), .A(n13973), .ZN(n10042) );
  OAI21_X1 U9380 ( .B1(n13973), .B2(n13972), .A(n13976), .ZN(n14179) );
  NAND2_X1 U9381 ( .A1(n15750), .A2(n15749), .ZN(n8037) );
  XNOR2_X1 U9382 ( .A(n15763), .B(n8034), .ZN(n15765) );
  INV_X1 U9383 ( .A(n15834), .ZN(n7967) );
  NAND2_X1 U9384 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7526), .ZN(n7525) );
  INV_X1 U9385 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7526) );
  NAND2_X1 U9386 ( .A1(n15734), .A2(n15735), .ZN(n7527) );
  OAI21_X1 U9387 ( .B1(n15791), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8040), .ZN(
        n8039) );
  XNOR2_X1 U9388 ( .A(n15807), .B(n8017), .ZN(n15809) );
  NAND3_X1 U9389 ( .A1(n8145), .A2(n7385), .A3(n7483), .ZN(n8144) );
  INV_X1 U9390 ( .A(n10641), .ZN(n10760) );
  NOR2_X1 U9391 ( .A1(n10696), .A2(n8173), .ZN(n8171) );
  NOR2_X1 U9392 ( .A1(n10707), .A2(n8159), .ZN(n8157) );
  NAND2_X1 U9393 ( .A1(n10650), .A2(n10649), .ZN(n10656) );
  NAND2_X1 U9394 ( .A1(n8122), .A2(n8119), .ZN(n10739) );
  NAND2_X1 U9395 ( .A1(n10730), .A2(n10729), .ZN(n8120) );
  AOI21_X1 U9396 ( .B1(n10632), .B2(n10631), .A(n10630), .ZN(n10633) );
  OR2_X1 U9397 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  INV_X1 U9398 ( .A(n8063), .ZN(n8062) );
  NAND2_X1 U9399 ( .A1(n10532), .A2(n10531), .ZN(n12661) );
  NAND2_X1 U9400 ( .A1(n14568), .A2(n14569), .ZN(n10545) );
  NAND2_X1 U9401 ( .A1(n10543), .A2(n10542), .ZN(n14568) );
  NAND2_X1 U9402 ( .A1(n7863), .A2(n10558), .ZN(n10560) );
  NAND2_X1 U9403 ( .A1(n12257), .A2(n10527), .ZN(n12422) );
  NAND2_X1 U9404 ( .A1(n7993), .A2(n7992), .ZN(n7991) );
  NAND2_X1 U9405 ( .A1(n9826), .A2(n9825), .ZN(n9647) );
  NAND2_X1 U9406 ( .A1(n10028), .A2(n9673), .ZN(n10030) );
  NAND2_X1 U9407 ( .A1(n7878), .A2(n7420), .ZN(n7877) );
  NAND2_X1 U9408 ( .A1(n15835), .A2(n11933), .ZN(n7966) );
  INV_X1 U9409 ( .A(n8039), .ZN(n15799) );
  NAND2_X1 U9410 ( .A1(n15809), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U9411 ( .A1(n15875), .A2(n15876), .ZN(n8032) );
  OAI21_X1 U9412 ( .B1(n15825), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7459), .ZN(
        n8030) );
  NOR2_X1 U9413 ( .A1(n15842), .A2(n15841), .ZN(n15843) );
  NAND2_X1 U9414 ( .A1(n10520), .A2(n10519), .ZN(n12098) );
  NAND2_X1 U9415 ( .A1(n15765), .A2(n15764), .ZN(n8033) );
  INV_X1 U9416 ( .A(n15792), .ZN(n8040) );
  OAI21_X1 U9417 ( .B1(n15802), .B2(n15801), .A(n15800), .ZN(n15807) );
  NAND2_X1 U9418 ( .A1(n8282), .A2(n11970), .ZN(n12067) );
  NOR2_X2 U9419 ( .A1(n7535), .A2(n7449), .ZN(n7646) );
  NAND2_X1 U9420 ( .A1(n15266), .A2(n7726), .ZN(n7654) );
  NAND2_X1 U9421 ( .A1(n15381), .A2(n13047), .ZN(n15363) );
  NAND2_X1 U9422 ( .A1(n10760), .A2(n16106), .ZN(n10568) );
  INV_X4 U9423 ( .A(n10747), .ZN(n10767) );
  AOI21_X1 U9424 ( .B1(n10746), .B2(n10745), .A(n10744), .ZN(n10754) );
  NAND2_X1 U9425 ( .A1(n14504), .A2(n14503), .ZN(n7944) );
  NAND2_X1 U9426 ( .A1(n7932), .A2(n16107), .ZN(n7929) );
  NAND2_X1 U9427 ( .A1(n14324), .A2(n14323), .ZN(n14325) );
  NAND2_X1 U9428 ( .A1(n9380), .A2(n9379), .ZN(n9394) );
  INV_X1 U9429 ( .A(n7547), .ZN(n9594) );
  NAND2_X1 U9430 ( .A1(n9468), .A2(n9469), .ZN(n7548) );
  OAI21_X1 U9431 ( .B1(n16143), .B2(n15143), .A(n9500), .ZN(n9058) );
  INV_X1 U9432 ( .A(n7650), .ZN(n7649) );
  INV_X1 U9433 ( .A(n7635), .ZN(n7634) );
  OR2_X1 U9434 ( .A1(n14358), .A2(n10846), .ZN(n10847) );
  NAND2_X1 U9435 ( .A1(n15281), .A2(n13058), .ZN(n15266) );
  NAND2_X1 U9436 ( .A1(n15260), .A2(n13061), .ZN(n13345) );
  NAND2_X2 U9437 ( .A1(n13051), .A2(n13050), .ZN(n15486) );
  NAND2_X1 U9438 ( .A1(n7544), .A2(n8323), .ZN(n9312) );
  NAND3_X1 U9439 ( .A1(n9282), .A2(n9281), .A3(n7472), .ZN(n7544) );
  NAND2_X1 U9440 ( .A1(n7545), .A2(n8308), .ZN(n9345) );
  NAND3_X1 U9441 ( .A1(n9317), .A2(n9316), .A3(n7474), .ZN(n7545) );
  NAND2_X1 U9442 ( .A1(n7546), .A2(n8321), .ZN(n9375) );
  NAND3_X1 U9443 ( .A1(n9350), .A2(n9349), .A3(n7475), .ZN(n7546) );
  NAND2_X1 U9444 ( .A1(n7549), .A2(n7548), .ZN(n7547) );
  NAND2_X1 U9445 ( .A1(n7551), .A2(n7550), .ZN(n7549) );
  NAND2_X1 U9446 ( .A1(n9467), .A2(n9466), .ZN(n7551) );
  CLKBUF_X3 U9447 ( .A(n9107), .Z(n9500) );
  NAND2_X1 U9448 ( .A1(n8779), .A2(n8599), .ZN(n8769) );
  INV_X1 U9449 ( .A(n14428), .ZN(n8064) );
  XNOR2_X1 U9450 ( .A(n8048), .B(n14372), .ZN(n14378) );
  OAI21_X2 U9451 ( .B1(n14099), .B2(n7898), .A(n7386), .ZN(n14053) );
  XNOR2_X1 U9452 ( .A(n10123), .B(n10122), .ZN(n7554) );
  NAND2_X1 U9453 ( .A1(n7554), .A2(n11413), .ZN(n11412) );
  NAND2_X1 U9454 ( .A1(n11412), .A2(n7553), .ZN(n11414) );
  OR2_X1 U9455 ( .A1(n11413), .A2(n7554), .ZN(n7553) );
  NAND2_X1 U9456 ( .A1(n10182), .A2(n7556), .ZN(n7555) );
  NAND2_X1 U9457 ( .A1(n7559), .A2(n7558), .ZN(n12755) );
  NAND2_X1 U9458 ( .A1(n7482), .A2(n11659), .ZN(n11728) );
  NAND2_X1 U9459 ( .A1(n7569), .A2(n7570), .ZN(n10171) );
  NAND2_X1 U9460 ( .A1(n12925), .A2(n7572), .ZN(n7569) );
  AND2_X1 U9461 ( .A1(n8376), .A2(n8338), .ZN(n8374) );
  NAND4_X1 U9462 ( .A1(n8361), .A2(n8376), .A3(n8338), .A4(n7576), .ZN(n8459)
         );
  XNOR2_X2 U9463 ( .A(n8461), .B(n8460), .ZN(n12984) );
  NAND2_X1 U9464 ( .A1(n7578), .A2(n13437), .ZN(n13363) );
  XNOR2_X1 U9465 ( .A(n7579), .B(n13358), .ZN(n7578) );
  NAND2_X1 U9466 ( .A1(n7580), .A2(n8197), .ZN(n7579) );
  NAND2_X1 U9467 ( .A1(n13388), .A2(n7411), .ZN(n7580) );
  CLKBUF_X1 U9468 ( .A(n7582), .Z(n7581) );
  NAND4_X1 U9469 ( .A1(n8182), .A2(n7582), .A3(n8406), .A4(n8346), .ZN(n8181)
         );
  NAND2_X1 U9470 ( .A1(n7581), .A2(n8406), .ZN(n8395) );
  NAND2_X1 U9471 ( .A1(n7581), .A2(n8346), .ZN(n8185) );
  NOR2_X1 U9472 ( .A1(n8405), .A2(n7581), .ZN(n7583) );
  NAND2_X1 U9473 ( .A1(n7588), .A2(n7587), .ZN(n13896) );
  INV_X1 U9474 ( .A(n7589), .ZN(n12800) );
  XNOR2_X1 U9475 ( .A(n8433), .B(n11019), .ZN(n12801) );
  OAI211_X1 U9476 ( .C1(n14435), .C2(n7606), .A(n7604), .B(n7603), .ZN(n14346)
         );
  NAND3_X1 U9477 ( .A1(n7611), .A2(n7417), .A3(n12789), .ZN(n7610) );
  NAND2_X1 U9478 ( .A1(n7624), .A2(n7622), .ZN(n12785) );
  NAND2_X1 U9479 ( .A1(n11429), .A2(n7628), .ZN(n11629) );
  NAND2_X2 U9480 ( .A1(n10845), .A2(n10844), .ZN(n10853) );
  NAND2_X2 U9481 ( .A1(n10825), .A2(n12739), .ZN(n10844) );
  NAND3_X1 U9482 ( .A1(n7629), .A2(n7846), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n7843) );
  NAND3_X1 U9483 ( .A1(n8070), .A2(n8069), .A3(n8071), .ZN(n8779) );
  NAND2_X1 U9484 ( .A1(n8612), .A2(n7633), .ZN(n7630) );
  NAND2_X1 U9485 ( .A1(n7630), .A2(n7436), .ZN(n8739) );
  NAND3_X1 U9486 ( .A1(n7642), .A2(n7641), .A3(n13057), .ZN(n15280) );
  NAND3_X1 U9487 ( .A1(n7642), .A2(n7641), .A3(n7639), .ZN(n15281) );
  INV_X1 U9488 ( .A(n13055), .ZN(n7644) );
  NAND2_X1 U9489 ( .A1(n7645), .A2(n7791), .ZN(n13056) );
  INV_X1 U9490 ( .A(n7647), .ZN(n8075) );
  NAND2_X1 U9491 ( .A1(n15259), .A2(n8290), .ZN(n8288) );
  MUX2_X1 U9492 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n10976), .Z(n7658) );
  NAND2_X1 U9493 ( .A1(n14983), .A2(n11487), .ZN(n11491) );
  NAND3_X1 U9494 ( .A1(n11476), .A2(n7659), .A3(n11475), .ZN(n14983) );
  NAND2_X1 U9495 ( .A1(n15095), .A2(n7667), .ZN(n7666) );
  NAND2_X1 U9496 ( .A1(n15095), .A2(n14961), .ZN(n14962) );
  OAI211_X1 U9497 ( .C1(n15095), .C2(n7484), .A(n7668), .B(n7666), .ZN(n15016)
         );
  NAND2_X1 U9498 ( .A1(n9190), .A2(n8999), .ZN(n9196) );
  NAND3_X1 U9499 ( .A1(n11963), .A2(n11962), .A3(n8344), .ZN(n7691) );
  NAND2_X1 U9500 ( .A1(n15398), .A2(n7692), .ZN(n15507) );
  INV_X2 U9501 ( .A(n9513), .ZN(n9359) );
  NAND2_X4 U9502 ( .A1(n9059), .A2(n10984), .ZN(n9513) );
  OR2_X1 U9503 ( .A1(n12457), .A2(n7702), .ZN(n7701) );
  NAND2_X1 U9504 ( .A1(n7701), .A2(n7699), .ZN(n12686) );
  NAND2_X1 U9505 ( .A1(n15331), .A2(n7456), .ZN(n7706) );
  NAND2_X1 U9506 ( .A1(n7706), .A2(n7429), .ZN(n7704) );
  NAND2_X1 U9507 ( .A1(n7704), .A2(n7462), .ZN(n15302) );
  INV_X1 U9508 ( .A(n7763), .ZN(n7709) );
  NAND4_X1 U9509 ( .A1(n7372), .A2(n7761), .A3(n7470), .A4(n7709), .ZN(n9596)
         );
  AND3_X1 U9510 ( .A1(n7372), .A2(n9004), .A3(n7761), .ZN(n7711) );
  NAND3_X1 U9511 ( .A1(n7711), .A2(n7713), .A3(n7712), .ZN(n9025) );
  NOR2_X1 U9512 ( .A1(n7722), .A2(n13344), .ZN(n7716) );
  OAI211_X1 U9513 ( .C1(n15277), .C2(n7461), .A(n7718), .B(n7715), .ZN(n13343)
         );
  NAND3_X1 U9514 ( .A1(n7719), .A2(n15277), .A3(n8258), .ZN(n7718) );
  NAND2_X1 U9515 ( .A1(n7370), .A2(n8499), .ZN(n7728) );
  OAI21_X1 U9516 ( .B1(n7370), .B2(n8499), .A(n7728), .ZN(n12004) );
  NAND2_X1 U9517 ( .A1(n12005), .A2(n12004), .ZN(n12009) );
  NAND2_X1 U9518 ( .A1(n12009), .A2(n8469), .ZN(n8470) );
  INV_X2 U9519 ( .A(n16214), .ZN(n16225) );
  AND2_X2 U9520 ( .A1(n8812), .A2(n8813), .ZN(n16214) );
  AND2_X2 U9521 ( .A1(n8767), .A2(n8766), .ZN(n16360) );
  INV_X1 U9522 ( .A(n7746), .ZN(n14633) );
  NAND3_X1 U9523 ( .A1(n7747), .A2(n7749), .A3(n12213), .ZN(n12662) );
  NAND3_X1 U9524 ( .A1(n7753), .A2(n14521), .A3(n14511), .ZN(n7750) );
  NAND4_X1 U9525 ( .A1(n7372), .A2(n7757), .A3(n7761), .A4(n7756), .ZN(n7755)
         );
  NOR2_X2 U9526 ( .A1(n7762), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n7761) );
  NAND3_X1 U9527 ( .A1(n8996), .A2(n8995), .A3(n8998), .ZN(n7759) );
  NAND4_X1 U9528 ( .A1(n13875), .A2(n7689), .A3(n9036), .A4(n9039), .ZN(n7762)
         );
  NAND2_X1 U9529 ( .A1(n7466), .A2(n12676), .ZN(n15404) );
  OR3_X1 U9530 ( .A1(n15284), .A2(n15274), .A3(n15436), .ZN(n15251) );
  NOR2_X1 U9531 ( .A1(n15284), .A2(n15274), .ZN(n15268) );
  AND2_X2 U9532 ( .A1(n12714), .A2(n12713), .ZN(n12717) );
  NAND2_X1 U9533 ( .A1(n9009), .A2(n7777), .ZN(n7776) );
  OAI21_X1 U9534 ( .B1(n15395), .B2(n7784), .A(n7479), .ZN(n15381) );
  INV_X1 U9535 ( .A(n13056), .ZN(n15292) );
  NAND2_X2 U9536 ( .A1(n13346), .A2(n13347), .ZN(n15431) );
  NAND3_X1 U9537 ( .A1(n7837), .A2(n8593), .A3(n8592), .ZN(n8807) );
  NAND2_X1 U9538 ( .A1(n7837), .A2(n8593), .ZN(n8805) );
  NAND2_X1 U9539 ( .A1(n8589), .A2(n10969), .ZN(n7837) );
  INV_X1 U9540 ( .A(n7846), .ZN(n7841) );
  NAND3_X1 U9541 ( .A1(n7840), .A2(n7842), .A3(n7843), .ZN(n7838) );
  NAND4_X1 U9542 ( .A1(n7843), .A2(n7842), .A3(n7840), .A4(n7839), .ZN(n7845)
         );
  NAND2_X1 U9543 ( .A1(n7480), .A2(n12081), .ZN(n11890) );
  NAND2_X1 U9544 ( .A1(n10547), .A2(n10546), .ZN(n14539) );
  NOR2_X1 U9545 ( .A1(n10549), .A2(n7851), .ZN(n7850) );
  INV_X1 U9546 ( .A(n10546), .ZN(n7851) );
  OAI21_X1 U9547 ( .B1(n14605), .B2(n7854), .A(n7477), .ZN(n10543) );
  NAND2_X1 U9548 ( .A1(n14514), .A2(n14513), .ZN(n14512) );
  AOI21_X2 U9549 ( .B1(n14036), .B2(n14038), .A(n7876), .ZN(n8339) );
  OR2_X1 U9550 ( .A1(n7908), .A2(n7881), .ZN(n8411) );
  NAND2_X1 U9551 ( .A1(n8345), .A2(n8406), .ZN(n7882) );
  NAND2_X1 U9552 ( .A1(n7468), .A2(n7908), .ZN(n7883) );
  OR2_X1 U9553 ( .A1(n7908), .A2(n7886), .ZN(n7885) );
  NAND2_X1 U9554 ( .A1(n7890), .A2(n7891), .ZN(n13034) );
  NAND2_X1 U9555 ( .A1(n12919), .A2(n7893), .ZN(n7890) );
  AND3_X1 U9556 ( .A1(n13145), .A2(n13146), .A3(n13137), .ZN(n7901) );
  NAND2_X1 U9557 ( .A1(n16174), .A2(n13146), .ZN(n12117) );
  NAND2_X1 U9558 ( .A1(n13145), .A2(n13146), .ZN(n16177) );
  NAND2_X1 U9559 ( .A1(n10065), .A2(n13137), .ZN(n16176) );
  OAI21_X1 U9560 ( .B1(n14017), .B2(n7906), .A(n7902), .ZN(n13978) );
  NAND2_X1 U9561 ( .A1(n8364), .A2(n8243), .ZN(n8457) );
  INV_X1 U9562 ( .A(n9614), .ZN(n9617) );
  NAND2_X1 U9563 ( .A1(n9614), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U9564 ( .A1(n13937), .A2(n7910), .ZN(n7909) );
  OAI211_X1 U9565 ( .C1(n13937), .C2(n7911), .A(n7909), .B(n8330), .ZN(
        P3_U3201) );
  INV_X1 U9566 ( .A(n8575), .ZN(n7915) );
  NAND2_X1 U9567 ( .A1(n7920), .A2(n7921), .ZN(n8433) );
  NAND2_X1 U9568 ( .A1(n12229), .A2(n8552), .ZN(n7920) );
  NAND2_X1 U9569 ( .A1(n12082), .A2(n12088), .ZN(n12081) );
  NAND2_X1 U9570 ( .A1(n7369), .A2(n8670), .ZN(n8677) );
  MUX2_X2 U9571 ( .A(n10244), .B(n10243), .S(n16473), .Z(n10245) );
  OAI211_X2 U9572 ( .C1(n9781), .C2(n10972), .A(n9754), .B(n9753), .ZN(n16333)
         );
  AND3_X2 U9573 ( .A1(n9065), .A2(n9063), .A3(n9064), .ZN(n16155) );
  NAND2_X2 U9574 ( .A1(n8957), .A2(n14808), .ZN(n8827) );
  NAND2_X1 U9575 ( .A1(n10295), .A2(n7923), .ZN(n16215) );
  NAND2_X1 U9576 ( .A1(n11740), .A2(n11757), .ZN(n7923) );
  XNOR2_X2 U9577 ( .A(n10571), .B(n11752), .ZN(n11757) );
  NAND4_X1 U9578 ( .A1(n10294), .A2(n10291), .A3(n10292), .A4(n10293), .ZN(
        n10571) );
  NAND2_X1 U9579 ( .A1(n8862), .A2(n7925), .ZN(n7924) );
  XNOR2_X1 U9580 ( .A(n10503), .B(n10552), .ZN(n7932) );
  NAND3_X1 U9581 ( .A1(n7929), .A2(n7927), .A3(n7926), .ZN(n10563) );
  NAND2_X1 U9582 ( .A1(n12665), .A2(n7936), .ZN(n7935) );
  NAND2_X1 U9583 ( .A1(n7944), .A2(n7942), .ZN(n14488) );
  NAND2_X1 U9584 ( .A1(n11457), .A2(n11456), .ZN(n11455) );
  NAND2_X1 U9585 ( .A1(n7945), .A2(n7946), .ZN(n10469) );
  NAND2_X1 U9586 ( .A1(n14556), .A2(n10457), .ZN(n7945) );
  OAI21_X1 U9587 ( .B1(n10359), .B2(n7956), .A(n7953), .ZN(n10380) );
  OR2_X2 U9588 ( .A1(n7965), .A2(n15843), .ZN(n7964) );
  NAND2_X1 U9589 ( .A1(n7968), .A2(n7972), .ZN(n9643) );
  NAND2_X1 U9590 ( .A1(n9640), .A2(n7969), .ZN(n7968) );
  NAND2_X1 U9591 ( .A1(n9802), .A2(n7977), .ZN(n7975) );
  NAND3_X1 U9592 ( .A1(n13287), .A2(n13289), .A3(n7984), .ZN(n7980) );
  NAND2_X1 U9593 ( .A1(n7984), .A2(n7983), .ZN(n7987) );
  NAND2_X1 U9594 ( .A1(n9867), .A2(n7999), .ZN(n7996) );
  NAND2_X1 U9595 ( .A1(n7996), .A2(n7997), .ZN(n9895) );
  NAND2_X1 U9596 ( .A1(n9699), .A2(n7457), .ZN(n8002) );
  NAND2_X1 U9597 ( .A1(n9699), .A2(n9697), .ZN(n8005) );
  NAND2_X1 U9598 ( .A1(n8002), .A2(n8003), .ZN(n9724) );
  NOR2_X1 U9599 ( .A1(n13235), .A2(n8006), .ZN(n13236) );
  NAND2_X1 U9600 ( .A1(n8007), .A2(n13295), .ZN(n8006) );
  NAND2_X1 U9601 ( .A1(n8009), .A2(n8010), .ZN(n8007) );
  INV_X1 U9602 ( .A(n13126), .ZN(n8009) );
  NOR2_X1 U9603 ( .A1(n13126), .A2(n13125), .ZN(n13240) );
  NAND2_X1 U9604 ( .A1(n9934), .A2(n7501), .ZN(n8021) );
  NAND2_X1 U9605 ( .A1(n8673), .A2(n8672), .ZN(n8952) );
  NAND2_X1 U9606 ( .A1(n8673), .A2(n8066), .ZN(n14796) );
  NAND2_X1 U9607 ( .A1(n8590), .A2(SI_2_), .ZN(n8593) );
  NAND2_X1 U9608 ( .A1(n8726), .A2(n8725), .ZN(n8068) );
  NAND2_X1 U9609 ( .A1(n8068), .A2(n8067), .ZN(n8631) );
  NAND2_X1 U9610 ( .A1(n8797), .A2(n8596), .ZN(n8788) );
  AOI21_X1 U9611 ( .B1(n8697), .B2(n8084), .A(n8081), .ZN(n8078) );
  OAI21_X1 U9612 ( .B1(n8697), .B2(n8698), .A(n8638), .ZN(n8694) );
  NAND2_X1 U9613 ( .A1(n8613), .A2(n8750), .ZN(n8835) );
  NAND3_X1 U9614 ( .A1(n8613), .A2(n8096), .A3(n8750), .ZN(n8088) );
  NAND3_X1 U9615 ( .A1(n8613), .A2(n8750), .A3(n8090), .ZN(n8089) );
  NAND2_X1 U9616 ( .A1(n8646), .A2(n8645), .ZN(n9405) );
  NAND2_X1 U9617 ( .A1(n8645), .A2(n8104), .ZN(n8103) );
  NAND2_X1 U9618 ( .A1(n11037), .A2(n11565), .ZN(n8106) );
  NAND2_X1 U9619 ( .A1(n11041), .A2(n8107), .ZN(n11084) );
  INV_X1 U9620 ( .A(n8109), .ZN(n8108) );
  OAI22_X1 U9621 ( .A1(n15000), .A2(n16142), .B1(n11039), .B2(n11496), .ZN(
        n8109) );
  NAND2_X1 U9622 ( .A1(n12649), .A2(n8112), .ZN(n8111) );
  NAND3_X1 U9623 ( .A1(n8121), .A2(n8120), .A3(n8127), .ZN(n8119) );
  NAND2_X1 U9624 ( .A1(n10726), .A2(n10725), .ZN(n8121) );
  NAND3_X1 U9625 ( .A1(n8124), .A2(n8123), .A3(n8128), .ZN(n8122) );
  NAND2_X1 U9626 ( .A1(n10726), .A2(n8126), .ZN(n8124) );
  NAND2_X1 U9627 ( .A1(n7369), .A2(n8335), .ZN(n8941) );
  NAND2_X1 U9628 ( .A1(n10741), .A2(n10740), .ZN(n8145) );
  NAND2_X1 U9629 ( .A1(n8144), .A2(n8146), .ZN(n10746) );
  NAND2_X1 U9630 ( .A1(n8149), .A2(n8152), .ZN(n8148) );
  AOI21_X1 U9631 ( .B1(n14917), .B2(n8151), .A(n8150), .ZN(n8149) );
  OAI211_X1 U9632 ( .C1(n7437), .C2(n10627), .A(n10622), .B(n10623), .ZN(n8154) );
  NAND2_X1 U9633 ( .A1(n8154), .A2(n8153), .ZN(n10632) );
  NAND2_X1 U9634 ( .A1(n8156), .A2(n8155), .ZN(n10719) );
  NAND2_X1 U9635 ( .A1(n8158), .A2(n8157), .ZN(n8156) );
  INV_X1 U9636 ( .A(n10708), .ZN(n8158) );
  NAND3_X1 U9637 ( .A1(n10657), .A2(n7463), .A3(n7383), .ZN(n8162) );
  NAND2_X1 U9638 ( .A1(n8162), .A2(n7478), .ZN(n10669) );
  NAND3_X1 U9639 ( .A1(n8165), .A2(n7448), .A3(n8164), .ZN(n8167) );
  INV_X1 U9640 ( .A(n10633), .ZN(n8165) );
  NAND2_X1 U9641 ( .A1(n8167), .A2(n8166), .ZN(n10645) );
  NAND2_X1 U9642 ( .A1(n8168), .A2(n10637), .ZN(n8166) );
  NAND2_X1 U9643 ( .A1(n8169), .A2(n8172), .ZN(n10706) );
  NAND2_X1 U9644 ( .A1(n8171), .A2(n8170), .ZN(n8169) );
  NAND2_X1 U9645 ( .A1(n8174), .A2(n8175), .ZN(n10685) );
  NAND3_X1 U9646 ( .A1(n10674), .A2(n7464), .A3(n10673), .ZN(n8174) );
  NAND3_X1 U9647 ( .A1(n8178), .A2(n8177), .A3(n8176), .ZN(n10612) );
  OR2_X1 U9648 ( .A1(n10605), .A2(n10606), .ZN(n8177) );
  NAND3_X1 U9649 ( .A1(n8179), .A2(n10598), .A3(n10599), .ZN(n8178) );
  NAND2_X1 U9650 ( .A1(n10605), .A2(n10606), .ZN(n8179) );
  NOR2_X2 U9651 ( .A1(n8181), .A2(n8186), .ZN(n8376) );
  NAND4_X1 U9652 ( .A1(n8345), .A2(n8401), .A3(n8406), .A4(n8403), .ZN(n8184)
         );
  NAND3_X1 U9653 ( .A1(n8401), .A2(n8403), .A3(n8347), .ZN(n8186) );
  OAI21_X1 U9654 ( .B1(n13412), .B2(n10196), .A(n10195), .ZN(n13388) );
  OAI21_X1 U9655 ( .B1(n13412), .B2(n8192), .A(n8191), .ZN(n8190) );
  NAND2_X1 U9656 ( .A1(n13405), .A2(n8205), .ZN(n8202) );
  INV_X1 U9657 ( .A(n12999), .ZN(n8211) );
  NAND2_X1 U9658 ( .A1(n8218), .A2(n8217), .ZN(n11994) );
  NAND2_X1 U9659 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  NAND2_X1 U9660 ( .A1(n13025), .A2(n8222), .ZN(n8219) );
  NAND2_X1 U9661 ( .A1(n8219), .A2(n8220), .ZN(n14143) );
  NAND2_X1 U9662 ( .A1(n8225), .A2(n7471), .ZN(n12325) );
  OAI211_X1 U9663 ( .C1(n9691), .C2(n13143), .A(n16181), .B(n8226), .ZN(n9703)
         );
  NAND2_X1 U9664 ( .A1(n8228), .A2(n8227), .ZN(n16182) );
  NAND2_X1 U9665 ( .A1(n13143), .A2(n13137), .ZN(n8228) );
  AND2_X1 U9666 ( .A1(n8364), .A2(n8362), .ZN(n8455) );
  NAND2_X1 U9667 ( .A1(n14006), .A2(n13108), .ZN(n13110) );
  INV_X1 U9668 ( .A(n11586), .ZN(n8253) );
  OAI21_X1 U9669 ( .B1(n11808), .B2(n8251), .A(n8248), .ZN(n11956) );
  NAND2_X1 U9670 ( .A1(n11956), .A2(n11955), .ZN(n11958) );
  NAND2_X1 U9671 ( .A1(n12955), .A2(n8260), .ZN(n15398) );
  NAND2_X1 U9672 ( .A1(n8264), .A2(n7644), .ZN(n8266) );
  INV_X1 U9673 ( .A(n15302), .ZN(n8264) );
  NOR2_X1 U9674 ( .A1(n15301), .A2(n8336), .ZN(n15278) );
  INV_X1 U9675 ( .A(n8343), .ZN(n8271) );
  NAND2_X2 U9676 ( .A1(n8272), .A2(n9547), .ZN(n16139) );
  OR2_X1 U9677 ( .A1(n16155), .A2(n15143), .ZN(n8272) );
  NAND3_X1 U9678 ( .A1(n12345), .A2(n12346), .A3(n12344), .ZN(n12457) );
  XNOR2_X2 U9679 ( .A(n8273), .B(n9028), .ZN(n15689) );
  AND2_X2 U9680 ( .A1(n13090), .A2(n9015), .ZN(n9075) );
  OR2_X1 U9681 ( .A1(n9015), .A2(P1_U3086), .ZN(n8274) );
  OAI21_X1 U9682 ( .B1(n15333), .B2(n8294), .A(n15332), .ZN(n15479) );
  OAI22_X2 U9683 ( .A1(n9181), .A2(n8296), .B1(n9182), .B2(n8295), .ZN(n9208)
         );
  NAND2_X1 U9684 ( .A1(n9208), .A2(n9207), .ZN(n9195) );
  OAI211_X1 U9685 ( .C1(n8306), .C2(n8304), .A(n8301), .B(n8300), .ZN(P1_U3242) );
  NAND2_X1 U9686 ( .A1(n9594), .A2(n8302), .ZN(n8300) );
  NAND2_X1 U9687 ( .A1(n7547), .A2(n8303), .ZN(n8301) );
  NAND3_X1 U9688 ( .A1(n9135), .A2(n9134), .A3(n8311), .ZN(n8310) );
  NAND3_X1 U9689 ( .A1(n9452), .A2(n9451), .A3(n7473), .ZN(n8312) );
  NAND3_X1 U9690 ( .A1(n9228), .A2(n9227), .A3(n7476), .ZN(n8315) );
  NAND2_X1 U9691 ( .A1(n8315), .A2(n8316), .ZN(n9256) );
  NAND2_X1 U9692 ( .A1(n8318), .A2(n8319), .ZN(n9447) );
  NAND3_X1 U9693 ( .A1(n9426), .A2(n7481), .A3(n9425), .ZN(n8318) );
  NAND2_X1 U9694 ( .A1(n8325), .A2(n8327), .ZN(n9421) );
  NAND3_X1 U9695 ( .A1(n9399), .A2(n9398), .A3(n8326), .ZN(n8325) );
  NAND2_X1 U9696 ( .A1(n8631), .A2(n8630), .ZN(n8861) );
  AOI21_X2 U9697 ( .B1(n15854), .B2(n15853), .A(n7394), .ZN(n15866) );
  INV_X1 U9698 ( .A(n14480), .ZN(n8927) );
  INV_X1 U9699 ( .A(n10455), .ZN(n14772) );
  NAND2_X1 U9700 ( .A1(n14685), .A2(n16516), .ZN(n8994) );
  NAND2_X1 U9701 ( .A1(n14817), .A2(n9512), .ZN(n9434) );
  INV_X1 U9702 ( .A(n10594), .ZN(n10597) );
  OAI21_X1 U9703 ( .B1(n15431), .B2(n16485), .A(n15430), .ZN(n15432) );
  AND2_X1 U9704 ( .A1(n16469), .A2(n13965), .ZN(n10084) );
  OR2_X1 U9705 ( .A1(n11987), .A2(n16202), .ZN(n9694) );
  OR2_X1 U9706 ( .A1(n10986), .A2(n9481), .ZN(n9093) );
  AOI22_X1 U9707 ( .A1(n9359), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9358), .B2(
        n15163), .ZN(n9092) );
  AOI21_X1 U9708 ( .B1(n14509), .B2(n10483), .A(n10482), .ZN(n14440) );
  INV_X1 U9709 ( .A(n10483), .ZN(n10496) );
  NAND2_X2 U9710 ( .A1(n9621), .A2(n14317), .ZN(n11987) );
  OAI21_X1 U9711 ( .B1(n9110), .B2(n9109), .A(n9106), .ZN(n9115) );
  OAI21_X2 U9712 ( .B1(n9115), .B2(n9114), .A(n9113), .ZN(n9130) );
  NOR2_X1 U9713 ( .A1(n13701), .A2(n13700), .ZN(n8329) );
  INV_X2 U9714 ( .A(n13471), .ZN(P3_U3897) );
  AND2_X1 U9715 ( .A1(n10772), .A2(n10771), .ZN(n8331) );
  AND2_X1 U9716 ( .A1(n10796), .A2(n10795), .ZN(n8332) );
  AND2_X1 U9717 ( .A1(n14788), .A2(n14626), .ZN(n8333) );
  INV_X1 U9718 ( .A(n14721), .ZN(n8873) );
  AND2_X2 U9719 ( .A1(n10556), .A2(n10924), .ZN(n16512) );
  AND2_X2 U9720 ( .A1(n10556), .A2(n15570), .ZN(n16516) );
  INV_X1 U9721 ( .A(n16516), .ZN(n16513) );
  NOR2_X1 U9722 ( .A1(n10930), .A2(n12843), .ZN(n8334) );
  AND4_X1 U9723 ( .A1(n8939), .A2(n8945), .A3(n8938), .A4(n8937), .ZN(n8335)
         );
  AND2_X1 U9724 ( .A1(n15299), .A2(n15122), .ZN(n8336) );
  INV_X1 U9725 ( .A(n16495), .ZN(n15501) );
  AND2_X2 U9726 ( .A1(n13079), .A2(n16104), .ZN(n16153) );
  OR2_X1 U9727 ( .A1(n11600), .A2(n11599), .ZN(n16540) );
  OR2_X1 U9728 ( .A1(n11600), .A2(n11789), .ZN(n16537) );
  OR2_X1 U9729 ( .A1(n13963), .A2(n14227), .ZN(n8337) );
  INV_X1 U9730 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14795) );
  NAND2_X2 U9731 ( .A1(n16194), .A2(n11924), .ZN(n14169) );
  INV_X1 U9732 ( .A(n9980), .ZN(n9670) );
  INV_X1 U9733 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n12180) );
  INV_X1 U9734 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8585) );
  INV_X1 U9735 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12740) );
  INV_X1 U9736 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n12338) );
  INV_X1 U9737 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n12024) );
  AND4_X1 U9738 ( .A1(n8349), .A2(n8348), .A3(n8378), .A4(n8388), .ZN(n8338)
         );
  INV_X1 U9739 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13015) );
  INV_X1 U9740 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12558) );
  INV_X1 U9741 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12771) );
  AND2_X1 U9742 ( .A1(n15932), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8340) );
  AND2_X1 U9743 ( .A1(n10780), .A2(n8331), .ZN(n8341) );
  CLKBUF_X3 U9744 ( .A(n10157), .Z(n10199) );
  NAND2_X1 U9745 ( .A1(n10120), .A2(n10119), .ZN(n10157) );
  INV_X1 U9746 ( .A(n13313), .ZN(n12759) );
  AND2_X1 U9747 ( .A1(n10164), .A2(n14160), .ZN(n8342) );
  AND2_X1 U9748 ( .A1(n15370), .A2(n15088), .ZN(n8343) );
  OR2_X1 U9749 ( .A1(n16388), .A2(n12365), .ZN(n8344) );
  BUF_X4 U9750 ( .A(n9692), .Z(n10035) );
  INV_X1 U9751 ( .A(n11807), .ZN(n9106) );
  AOI21_X1 U9752 ( .B1(n9110), .B2(n9109), .A(n9108), .ZN(n9114) );
  INV_X1 U9753 ( .A(n10595), .ZN(n10596) );
  AOI21_X1 U9754 ( .B1(n12101), .B2(n10759), .A(n10602), .ZN(n10608) );
  NAND2_X1 U9755 ( .A1(n9169), .A2(n9168), .ZN(n9181) );
  XNOR2_X1 U9756 ( .A(SI_19_), .B(keyinput_13), .ZN(n13684) );
  OAI21_X1 U9757 ( .B1(n12247), .B2(n10789), .A(n10642), .ZN(n10643) );
  NAND2_X1 U9758 ( .A1(n9261), .A2(n9260), .ZN(n9277) );
  NAND2_X1 U9759 ( .A1(n13704), .A2(n13703), .ZN(n13710) );
  INV_X1 U9760 ( .A(n10670), .ZN(n10671) );
  OAI22_X1 U9761 ( .A1(n13723), .A2(keyinput_36), .B1(n13722), .B2(
        P3_REG3_REG_27__SCAN_IN), .ZN(n13724) );
  INV_X1 U9762 ( .A(n13724), .ZN(n13725) );
  NAND2_X1 U9763 ( .A1(n13721), .A2(n13720), .ZN(n13726) );
  XNOR2_X1 U9764 ( .A(keyinput_39), .B(P3_REG3_REG_10__SCAN_IN), .ZN(n13729)
         );
  NAND2_X1 U9765 ( .A1(n10683), .A2(n10682), .ZN(n10690) );
  OAI22_X1 U9766 ( .A1(n13751), .A2(keyinput_51), .B1(n13750), .B2(
        P3_REG3_REG_24__SCAN_IN), .ZN(n13752) );
  OAI22_X1 U9767 ( .A1(n13756), .A2(n13755), .B1(P3_REG3_REG_4__SCAN_IN), .B2(
        keyinput_52), .ZN(n13757) );
  INV_X1 U9768 ( .A(n13757), .ZN(n13758) );
  NAND2_X1 U9769 ( .A1(n13759), .A2(n13758), .ZN(n13765) );
  INV_X1 U9770 ( .A(keyinput_76), .ZN(n13797) );
  NAND2_X1 U9771 ( .A1(n13798), .A2(n13797), .ZN(n13800) );
  AND2_X1 U9772 ( .A1(n13800), .A2(n13799), .ZN(n13801) );
  XNOR2_X1 U9773 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n13813)
         );
  NOR2_X1 U9774 ( .A1(n13814), .A2(n13813), .ZN(n13815) );
  NOR3_X1 U9775 ( .A1(n13328), .A2(n13239), .A3(n13238), .ZN(n13244) );
  INV_X1 U9776 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8355) );
  AOI211_X1 U9777 ( .C1(n13851), .C2(n13850), .A(n13849), .B(n13848), .ZN(
        n13854) );
  NAND2_X1 U9778 ( .A1(n13295), .A2(n13291), .ZN(n13126) );
  INV_X1 U9779 ( .A(n14144), .ZN(n9877) );
  INV_X1 U9780 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9665) );
  INV_X1 U9781 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8580) );
  OR4_X1 U9782 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8982) );
  OR2_X1 U9783 ( .A1(n16155), .A2(n15000), .ZN(n11078) );
  INV_X1 U9784 ( .A(n12452), .ZN(n12346) );
  OR4_X1 U9785 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n11048) );
  INV_X1 U9786 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8999) );
  INV_X1 U9787 ( .A(n13287), .ZN(n13288) );
  INV_X1 U9788 ( .A(n14317), .ZN(n9622) );
  INV_X1 U9789 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13748) );
  OAI22_X1 U9790 ( .A1(n14058), .A2(n9955), .B1(n14041), .B2(n14199), .ZN(
        n14037) );
  INV_X1 U9791 ( .A(n13302), .ZN(n9743) );
  INV_X1 U9792 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8362) );
  INV_X1 U9793 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9656) );
  INV_X1 U9794 ( .A(n10424), .ZN(n10254) );
  AND2_X1 U9795 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10309) );
  INV_X1 U9796 ( .A(n10369), .ZN(n10249) );
  INV_X1 U9797 ( .A(n14529), .ZN(n10820) );
  NOR2_X1 U9798 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  INV_X1 U9799 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9233) );
  OR2_X1 U9800 ( .A1(n15334), .A2(n13070), .ZN(n13071) );
  INV_X1 U9801 ( .A(n15397), .ZN(n12956) );
  INV_X1 U9802 ( .A(SI_22_), .ZN(n8644) );
  NOR2_X1 U9803 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9291) );
  INV_X1 U9804 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9144) );
  INV_X1 U9805 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9870) );
  AND2_X1 U9806 ( .A1(n15548), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9671) );
  INV_X1 U9807 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9646) );
  AND2_X1 U9808 ( .A1(n10786), .A2(n10785), .ZN(n10787) );
  OR2_X1 U9809 ( .A1(n10470), .A2(n14441), .ZN(n10487) );
  NAND2_X1 U9810 ( .A1(n10254), .A2(n10253), .ZN(n10435) );
  OR2_X1 U9811 ( .A1(n10422), .A2(n10421), .ZN(n10424) );
  INV_X1 U9812 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10381) );
  INV_X1 U9813 ( .A(n16512), .ZN(n14686) );
  OR2_X1 U9814 ( .A1(n12987), .A2(n12877), .ZN(n10831) );
  INV_X1 U9815 ( .A(n9427), .ZN(n9438) );
  INV_X1 U9816 ( .A(n9411), .ZN(n9428) );
  AND2_X1 U9817 ( .A1(n9519), .A2(n9540), .ZN(n9518) );
  AND2_X1 U9818 ( .A1(n9351), .A2(n9016), .ZN(n9365) );
  NAND2_X1 U9819 ( .A1(n15428), .A2(n15119), .ZN(n13062) );
  INV_X1 U9820 ( .A(n16493), .ZN(n12677) );
  OR2_X1 U9821 ( .A1(n12273), .A2(n16421), .ZN(n12350) );
  INV_X1 U9822 ( .A(n8895), .ZN(n8883) );
  NAND2_X1 U9823 ( .A1(n8629), .A2(SI_16_), .ZN(n8630) );
  INV_X1 U9824 ( .A(n8804), .ZN(n8592) );
  AND2_X1 U9825 ( .A1(n9769), .A2(n13737), .ZN(n9783) );
  INV_X1 U9826 ( .A(n14042), .ZN(n14009) );
  AND2_X1 U9827 ( .A1(n9871), .A2(n9870), .ZN(n9886) );
  NOR2_X1 U9828 ( .A1(n9969), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U9829 ( .A1(n9833), .A2(n13555), .ZN(n9846) );
  OR2_X1 U9830 ( .A1(n9899), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9911) );
  AND2_X1 U9831 ( .A1(n10104), .A2(n11932), .ZN(n13332) );
  AND3_X1 U9832 ( .A1(n12880), .A2(n12633), .A3(n10087), .ZN(n8463) );
  INV_X1 U9833 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15733) );
  OAI21_X1 U9834 ( .B1(n7370), .B2(n16202), .A(n8407), .ZN(n12003) );
  INV_X1 U9835 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n13745) );
  AND2_X1 U9836 ( .A1(n8490), .A2(n8491), .ZN(n8488) );
  INV_X1 U9837 ( .A(n13463), .ZN(n14027) );
  NAND2_X1 U9838 ( .A1(n9937), .A2(n13740), .ZN(n9948) );
  AND4_X1 U9839 ( .A1(n9904), .A2(n9903), .A3(n9902), .A4(n9901), .ZN(n14108)
         );
  AND2_X1 U9840 ( .A1(n9892), .A2(n10077), .ZN(n13321) );
  AND4_X1 U9841 ( .A1(n9864), .A2(n9863), .A3(n9862), .A4(n9861), .ZN(n14146)
         );
  INV_X1 U9842 ( .A(n14163), .ZN(n16194) );
  INV_X1 U9843 ( .A(n14305), .ZN(n11917) );
  INV_X1 U9844 ( .A(n10108), .ZN(n10236) );
  INV_X1 U9845 ( .A(n13997), .ZN(n13993) );
  INV_X1 U9846 ( .A(n13318), .ZN(n12918) );
  AND2_X1 U9847 ( .A1(n10106), .A2(n10047), .ZN(n14156) );
  AND2_X1 U9848 ( .A1(n13336), .A2(n10214), .ZN(n10110) );
  INV_X1 U9849 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8353) );
  INV_X1 U9850 ( .A(n9979), .ZN(n9981) );
  OAI21_X1 U9851 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(n11403), .A(n9647), .ZN(
        n9648) );
  OR2_X1 U9852 ( .A1(n10437), .A2(n10255), .ZN(n10448) );
  INV_X1 U9853 ( .A(n14626), .ZN(n14360) );
  INV_X1 U9854 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n11509) );
  INV_X1 U9855 ( .A(n14652), .ZN(n14627) );
  OR2_X1 U9856 ( .A1(n14495), .A2(n10496), .ZN(n10493) );
  OR2_X1 U9857 ( .A1(n11247), .A2(n11246), .ZN(n11540) );
  OR2_X1 U9858 ( .A1(n11939), .A2(n11938), .ZN(n12815) );
  OR2_X1 U9859 ( .A1(n11124), .A2(n11102), .ZN(n15645) );
  INV_X1 U9860 ( .A(n14691), .ZN(n8926) );
  INV_X1 U9861 ( .A(n14513), .ZN(n14503) );
  INV_X1 U9862 ( .A(n12935), .ZN(n14644) );
  OR3_X1 U9863 ( .A1(n10383), .A2(n10382), .A3(n10381), .ZN(n10394) );
  INV_X1 U9864 ( .A(n16399), .ZN(n14648) );
  NAND2_X1 U9865 ( .A1(n16513), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8990) );
  INV_X1 U9866 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10561) );
  NAND2_X1 U9867 ( .A1(n10842), .A2(n12739), .ZN(n10835) );
  INV_X1 U9868 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8974) );
  INV_X1 U9869 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8752) );
  INV_X1 U9870 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n12174) );
  AND2_X1 U9871 ( .A1(n9017), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9412) );
  OR2_X1 U9872 ( .A1(n11065), .A2(n11062), .ZN(n15102) );
  OR2_X1 U9873 ( .A1(n11005), .A2(n9610), .ZN(n11554) );
  AND2_X1 U9874 ( .A1(n9365), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9381) );
  OR2_X1 U9875 ( .A1(n11668), .A2(n11667), .ZN(n11665) );
  INV_X1 U9876 ( .A(n15119), .ZN(n15004) );
  AND2_X1 U9877 ( .A1(n15001), .A2(n11581), .ZN(n11805) );
  INV_X1 U9878 ( .A(n15099), .ZN(n15401) );
  INV_X1 U9879 ( .A(n11068), .ZN(n16495) );
  XNOR2_X1 U9880 ( .A(n8632), .B(SI_17_), .ZN(n8860) );
  XNOR2_X1 U9881 ( .A(n8619), .B(n13699), .ZN(n8850) );
  INV_X1 U9882 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15749) );
  AOI21_X1 U9883 ( .B1(n11643), .B2(n11644), .A(n10128), .ZN(n11661) );
  AND3_X1 U9884 ( .A1(n9829), .A2(n9828), .A3(n9827), .ZN(n12782) );
  INV_X1 U9885 ( .A(n13447), .ZN(n13455) );
  NOR2_X1 U9886 ( .A1(n13337), .A2(n16467), .ZN(n11923) );
  INV_X1 U9887 ( .A(n14108), .ZN(n14132) );
  OAI21_X1 U9888 ( .B1(n13884), .B2(n13883), .A(n13882), .ZN(n13890) );
  INV_X1 U9889 ( .A(n16076), .ZN(n16043) );
  AND2_X1 U9890 ( .A1(n8488), .A2(n8466), .ZN(n16054) );
  INV_X1 U9891 ( .A(n13321), .ZN(n14130) );
  AND2_X1 U9892 ( .A1(n14169), .A2(n12414), .ZN(n14100) );
  AND2_X2 U9893 ( .A1(n11923), .A2(n13289), .ZN(n14163) );
  NOR2_X1 U9894 ( .A1(n13337), .A2(n10236), .ZN(n11920) );
  NAND2_X1 U9895 ( .A1(n10064), .A2(n10238), .ZN(n16475) );
  OR2_X1 U9896 ( .A1(n16475), .A2(n16382), .ZN(n16469) );
  INV_X1 U9897 ( .A(n16413), .ZN(n16382) );
  XNOR2_X1 U9898 ( .A(n8451), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13338) );
  INV_X1 U9899 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8448) );
  OR2_X1 U9900 ( .A1(n8385), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8434) );
  INV_X1 U9901 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8388) );
  INV_X1 U9902 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8401) );
  INV_X1 U9903 ( .A(n14442), .ZN(n14420) );
  AND2_X1 U9904 ( .A1(n10940), .A2(n10939), .ZN(n14445) );
  AND2_X1 U9905 ( .A1(n10502), .A2(n10501), .ZN(n14373) );
  INV_X1 U9906 ( .A(n10506), .ZN(n10499) );
  INV_X1 U9907 ( .A(n15681), .ZN(n15668) );
  NOR2_X1 U9908 ( .A1(n15645), .A2(P2_U3088), .ZN(n15678) );
  NAND2_X1 U9909 ( .A1(n8927), .A2(n8926), .ZN(n14481) );
  XNOR2_X1 U9910 ( .A(n11853), .B(n14470), .ZN(n11856) );
  INV_X1 U9911 ( .A(n16117), .ZN(n16397) );
  INV_X1 U9912 ( .A(n14750), .ZN(n14757) );
  NAND2_X1 U9913 ( .A1(n16513), .A2(n10561), .ZN(n10562) );
  AND2_X1 U9914 ( .A1(n16105), .A2(n10835), .ZN(n16265) );
  INV_X1 U9915 ( .A(n14787), .ZN(n14792) );
  INV_X1 U9916 ( .A(n16430), .ZN(n16509) );
  INV_X1 U9917 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8962) );
  OR2_X1 U9918 ( .A1(n8943), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8950) );
  INV_X1 U9919 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8763) );
  AND4_X1 U9920 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(n9565)
         );
  AND2_X1 U9921 ( .A1(n9357), .A2(n9356), .ZN(n15088) );
  INV_X1 U9922 ( .A(n15227), .ZN(n15720) );
  OR2_X1 U9923 ( .A1(n11059), .A2(n12770), .ZN(n11798) );
  AND2_X1 U9924 ( .A1(n15349), .A2(n15348), .ZN(n15487) );
  INV_X1 U9925 ( .A(n16099), .ZN(n15387) );
  INV_X1 U9926 ( .A(n15412), .ZN(n15393) );
  INV_X1 U9927 ( .A(n16153), .ZN(n15356) );
  NAND2_X1 U9928 ( .A1(n11057), .A2(n15541), .ZN(n11789) );
  INV_X1 U9929 ( .A(n15432), .ZN(n15433) );
  AND2_X1 U9930 ( .A1(n16085), .A2(n16485), .ZN(n16243) );
  INV_X1 U9931 ( .A(n16248), .ZN(n16532) );
  INV_X1 U9932 ( .A(n16243), .ZN(n16536) );
  INV_X1 U9933 ( .A(n11789), .ZN(n11599) );
  NAND2_X1 U9934 ( .A1(n10995), .A2(n10994), .ZN(n11557) );
  AND2_X1 U9935 ( .A1(n8492), .A2(n8491), .ZN(n16073) );
  INV_X1 U9936 ( .A(n10231), .ZN(n10232) );
  INV_X1 U9937 ( .A(n13454), .ZN(n12702) );
  NAND2_X1 U9938 ( .A1(n9991), .A2(n9990), .ZN(n13463) );
  INV_X1 U9939 ( .A(n14160), .ZN(n13465) );
  INV_X1 U9940 ( .A(n16073), .ZN(n15981) );
  INV_X1 U9941 ( .A(n16054), .ZN(n16082) );
  INV_X1 U9942 ( .A(n14100), .ZN(n14171) );
  NAND2_X1 U9943 ( .A1(n16473), .A2(n16410), .ZN(n14227) );
  AND4_X2 U9944 ( .A1(n11921), .A2(n11920), .A3(n10242), .A4(n10241), .ZN(
        n16473) );
  NAND2_X1 U9945 ( .A1(n16447), .A2(n16410), .ZN(n14296) );
  AND2_X1 U9946 ( .A1(n16385), .A2(n16384), .ZN(n16387) );
  AND2_X2 U9947 ( .A1(n10111), .A2(n10208), .ZN(n16447) );
  NAND2_X1 U9948 ( .A1(n11410), .A2(n11024), .ZN(n11025) );
  INV_X1 U9949 ( .A(SI_14_), .ZN(n11032) );
  INV_X1 U9950 ( .A(SI_11_), .ZN(n13698) );
  INV_X1 U9951 ( .A(n14437), .ZN(n14427) );
  INV_X1 U9952 ( .A(n14437), .ZN(n14408) );
  INV_X1 U9953 ( .A(n14373), .ZN(n14450) );
  INV_X1 U9954 ( .A(n14439), .ZN(n14559) );
  OR2_X1 U9955 ( .A1(n10397), .A2(n10396), .ZN(n14461) );
  INV_X1 U9956 ( .A(n15678), .ZN(n15626) );
  OR2_X1 U9957 ( .A1(n11124), .A2(n11123), .ZN(n15686) );
  INV_X1 U9958 ( .A(n14678), .ZN(n14620) );
  NAND2_X1 U9959 ( .A1(n13098), .A2(n14757), .ZN(n10559) );
  INV_X1 U9960 ( .A(n16512), .ZN(n16510) );
  NAND2_X1 U9961 ( .A1(n16516), .A2(n16265), .ZN(n14787) );
  AND4_X1 U9962 ( .A1(n16277), .A2(n16272), .A3(n16267), .A4(n16266), .ZN(
        n16269) );
  OR2_X1 U9963 ( .A1(n15568), .A2(n15566), .ZN(n15567) );
  INV_X1 U9964 ( .A(n15571), .ZN(n15568) );
  XNOR2_X1 U9965 ( .A(n8963), .B(n8962), .ZN(n14813) );
  INV_X1 U9966 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11403) );
  INV_X1 U9967 ( .A(n12071), .ZN(n16351) );
  AND2_X1 U9968 ( .A1(n11499), .A2(n13013), .ZN(n16555) );
  INV_X1 U9969 ( .A(n11802), .ZN(n16204) );
  OR2_X1 U9970 ( .A1(n11065), .A2(n11061), .ZN(n15115) );
  INV_X1 U9971 ( .A(n15056), .ZN(n15121) );
  OR2_X1 U9972 ( .A1(n9288), .A2(n9287), .ZN(n15131) );
  INV_X1 U9973 ( .A(n12640), .ZN(n15135) );
  OR2_X1 U9974 ( .A1(n15699), .A2(n11296), .ZN(n15227) );
  INV_X1 U9975 ( .A(n15696), .ZN(n15728) );
  OR2_X1 U9976 ( .A1(n16153), .A2(n11798), .ZN(n16156) );
  AND2_X1 U9977 ( .A1(n15380), .A2(n15379), .ZN(n15504) );
  OR2_X1 U9978 ( .A1(n16153), .A2(n12276), .ZN(n15412) );
  AND2_X1 U9979 ( .A1(n16394), .A2(n16393), .ZN(n16396) );
  AND2_X1 U9980 ( .A1(n9609), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10996) );
  INV_X1 U9981 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15553) );
  INV_X1 U9982 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11401) );
  AND2_X1 U9983 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10840), .ZN(P2_U3947) );
  NAND2_X1 U9984 ( .A1(n8994), .A2(n8993), .ZN(P2_U3498) );
  INV_X2 U9985 ( .A(n15142), .ZN(P1_U4016) );
  NAND2_X1 U9986 ( .A1(n8374), .A2(n8360), .ZN(n8372) );
  INV_X1 U9987 ( .A(n8372), .ZN(n8350) );
  NAND2_X1 U9988 ( .A1(n8350), .A2(n8359), .ZN(n8443) );
  NAND2_X1 U9989 ( .A1(n10043), .A2(n10045), .ZN(n8452) );
  NOR2_X1 U9990 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n8358) );
  NOR2_X1 U9991 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8357) );
  AND2_X2 U9992 ( .A1(n7447), .A2(n8360), .ZN(n8361) );
  INV_X1 U9993 ( .A(n8455), .ZN(n8366) );
  NAND2_X1 U9994 ( .A1(n8366), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8363) );
  MUX2_X1 U9995 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8365), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8367) );
  NAND2_X1 U9996 ( .A1(n8368), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8369) );
  MUX2_X1 U9997 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8369), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8371) );
  INV_X1 U9998 ( .A(n12537), .ZN(n10087) );
  INV_X1 U9999 ( .A(n8463), .ZN(n10217) );
  NAND2_X1 U10000 ( .A1(n8372), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8373) );
  XNOR2_X1 U10001 ( .A(n8373), .B(P3_IR_REG_17__SCAN_IN), .ZN(n9883) );
  INV_X1 U10002 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8405) );
  OR2_X1 U10003 ( .A1(n8374), .A2(n8405), .ZN(n8375) );
  XNOR2_X1 U10004 ( .A(n8375), .B(P3_IR_REG_16__SCAN_IN), .ZN(n16042) );
  INV_X1 U10005 ( .A(n16042), .ZN(n11136) );
  OR2_X1 U10006 ( .A1(n8425), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10007 ( .A1(n8382), .A2(n8378), .ZN(n8385) );
  OAI21_X1 U10008 ( .B1(n8434), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8379) );
  XNOR2_X1 U10009 ( .A(n8379), .B(P3_IR_REG_15__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U10010 ( .A1(n8385), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8380) );
  MUX2_X1 U10011 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8380), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8381) );
  NAND2_X1 U10012 ( .A1(n8381), .A2(n8434), .ZN(n11019) );
  NOR2_X1 U10013 ( .A1(n8382), .A2(n8405), .ZN(n8383) );
  MUX2_X1 U10014 ( .A(n8405), .B(n8383), .S(P3_IR_REG_12__SCAN_IN), .Z(n8384)
         );
  INV_X1 U10015 ( .A(n8384), .ZN(n8386) );
  NAND2_X1 U10016 ( .A1(n8386), .A2(n8385), .ZN(n12524) );
  NAND2_X1 U10017 ( .A1(n12524), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U10018 ( .A1(n8387), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8389) );
  XNOR2_X1 U10019 ( .A(n8389), .B(n8388), .ZN(n12238) );
  INV_X1 U10020 ( .A(n12238), .ZN(n8550) );
  NAND2_X1 U10021 ( .A1(n8390), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8391) );
  MUX2_X1 U10022 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8391), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8392) );
  NAND2_X1 U10023 ( .A1(n8392), .A2(n8425), .ZN(n16032) );
  INV_X1 U10024 ( .A(n16032), .ZN(n8537) );
  OR2_X1 U10025 ( .A1(n8393), .A2(n8405), .ZN(n8394) );
  XNOR2_X1 U10026 ( .A(n8394), .B(P3_IR_REG_8__SCAN_IN), .ZN(n9778) );
  NOR2_X1 U10027 ( .A1(n8395), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8414) );
  INV_X1 U10028 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10029 ( .A1(n8414), .A2(n8396), .ZN(n8417) );
  OAI21_X1 U10030 ( .B1(n8399), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8398) );
  INV_X1 U10031 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8397) );
  XNOR2_X1 U10032 ( .A(n8398), .B(n8397), .ZN(n15992) );
  NAND2_X1 U10033 ( .A1(n8399), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8400) );
  XNOR2_X1 U10034 ( .A(n8400), .B(P3_IR_REG_6__SCAN_IN), .ZN(n15978) );
  INV_X1 U10035 ( .A(n15978), .ZN(n10973) );
  NAND2_X1 U10036 ( .A1(n8417), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8402) );
  XNOR2_X1 U10037 ( .A(n8402), .B(n8401), .ZN(n15952) );
  NAND2_X1 U10038 ( .A1(n8395), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8404) );
  XNOR2_X1 U10039 ( .A(n8404), .B(n8403), .ZN(n10965) );
  INV_X1 U10040 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n16202) );
  NAND2_X1 U10041 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8408) );
  XNOR2_X1 U10042 ( .A(n8408), .B(P3_IR_REG_1__SCAN_IN), .ZN(n11784) );
  INV_X1 U10043 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10960) );
  NAND2_X1 U10044 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n10960), .ZN(n8409) );
  NAND2_X1 U10045 ( .A1(n11784), .A2(n8409), .ZN(n8410) );
  NAND2_X1 U10046 ( .A1(n8410), .A2(n8411), .ZN(n11778) );
  INV_X1 U10047 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n16137) );
  OR2_X1 U10048 ( .A1(n11778), .A2(n16137), .ZN(n11780) );
  NAND2_X1 U10049 ( .A1(n11780), .A2(n8411), .ZN(n12002) );
  NAND2_X1 U10050 ( .A1(n12003), .A2(n12002), .ZN(n12001) );
  NAND2_X1 U10051 ( .A1(n7370), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8412) );
  INV_X1 U10052 ( .A(n10965), .ZN(n15917) );
  INV_X1 U10053 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n8511) );
  INV_X1 U10054 ( .A(n8414), .ZN(n8415) );
  NAND2_X1 U10055 ( .A1(n8415), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8416) );
  MUX2_X1 U10056 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8416), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8418) );
  NAND2_X1 U10057 ( .A1(n8418), .A2(n8417), .ZN(n15932) );
  MUX2_X1 U10058 ( .A(n8511), .B(P3_REG2_REG_4__SCAN_IN), .S(n15932), .Z(
        n15924) );
  NOR2_X1 U10059 ( .A1(n7735), .A2(n8419), .ZN(n8420) );
  INV_X1 U10060 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15945) );
  INV_X1 U10061 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n8522) );
  MUX2_X1 U10062 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n8522), .S(n15978), .Z(
        n15966) );
  NOR2_X1 U10063 ( .A1(n7737), .A2(n8421), .ZN(n8422) );
  INV_X1 U10064 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15985) );
  INV_X1 U10065 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U10066 ( .A1(n9778), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n12418), .B2(
        n16011), .ZN(n16003) );
  NOR2_X1 U10067 ( .A1(n8537), .A2(n8423), .ZN(n8424) );
  INV_X1 U10068 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n16024) );
  NAND2_X1 U10069 ( .A1(n8425), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8427) );
  INV_X1 U10070 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8426) );
  XNOR2_X1 U10071 ( .A(n8427), .B(n8426), .ZN(n12547) );
  NAND2_X1 U10072 ( .A1(n12547), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8429) );
  OR2_X1 U10073 ( .A1(n12547), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10074 ( .A1(n8429), .A2(n8428), .ZN(n12542) );
  NOR2_X1 U10075 ( .A1(n8550), .A2(n8430), .ZN(n8431) );
  INV_X1 U10076 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12991) );
  NOR2_X1 U10077 ( .A1(n12991), .A2(n12230), .ZN(n12229) );
  OR2_X1 U10078 ( .A1(n12524), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U10079 ( .A1(n8555), .A2(n8432), .ZN(n12518) );
  INV_X1 U10080 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12802) );
  NAND2_X1 U10081 ( .A1(n8434), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8436) );
  INV_X1 U10082 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8435) );
  XNOR2_X1 U10083 ( .A(n8436), .B(n8435), .ZN(n11031) );
  NAND2_X1 U10084 ( .A1(n11031), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8438) );
  OR2_X1 U10085 ( .A1(n11031), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10086 ( .A1(n8438), .A2(n8437), .ZN(n13898) );
  NOR2_X1 U10087 ( .A1(n11075), .A2(n8439), .ZN(n8440) );
  INV_X1 U10088 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13919) );
  INV_X1 U10089 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n8441) );
  AOI22_X1 U10090 ( .A1(n16042), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n8441), 
        .B2(n11136), .ZN(n16055) );
  AOI21_X1 U10091 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n11136), .A(n16056), 
        .ZN(n8442) );
  XNOR2_X1 U10092 ( .A(n9883), .B(n8442), .ZN(n16063) );
  INV_X1 U10093 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n16064) );
  OR2_X1 U10094 ( .A1(n8442), .A2(n9883), .ZN(n13935) );
  NAND2_X1 U10095 ( .A1(n8443), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8444) );
  XNOR2_X1 U10096 ( .A(n8444), .B(P3_IR_REG_18__SCAN_IN), .ZN(n9896) );
  INV_X1 U10097 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8571) );
  OR2_X1 U10098 ( .A1(n9896), .A2(n8571), .ZN(n8446) );
  NAND2_X1 U10099 ( .A1(n9896), .A2(n8571), .ZN(n8445) );
  NAND2_X1 U10100 ( .A1(n8446), .A2(n8445), .ZN(n13934) );
  INV_X1 U10101 ( .A(n8446), .ZN(n8447) );
  NAND2_X1 U10102 ( .A1(n8351), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8449) );
  XNOR2_X1 U10103 ( .A(n11452), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10104 ( .A1(n8450), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10105 ( .A1(n8452), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10106 ( .A1(n13207), .A2(n8464), .ZN(n8462) );
  NAND2_X1 U10107 ( .A1(n8457), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10108 ( .A1(n8459), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8461) );
  AND2_X1 U10109 ( .A1(n8462), .A2(n10054), .ZN(n8490) );
  INV_X1 U10110 ( .A(n8464), .ZN(n8465) );
  NAND2_X1 U10111 ( .A1(n8465), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13341) );
  NAND2_X1 U10112 ( .A1(n13337), .A2(n13341), .ZN(n8491) );
  INV_X1 U10113 ( .A(n13335), .ZN(n10056) );
  NAND2_X1 U10114 ( .A1(n10056), .A2(n13334), .ZN(n10055) );
  INV_X1 U10115 ( .A(n10055), .ZN(n8466) );
  INV_X1 U10116 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n14217) );
  INV_X1 U10117 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n14225) );
  AOI22_X1 U10118 ( .A1(n16042), .A2(n14225), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n11136), .ZN(n16046) );
  INV_X1 U10119 ( .A(n11075), .ZN(n13929) );
  NAND2_X1 U10120 ( .A1(n12524), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8554) );
  OR2_X1 U10121 ( .A1(n12524), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8467) );
  AND2_X1 U10122 ( .A1(n8554), .A2(n8467), .ZN(n12521) );
  NAND2_X1 U10123 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n12547), .ZN(n8478) );
  INV_X1 U10124 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8542) );
  MUX2_X1 U10125 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n8542), .S(n12547), .Z(
        n12539) );
  INV_X1 U10126 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n16371) );
  AOI22_X1 U10127 ( .A1(n9778), .A2(n16371), .B1(P3_REG1_REG_8__SCAN_IN), .B2(
        n16011), .ZN(n16016) );
  INV_X1 U10128 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n16334) );
  INV_X1 U10129 ( .A(n15932), .ZN(n8512) );
  INV_X1 U10130 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n16282) );
  INV_X1 U10131 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U10132 ( .A1(n11777), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10133 ( .A1(n8468), .A2(n7885), .ZN(n12005) );
  NAND2_X1 U10134 ( .A1(n7370), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8469) );
  XNOR2_X1 U10135 ( .A(n8470), .B(n15917), .ZN(n15918) );
  AND2_X1 U10136 ( .A1(n8470), .A2(n10965), .ZN(n8471) );
  AOI21_X1 U10137 ( .B1(n15918), .B2(P3_REG1_REG_3__SCAN_IN), .A(n8471), .ZN(
        n15938) );
  MUX2_X1 U10138 ( .A(n16282), .B(P3_REG1_REG_4__SCAN_IN), .S(n15932), .Z(
        n15937) );
  NAND2_X1 U10139 ( .A1(n15952), .A2(n8472), .ZN(n8473) );
  NAND2_X1 U10140 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15957), .ZN(n15956) );
  AND2_X1 U10141 ( .A1(n8473), .A2(n15956), .ZN(n15964) );
  MUX2_X1 U10142 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n16334), .S(n15978), .Z(
        n15963) );
  NAND2_X1 U10143 ( .A1(n15992), .A2(n8474), .ZN(n8475) );
  NAND2_X1 U10144 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15997), .ZN(n15996) );
  NAND2_X1 U10145 ( .A1(n8475), .A2(n15996), .ZN(n16017) );
  NAND2_X1 U10146 ( .A1(n16016), .A2(n16017), .ZN(n16015) );
  OAI21_X1 U10147 ( .B1(n9778), .B2(n16371), .A(n16015), .ZN(n8476) );
  NAND2_X1 U10148 ( .A1(n16032), .A2(n8476), .ZN(n8477) );
  XNOR2_X1 U10149 ( .A(n8476), .B(n8537), .ZN(n16037) );
  NAND2_X1 U10150 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n16037), .ZN(n16036) );
  NAND2_X1 U10151 ( .A1(n12238), .A2(n8479), .ZN(n8480) );
  NAND2_X1 U10152 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n12234), .ZN(n12233) );
  NAND2_X1 U10153 ( .A1(n8480), .A2(n12233), .ZN(n12522) );
  NAND2_X1 U10154 ( .A1(n12521), .A2(n12522), .ZN(n12520) );
  NAND2_X1 U10155 ( .A1(n11019), .A2(n8481), .ZN(n8482) );
  INV_X1 U10156 ( .A(n11031), .ZN(n13909) );
  XNOR2_X1 U10157 ( .A(n13909), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U10158 ( .A1(n13901), .A2(n13900), .B1(P3_REG1_REG_14__SCAN_IN), 
        .B2(n11031), .ZN(n8483) );
  NAND2_X1 U10159 ( .A1(n13929), .A2(n8484), .ZN(n8485) );
  NAND2_X1 U10160 ( .A1(n16046), .A2(n16045), .ZN(n16044) );
  OAI21_X1 U10161 ( .B1(n16042), .B2(n14225), .A(n16044), .ZN(n8486) );
  INV_X1 U10162 ( .A(n9883), .ZN(n16075) );
  NAND2_X1 U10163 ( .A1(n8486), .A2(n16075), .ZN(n13946) );
  XNOR2_X1 U10164 ( .A(n8486), .B(n9883), .ZN(n16066) );
  NAND2_X1 U10165 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n16066), .ZN(n16065) );
  NAND2_X1 U10166 ( .A1(n13946), .A2(n16065), .ZN(n8487) );
  XNOR2_X1 U10167 ( .A(n9896), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n13944) );
  NAND2_X1 U10168 ( .A1(n8487), .A2(n13944), .ZN(n13948) );
  INV_X1 U10169 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n14213) );
  XNOR2_X1 U10170 ( .A(n11452), .B(n14213), .ZN(n8573) );
  INV_X1 U10171 ( .A(n8488), .ZN(n8489) );
  MUX2_X1 U10172 ( .A(n8489), .B(n13471), .S(n10056), .Z(n16076) );
  INV_X1 U10173 ( .A(n8490), .ZN(n8492) );
  AND2_X1 U10174 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13373) );
  AOI21_X1 U10175 ( .B1(n16073), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n13373), 
        .ZN(n8493) );
  OAI21_X1 U10176 ( .B1(n16076), .B2(n11452), .A(n8493), .ZN(n8494) );
  INV_X1 U10177 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8495) );
  MUX2_X1 U10178 ( .A(n16137), .B(n8495), .S(n8565), .Z(n8496) );
  NAND2_X1 U10179 ( .A1(n8496), .A2(n11784), .ZN(n12013) );
  INV_X1 U10180 ( .A(n8496), .ZN(n8497) );
  NAND2_X1 U10181 ( .A1(n8497), .A2(n7889), .ZN(n8498) );
  NAND2_X1 U10182 ( .A1(n12013), .A2(n8498), .ZN(n11776) );
  MUX2_X1 U10183 ( .A(n7881), .B(n7886), .S(n8565), .Z(n15899) );
  NAND2_X1 U10184 ( .A1(n15899), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15898) );
  OR2_X1 U10185 ( .A1(n11776), .A2(n15898), .ZN(n11775) );
  NAND2_X1 U10186 ( .A1(n11775), .A2(n12013), .ZN(n8504) );
  MUX2_X1 U10187 ( .A(n16202), .B(n8499), .S(n8565), .Z(n8501) );
  INV_X1 U10188 ( .A(n7370), .ZN(n8500) );
  NAND2_X1 U10189 ( .A1(n8501), .A2(n8500), .ZN(n15912) );
  INV_X1 U10190 ( .A(n8501), .ZN(n8502) );
  NAND2_X1 U10191 ( .A1(n8502), .A2(n7370), .ZN(n8503) );
  AND2_X1 U10192 ( .A1(n15912), .A2(n8503), .ZN(n12014) );
  NAND2_X1 U10193 ( .A1(n8504), .A2(n12014), .ZN(n15913) );
  NAND2_X1 U10194 ( .A1(n15913), .A2(n15912), .ZN(n8510) );
  INV_X1 U10195 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n8506) );
  INV_X1 U10196 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n8505) );
  MUX2_X1 U10197 ( .A(n8506), .B(n8505), .S(n8565), .Z(n8507) );
  NAND2_X1 U10198 ( .A1(n8507), .A2(n15917), .ZN(n15926) );
  INV_X1 U10199 ( .A(n8507), .ZN(n8508) );
  NAND2_X1 U10200 ( .A1(n8508), .A2(n10965), .ZN(n8509) );
  AND2_X1 U10201 ( .A1(n15926), .A2(n8509), .ZN(n15910) );
  NAND2_X1 U10202 ( .A1(n8510), .A2(n15910), .ZN(n15930) );
  NAND2_X1 U10203 ( .A1(n15930), .A2(n15926), .ZN(n8516) );
  MUX2_X1 U10204 ( .A(n8511), .B(n16282), .S(n8565), .Z(n8513) );
  NAND2_X1 U10205 ( .A1(n8513), .A2(n8512), .ZN(n15946) );
  INV_X1 U10206 ( .A(n8513), .ZN(n8514) );
  NAND2_X1 U10207 ( .A1(n8514), .A2(n15932), .ZN(n8515) );
  AND2_X1 U10208 ( .A1(n15946), .A2(n8515), .ZN(n15928) );
  NAND2_X1 U10209 ( .A1(n8516), .A2(n15928), .ZN(n15950) );
  NAND2_X1 U10210 ( .A1(n15950), .A2(n15946), .ZN(n8521) );
  INV_X1 U10211 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n8517) );
  MUX2_X1 U10212 ( .A(n15945), .B(n8517), .S(n8565), .Z(n8518) );
  NAND2_X1 U10213 ( .A1(n8518), .A2(n7735), .ZN(n15973) );
  INV_X1 U10214 ( .A(n8518), .ZN(n8519) );
  NAND2_X1 U10215 ( .A1(n8519), .A2(n15952), .ZN(n8520) );
  AND2_X1 U10216 ( .A1(n15973), .A2(n8520), .ZN(n15948) );
  NAND2_X1 U10217 ( .A1(n8521), .A2(n15948), .ZN(n15974) );
  NAND2_X1 U10218 ( .A1(n15974), .A2(n15973), .ZN(n8526) );
  MUX2_X1 U10219 ( .A(n8522), .B(n16334), .S(n8565), .Z(n8523) );
  NAND2_X1 U10220 ( .A1(n8523), .A2(n15978), .ZN(n15986) );
  INV_X1 U10221 ( .A(n8523), .ZN(n8524) );
  NAND2_X1 U10222 ( .A1(n8524), .A2(n10973), .ZN(n8525) );
  AND2_X1 U10223 ( .A1(n15986), .A2(n8525), .ZN(n15971) );
  NAND2_X1 U10224 ( .A1(n8526), .A2(n15971), .ZN(n15990) );
  NAND2_X1 U10225 ( .A1(n15990), .A2(n15986), .ZN(n8531) );
  INV_X1 U10226 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8527) );
  MUX2_X1 U10227 ( .A(n15985), .B(n8527), .S(n8565), .Z(n8528) );
  NAND2_X1 U10228 ( .A1(n8528), .A2(n7737), .ZN(n16005) );
  INV_X1 U10229 ( .A(n8528), .ZN(n8529) );
  NAND2_X1 U10230 ( .A1(n8529), .A2(n15992), .ZN(n8530) );
  AND2_X1 U10231 ( .A1(n16005), .A2(n8530), .ZN(n15988) );
  NAND2_X1 U10232 ( .A1(n8531), .A2(n15988), .ZN(n16009) );
  NAND2_X1 U10233 ( .A1(n16009), .A2(n16005), .ZN(n8535) );
  MUX2_X1 U10234 ( .A(n12418), .B(n16371), .S(n8565), .Z(n8532) );
  NAND2_X1 U10235 ( .A1(n8532), .A2(n9778), .ZN(n16025) );
  INV_X1 U10236 ( .A(n8532), .ZN(n8533) );
  NAND2_X1 U10237 ( .A1(n8533), .A2(n16011), .ZN(n8534) );
  AND2_X1 U10238 ( .A1(n16025), .A2(n8534), .ZN(n16007) );
  NAND2_X1 U10239 ( .A1(n8535), .A2(n16007), .ZN(n16030) );
  NAND2_X1 U10240 ( .A1(n16030), .A2(n16025), .ZN(n8541) );
  INV_X1 U10241 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n8536) );
  MUX2_X1 U10242 ( .A(n16024), .B(n8536), .S(n8565), .Z(n8538) );
  NAND2_X1 U10243 ( .A1(n8538), .A2(n8537), .ZN(n12550) );
  INV_X1 U10244 ( .A(n8538), .ZN(n8539) );
  NAND2_X1 U10245 ( .A1(n8539), .A2(n16032), .ZN(n8540) );
  AND2_X1 U10246 ( .A1(n12550), .A2(n8540), .ZN(n16027) );
  NAND2_X1 U10247 ( .A1(n8541), .A2(n16027), .ZN(n16028) );
  NAND2_X1 U10248 ( .A1(n16028), .A2(n12550), .ZN(n8547) );
  INV_X1 U10249 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12765) );
  MUX2_X1 U10250 ( .A(n12765), .B(n8542), .S(n12984), .Z(n8544) );
  INV_X1 U10251 ( .A(n12547), .ZN(n8543) );
  NAND2_X1 U10252 ( .A1(n8544), .A2(n8543), .ZN(n8548) );
  INV_X1 U10253 ( .A(n8544), .ZN(n8545) );
  NAND2_X1 U10254 ( .A1(n8545), .A2(n12547), .ZN(n8546) );
  AND2_X1 U10255 ( .A1(n8548), .A2(n8546), .ZN(n12548) );
  NAND2_X1 U10256 ( .A1(n8547), .A2(n12548), .ZN(n12552) );
  NAND2_X1 U10257 ( .A1(n12552), .A2(n8548), .ZN(n12232) );
  MUX2_X1 U10258 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12984), .Z(n8549) );
  XNOR2_X1 U10259 ( .A(n8549), .B(n8550), .ZN(n12231) );
  NAND2_X1 U10260 ( .A1(n12232), .A2(n12231), .ZN(n12528) );
  INV_X1 U10261 ( .A(n8549), .ZN(n8551) );
  NAND2_X1 U10262 ( .A1(n8551), .A2(n8550), .ZN(n12527) );
  INV_X1 U10263 ( .A(n12518), .ZN(n8552) );
  MUX2_X1 U10264 ( .A(n8552), .B(n12521), .S(n12984), .Z(n12530) );
  AND2_X1 U10265 ( .A1(n12527), .A2(n12530), .ZN(n8553) );
  NAND2_X1 U10266 ( .A1(n12528), .A2(n8553), .ZN(n12529) );
  MUX2_X1 U10267 ( .A(n8555), .B(n8554), .S(n8565), .Z(n8556) );
  NAND2_X1 U10268 ( .A1(n12529), .A2(n8556), .ZN(n12806) );
  MUX2_X1 U10269 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12984), .Z(n8557) );
  XNOR2_X1 U10270 ( .A(n8557), .B(n11019), .ZN(n12807) );
  MUX2_X1 U10271 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n12984), .Z(n8560) );
  XNOR2_X1 U10272 ( .A(n8560), .B(n13909), .ZN(n13903) );
  INV_X1 U10273 ( .A(n8557), .ZN(n8558) );
  NAND2_X1 U10274 ( .A1(n8558), .A2(n7734), .ZN(n13904) );
  AND2_X1 U10275 ( .A1(n13903), .A2(n13904), .ZN(n8559) );
  NAND2_X1 U10276 ( .A1(n13905), .A2(n8559), .ZN(n13902) );
  NAND2_X1 U10277 ( .A1(n8560), .A2(n11031), .ZN(n8561) );
  NAND2_X1 U10278 ( .A1(n13902), .A2(n8561), .ZN(n8563) );
  XNOR2_X1 U10279 ( .A(n8563), .B(n11075), .ZN(n13922) );
  INV_X1 U10280 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n8562) );
  MUX2_X1 U10281 ( .A(n13919), .B(n8562), .S(n8565), .Z(n13921) );
  NAND2_X1 U10282 ( .A1(n13922), .A2(n13921), .ZN(n13920) );
  OR2_X1 U10283 ( .A1(n8563), .A2(n13929), .ZN(n8564) );
  NAND2_X1 U10284 ( .A1(n13920), .A2(n8564), .ZN(n16049) );
  MUX2_X1 U10285 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n8565), .Z(n8566) );
  NAND2_X1 U10286 ( .A1(n8566), .A2(n11136), .ZN(n16047) );
  NAND2_X1 U10287 ( .A1(n16049), .A2(n16047), .ZN(n8568) );
  INV_X1 U10288 ( .A(n8566), .ZN(n8567) );
  NAND2_X1 U10289 ( .A1(n8567), .A2(n16042), .ZN(n16048) );
  NAND2_X1 U10290 ( .A1(n8568), .A2(n16048), .ZN(n16070) );
  MUX2_X1 U10291 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12984), .Z(n8569) );
  XNOR2_X1 U10292 ( .A(n8569), .B(n16075), .ZN(n16071) );
  NAND2_X1 U10293 ( .A1(n8569), .A2(n16075), .ZN(n8570) );
  NAND2_X1 U10294 ( .A1(n16067), .A2(n8570), .ZN(n8572) );
  INV_X1 U10295 ( .A(n9896), .ZN(n13943) );
  XNOR2_X1 U10296 ( .A(n8572), .B(n9896), .ZN(n13940) );
  MUX2_X1 U10297 ( .A(n8571), .B(n14217), .S(n12984), .Z(n13939) );
  NAND2_X1 U10298 ( .A1(n13940), .A2(n13939), .ZN(n13938) );
  OAI21_X1 U10299 ( .B1(n8572), .B2(n13943), .A(n13938), .ZN(n8577) );
  INV_X1 U10300 ( .A(n8573), .ZN(n8574) );
  MUX2_X1 U10301 ( .A(n8575), .B(n8574), .S(n12984), .Z(n8576) );
  NAND2_X1 U10302 ( .A1(P3_U3897), .A2(n13335), .ZN(n16069) );
  NAND2_X1 U10303 ( .A1(n7427), .A2(n16052), .ZN(n8578) );
  INV_X1 U10304 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8579) );
  NAND3_X1 U10305 ( .A1(n8580), .A2(n8579), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n8582) );
  INV_X1 U10306 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8583) );
  NAND3_X1 U10307 ( .A1(n15886), .A2(n8583), .A3(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8584) );
  INV_X1 U10308 ( .A(n8815), .ZN(n8587) );
  INV_X1 U10309 ( .A(SI_0_), .ZN(n13718) );
  NOR2_X1 U10310 ( .A1(n8586), .A2(n13718), .ZN(n8816) );
  NAND2_X1 U10311 ( .A1(n8587), .A2(n8816), .ZN(n8814) );
  INV_X1 U10312 ( .A(n8590), .ZN(n8589) );
  INV_X1 U10313 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10980) );
  NAND2_X1 U10314 ( .A1(n8807), .A2(n8593), .ZN(n8796) );
  NAND2_X1 U10315 ( .A1(n8594), .A2(SI_3_), .ZN(n8596) );
  OAI21_X1 U10316 ( .B1(SI_3_), .B2(n8594), .A(n8596), .ZN(n8595) );
  INV_X1 U10317 ( .A(n8595), .ZN(n8798) );
  NAND2_X1 U10318 ( .A1(n8796), .A2(n8798), .ZN(n8797) );
  MUX2_X1 U10319 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10984), .Z(n8598) );
  NAND2_X1 U10320 ( .A1(n8598), .A2(SI_5_), .ZN(n8599) );
  OAI21_X1 U10321 ( .B1(SI_5_), .B2(n8598), .A(n8599), .ZN(n8777) );
  MUX2_X1 U10322 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10984), .Z(n8600) );
  NAND2_X1 U10323 ( .A1(n8600), .A2(SI_6_), .ZN(n8602) );
  OAI21_X1 U10324 ( .B1(n8600), .B2(SI_6_), .A(n8602), .ZN(n8601) );
  INV_X1 U10325 ( .A(n8601), .ZN(n8768) );
  NAND2_X1 U10326 ( .A1(n8769), .A2(n8768), .ZN(n8771) );
  MUX2_X1 U10327 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10984), .Z(n8603) );
  NAND2_X1 U10328 ( .A1(n8603), .A2(SI_7_), .ZN(n8605) );
  OAI21_X1 U10329 ( .B1(SI_7_), .B2(n8603), .A(n8605), .ZN(n8604) );
  INV_X1 U10330 ( .A(n8604), .ZN(n8758) );
  MUX2_X1 U10331 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10983), .Z(n8606) );
  XNOR2_X1 U10332 ( .A(n8606), .B(SI_8_), .ZN(n8828) );
  INV_X1 U10333 ( .A(n8606), .ZN(n8607) );
  NAND2_X1 U10334 ( .A1(n8607), .A2(n13705), .ZN(n8610) );
  MUX2_X1 U10335 ( .A(n11132), .B(n11134), .S(n10984), .Z(n8608) );
  MUX2_X1 U10336 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10984), .Z(n8609) );
  MUX2_X1 U10337 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10984), .Z(n8614) );
  OAI21_X1 U10338 ( .B1(n8614), .B2(SI_10_), .A(n8615), .ZN(n8834) );
  MUX2_X1 U10339 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10984), .Z(n8616) );
  XNOR2_X1 U10340 ( .A(n8616), .B(SI_11_), .ZN(n8841) );
  INV_X1 U10341 ( .A(n8616), .ZN(n8617) );
  NAND2_X1 U10342 ( .A1(n8617), .A2(n13698), .ZN(n8618) );
  MUX2_X1 U10343 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n10983), .Z(n8619) );
  MUX2_X1 U10344 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10984), .Z(n8620) );
  NAND2_X1 U10345 ( .A1(n8620), .A2(SI_13_), .ZN(n8622) );
  OAI21_X1 U10346 ( .B1(SI_13_), .B2(n8620), .A(n8622), .ZN(n8740) );
  INV_X1 U10347 ( .A(n8740), .ZN(n8621) );
  NAND2_X1 U10348 ( .A1(n8739), .A2(n8621), .ZN(n8743) );
  NAND2_X1 U10349 ( .A1(n8743), .A2(n8622), .ZN(n8733) );
  MUX2_X1 U10350 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10984), .Z(n8623) );
  XNOR2_X1 U10351 ( .A(n8623), .B(SI_14_), .ZN(n8732) );
  INV_X1 U10352 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U10353 ( .A1(n8624), .A2(n11032), .ZN(n8625) );
  MUX2_X1 U10354 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10984), .Z(n8626) );
  XNOR2_X1 U10355 ( .A(n8626), .B(n13692), .ZN(n8725) );
  INV_X1 U10356 ( .A(n8626), .ZN(n8627) );
  NAND2_X1 U10357 ( .A1(n8627), .A2(n13692), .ZN(n8628) );
  MUX2_X1 U10358 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n10984), .Z(n8629) );
  OAI21_X1 U10359 ( .B1(n8629), .B2(SI_16_), .A(n8630), .ZN(n8713) );
  MUX2_X1 U10360 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10983), .Z(n8632) );
  MUX2_X1 U10361 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10984), .Z(n8706) );
  MUX2_X1 U10362 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10984), .Z(n8636) );
  XNOR2_X1 U10363 ( .A(n8636), .B(SI_19_), .ZN(n8698) );
  INV_X1 U10364 ( .A(n8636), .ZN(n8637) );
  INV_X1 U10365 ( .A(SI_19_), .ZN(n11451) );
  NAND2_X1 U10366 ( .A1(n8637), .A2(n11451), .ZN(n8638) );
  MUX2_X1 U10367 ( .A(n12771), .B(n12740), .S(n10984), .Z(n8692) );
  INV_X1 U10368 ( .A(n8692), .ZN(n8639) );
  MUX2_X1 U10369 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10984), .Z(n8642) );
  XNOR2_X1 U10370 ( .A(n8642), .B(SI_21_), .ZN(n8689) );
  INV_X1 U10371 ( .A(n8689), .ZN(n8641) );
  NAND2_X1 U10372 ( .A1(n8642), .A2(SI_21_), .ZN(n8643) );
  NAND2_X1 U10373 ( .A1(n7647), .A2(SI_22_), .ZN(n8645) );
  MUX2_X1 U10374 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10984), .Z(n8868) );
  MUX2_X1 U10375 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10983), .Z(n8647) );
  XNOR2_X1 U10376 ( .A(n8647), .B(n12149), .ZN(n8684) );
  INV_X1 U10377 ( .A(n8684), .ZN(n8648) );
  INV_X1 U10378 ( .A(n8681), .ZN(n8649) );
  MUX2_X1 U10379 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10984), .Z(n8875) );
  NAND2_X1 U10380 ( .A1(n8649), .A2(n8875), .ZN(n8651) );
  NAND2_X1 U10381 ( .A1(n8882), .A2(SI_24_), .ZN(n8650) );
  NAND2_X1 U10382 ( .A1(n8651), .A2(n8650), .ZN(n8655) );
  MUX2_X1 U10383 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10984), .Z(n8652) );
  NAND2_X1 U10384 ( .A1(n8652), .A2(SI_25_), .ZN(n8878) );
  INV_X1 U10385 ( .A(n8652), .ZN(n8653) );
  NAND2_X1 U10386 ( .A1(n8653), .A2(n13680), .ZN(n8876) );
  NAND2_X1 U10387 ( .A1(n8878), .A2(n8876), .ZN(n8654) );
  NAND4_X1 U10388 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8752), .ZN(n8716)
         );
  INV_X1 U10389 ( .A(n8716), .ZN(n8666) );
  NAND3_X1 U10390 ( .A1(n8772), .A2(n8836), .A3(n8843), .ZN(n8718) );
  INV_X1 U10391 ( .A(n8718), .ZN(n8664) );
  NOR2_X1 U10392 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n8663) );
  NOR2_X1 U10393 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n8662) );
  NAND4_X1 U10394 ( .A1(n8666), .A2(n8665), .A3(n8664), .A4(n8719), .ZN(n8699)
         );
  NOR2_X1 U10395 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8667) );
  NAND4_X1 U10396 ( .A1(n8944), .A2(n8667), .A3(n8965), .A4(n8967), .ZN(n8669)
         );
  NAND4_X1 U10397 ( .A1(n8942), .A2(n8939), .A3(n8945), .A4(n8962), .ZN(n8668)
         );
  INV_X1 U10398 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U10399 ( .A1(n8674), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8675) );
  XNOR2_X2 U10400 ( .A(n8678), .B(n8671), .ZN(n14808) );
  NAND2_X2 U10401 ( .A1(n8827), .A2(n10984), .ZN(n8923) );
  INV_X2 U10402 ( .A(n8923), .ZN(n8862) );
  NAND2_X1 U10403 ( .A1(n14814), .A2(n8933), .ZN(n8680) );
  NAND2_X1 U10404 ( .A1(n8934), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U10405 ( .A1(n14817), .A2(n8933), .ZN(n8683) );
  NAND2_X1 U10406 ( .A1(n8934), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8682) );
  XNOR2_X1 U10407 ( .A(n8685), .B(n8684), .ZN(n13009) );
  NAND2_X1 U10408 ( .A1(n13009), .A2(n8933), .ZN(n8687) );
  NAND2_X1 U10409 ( .A1(n8934), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U10410 ( .A1(n12874), .A2(n8933), .ZN(n8691) );
  NAND2_X1 U10411 ( .A1(n8934), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8690) );
  XNOR2_X1 U10412 ( .A(n8692), .B(SI_20_), .ZN(n8693) );
  XNOR2_X1 U10413 ( .A(n8694), .B(n8693), .ZN(n12738) );
  NAND2_X1 U10414 ( .A1(n12738), .A2(n8933), .ZN(n8696) );
  NAND2_X1 U10415 ( .A1(n8934), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8695) );
  INV_X1 U10416 ( .A(n14739), .ZN(n14782) );
  NAND2_X1 U10417 ( .A1(n12557), .A2(n8933), .ZN(n8705) );
  NAND2_X1 U10418 ( .A1(n8863), .A2(n8945), .ZN(n8700) );
  NAND2_X1 U10419 ( .A1(n8709), .A2(n8938), .ZN(n8701) );
  OAI22_X1 U10420 ( .A1(n8864), .A2(n12558), .B1(n10830), .B2(n12843), .ZN(
        n8703) );
  INV_X1 U10421 ( .A(n8703), .ZN(n8704) );
  INV_X1 U10422 ( .A(n8706), .ZN(n8707) );
  XNOR2_X1 U10423 ( .A(n8709), .B(n8938), .ZN(n12841) );
  OAI22_X1 U10424 ( .A1(n8864), .A2(n12338), .B1(n10830), .B2(n12841), .ZN(
        n8710) );
  INV_X1 U10425 ( .A(n8710), .ZN(n8711) );
  INV_X1 U10426 ( .A(n8713), .ZN(n8714) );
  XNOR2_X1 U10427 ( .A(n8715), .B(n8714), .ZN(n12022) );
  NAND2_X1 U10428 ( .A1(n12022), .A2(n8862), .ZN(n8724) );
  INV_X1 U10429 ( .A(n8821), .ZN(n8808) );
  INV_X2 U10430 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8809) );
  AND2_X1 U10431 ( .A1(n8808), .A2(n8809), .ZN(n8799) );
  NOR2_X1 U10432 ( .A1(n8717), .A2(n8718), .ZN(n8727) );
  NAND3_X1 U10433 ( .A1(n8801), .A2(n8719), .A3(n8727), .ZN(n8720) );
  NAND2_X1 U10434 ( .A1(n8720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8721) );
  XNOR2_X1 U10435 ( .A(n8721), .B(P2_IR_REG_16__SCAN_IN), .ZN(n12829) );
  INV_X1 U10436 ( .A(n12829), .ZN(n15644) );
  OAI22_X1 U10437 ( .A1(n8864), .A2(n12024), .B1(n10830), .B2(n15644), .ZN(
        n8722) );
  INV_X1 U10438 ( .A(n8722), .ZN(n8723) );
  INV_X1 U10439 ( .A(n12795), .ZN(n12886) );
  XNOR2_X1 U10440 ( .A(n8726), .B(n8725), .ZN(n11863) );
  NAND2_X1 U10441 ( .A1(n11863), .A2(n8862), .ZN(n8731) );
  NAND2_X1 U10442 ( .A1(n8801), .A2(n8727), .ZN(n8853) );
  NOR2_X1 U10443 ( .A1(n8853), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8852) );
  INV_X1 U10444 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U10445 ( .A1(n8852), .A2(n8728), .ZN(n8745) );
  OAI21_X1 U10446 ( .B1(n8745), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8729) );
  XNOR2_X1 U10447 ( .A(n8729), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15637) );
  INV_X1 U10448 ( .A(n8827), .ZN(n8847) );
  AOI22_X1 U10449 ( .A1(n8934), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n15637), 
        .B2(n8847), .ZN(n8730) );
  XNOR2_X1 U10450 ( .A(n8733), .B(n8732), .ZN(n11515) );
  NAND2_X1 U10451 ( .A1(n11515), .A2(n8862), .ZN(n8738) );
  INV_X1 U10452 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11605) );
  NAND2_X1 U10453 ( .A1(n8745), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8735) );
  INV_X1 U10454 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8734) );
  XNOR2_X1 U10455 ( .A(n8735), .B(n8734), .ZN(n15625) );
  OAI22_X1 U10456 ( .A1(n8864), .A2(n11605), .B1(n10830), .B2(n15625), .ZN(
        n8736) );
  INV_X1 U10457 ( .A(n8736), .ZN(n8737) );
  INV_X1 U10458 ( .A(n8739), .ZN(n8741) );
  NAND2_X1 U10459 ( .A1(n8741), .A2(n8740), .ZN(n8742) );
  NAND2_X1 U10460 ( .A1(n8743), .A2(n8742), .ZN(n11400) );
  OR2_X1 U10461 ( .A1(n8852), .A2(n14795), .ZN(n8744) );
  MUX2_X1 U10462 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8744), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8746) );
  AND2_X1 U10463 ( .A1(n8746), .A2(n8745), .ZN(n11950) );
  AOI22_X1 U10464 ( .A1(n8934), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8847), 
        .B2(n11950), .ZN(n8747) );
  INV_X1 U10465 ( .A(n12504), .ZN(n16505) );
  NAND2_X1 U10466 ( .A1(n8750), .A2(n8749), .ZN(n8751) );
  XNOR2_X1 U10467 ( .A(n8751), .B(SI_9_), .ZN(n11131) );
  NAND2_X1 U10468 ( .A1(n11131), .A2(n8933), .ZN(n8757) );
  NAND2_X1 U10469 ( .A1(n8801), .A2(n8752), .ZN(n8791) );
  INV_X1 U10470 ( .A(n8782), .ZN(n8753) );
  NAND2_X1 U10471 ( .A1(n8753), .A2(n8772), .ZN(n8762) );
  INV_X1 U10472 ( .A(n8762), .ZN(n8754) );
  NAND2_X1 U10473 ( .A1(n8754), .A2(n8763), .ZN(n8830) );
  NAND2_X1 U10474 ( .A1(n8755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8837) );
  XNOR2_X1 U10475 ( .A(n8837), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U10476 ( .A1(n8847), .A2(n11258), .B1(n8934), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n8756) );
  NAND2_X2 U10477 ( .A1(n8757), .A2(n8756), .ZN(n16400) );
  NAND2_X1 U10478 ( .A1(n8761), .A2(n8760), .ZN(n11014) );
  INV_X1 U10479 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n11015) );
  NAND2_X1 U10480 ( .A1(n8762), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8764) );
  XNOR2_X1 U10481 ( .A(n8764), .B(n8763), .ZN(n11236) );
  OAI22_X1 U10482 ( .A1(n8864), .A2(n11015), .B1(n10830), .B2(n11236), .ZN(
        n8765) );
  INV_X1 U10483 ( .A(n8765), .ZN(n8766) );
  OR2_X1 U10484 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  AND2_X1 U10485 ( .A1(n8771), .A2(n8770), .ZN(n11009) );
  NAND2_X1 U10486 ( .A1(n11009), .A2(n8933), .ZN(n8776) );
  NAND2_X1 U10487 ( .A1(n8782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8773) );
  XNOR2_X1 U10488 ( .A(n8773), .B(n8772), .ZN(n11117) );
  OAI22_X1 U10489 ( .A1(n8864), .A2(n11010), .B1(n10830), .B2(n11117), .ZN(
        n8774) );
  INV_X1 U10490 ( .A(n8774), .ZN(n8775) );
  NAND2_X1 U10491 ( .A1(n8776), .A2(n8775), .ZN(n11906) );
  NAND2_X1 U10492 ( .A1(n8778), .A2(n8777), .ZN(n8780) );
  NAND2_X1 U10493 ( .A1(n8780), .A2(n8779), .ZN(n11001) );
  OR2_X1 U10494 ( .A1(n11001), .A2(n8923), .ZN(n8786) );
  NAND2_X1 U10495 ( .A1(n8791), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8781) );
  MUX2_X1 U10496 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8781), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8783) );
  NAND2_X1 U10497 ( .A1(n8783), .A2(n8782), .ZN(n11162) );
  OAI22_X1 U10498 ( .A1(n8864), .A2(n11002), .B1(n10830), .B2(n11162), .ZN(
        n8784) );
  INV_X1 U10499 ( .A(n8784), .ZN(n8785) );
  XNOR2_X1 U10500 ( .A(n8788), .B(n8787), .ZN(n10998) );
  NAND2_X1 U10501 ( .A1(n10998), .A2(n8862), .ZN(n8795) );
  NOR2_X1 U10502 ( .A1(n8801), .A2(n14795), .ZN(n8789) );
  MUX2_X1 U10503 ( .A(n14795), .B(n8789), .S(P2_IR_REG_4__SCAN_IN), .Z(n8790)
         );
  INV_X1 U10504 ( .A(n8790), .ZN(n8792) );
  NAND2_X1 U10505 ( .A1(n8792), .A2(n8791), .ZN(n11205) );
  OAI22_X1 U10506 ( .A1(n8864), .A2(n11016), .B1(n10830), .B2(n11205), .ZN(
        n8793) );
  INV_X1 U10507 ( .A(n8793), .ZN(n8794) );
  NAND2_X1 U10508 ( .A1(n8795), .A2(n8794), .ZN(n11853) );
  INV_X1 U10509 ( .A(n11853), .ZN(n16298) );
  NOR2_X1 U10510 ( .A1(n8799), .A2(n14795), .ZN(n8800) );
  MUX2_X1 U10511 ( .A(n14795), .B(n8800), .S(P2_IR_REG_3__SCAN_IN), .Z(n8802)
         );
  NOR2_X1 U10512 ( .A1(n8802), .A2(n8801), .ZN(n15572) );
  AOI22_X1 U10513 ( .A1(n8819), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8847), .B2(
        n15572), .ZN(n8803) );
  NAND2_X1 U10514 ( .A1(n8805), .A2(n8804), .ZN(n8806) );
  AND2_X1 U10515 ( .A1(n8807), .A2(n8806), .ZN(n10978) );
  NAND2_X1 U10516 ( .A1(n10978), .A2(n8862), .ZN(n8813) );
  OR2_X1 U10517 ( .A1(n8808), .A2(n14795), .ZN(n8810) );
  XNOR2_X1 U10518 ( .A(n8810), .B(n8809), .ZN(n11220) );
  OAI22_X1 U10519 ( .A1(n8864), .A2(n10989), .B1(n10830), .B2(n11220), .ZN(
        n8811) );
  INV_X1 U10520 ( .A(n8811), .ZN(n8812) );
  INV_X1 U10521 ( .A(n8816), .ZN(n8817) );
  NAND2_X1 U10522 ( .A1(n8815), .A2(n8817), .ZN(n8818) );
  NAND2_X1 U10523 ( .A1(n8814), .A2(n8818), .ZN(n10988) );
  NAND2_X1 U10524 ( .A1(n8819), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U10525 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8820) );
  MUX2_X1 U10526 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8820), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8822) );
  NAND2_X1 U10527 ( .A1(n8822), .A2(n8821), .ZN(n11191) );
  INV_X1 U10528 ( .A(n11191), .ZN(n8823) );
  NAND2_X1 U10529 ( .A1(n8847), .A2(n8823), .ZN(n8824) );
  INV_X1 U10530 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U10531 ( .A1(n10984), .A2(SI_0_), .ZN(n8826) );
  XNOR2_X1 U10532 ( .A(n8826), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14822) );
  MUX2_X1 U10533 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14822), .S(n8827), .Z(n16106)
         );
  XNOR2_X1 U10534 ( .A(n8829), .B(n8828), .ZN(n11022) );
  NAND2_X1 U10535 ( .A1(n11022), .A2(n8933), .ZN(n8833) );
  NAND2_X1 U10536 ( .A1(n8830), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8831) );
  XNOR2_X1 U10537 ( .A(n8831), .B(P2_IR_REG_8__SCAN_IN), .ZN(n15594) );
  AOI22_X1 U10538 ( .A1(n8934), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n15594), 
        .B2(n8847), .ZN(n8832) );
  XNOR2_X1 U10539 ( .A(n8835), .B(n8096), .ZN(n11091) );
  NAND2_X1 U10540 ( .A1(n11091), .A2(n8933), .ZN(n8840) );
  NAND2_X1 U10541 ( .A1(n8837), .A2(n8836), .ZN(n8838) );
  NAND2_X1 U10542 ( .A1(n8838), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8844) );
  XNOR2_X1 U10543 ( .A(n8844), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U10544 ( .A1(n11538), .A2(n8847), .B1(n8934), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8839) );
  INV_X1 U10545 ( .A(n12037), .ZN(n16434) );
  XNOR2_X1 U10546 ( .A(n8842), .B(n8841), .ZN(n11206) );
  NAND2_X1 U10547 ( .A1(n11206), .A2(n8862), .ZN(n8849) );
  NAND2_X1 U10548 ( .A1(n8844), .A2(n8843), .ZN(n8845) );
  NAND2_X1 U10549 ( .A1(n8845), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8846) );
  XNOR2_X1 U10550 ( .A(n8846), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U10551 ( .A1(n11541), .A2(n8847), .B1(n8934), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8848) );
  XNOR2_X1 U10552 ( .A(n8851), .B(n8850), .ZN(n11371) );
  NAND2_X1 U10553 ( .A1(n11371), .A2(n8862), .ZN(n8859) );
  INV_X1 U10554 ( .A(n8852), .ZN(n8856) );
  NAND2_X1 U10555 ( .A1(n8853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8854) );
  MUX2_X1 U10556 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8854), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8855) );
  NAND2_X1 U10557 ( .A1(n8856), .A2(n8855), .ZN(n11943) );
  OAI22_X1 U10558 ( .A1(n8864), .A2(n11403), .B1(n10830), .B2(n11943), .ZN(
        n8857) );
  INV_X1 U10559 ( .A(n8857), .ZN(n8858) );
  NAND2_X1 U10560 ( .A1(n12886), .A2(n12748), .ZN(n12936) );
  XNOR2_X1 U10561 ( .A(n8861), .B(n8860), .ZN(n12178) );
  NAND2_X1 U10562 ( .A1(n12178), .A2(n8933), .ZN(n8867) );
  XNOR2_X1 U10563 ( .A(n8863), .B(n8945), .ZN(n15658) );
  OAI22_X1 U10564 ( .A1(n8864), .A2(n12180), .B1(n10830), .B2(n15658), .ZN(
        n8865) );
  INV_X1 U10565 ( .A(n8865), .ZN(n8866) );
  XNOR2_X1 U10566 ( .A(n9405), .B(n8868), .ZN(n12985) );
  NAND2_X1 U10567 ( .A1(n12985), .A2(n8933), .ZN(n8870) );
  NAND2_X1 U10568 ( .A1(n8934), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8869) );
  INV_X1 U10569 ( .A(n8875), .ZN(n8874) );
  OAI21_X1 U10570 ( .B1(n8874), .B2(n13681), .A(n8878), .ZN(n8881) );
  NOR2_X1 U10571 ( .A1(n8875), .A2(SI_24_), .ZN(n8879) );
  INV_X1 U10572 ( .A(n8876), .ZN(n8877) );
  AOI21_X1 U10573 ( .B1(n8879), .B2(n8878), .A(n8877), .ZN(n8880) );
  MUX2_X1 U10574 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10983), .Z(n8895) );
  NAND2_X1 U10575 ( .A1(n14811), .A2(n8933), .ZN(n8885) );
  NAND2_X1 U10576 ( .A1(n8934), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8884) );
  INV_X1 U10577 ( .A(n14705), .ZN(n14521) );
  NAND2_X1 U10578 ( .A1(n8886), .A2(n8895), .ZN(n8889) );
  INV_X1 U10579 ( .A(n8901), .ZN(n8887) );
  NAND2_X1 U10580 ( .A1(n8887), .A2(SI_26_), .ZN(n8888) );
  MUX2_X1 U10581 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10984), .Z(n8896) );
  XNOR2_X1 U10582 ( .A(n8896), .B(SI_27_), .ZN(n8890) );
  NAND2_X1 U10583 ( .A1(n13086), .A2(n8933), .ZN(n8893) );
  NAND2_X1 U10584 ( .A1(n8934), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8892) );
  INV_X1 U10585 ( .A(n8896), .ZN(n8894) );
  INV_X1 U10586 ( .A(SI_27_), .ZN(n12983) );
  NAND2_X1 U10587 ( .A1(n8894), .A2(n12983), .ZN(n8897) );
  OAI21_X1 U10588 ( .B1(n8895), .B2(SI_26_), .A(n8897), .ZN(n8900) );
  INV_X1 U10589 ( .A(SI_26_), .ZN(n13677) );
  NOR2_X1 U10590 ( .A1(n8883), .A2(n13677), .ZN(n8898) );
  AOI22_X1 U10591 ( .A1(n8898), .A2(n8897), .B1(n8896), .B2(SI_27_), .ZN(n8899) );
  MUX2_X1 U10592 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10984), .Z(n8906) );
  XNOR2_X1 U10593 ( .A(n8906), .B(SI_28_), .ZN(n8904) );
  NAND2_X1 U10594 ( .A1(n14804), .A2(n8933), .ZN(n8903) );
  NAND2_X1 U10595 ( .A1(n8934), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U10596 ( .A1(n14507), .A2(n14493), .ZN(n14490) );
  INV_X1 U10597 ( .A(n8906), .ZN(n8907) );
  INV_X1 U10598 ( .A(SI_28_), .ZN(n13120) );
  NAND2_X1 U10599 ( .A1(n8907), .A2(n13120), .ZN(n8908) );
  MUX2_X1 U10600 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n10984), .Z(n8913) );
  INV_X1 U10601 ( .A(SI_29_), .ZN(n14316) );
  XNOR2_X1 U10602 ( .A(n8913), .B(n14316), .ZN(n8915) );
  NAND2_X1 U10603 ( .A1(n13088), .A2(n8933), .ZN(n8911) );
  NAND2_X1 U10604 ( .A1(n8934), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8910) );
  NOR2_X1 U10605 ( .A1(n8913), .A2(SI_29_), .ZN(n8914) );
  MUX2_X1 U10606 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10984), .Z(n8917) );
  NAND2_X1 U10607 ( .A1(n8917), .A2(SI_30_), .ZN(n8928) );
  OAI21_X1 U10608 ( .B1(SI_30_), .B2(n8917), .A(n8928), .ZN(n8920) );
  INV_X1 U10609 ( .A(n8920), .ZN(n8918) );
  INV_X1 U10610 ( .A(n8919), .ZN(n8921) );
  NAND2_X1 U10611 ( .A1(n8921), .A2(n8920), .ZN(n8922) );
  NAND2_X1 U10612 ( .A1(n8929), .A2(n8922), .ZN(n13122) );
  OR2_X1 U10613 ( .A1(n13122), .A2(n8923), .ZN(n8925) );
  NAND2_X1 U10614 ( .A1(n8934), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U10615 ( .A1(n8929), .A2(n8928), .ZN(n8932) );
  MUX2_X1 U10616 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10983), .Z(n8930) );
  XNOR2_X1 U10617 ( .A(n8930), .B(SI_31_), .ZN(n8931) );
  NAND2_X1 U10618 ( .A1(n14794), .A2(n8933), .ZN(n8936) );
  NAND2_X1 U10619 ( .A1(n8934), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8935) );
  XNOR2_X1 U10620 ( .A(n14481), .B(n8991), .ZN(n8951) );
  NAND2_X1 U10621 ( .A1(n8941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8943) );
  INV_X1 U10622 ( .A(n8944), .ZN(n8947) );
  NAND2_X1 U10623 ( .A1(n8945), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8946) );
  NOR2_X1 U10624 ( .A1(n8947), .A2(n8946), .ZN(n8948) );
  AOI22_X1 U10625 ( .A1(n8863), .A2(n8948), .B1(P2_IR_REG_20__SCAN_IN), .B2(
        n14795), .ZN(n8949) );
  AND2_X2 U10626 ( .A1(n16105), .A2(n12739), .ZN(n16261) );
  NAND2_X1 U10627 ( .A1(n8951), .A2(n16261), .ZN(n14479) );
  XNOR2_X2 U10628 ( .A(n8953), .B(P2_IR_REG_30__SCAN_IN), .ZN(n10259) );
  AND2_X4 U10629 ( .A1(n14802), .A2(n10259), .ZN(n10506) );
  INV_X1 U10630 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n14476) );
  NAND2_X1 U10631 ( .A1(n10505), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8956) );
  AND2_X2 U10632 ( .A1(n13091), .A2(n14802), .ZN(n10302) );
  NAND2_X1 U10633 ( .A1(n10507), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8955) );
  OAI211_X1 U10634 ( .C1(n10499), .C2(n14476), .A(n8956), .B(n8955), .ZN(
        n11026) );
  NOR2_X2 U10635 ( .A1(n10831), .A2(n11102), .ZN(n14628) );
  INV_X1 U10636 ( .A(n14808), .ZN(n11121) );
  NAND2_X1 U10637 ( .A1(n11121), .A2(P2_B_REG_SCAN_IN), .ZN(n8958) );
  NAND2_X1 U10638 ( .A1(n14628), .A2(n8958), .ZN(n10511) );
  INV_X1 U10639 ( .A(n10511), .ZN(n8959) );
  NAND2_X1 U10640 ( .A1(n11026), .A2(n8959), .ZN(n14688) );
  NAND2_X1 U10641 ( .A1(n14479), .A2(n14688), .ZN(n14685) );
  NAND2_X1 U10642 ( .A1(n8968), .A2(n8967), .ZN(n8961) );
  INV_X1 U10643 ( .A(P2_B_REG_SCAN_IN), .ZN(n8969) );
  XOR2_X1 U10644 ( .A(n14818), .B(n8969), .Z(n8970) );
  AND2_X1 U10645 ( .A1(n14815), .A2(n8970), .ZN(n8971) );
  NAND2_X1 U10646 ( .A1(n14813), .A2(n14815), .ZN(n8972) );
  OAI21_X1 U10647 ( .B1(n8989), .B2(P2_D_REG_1__SCAN_IN), .A(n8972), .ZN(
        n10923) );
  NAND2_X1 U10648 ( .A1(n8973), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8975) );
  INV_X1 U10649 ( .A(n10829), .ZN(n10934) );
  AND2_X1 U10650 ( .A1(n10923), .A2(n15571), .ZN(n15564) );
  NOR4_X1 U10651 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n8985) );
  NOR4_X1 U10652 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8980) );
  NOR4_X1 U10653 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8979) );
  NOR4_X1 U10654 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8978) );
  NOR4_X1 U10655 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8977) );
  NAND4_X1 U10656 ( .A1(n8980), .A2(n8979), .A3(n8978), .A4(n8977), .ZN(n8981)
         );
  NOR4_X1 U10657 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        n8982), .A4(n8981), .ZN(n8984) );
  NOR4_X1 U10658 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8983) );
  NAND3_X1 U10659 ( .A1(n8985), .A2(n8984), .A3(n8983), .ZN(n8986) );
  INV_X1 U10660 ( .A(n8989), .ZN(n15566) );
  NAND2_X1 U10661 ( .A1(n8986), .A2(n15566), .ZN(n11739) );
  NAND2_X1 U10662 ( .A1(n16261), .A2(n12849), .ZN(n10932) );
  INV_X1 U10663 ( .A(n10831), .ZN(n10925) );
  NAND2_X1 U10664 ( .A1(n10925), .A2(n10835), .ZN(n11736) );
  AND2_X1 U10665 ( .A1(n10932), .A2(n11736), .ZN(n8987) );
  NAND2_X1 U10666 ( .A1(n14813), .A2(n14818), .ZN(n8988) );
  INV_X1 U10667 ( .A(n8992), .ZN(n8993) );
  NOR2_X2 U10668 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n8996) );
  NOR2_X1 U10669 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .ZN(n9003) );
  NOR2_X1 U10670 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .ZN(n9002) );
  NAND4_X1 U10671 ( .A1(n9599), .A2(n9006), .A3(n9005), .A4(n9602), .ZN(n9007)
         );
  INV_X1 U10672 ( .A(n9015), .ZN(n9013) );
  INV_X2 U10673 ( .A(n9386), .ZN(n9410) );
  NAND2_X1 U10674 ( .A1(n9410), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9024) );
  INV_X1 U10675 ( .A(n9075), .ZN(n9122) );
  NAND2_X1 U10676 ( .A1(n9456), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U10677 ( .A1(n7366), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9022) );
  AND2_X1 U10678 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9123) );
  NAND2_X1 U10679 ( .A1(n9123), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9137) );
  INV_X1 U10680 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9136) );
  NOR2_X1 U10681 ( .A1(n9137), .A2(n9136), .ZN(n9156) );
  NAND2_X1 U10682 ( .A1(n9156), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9170) );
  INV_X1 U10683 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9246) );
  INV_X1 U10684 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U10685 ( .A1(n9283), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9303) );
  INV_X1 U10686 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9302) );
  INV_X1 U10687 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9318) );
  AND2_X1 U10688 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n9016) );
  NAND2_X1 U10689 ( .A1(n9428), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U10690 ( .A1(n9438), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U10691 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n9454), .ZN(n9453) );
  INV_X1 U10692 ( .A(n9453), .ZN(n9018) );
  NAND2_X1 U10693 ( .A1(n9018), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9505) );
  INV_X1 U10694 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U10695 ( .A1(n9453), .A2(n9019), .ZN(n9020) );
  NAND2_X1 U10696 ( .A1(n9505), .A2(n9020), .ZN(n15254) );
  OR2_X1 U10697 ( .A1(n9455), .A2(n15254), .ZN(n9021) );
  XNOR2_X2 U10698 ( .A(n9027), .B(n9026), .ZN(n9598) );
  NAND2_X2 U10699 ( .A1(n9059), .A2(n10976), .ZN(n9481) );
  OR2_X1 U10700 ( .A1(n9513), .A2(n13087), .ZN(n9029) );
  INV_X1 U10701 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U10702 ( .A1(n9033), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9034) );
  MUX2_X1 U10703 ( .A(n9034), .B(P1_IR_REG_31__SCAN_IN), .S(n13875), .Z(n9035)
         );
  NAND2_X1 U10704 ( .A1(n9038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U10705 ( .A1(n9489), .A2(n15311), .ZN(n9042) );
  NAND2_X1 U10706 ( .A1(n11580), .A2(n9042), .ZN(n9479) );
  MUX2_X1 U10707 ( .A(n7690), .B(n12875), .S(n9479), .Z(n9107) );
  MUX2_X1 U10708 ( .A(n8086), .B(n15436), .S(n9500), .Z(n9466) );
  INV_X1 U10709 ( .A(n9466), .ZN(n9469) );
  NAND2_X1 U10710 ( .A1(n9075), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9045) );
  INV_X1 U10711 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9043) );
  INV_X1 U10712 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15691) );
  NOR2_X1 U10713 ( .A1(n10983), .A2(n13718), .ZN(n9046) );
  XNOR2_X1 U10714 ( .A(n9046), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15561) );
  MUX2_X1 U10715 ( .A(n15691), .B(n15561), .S(n9059), .Z(n16142) );
  INV_X1 U10716 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U10717 ( .A1(n9075), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U10718 ( .A1(n9049), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U10719 ( .A1(n9050), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9051) );
  AND2_X1 U10720 ( .A1(n16142), .A2(n11579), .ZN(n9067) );
  OR2_X1 U10721 ( .A1(n16142), .A2(n11579), .ZN(n9068) );
  OAI211_X1 U10722 ( .C1(n11565), .C2(n9067), .A(n15143), .B(n9068), .ZN(n9056) );
  INV_X2 U10723 ( .A(n9107), .ZN(n9253) );
  NAND2_X1 U10724 ( .A1(n9056), .A2(n9253), .ZN(n9057) );
  NAND2_X1 U10725 ( .A1(n9058), .A2(n9057), .ZN(n9074) );
  NAND2_X1 U10726 ( .A1(n16143), .A2(n15143), .ZN(n9066) );
  OR2_X1 U10727 ( .A1(n9513), .A2(n8585), .ZN(n9065) );
  OR2_X1 U10728 ( .A1(n9481), .A2(n10988), .ZN(n9064) );
  NAND2_X1 U10729 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9060) );
  MUX2_X1 U10730 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9060), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9062) );
  NOR2_X1 U10731 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9080) );
  INV_X1 U10732 ( .A(n9080), .ZN(n9061) );
  NAND2_X1 U10733 ( .A1(n9062), .A2(n9061), .ZN(n11288) );
  OR2_X1 U10734 ( .A1(n9059), .A2(n11288), .ZN(n9063) );
  INV_X1 U10735 ( .A(n16155), .ZN(n11566) );
  NAND3_X1 U10736 ( .A1(n9066), .A2(n11566), .A3(n9500), .ZN(n9073) );
  INV_X1 U10737 ( .A(n15143), .ZN(n11064) );
  INV_X1 U10738 ( .A(n9067), .ZN(n9070) );
  NAND2_X1 U10739 ( .A1(n11565), .A2(n9068), .ZN(n9069) );
  NAND3_X1 U10740 ( .A1(n11064), .A2(n9070), .A3(n9069), .ZN(n9071) );
  NAND3_X1 U10741 ( .A1(n9071), .A2(n9253), .A3(n16155), .ZN(n9072) );
  NAND3_X1 U10742 ( .A1(n9074), .A2(n9073), .A3(n9072), .ZN(n9088) );
  NAND2_X1 U10743 ( .A1(n9410), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U10744 ( .A1(n9075), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U10745 ( .A1(n9050), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U10746 ( .A1(n9507), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9076) );
  NAND4_X2 U10747 ( .A1(n9079), .A2(n9078), .A3(n9077), .A4(n9076), .ZN(n11171) );
  INV_X1 U10748 ( .A(n9513), .ZN(n9083) );
  NOR2_X1 U10749 ( .A1(n9080), .A2(n15542), .ZN(n9081) );
  MUX2_X1 U10750 ( .A(n15542), .B(n9081), .S(P1_IR_REG_2__SCAN_IN), .Z(n9082)
         );
  AOI22_X1 U10751 ( .A1(n9083), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9358), .B2(
        n11386), .ZN(n9085) );
  NAND2_X1 U10752 ( .A1(n10978), .A2(n7368), .ZN(n9084) );
  OR2_X1 U10753 ( .A1(n11171), .A2(n11802), .ZN(n11570) );
  INV_X1 U10754 ( .A(n11171), .ZN(n11582) );
  MUX2_X1 U10755 ( .A(n11582), .B(n16204), .S(n9253), .Z(n9086) );
  OAI21_X1 U10756 ( .B1(n9088), .B2(n11570), .A(n9086), .ZN(n9090) );
  NAND2_X1 U10757 ( .A1(n11171), .A2(n11802), .ZN(n9549) );
  INV_X1 U10758 ( .A(n9549), .ZN(n9087) );
  NAND2_X1 U10759 ( .A1(n9088), .A2(n9087), .ZN(n9089) );
  NAND2_X1 U10760 ( .A1(n9090), .A2(n9089), .ZN(n9110) );
  NAND2_X1 U10761 ( .A1(n7537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9091) );
  XNOR2_X1 U10762 ( .A(n9091), .B(P1_IR_REG_3__SCAN_IN), .ZN(n15163) );
  NAND2_X1 U10763 ( .A1(n9504), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U10764 ( .A1(n9075), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9096) );
  NAND2_X1 U10765 ( .A1(n7366), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9095) );
  INV_X1 U10766 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14987) );
  NAND2_X1 U10767 ( .A1(n9507), .A2(n14987), .ZN(n9094) );
  MUX2_X1 U10768 ( .A(n14985), .B(n15141), .S(n9253), .Z(n9109) );
  NAND2_X1 U10769 ( .A1(n10998), .A2(n7368), .ZN(n9100) );
  OR2_X1 U10770 ( .A1(n7537), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U10771 ( .A1(n9116), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9099) );
  XNOR2_X1 U10772 ( .A(n9099), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15172) );
  NAND2_X1 U10773 ( .A1(n9504), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U10774 ( .A1(n9456), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9104) );
  NOR2_X1 U10775 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9101) );
  NOR2_X1 U10776 ( .A1(n9123), .A2(n9101), .ZN(n11811) );
  NAND2_X1 U10777 ( .A1(n9507), .A2(n11811), .ZN(n9103) );
  NAND2_X1 U10778 ( .A1(n7366), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9102) );
  XNOR2_X1 U10779 ( .A(n11816), .B(n12048), .ZN(n11807) );
  INV_X1 U10780 ( .A(n14985), .ZN(n16242) );
  INV_X1 U10781 ( .A(n15141), .ZN(n11573) );
  MUX2_X1 U10782 ( .A(n16242), .B(n11573), .S(n9530), .Z(n9108) );
  NOR2_X1 U10783 ( .A1(n12048), .A2(n9530), .ZN(n9112) );
  INV_X1 U10784 ( .A(n12048), .ZN(n11576) );
  OAI21_X1 U10785 ( .B1(n11576), .B2(n9529), .A(n11816), .ZN(n9111) );
  OAI21_X1 U10786 ( .B1(n9112), .B2(n11816), .A(n9111), .ZN(n9113) );
  OR2_X1 U10787 ( .A1(n11001), .A2(n9481), .ZN(n9121) );
  INV_X1 U10788 ( .A(n9116), .ZN(n9118) );
  INV_X1 U10789 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U10790 ( .A1(n9118), .A2(n9117), .ZN(n9143) );
  NAND2_X1 U10791 ( .A1(n9143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9119) );
  XNOR2_X1 U10792 ( .A(n9119), .B(P1_IR_REG_5__SCAN_IN), .ZN(n11293) );
  AOI22_X1 U10793 ( .A1(n9359), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7365), .B2(
        n11293), .ZN(n9120) );
  NAND2_X1 U10794 ( .A1(n9121), .A2(n9120), .ZN(n16314) );
  NAND2_X1 U10795 ( .A1(n9410), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U10796 ( .A1(n9456), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U10797 ( .A1(n7366), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9125) );
  OAI21_X1 U10798 ( .B1(n9123), .B2(P1_REG3_REG_5__SCAN_IN), .A(n9137), .ZN(
        n11526) );
  OR2_X1 U10799 ( .A1(n9455), .A2(n11526), .ZN(n9124) );
  INV_X1 U10800 ( .A(n11823), .ZN(n15140) );
  MUX2_X1 U10801 ( .A(n16314), .B(n15140), .S(n9253), .Z(n9131) );
  NAND2_X1 U10802 ( .A1(n9130), .A2(n9131), .ZN(n9129) );
  MUX2_X1 U10803 ( .A(n16314), .B(n15140), .S(n9500), .Z(n9128) );
  NAND2_X1 U10804 ( .A1(n9129), .A2(n9128), .ZN(n9135) );
  INV_X1 U10805 ( .A(n9130), .ZN(n9133) );
  INV_X1 U10806 ( .A(n9131), .ZN(n9132) );
  NAND2_X1 U10807 ( .A1(n9133), .A2(n9132), .ZN(n9134) );
  NAND2_X1 U10808 ( .A1(n9456), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U10809 ( .A1(n9504), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9141) );
  AND2_X1 U10810 ( .A1(n9137), .A2(n9136), .ZN(n9138) );
  NOR2_X1 U10811 ( .A1(n9156), .A2(n9138), .ZN(n11831) );
  NAND2_X1 U10812 ( .A1(n9507), .A2(n11831), .ZN(n9140) );
  NAND2_X1 U10813 ( .A1(n7366), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9139) );
  NAND4_X1 U10814 ( .A1(n9142), .A2(n9141), .A3(n9140), .A4(n9139), .ZN(n15139) );
  NAND2_X1 U10815 ( .A1(n11009), .A2(n9512), .ZN(n9148) );
  INV_X1 U10816 ( .A(n9143), .ZN(n9145) );
  NAND2_X1 U10817 ( .A1(n9145), .A2(n9144), .ZN(n9152) );
  NAND2_X1 U10818 ( .A1(n9152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9146) );
  XNOR2_X1 U10819 ( .A(n9146), .B(P1_IR_REG_6__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U10820 ( .A1(n9359), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7365), .B2(
        n11434), .ZN(n9147) );
  NAND2_X1 U10821 ( .A1(n9148), .A2(n9147), .ZN(n11838) );
  MUX2_X1 U10822 ( .A(n15139), .B(n11838), .S(n9253), .Z(n9150) );
  MUX2_X1 U10823 ( .A(n11838), .B(n15139), .S(n9253), .Z(n9149) );
  INV_X1 U10824 ( .A(n9150), .ZN(n9151) );
  OR2_X1 U10825 ( .A1(n11014), .A2(n9481), .ZN(n9155) );
  NAND2_X1 U10826 ( .A1(n9176), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9153) );
  XNOR2_X1 U10827 ( .A(n9153), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U10828 ( .A1(n9359), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7365), .B2(
        n11322), .ZN(n9154) );
  NAND2_X1 U10829 ( .A1(n9155), .A2(n9154), .ZN(n12071) );
  NAND2_X1 U10830 ( .A1(n9504), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U10831 ( .A1(n9456), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9160) );
  OR2_X1 U10832 ( .A1(n9156), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9157) );
  AND2_X1 U10833 ( .A1(n9170), .A2(n9157), .ZN(n12070) );
  NAND2_X1 U10834 ( .A1(n9507), .A2(n12070), .ZN(n9159) );
  NAND2_X1 U10835 ( .A1(n7366), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9158) );
  NAND4_X1 U10836 ( .A1(n9161), .A2(n9160), .A3(n9159), .A4(n9158), .ZN(n15138) );
  MUX2_X1 U10837 ( .A(n12071), .B(n15138), .S(n9253), .Z(n9165) );
  NAND2_X1 U10838 ( .A1(n9164), .A2(n9165), .ZN(n9163) );
  MUX2_X1 U10839 ( .A(n12071), .B(n15138), .S(n9500), .Z(n9162) );
  NAND2_X1 U10840 ( .A1(n9163), .A2(n9162), .ZN(n9169) );
  INV_X1 U10841 ( .A(n9164), .ZN(n9167) );
  INV_X1 U10842 ( .A(n9165), .ZN(n9166) );
  NAND2_X1 U10843 ( .A1(n9167), .A2(n9166), .ZN(n9168) );
  NAND2_X1 U10844 ( .A1(n9456), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U10845 ( .A1(n7366), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U10846 ( .A1(n9170), .A2(n12174), .ZN(n9171) );
  AND2_X1 U10847 ( .A1(n9184), .A2(n9171), .ZN(n12185) );
  NAND2_X1 U10848 ( .A1(n9507), .A2(n12185), .ZN(n9173) );
  NAND2_X1 U10849 ( .A1(n9410), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9172) );
  NAND4_X1 U10850 ( .A1(n9175), .A2(n9174), .A3(n9173), .A4(n9172), .ZN(n15137) );
  NAND2_X1 U10851 ( .A1(n11022), .A2(n9512), .ZN(n9179) );
  OAI21_X1 U10852 ( .B1(n9176), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9177) );
  XNOR2_X1 U10853 ( .A(n9177), .B(P1_IR_REG_8__SCAN_IN), .ZN(n15196) );
  AOI22_X1 U10854 ( .A1(n9359), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7365), .B2(
        n15196), .ZN(n9178) );
  NAND2_X1 U10855 ( .A1(n9179), .A2(n9178), .ZN(n12186) );
  MUX2_X1 U10856 ( .A(n15137), .B(n12186), .S(n9253), .Z(n9182) );
  MUX2_X1 U10857 ( .A(n15137), .B(n12186), .S(n9500), .Z(n9180) );
  NAND2_X1 U10858 ( .A1(n9504), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9189) );
  NAND2_X1 U10859 ( .A1(n9456), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9188) );
  AND2_X1 U10860 ( .A1(n9184), .A2(n9183), .ZN(n9185) );
  NOR2_X1 U10861 ( .A1(n9200), .A2(n9185), .ZN(n12369) );
  NAND2_X1 U10862 ( .A1(n9507), .A2(n12369), .ZN(n9187) );
  NAND2_X1 U10863 ( .A1(n7366), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9186) );
  INV_X1 U10864 ( .A(n12365), .ZN(n12270) );
  NAND2_X1 U10865 ( .A1(n11131), .A2(n9512), .ZN(n9193) );
  OR2_X1 U10866 ( .A1(n9190), .A2(n15542), .ZN(n9191) );
  XNOR2_X1 U10867 ( .A(n9191), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U10868 ( .A1(n9359), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7365), .B2(
        n11356), .ZN(n9192) );
  NAND2_X2 U10869 ( .A1(n9193), .A2(n9192), .ZN(n16388) );
  MUX2_X1 U10870 ( .A(n12270), .B(n16388), .S(n9500), .Z(n9207) );
  MUX2_X1 U10871 ( .A(n12270), .B(n16388), .S(n9253), .Z(n9194) );
  NAND2_X1 U10872 ( .A1(n9195), .A2(n9194), .ZN(n9206) );
  NAND2_X1 U10873 ( .A1(n11091), .A2(n9512), .ZN(n9199) );
  NAND2_X1 U10874 ( .A1(n9196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9197) );
  XNOR2_X1 U10875 ( .A(n9197), .B(P1_IR_REG_10__SCAN_IN), .ZN(n15212) );
  AOI22_X1 U10876 ( .A1(n9359), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7365), 
        .B2(n15212), .ZN(n9198) );
  NAND2_X1 U10877 ( .A1(n9504), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U10878 ( .A1(n9456), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U10879 ( .A1(n7366), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9203) );
  NOR2_X1 U10880 ( .A1(n9200), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9201) );
  OR2_X1 U10881 ( .A1(n9213), .A2(n9201), .ZN(n12488) );
  OR2_X1 U10882 ( .A1(n9455), .A2(n12488), .ZN(n9202) );
  XNOR2_X1 U10883 ( .A(n16421), .B(n12343), .ZN(n12339) );
  OAI211_X1 U10884 ( .C1(n9208), .C2(n9207), .A(n9206), .B(n12268), .ZN(n9212)
         );
  NOR2_X1 U10885 ( .A1(n12343), .A2(n9530), .ZN(n9210) );
  OAI21_X1 U10886 ( .B1(n9529), .B2(n15136), .A(n16421), .ZN(n9209) );
  OAI21_X1 U10887 ( .B1(n9210), .B2(n16421), .A(n9209), .ZN(n9211) );
  NAND2_X1 U10888 ( .A1(n9212), .A2(n9211), .ZN(n9223) );
  NAND2_X1 U10889 ( .A1(n9410), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U10890 ( .A1(n9456), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U10891 ( .A1(n7366), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9216) );
  OR2_X1 U10892 ( .A1(n9213), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U10893 ( .A1(n9234), .A2(n9214), .ZN(n12352) );
  OR2_X1 U10894 ( .A1(n9455), .A2(n12352), .ZN(n9215) );
  NAND2_X1 U10895 ( .A1(n11206), .A2(n9512), .ZN(n9220) );
  OR2_X1 U10896 ( .A1(n9196), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U10897 ( .A1(n9293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9229) );
  XNOR2_X1 U10898 ( .A(n9229), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U10899 ( .A1(n9359), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7365), 
        .B2(n11614), .ZN(n9219) );
  MUX2_X1 U10900 ( .A(n15135), .B(n12642), .S(n9530), .Z(n9224) );
  NAND2_X1 U10901 ( .A1(n9223), .A2(n9224), .ZN(n9222) );
  MUX2_X1 U10902 ( .A(n15135), .B(n12642), .S(n9253), .Z(n9221) );
  NAND2_X1 U10903 ( .A1(n9222), .A2(n9221), .ZN(n9228) );
  INV_X1 U10904 ( .A(n9223), .ZN(n9226) );
  INV_X1 U10905 ( .A(n9224), .ZN(n9225) );
  NAND2_X1 U10906 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  NAND2_X1 U10907 ( .A1(n11371), .A2(n9512), .ZN(n9232) );
  INV_X1 U10908 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n13862) );
  NAND2_X1 U10909 ( .A1(n9229), .A2(n13862), .ZN(n9230) );
  NAND2_X1 U10910 ( .A1(n9230), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9242) );
  XNOR2_X1 U10911 ( .A(n9242), .B(P1_IR_REG_12__SCAN_IN), .ZN(n15723) );
  AOI22_X1 U10912 ( .A1(n9359), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7365), 
        .B2(n15723), .ZN(n9231) );
  NAND2_X1 U10913 ( .A1(n9456), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U10914 ( .A1(n9504), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U10915 ( .A1(n9234), .A2(n9233), .ZN(n9235) );
  AND2_X1 U10916 ( .A1(n9247), .A2(n9235), .ZN(n12732) );
  NAND2_X1 U10917 ( .A1(n9507), .A2(n12732), .ZN(n9237) );
  NAND2_X1 U10918 ( .A1(n7366), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9236) );
  NAND4_X1 U10919 ( .A1(n9239), .A2(n9238), .A3(n9237), .A4(n9236), .ZN(n15134) );
  MUX2_X1 U10920 ( .A(n16482), .B(n15134), .S(n9530), .Z(n9241) );
  MUX2_X1 U10921 ( .A(n16482), .B(n15134), .S(n9253), .Z(n9240) );
  OR2_X1 U10922 ( .A1(n11400), .A2(n9481), .ZN(n9245) );
  INV_X1 U10923 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U10924 ( .A1(n9242), .A2(n9289), .ZN(n9243) );
  NAND2_X1 U10925 ( .A1(n9243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9270) );
  XNOR2_X1 U10926 ( .A(n9270), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U10927 ( .A1(n9359), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7365), 
        .B2(n11617), .ZN(n9244) );
  NAND2_X1 U10928 ( .A1(n9456), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U10929 ( .A1(n7366), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U10930 ( .A1(n9247), .A2(n9246), .ZN(n9248) );
  AND2_X1 U10931 ( .A1(n9263), .A2(n9248), .ZN(n12868) );
  NAND2_X1 U10932 ( .A1(n9507), .A2(n12868), .ZN(n9250) );
  NAND2_X1 U10933 ( .A1(n9410), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9249) );
  NAND4_X1 U10934 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(n15133) );
  MUX2_X1 U10935 ( .A(n16493), .B(n15133), .S(n9253), .Z(n9257) );
  NAND2_X1 U10936 ( .A1(n9256), .A2(n9257), .ZN(n9255) );
  MUX2_X1 U10937 ( .A(n15133), .B(n16493), .S(n9529), .Z(n9254) );
  NAND2_X1 U10938 ( .A1(n9255), .A2(n9254), .ZN(n9261) );
  INV_X1 U10939 ( .A(n9256), .ZN(n9259) );
  INV_X1 U10940 ( .A(n9257), .ZN(n9258) );
  NAND2_X1 U10941 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  AND2_X1 U10942 ( .A1(n9263), .A2(n9262), .ZN(n9264) );
  OR2_X1 U10943 ( .A1(n9264), .A2(n9283), .ZN(n16526) );
  INV_X1 U10944 ( .A(n16526), .ZN(n9265) );
  NAND2_X1 U10945 ( .A1(n9265), .A2(n9507), .ZN(n9269) );
  NAND2_X1 U10946 ( .A1(n9504), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U10947 ( .A1(n9456), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U10948 ( .A1(n7366), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9266) );
  NAND4_X1 U10949 ( .A1(n9269), .A2(n9268), .A3(n9267), .A4(n9266), .ZN(n15132) );
  NAND2_X1 U10950 ( .A1(n11515), .A2(n9512), .ZN(n9274) );
  INV_X1 U10951 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U10952 ( .A1(n9270), .A2(n13868), .ZN(n9271) );
  NAND2_X1 U10953 ( .A1(n9271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9272) );
  XNOR2_X1 U10954 ( .A(n9272), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U10955 ( .A1(n9359), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n12311), 
        .B2(n7365), .ZN(n9273) );
  MUX2_X1 U10956 ( .A(n15132), .B(n16523), .S(n9529), .Z(n9278) );
  NAND2_X1 U10957 ( .A1(n9277), .A2(n9278), .ZN(n9276) );
  MUX2_X1 U10958 ( .A(n15132), .B(n16523), .S(n9530), .Z(n9275) );
  NAND2_X1 U10959 ( .A1(n9276), .A2(n9275), .ZN(n9282) );
  INV_X1 U10960 ( .A(n9277), .ZN(n9280) );
  INV_X1 U10961 ( .A(n9278), .ZN(n9279) );
  NAND2_X1 U10962 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  OR2_X1 U10963 ( .A1(n9283), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U10964 ( .A1(n9303), .A2(n9284), .ZN(n15112) );
  NAND2_X1 U10965 ( .A1(n7366), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9285) );
  OAI21_X1 U10966 ( .B1(n15112), .B2(n9455), .A(n9285), .ZN(n9288) );
  INV_X1 U10967 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12709) );
  NAND2_X1 U10968 ( .A1(n9456), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9286) );
  OAI21_X1 U10969 ( .B1(n12709), .B2(n9386), .A(n9286), .ZN(n9287) );
  NAND2_X1 U10970 ( .A1(n11863), .A2(n9512), .ZN(n9299) );
  INV_X1 U10971 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9290) );
  NAND3_X1 U10972 ( .A1(n9291), .A2(n9290), .A3(n9289), .ZN(n9292) );
  NOR2_X1 U10973 ( .A1(n9293), .A2(n9292), .ZN(n9295) );
  OR2_X1 U10974 ( .A1(n9295), .A2(n15542), .ZN(n9294) );
  MUX2_X1 U10975 ( .A(n9294), .B(P1_IR_REG_31__SCAN_IN), .S(n13871), .Z(n9296)
         );
  NAND2_X1 U10976 ( .A1(n9295), .A2(n13871), .ZN(n9323) );
  NAND2_X1 U10977 ( .A1(n9296), .A2(n9323), .ZN(n15705) );
  INV_X1 U10978 ( .A(n15705), .ZN(n9297) );
  AOI22_X1 U10979 ( .A1(n9359), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7365), 
        .B2(n9297), .ZN(n9298) );
  MUX2_X1 U10980 ( .A(n15131), .B(n16529), .S(n9530), .Z(n9301) );
  MUX2_X1 U10981 ( .A(n15131), .B(n16529), .S(n9529), .Z(n9300) );
  NAND2_X1 U10982 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  NAND2_X1 U10983 ( .A1(n9319), .A2(n9304), .ZN(n16554) );
  AOI22_X1 U10984 ( .A1(n9410), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9456), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n9306) );
  NAND2_X1 U10985 ( .A1(n7366), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9305) );
  OAI211_X1 U10986 ( .C1(n16554), .C2(n9455), .A(n9306), .B(n9305), .ZN(n15130) );
  NAND2_X1 U10987 ( .A1(n12022), .A2(n9512), .ZN(n9309) );
  NAND2_X1 U10988 ( .A1(n9323), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9307) );
  XNOR2_X1 U10989 ( .A(n9307), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U10990 ( .A1(n9359), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7365), 
        .B2(n12609), .ZN(n9308) );
  MUX2_X1 U10991 ( .A(n15130), .B(n16550), .S(n9529), .Z(n9313) );
  NAND2_X1 U10992 ( .A1(n9312), .A2(n9313), .ZN(n9311) );
  MUX2_X1 U10993 ( .A(n15130), .B(n16550), .S(n9530), .Z(n9310) );
  NAND2_X1 U10994 ( .A1(n9311), .A2(n9310), .ZN(n9317) );
  INV_X1 U10995 ( .A(n9312), .ZN(n9315) );
  INV_X1 U10996 ( .A(n9313), .ZN(n9314) );
  NAND2_X1 U10997 ( .A1(n9315), .A2(n9314), .ZN(n9316) );
  AND2_X1 U10998 ( .A1(n9319), .A2(n9318), .ZN(n9320) );
  OR2_X1 U10999 ( .A1(n9320), .A2(n9351), .ZN(n15044) );
  AOI22_X1 U11000 ( .A1(n9410), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9456), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U11001 ( .A1(n7366), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9321) );
  OAI211_X1 U11002 ( .C1(n15044), .C2(n9455), .A(n9322), .B(n9321), .ZN(n15129) );
  NAND2_X1 U11003 ( .A1(n12178), .A2(n9512), .ZN(n9328) );
  OR2_X1 U11004 ( .A1(n9323), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U11005 ( .A1(n9324), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11006 ( .A1(n9325), .A2(n13878), .ZN(n9339) );
  OR2_X1 U11007 ( .A1(n9325), .A2(n13878), .ZN(n9326) );
  AND2_X1 U11008 ( .A1(n9339), .A2(n9326), .ZN(n12970) );
  AOI22_X1 U11009 ( .A1(n9359), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7365), 
        .B2(n12970), .ZN(n9327) );
  MUX2_X1 U11010 ( .A(n15129), .B(n15508), .S(n9500), .Z(n9330) );
  MUX2_X1 U11011 ( .A(n15129), .B(n15508), .S(n9529), .Z(n9329) );
  INV_X1 U11012 ( .A(n9330), .ZN(n9331) );
  INV_X1 U11013 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9332) );
  XNOR2_X1 U11014 ( .A(n9351), .B(n9332), .ZN(n15388) );
  NAND2_X1 U11015 ( .A1(n15388), .A2(n9507), .ZN(n9338) );
  INV_X1 U11016 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n12971) );
  NAND2_X1 U11017 ( .A1(n9504), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11018 ( .A1(n9456), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9333) );
  OAI211_X1 U11019 ( .C1(n12971), .C2(n9335), .A(n9334), .B(n9333), .ZN(n9336)
         );
  INV_X1 U11020 ( .A(n9336), .ZN(n9337) );
  NAND2_X1 U11021 ( .A1(n9338), .A2(n9337), .ZN(n15128) );
  NAND2_X1 U11022 ( .A1(n9339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9340) );
  XNOR2_X1 U11023 ( .A(n9340), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15222) );
  AOI22_X1 U11024 ( .A1(n15222), .A2(n7365), .B1(n9359), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n9341) );
  MUX2_X1 U11025 ( .A(n15128), .B(n15500), .S(n9529), .Z(n9346) );
  NAND2_X1 U11026 ( .A1(n9345), .A2(n9346), .ZN(n9344) );
  MUX2_X1 U11027 ( .A(n15500), .B(n15128), .S(n9529), .Z(n9343) );
  NAND2_X1 U11028 ( .A1(n9344), .A2(n9343), .ZN(n9350) );
  INV_X1 U11029 ( .A(n9345), .ZN(n9348) );
  INV_X1 U11030 ( .A(n9346), .ZN(n9347) );
  NAND2_X1 U11031 ( .A1(n9348), .A2(n9347), .ZN(n9349) );
  AOI21_X1 U11032 ( .B1(n9351), .B2(P1_REG3_REG_18__SCAN_IN), .A(
        P1_REG3_REG_19__SCAN_IN), .ZN(n9352) );
  OR2_X1 U11033 ( .A1(n9365), .A2(n9352), .ZN(n15367) );
  INV_X1 U11034 ( .A(n15367), .ZN(n14995) );
  NAND2_X1 U11035 ( .A1(n14995), .A2(n9507), .ZN(n9357) );
  INV_X1 U11036 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15366) );
  NAND2_X1 U11037 ( .A1(n7366), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U11038 ( .A1(n9456), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9353) );
  OAI211_X1 U11039 ( .C1(n9386), .C2(n15366), .A(n9354), .B(n9353), .ZN(n9355)
         );
  INV_X1 U11040 ( .A(n9355), .ZN(n9356) );
  INV_X1 U11041 ( .A(n15088), .ZN(n15127) );
  NAND2_X1 U11042 ( .A1(n12557), .A2(n9512), .ZN(n9361) );
  AOI22_X1 U11043 ( .A1(n9359), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7363), 
        .B2(n7365), .ZN(n9360) );
  MUX2_X1 U11044 ( .A(n15127), .B(n15370), .S(n9500), .Z(n9363) );
  MUX2_X1 U11045 ( .A(n15127), .B(n15370), .S(n9529), .Z(n9362) );
  INV_X1 U11046 ( .A(n9363), .ZN(n9364) );
  NOR2_X1 U11047 ( .A1(n9365), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9366) );
  OR2_X1 U11048 ( .A1(n9381), .A2(n9366), .ZN(n15350) );
  INV_X1 U11049 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15355) );
  NAND2_X1 U11050 ( .A1(n9456), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11051 ( .A1(n7366), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9367) );
  OAI211_X1 U11052 ( .C1(n9386), .C2(n15355), .A(n9368), .B(n9367), .ZN(n9369)
         );
  INV_X1 U11053 ( .A(n9369), .ZN(n9370) );
  OAI21_X1 U11054 ( .B1(n15350), .B2(n9455), .A(n9370), .ZN(n15126) );
  NAND2_X1 U11055 ( .A1(n12738), .A2(n9512), .ZN(n9372) );
  OR2_X1 U11056 ( .A1(n9513), .A2(n12771), .ZN(n9371) );
  MUX2_X1 U11057 ( .A(n15126), .B(n15484), .S(n9529), .Z(n9376) );
  NAND2_X1 U11058 ( .A1(n9375), .A2(n9376), .ZN(n9374) );
  MUX2_X1 U11059 ( .A(n15484), .B(n15126), .S(n9529), .Z(n9373) );
  NAND2_X1 U11060 ( .A1(n9374), .A2(n9373), .ZN(n9380) );
  INV_X1 U11061 ( .A(n9375), .ZN(n9378) );
  INV_X1 U11062 ( .A(n9376), .ZN(n9377) );
  NAND2_X1 U11063 ( .A1(n9378), .A2(n9377), .ZN(n9379) );
  OR2_X1 U11064 ( .A1(n9381), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9382) );
  AND2_X1 U11065 ( .A1(n9382), .A2(n9400), .ZN(n15338) );
  NAND2_X1 U11066 ( .A1(n15338), .A2(n9507), .ZN(n9389) );
  INV_X1 U11067 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U11068 ( .A1(n7366), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11069 ( .A1(n9456), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9383) );
  OAI211_X1 U11070 ( .C1(n9386), .C2(n9385), .A(n9384), .B(n9383), .ZN(n9387)
         );
  INV_X1 U11071 ( .A(n9387), .ZN(n9388) );
  NAND2_X1 U11072 ( .A1(n9389), .A2(n9388), .ZN(n15125) );
  NAND2_X1 U11073 ( .A1(n12874), .A2(n9512), .ZN(n9391) );
  OR2_X1 U11074 ( .A1(n9513), .A2(n12876), .ZN(n9390) );
  MUX2_X1 U11075 ( .A(n15125), .B(n15334), .S(n9500), .Z(n9395) );
  NAND2_X1 U11076 ( .A1(n9394), .A2(n9395), .ZN(n9393) );
  MUX2_X1 U11077 ( .A(n15125), .B(n15334), .S(n9529), .Z(n9392) );
  NAND2_X1 U11078 ( .A1(n9393), .A2(n9392), .ZN(n9399) );
  INV_X1 U11079 ( .A(n9394), .ZN(n9397) );
  INV_X1 U11080 ( .A(n9395), .ZN(n9396) );
  NAND2_X1 U11081 ( .A1(n9397), .A2(n9396), .ZN(n9398) );
  NAND2_X1 U11082 ( .A1(n9504), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U11083 ( .A1(n9456), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9403) );
  INV_X1 U11084 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15077) );
  AOI21_X1 U11085 ( .B1(n15077), .B2(n9400), .A(n9412), .ZN(n15323) );
  NAND2_X1 U11086 ( .A1(n9507), .A2(n15323), .ZN(n9402) );
  NAND2_X1 U11087 ( .A1(n7366), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9401) );
  NAND4_X1 U11088 ( .A1(n9404), .A2(n9403), .A3(n9402), .A4(n9401), .ZN(n15124) );
  OR2_X1 U11089 ( .A1(n9405), .A2(n10984), .ZN(n9406) );
  MUX2_X1 U11090 ( .A(n15124), .B(n15470), .S(n9529), .Z(n9408) );
  MUX2_X1 U11091 ( .A(n15470), .B(n15124), .S(n9529), .Z(n9407) );
  INV_X1 U11092 ( .A(n9408), .ZN(n9409) );
  NAND2_X1 U11093 ( .A1(n9410), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U11094 ( .A1(n9456), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U11095 ( .A1(n7366), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9414) );
  OAI21_X1 U11096 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9412), .A(n9411), .ZN(
        n14976) );
  OR2_X1 U11097 ( .A1(n9455), .A2(n14976), .ZN(n9413) );
  NAND2_X1 U11098 ( .A1(n13009), .A2(n9512), .ZN(n9418) );
  OR2_X1 U11099 ( .A1(n9513), .A2(n13015), .ZN(n9417) );
  MUX2_X1 U11100 ( .A(n15123), .B(n14928), .S(n9500), .Z(n9422) );
  NAND2_X1 U11101 ( .A1(n9421), .A2(n9422), .ZN(n9420) );
  MUX2_X1 U11102 ( .A(n15123), .B(n14928), .S(n9529), .Z(n9419) );
  NAND2_X1 U11103 ( .A1(n9420), .A2(n9419), .ZN(n9426) );
  INV_X1 U11104 ( .A(n9421), .ZN(n9424) );
  INV_X1 U11105 ( .A(n9422), .ZN(n9423) );
  NAND2_X1 U11106 ( .A1(n9424), .A2(n9423), .ZN(n9425) );
  NAND2_X1 U11107 ( .A1(n9456), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11108 ( .A1(n7366), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U11109 ( .A1(n9410), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9430) );
  OAI21_X1 U11110 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9428), .A(n9427), .ZN(
        n15295) );
  OR2_X1 U11111 ( .A1(n9455), .A2(n15295), .ZN(n9429) );
  INV_X1 U11112 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15557) );
  OR2_X1 U11113 ( .A1(n9513), .A2(n15557), .ZN(n9433) );
  MUX2_X1 U11114 ( .A(n15122), .B(n15457), .S(n9529), .Z(n9436) );
  MUX2_X1 U11115 ( .A(n15122), .B(n15457), .S(n9500), .Z(n9435) );
  NAND2_X1 U11116 ( .A1(n9410), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U11117 ( .A1(n9456), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U11118 ( .A1(n7366), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9440) );
  OAI21_X1 U11119 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9438), .A(n9437), .ZN(
        n15031) );
  OR2_X1 U11120 ( .A1(n9455), .A2(n15031), .ZN(n9439) );
  OR2_X1 U11121 ( .A1(n9513), .A2(n15553), .ZN(n9443) );
  MUX2_X1 U11122 ( .A(n15121), .B(n9544), .S(n9500), .Z(n9448) );
  NAND2_X1 U11123 ( .A1(n9447), .A2(n9448), .ZN(n9446) );
  MUX2_X1 U11124 ( .A(n15121), .B(n9544), .S(n9529), .Z(n9445) );
  NAND2_X1 U11125 ( .A1(n9446), .A2(n9445), .ZN(n9452) );
  INV_X1 U11126 ( .A(n9447), .ZN(n9450) );
  INV_X1 U11127 ( .A(n9448), .ZN(n9449) );
  NAND2_X1 U11128 ( .A1(n9450), .A2(n9449), .ZN(n9451) );
  OAI21_X1 U11129 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n9454), .A(n9453), .ZN(
        n15270) );
  OR2_X1 U11130 ( .A1(n9455), .A2(n15270), .ZN(n9460) );
  NAND2_X1 U11131 ( .A1(n9504), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9459) );
  NAND2_X1 U11132 ( .A1(n9456), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9458) );
  NAND2_X1 U11133 ( .A1(n7366), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9457) );
  NAND4_X1 U11134 ( .A1(n9460), .A2(n9459), .A3(n9458), .A4(n9457), .ZN(n15120) );
  NAND2_X1 U11135 ( .A1(n14811), .A2(n9512), .ZN(n9462) );
  INV_X1 U11136 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15548) );
  OR2_X1 U11137 ( .A1(n9513), .A2(n15548), .ZN(n9461) );
  MUX2_X1 U11138 ( .A(n15120), .B(n15274), .S(n9529), .Z(n9464) );
  MUX2_X1 U11139 ( .A(n15274), .B(n15120), .S(n9529), .Z(n9463) );
  INV_X1 U11140 ( .A(n9467), .ZN(n9468) );
  INV_X1 U11141 ( .A(n15436), .ZN(n15257) );
  MUX2_X1 U11142 ( .A(n9565), .B(n15257), .S(n9529), .Z(n9465) );
  NAND2_X1 U11143 ( .A1(n14794), .A2(n9512), .ZN(n9472) );
  INV_X1 U11144 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9470) );
  OR2_X1 U11145 ( .A1(n9513), .A2(n9470), .ZN(n9471) );
  NAND2_X1 U11146 ( .A1(n7366), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U11147 ( .A1(n9504), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U11148 ( .A1(n9456), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9473) );
  NAND3_X1 U11149 ( .A1(n9475), .A2(n9474), .A3(n9473), .ZN(n15238) );
  XNOR2_X1 U11150 ( .A(n9583), .B(n15238), .ZN(n9567) );
  NAND2_X1 U11151 ( .A1(n7366), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9478) );
  NAND2_X1 U11152 ( .A1(n9410), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U11153 ( .A1(n9456), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9476) );
  NAND3_X1 U11154 ( .A1(n9478), .A2(n9477), .A3(n9476), .ZN(n15117) );
  OAI21_X1 U11155 ( .B1(n15238), .B2(n9479), .A(n15117), .ZN(n9480) );
  INV_X1 U11156 ( .A(n9480), .ZN(n9484) );
  OR2_X1 U11157 ( .A1(n13122), .A2(n9481), .ZN(n9483) );
  INV_X1 U11158 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13268) );
  OR2_X1 U11159 ( .A1(n9513), .A2(n13268), .ZN(n9482) );
  MUX2_X1 U11160 ( .A(n9484), .B(n15241), .S(n9529), .Z(n9524) );
  INV_X1 U11161 ( .A(n9524), .ZN(n9487) );
  OAI21_X1 U11162 ( .B1(n15238), .B2(n12770), .A(n15117), .ZN(n9485) );
  INV_X1 U11163 ( .A(n9485), .ZN(n9486) );
  MUX2_X1 U11164 ( .A(n15241), .B(n9486), .S(n9529), .Z(n9523) );
  NAND2_X1 U11165 ( .A1(n9487), .A2(n9523), .ZN(n9569) );
  NAND2_X1 U11166 ( .A1(n15559), .A2(n11588), .ZN(n11005) );
  NAND2_X1 U11167 ( .A1(n11564), .A2(n12770), .ZN(n9490) );
  NAND2_X1 U11168 ( .A1(n11005), .A2(n9490), .ZN(n9491) );
  OR2_X1 U11169 ( .A1(n11579), .A2(n12559), .ZN(n16093) );
  NAND2_X1 U11170 ( .A1(n9491), .A2(n16093), .ZN(n9581) );
  INV_X1 U11171 ( .A(n9581), .ZN(n9492) );
  NAND3_X1 U11172 ( .A1(n9567), .A2(n9569), .A3(n9492), .ZN(n9531) );
  INV_X1 U11173 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13089) );
  NOR2_X1 U11174 ( .A1(n9513), .A2(n13089), .ZN(n9493) );
  NAND2_X1 U11175 ( .A1(n9504), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U11176 ( .A1(n9456), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9498) );
  INV_X1 U11177 ( .A(n9505), .ZN(n9494) );
  NAND2_X1 U11178 ( .A1(n9494), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13078) );
  INV_X1 U11179 ( .A(n13078), .ZN(n9495) );
  NAND2_X1 U11180 ( .A1(n9507), .A2(n9495), .ZN(n9497) );
  NAND2_X1 U11181 ( .A1(n7366), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9496) );
  NAND4_X1 U11182 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n15118) );
  MUX2_X1 U11183 ( .A(n13075), .B(n15118), .S(n9530), .Z(n9526) );
  INV_X1 U11184 ( .A(n9526), .ZN(n9503) );
  INV_X1 U11185 ( .A(n15118), .ZN(n9501) );
  MUX2_X1 U11186 ( .A(n9501), .B(n15422), .S(n9500), .Z(n9527) );
  INV_X1 U11187 ( .A(n9527), .ZN(n9502) );
  AND2_X1 U11188 ( .A1(n9503), .A2(n9502), .ZN(n9536) );
  NOR2_X1 U11189 ( .A1(n9531), .A2(n9536), .ZN(n9519) );
  NAND2_X1 U11190 ( .A1(n9456), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U11191 ( .A1(n9504), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9510) );
  INV_X1 U11192 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n15010) );
  NAND2_X1 U11193 ( .A1(n9505), .A2(n15010), .ZN(n9506) );
  NAND2_X1 U11194 ( .A1(n9507), .A2(n15013), .ZN(n9509) );
  NAND2_X1 U11195 ( .A1(n7366), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9508) );
  NAND4_X1 U11196 ( .A1(n9511), .A2(n9510), .A3(n9509), .A4(n9508), .ZN(n15119) );
  NAND2_X1 U11197 ( .A1(n14804), .A2(n9512), .ZN(n9515) );
  INV_X1 U11198 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13093) );
  OR2_X1 U11199 ( .A1(n9513), .A2(n13093), .ZN(n9514) );
  MUX2_X1 U11200 ( .A(n15119), .B(n15428), .S(n9529), .Z(n9520) );
  INV_X1 U11201 ( .A(n9520), .ZN(n9517) );
  MUX2_X1 U11202 ( .A(n15004), .B(n15006), .S(n9530), .Z(n9521) );
  INV_X1 U11203 ( .A(n9521), .ZN(n9516) );
  NAND2_X1 U11204 ( .A1(n9517), .A2(n9516), .ZN(n9540) );
  INV_X1 U11205 ( .A(n9519), .ZN(n9522) );
  NAND2_X1 U11206 ( .A1(n9521), .A2(n9520), .ZN(n9592) );
  NOR2_X1 U11207 ( .A1(n9522), .A2(n9592), .ZN(n9543) );
  INV_X1 U11208 ( .A(n9523), .ZN(n9525) );
  NAND2_X1 U11209 ( .A1(n9525), .A2(n9524), .ZN(n9535) );
  NAND2_X1 U11210 ( .A1(n9527), .A2(n9526), .ZN(n9528) );
  NAND2_X1 U11211 ( .A1(n9535), .A2(n9528), .ZN(n9532) );
  NAND2_X1 U11212 ( .A1(n9529), .A2(n15238), .ZN(n9574) );
  OR2_X1 U11213 ( .A1(n9583), .A2(n9574), .ZN(n9570) );
  INV_X1 U11214 ( .A(n15238), .ZN(n9578) );
  AND2_X1 U11215 ( .A1(n9578), .A2(n9530), .ZN(n9577) );
  NAND2_X1 U11216 ( .A1(n9583), .A2(n9577), .ZN(n9571) );
  NAND2_X1 U11217 ( .A1(n12875), .A2(n7690), .ZN(n9588) );
  NAND4_X1 U11218 ( .A1(n9570), .A2(n9571), .A3(n9581), .A4(n9588), .ZN(n9534)
         );
  NOR2_X1 U11219 ( .A1(n9532), .A2(n9534), .ZN(n9593) );
  INV_X1 U11220 ( .A(n9593), .ZN(n9541) );
  INV_X1 U11221 ( .A(n9531), .ZN(n9533) );
  NAND2_X1 U11222 ( .A1(n9533), .A2(n9532), .ZN(n9539) );
  INV_X1 U11223 ( .A(n9534), .ZN(n9537) );
  NAND3_X1 U11224 ( .A1(n9537), .A2(n9536), .A3(n9535), .ZN(n9538) );
  OAI211_X1 U11225 ( .C1(n9541), .C2(n9540), .A(n9539), .B(n9538), .ZN(n9542)
         );
  NOR2_X1 U11226 ( .A1(n9543), .A2(n9542), .ZN(n9591) );
  XNOR2_X1 U11227 ( .A(n15241), .B(n15117), .ZN(n9563) );
  NAND2_X1 U11228 ( .A1(n9544), .A2(n15056), .ZN(n13072) );
  XNOR2_X1 U11229 ( .A(n14928), .B(n15057), .ZN(n15305) );
  XNOR2_X1 U11230 ( .A(n15326), .B(n15124), .ZN(n15318) );
  INV_X1 U11231 ( .A(n15318), .ZN(n9559) );
  XNOR2_X1 U11232 ( .A(n15484), .B(n15126), .ZN(n15359) );
  INV_X1 U11233 ( .A(n15129), .ZN(n15402) );
  XNOR2_X1 U11234 ( .A(n15508), .B(n15402), .ZN(n12959) );
  INV_X1 U11235 ( .A(n15130), .ZN(n12957) );
  XNOR2_X1 U11236 ( .A(n16550), .B(n12957), .ZN(n15397) );
  XNOR2_X1 U11237 ( .A(n16529), .B(n15131), .ZN(n12715) );
  INV_X1 U11238 ( .A(n12715), .ZN(n12716) );
  XNOR2_X1 U11239 ( .A(n16523), .B(n15132), .ZN(n12582) );
  XNOR2_X1 U11240 ( .A(n12642), .B(n12640), .ZN(n12452) );
  XNOR2_X1 U11241 ( .A(n16388), .B(n12365), .ZN(n12262) );
  XNOR2_X1 U11242 ( .A(n12186), .B(n15137), .ZN(n12189) );
  INV_X1 U11243 ( .A(n12189), .ZN(n12182) );
  XNOR2_X1 U11244 ( .A(n12071), .B(n15138), .ZN(n12074) );
  XNOR2_X1 U11245 ( .A(n16314), .B(n11823), .ZN(n11587) );
  NAND2_X1 U11246 ( .A1(n16242), .A2(n15141), .ZN(n9546) );
  NAND2_X1 U11247 ( .A1(n11573), .A2(n14985), .ZN(n11584) );
  AND2_X2 U11248 ( .A1(n9546), .A2(n11584), .ZN(n12042) );
  NAND2_X1 U11249 ( .A1(n15143), .A2(n16155), .ZN(n9547) );
  INV_X1 U11250 ( .A(n16139), .ZN(n16144) );
  NAND2_X1 U11251 ( .A1(n11565), .A2(n16142), .ZN(n9548) );
  NAND2_X1 U11252 ( .A1(n16143), .A2(n9548), .ZN(n16094) );
  INV_X1 U11253 ( .A(n16094), .ZN(n16088) );
  NAND4_X1 U11254 ( .A1(n12042), .A2(n16144), .A3(n16088), .A4(n11793), .ZN(
        n9550) );
  NOR2_X1 U11255 ( .A1(n11587), .A2(n9550), .ZN(n9551) );
  XNOR2_X1 U11256 ( .A(n11838), .B(n15139), .ZN(n11955) );
  NAND4_X1 U11257 ( .A1(n12074), .A2(n9551), .A3(n11955), .A4(n9106), .ZN(
        n9552) );
  OR4_X1 U11258 ( .A1(n12339), .A2(n12262), .A3(n12182), .A4(n9552), .ZN(n9553) );
  NOR2_X1 U11259 ( .A1(n12452), .A2(n9553), .ZN(n9554) );
  XNOR2_X1 U11260 ( .A(n16493), .B(n15133), .ZN(n12687) );
  XNOR2_X1 U11261 ( .A(n16482), .B(n15134), .ZN(n12575) );
  NAND4_X1 U11262 ( .A1(n12582), .A2(n9554), .A3(n12687), .A4(n12575), .ZN(
        n9555) );
  OR3_X1 U11263 ( .A1(n15397), .A2(n12716), .A3(n9555), .ZN(n9556) );
  NOR2_X1 U11264 ( .A1(n12959), .A2(n9556), .ZN(n9557) );
  XNOR2_X1 U11265 ( .A(n15370), .B(n15088), .ZN(n13067) );
  INV_X1 U11266 ( .A(n13067), .ZN(n15364) );
  AND4_X1 U11267 ( .A1(n15359), .A2(n9557), .A3(n15364), .A4(n15378), .ZN(
        n9558) );
  XNOR2_X1 U11268 ( .A(n15334), .B(n15125), .ZN(n15330) );
  NAND3_X1 U11269 ( .A1(n9559), .A2(n9558), .A3(n15330), .ZN(n9560) );
  NOR2_X1 U11270 ( .A1(n15305), .A2(n9560), .ZN(n9561) );
  AND3_X1 U11271 ( .A1(n7380), .A2(n9561), .A3(n7644), .ZN(n9562) );
  XNOR2_X1 U11272 ( .A(n13075), .B(n15118), .ZN(n13074) );
  NAND4_X1 U11273 ( .A1(n9563), .A2(n9562), .A3(n13074), .A4(n13344), .ZN(
        n9564) );
  XNOR2_X1 U11274 ( .A(n15274), .B(n15120), .ZN(n13073) );
  NOR2_X1 U11275 ( .A1(n9564), .A2(n7726), .ZN(n9566) );
  NAND3_X1 U11276 ( .A1(n9567), .A2(n9566), .A3(n15262), .ZN(n9568) );
  XNOR2_X1 U11277 ( .A(n9568), .B(n7363), .ZN(n9589) );
  INV_X1 U11278 ( .A(n9569), .ZN(n9572) );
  NAND4_X1 U11279 ( .A1(n9572), .A2(n9571), .A3(n9570), .A4(n9581), .ZN(n9586)
         );
  NAND3_X1 U11280 ( .A1(n9574), .A2(n15238), .A3(n9581), .ZN(n9573) );
  OAI21_X1 U11281 ( .B1(n9581), .B2(n9574), .A(n9573), .ZN(n9576) );
  INV_X1 U11282 ( .A(n9588), .ZN(n9575) );
  AOI21_X1 U11283 ( .B1(n15415), .B2(n9576), .A(n9575), .ZN(n9585) );
  INV_X1 U11284 ( .A(n9577), .ZN(n9580) );
  NAND3_X1 U11285 ( .A1(n9580), .A2(n9578), .A3(n9581), .ZN(n9579) );
  OAI21_X1 U11286 ( .B1(n9581), .B2(n9580), .A(n9579), .ZN(n9582) );
  NAND2_X1 U11287 ( .A1(n9583), .A2(n9582), .ZN(n9584) );
  NAND3_X1 U11288 ( .A1(n9586), .A2(n9585), .A3(n9584), .ZN(n9587) );
  OAI21_X1 U11289 ( .B1(n9589), .B2(n9588), .A(n9587), .ZN(n9590) );
  XNOR2_X1 U11290 ( .A(n9597), .B(n9599), .ZN(n9609) );
  INV_X1 U11291 ( .A(n9609), .ZN(n11004) );
  NAND2_X1 U11292 ( .A1(n11004), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13013) );
  INV_X1 U11293 ( .A(n11005), .ZN(n11063) );
  INV_X1 U11294 ( .A(n9598), .ZN(n11285) );
  INV_X1 U11295 ( .A(n15689), .ZN(n11296) );
  NAND2_X1 U11296 ( .A1(n9600), .A2(n9599), .ZN(n9606) );
  INV_X1 U11297 ( .A(n9606), .ZN(n9601) );
  NAND2_X1 U11298 ( .A1(n9601), .A2(n9006), .ZN(n9604) );
  NAND2_X1 U11299 ( .A1(n9604), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9605) );
  XNOR2_X1 U11300 ( .A(n9605), .B(P1_IR_REG_25__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U11301 ( .A1(n9606), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9607) );
  NAND2_X1 U11302 ( .A1(n10992), .A2(n11056), .ZN(n9608) );
  AND2_X1 U11303 ( .A1(n12770), .A2(n12559), .ZN(n9610) );
  NAND4_X1 U11304 ( .A1(n15100), .A2(n11296), .A3(n11555), .A4(n11554), .ZN(
        n9611) );
  OAI211_X1 U11305 ( .C1(n15559), .C2(n13013), .A(n9611), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9612) );
  NOR2_X1 U11306 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9730) );
  NAND2_X1 U11307 ( .A1(n9730), .A2(n13745), .ZN(n9744) );
  NOR2_X2 U11308 ( .A1(n9819), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9833) );
  INV_X1 U11309 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n13556) );
  INV_X1 U11310 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n13541) );
  NAND2_X1 U11311 ( .A1(n9984), .A2(n13541), .ZN(n9998) );
  INV_X1 U11312 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13664) );
  NOR2_X1 U11313 ( .A1(n10011), .A2(n13664), .ZN(n9613) );
  OR2_X2 U11314 ( .A1(n13961), .A2(n9613), .ZN(n13981) );
  MUX2_X1 U11315 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9615), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n9619) );
  INV_X1 U11316 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9616) );
  XNOR2_X2 U11317 ( .A(n9620), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U11318 ( .A1(n13981), .A2(n10035), .ZN(n9628) );
  INV_X1 U11319 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9625) );
  INV_X1 U11320 ( .A(n9621), .ZN(n13356) );
  NAND2_X1 U11321 ( .A1(n10036), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U11322 ( .A1(n10048), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9623) );
  OAI211_X1 U11323 ( .C1(n9625), .C2(n11987), .A(n9624), .B(n9623), .ZN(n9626)
         );
  INV_X1 U11324 ( .A(n9626), .ZN(n9627) );
  INV_X1 U11325 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14820) );
  AOI22_X1 U11326 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n9665), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n13015), .ZN(n9957) );
  XNOR2_X1 U11327 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9825) );
  INV_X1 U11328 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U11329 ( .A1(n10987), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U11330 ( .A1(n9681), .A2(n9630), .ZN(n9699) );
  XNOR2_X1 U11331 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9697) );
  NAND2_X1 U11332 ( .A1(n10989), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9631) );
  INV_X1 U11333 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U11334 ( .A1(n9724), .A2(n9722), .ZN(n9634) );
  NAND2_X1 U11335 ( .A1(n11016), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U11336 ( .A1(n9634), .A2(n9633), .ZN(n9738) );
  NAND2_X1 U11337 ( .A1(n9738), .A2(n9736), .ZN(n9636) );
  NAND2_X1 U11338 ( .A1(n11002), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U11339 ( .A1(n9636), .A2(n9635), .ZN(n9752) );
  NAND2_X1 U11340 ( .A1(n11012), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U11341 ( .A1(n9763), .A2(n9762), .ZN(n9640) );
  NAND2_X1 U11342 ( .A1(n11013), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U11343 ( .A1(n11132), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U11344 ( .A1(n9643), .A2(n9642), .ZN(n9802) );
  XNOR2_X1 U11345 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9801) );
  NAND2_X1 U11346 ( .A1(n9644), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9645) );
  XNOR2_X1 U11347 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9813) );
  XNOR2_X1 U11348 ( .A(n9648), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U11349 ( .A1(n9830), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U11350 ( .A1(n11401), .A2(n9648), .ZN(n9649) );
  NAND2_X1 U11351 ( .A1(n9650), .A2(n9649), .ZN(n9843) );
  XNOR2_X1 U11352 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9842) );
  NAND2_X1 U11353 ( .A1(n9843), .A2(n9842), .ZN(n9653) );
  INV_X1 U11354 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U11355 ( .A1(n9651), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9652) );
  XNOR2_X1 U11356 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9854) );
  NAND2_X1 U11357 ( .A1(n9856), .A2(n9854), .ZN(n9654) );
  INV_X1 U11358 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U11359 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n12024), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n12023), .ZN(n9865) );
  AOI22_X1 U11360 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n12180), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9656), .ZN(n9880) );
  INV_X1 U11361 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U11362 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n12338), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n12336), .ZN(n9893) );
  NAND2_X1 U11363 ( .A1(n9895), .A2(n9893), .ZN(n9658) );
  INV_X1 U11364 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U11365 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n12558), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n12561), .ZN(n9906) );
  NAND2_X1 U11366 ( .A1(n9907), .A2(n9906), .ZN(n9660) );
  AOI22_X1 U11367 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n12740), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n12771), .ZN(n9918) );
  NAND2_X1 U11368 ( .A1(n9920), .A2(n9918), .ZN(n9662) );
  INV_X1 U11369 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12879) );
  NAND2_X1 U11370 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n12879), .ZN(n9663) );
  INV_X1 U11371 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U11372 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n12988), .B2(n9664), .ZN(n9944) );
  INV_X1 U11373 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14816) );
  AOI22_X1 U11374 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n14816), .B2(n15553), .ZN(n9980) );
  INV_X1 U11375 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14812) );
  AOI22_X1 U11376 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n14812), .B2(n15548), .ZN(n9992) );
  INV_X1 U11377 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14810) );
  AOI22_X1 U11378 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n14810), .B2(n13087), .ZN(n10006) );
  INV_X1 U11379 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14807) );
  AOI22_X1 U11380 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n14807), .B2(n13093), .ZN(n10027) );
  INV_X1 U11381 ( .A(n10027), .ZN(n9673) );
  XNOR2_X1 U11382 ( .A(n10026), .B(n9673), .ZN(n13119) );
  NAND2_X1 U11383 ( .A1(n13119), .A2(n10032), .ZN(n9675) );
  NAND2_X1 U11384 ( .A1(n13279), .A2(SI_28_), .ZN(n9674) );
  NAND2_X2 U11385 ( .A1(n9675), .A2(n9674), .ZN(n10022) );
  NAND2_X1 U11386 ( .A1(n7367), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U11387 ( .A1(n9746), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U11388 ( .A1(n9729), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U11389 ( .A1(n9692), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9676) );
  OAI21_X1 U11390 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n10966) );
  NAND2_X1 U11391 ( .A1(n9739), .A2(n10966), .ZN(n9685) );
  OAI211_X1 U11392 ( .C1(n9721), .C2(n7839), .A(n9685), .B(n9684), .ZN(n10121)
         );
  INV_X1 U11393 ( .A(n10121), .ZN(n16130) );
  NAND2_X1 U11394 ( .A1(n9729), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U11395 ( .A1(n7367), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U11396 ( .A1(n9692), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9687) );
  NAND2_X1 U11397 ( .A1(n9746), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9686) );
  XNOR2_X1 U11398 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .ZN(n9690) );
  MUX2_X1 U11399 ( .A(n9690), .B(n13718), .S(n10984), .Z(n10961) );
  MUX2_X1 U11400 ( .A(n10960), .B(n10961), .S(n10054), .Z(n11928) );
  INV_X1 U11401 ( .A(n11928), .ZN(n11883) );
  AND2_X1 U11402 ( .A1(n13893), .A2(n11883), .ZN(n9691) );
  NAND2_X1 U11403 ( .A1(n10122), .A2(n16130), .ZN(n16181) );
  NAND2_X1 U11404 ( .A1(n11983), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U11405 ( .A1(n9746), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U11406 ( .A1(n9692), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9693) );
  AND4_X2 U11407 ( .A1(n9696), .A2(n9695), .A3(n9694), .A4(n9693), .ZN(n12118)
         );
  INV_X1 U11408 ( .A(n12118), .ZN(n11310) );
  INV_X1 U11409 ( .A(n9697), .ZN(n9698) );
  XNOR2_X1 U11410 ( .A(n9699), .B(n9698), .ZN(n10970) );
  NAND2_X1 U11411 ( .A1(n9739), .A2(n10970), .ZN(n9701) );
  NAND2_X1 U11412 ( .A1(n9908), .A2(n7370), .ZN(n9700) );
  INV_X1 U11413 ( .A(n11645), .ZN(n16196) );
  NAND2_X1 U11414 ( .A1(n11310), .A2(n16196), .ZN(n13145) );
  NAND2_X1 U11415 ( .A1(n12118), .A2(n11645), .ZN(n13146) );
  NAND2_X1 U11416 ( .A1(n9703), .A2(n16177), .ZN(n12121) );
  INV_X1 U11417 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n13734) );
  NAND2_X1 U11418 ( .A1(n10035), .A2(n13734), .ZN(n9707) );
  NAND2_X1 U11419 ( .A1(n11983), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U11420 ( .A1(n9746), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U11421 ( .A1(n7367), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9704) );
  AND4_X2 U11422 ( .A1(n9707), .A2(n9706), .A3(n9705), .A4(n9704), .ZN(n12136)
         );
  INV_X1 U11423 ( .A(SI_3_), .ZN(n13715) );
  NAND2_X1 U11424 ( .A1(n13279), .A2(n13715), .ZN(n9713) );
  INV_X1 U11425 ( .A(n9708), .ZN(n9709) );
  XNOR2_X1 U11426 ( .A(n9710), .B(n9709), .ZN(n10964) );
  NAND2_X1 U11427 ( .A1(n9739), .A2(n10964), .ZN(n9712) );
  NAND2_X1 U11428 ( .A1(n9908), .A2(n10965), .ZN(n9711) );
  NAND2_X1 U11429 ( .A1(n12136), .A2(n12128), .ZN(n13153) );
  NAND2_X1 U11430 ( .A1(n16179), .A2(n16234), .ZN(n13154) );
  AND2_X1 U11431 ( .A1(n12118), .A2(n16196), .ZN(n12122) );
  NAND2_X1 U11432 ( .A1(n12121), .A2(n9714), .ZN(n12123) );
  NAND2_X1 U11433 ( .A1(n16179), .A2(n12128), .ZN(n9715) );
  NAND2_X1 U11434 ( .A1(n12123), .A2(n9715), .ZN(n12134) );
  NAND2_X1 U11435 ( .A1(n11983), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U11436 ( .A1(n7367), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9719) );
  AND2_X1 U11437 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9716) );
  OR2_X1 U11438 ( .A1(n9716), .A2(n9730), .ZN(n12140) );
  NAND2_X1 U11439 ( .A1(n10035), .A2(n12140), .ZN(n9718) );
  NAND2_X1 U11440 ( .A1(n10048), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9717) );
  AND4_X2 U11441 ( .A1(n9720), .A2(n9719), .A3(n9718), .A4(n9717), .ZN(n12119)
         );
  NAND2_X1 U11442 ( .A1(n9995), .A2(n7656), .ZN(n9727) );
  INV_X1 U11443 ( .A(n9722), .ZN(n9723) );
  XNOR2_X1 U11444 ( .A(n9724), .B(n9723), .ZN(n10974) );
  NAND2_X1 U11445 ( .A1(n9739), .A2(n10974), .ZN(n9726) );
  NAND2_X1 U11446 ( .A1(n9908), .A2(n15932), .ZN(n9725) );
  NAND2_X1 U11447 ( .A1(n12119), .A2(n12141), .ZN(n13157) );
  INV_X1 U11448 ( .A(n12119), .ZN(n13475) );
  INV_X1 U11449 ( .A(n12141), .ZN(n16278) );
  NAND2_X1 U11450 ( .A1(n13475), .A2(n16278), .ZN(n13158) );
  INV_X1 U11451 ( .A(n13306), .ZN(n12133) );
  NAND2_X1 U11452 ( .A1(n13475), .A2(n12141), .ZN(n9728) );
  NAND2_X1 U11453 ( .A1(n9729), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9735) );
  NAND2_X1 U11454 ( .A1(n9746), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9734) );
  OR2_X1 U11455 ( .A1(n13745), .A2(n9730), .ZN(n9731) );
  NAND2_X1 U11456 ( .A1(n9744), .A2(n9731), .ZN(n12332) );
  NAND2_X1 U11457 ( .A1(n10035), .A2(n12332), .ZN(n9733) );
  NAND2_X1 U11458 ( .A1(n7367), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9732) );
  INV_X1 U11459 ( .A(SI_5_), .ZN(n13666) );
  NAND2_X1 U11460 ( .A1(n13279), .A2(n13666), .ZN(n9742) );
  INV_X1 U11461 ( .A(n9736), .ZN(n9737) );
  XNOR2_X1 U11462 ( .A(n9738), .B(n9737), .ZN(n10968) );
  NAND2_X1 U11463 ( .A1(n9739), .A2(n10968), .ZN(n9741) );
  NAND2_X1 U11464 ( .A1(n9908), .A2(n15952), .ZN(n9740) );
  NAND2_X1 U11465 ( .A1(n12293), .A2(n12333), .ZN(n13162) );
  INV_X1 U11466 ( .A(n12293), .ZN(n13474) );
  INV_X1 U11467 ( .A(n12333), .ZN(n16305) );
  NAND2_X1 U11468 ( .A1(n13474), .A2(n16305), .ZN(n13161) );
  AND2_X2 U11469 ( .A1(n13162), .A2(n13161), .ZN(n13302) );
  NAND2_X1 U11470 ( .A1(n7367), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U11471 ( .A1(n11983), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U11472 ( .A1(n9744), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U11473 ( .A1(n9756), .A2(n9745), .ZN(n12301) );
  NAND2_X1 U11474 ( .A1(n10035), .A2(n12301), .ZN(n9748) );
  NAND2_X1 U11475 ( .A1(n9746), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9747) );
  NAND4_X2 U11476 ( .A1(n9750), .A2(n9749), .A3(n9748), .A4(n9747), .ZN(n13472) );
  XNOR2_X1 U11477 ( .A(n11010), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9751) );
  XNOR2_X1 U11478 ( .A(n9752), .B(n9751), .ZN(n10972) );
  NAND2_X1 U11479 ( .A1(n13279), .A2(SI_6_), .ZN(n9754) );
  NAND2_X1 U11480 ( .A1(n9908), .A2(n15978), .ZN(n9753) );
  AND2_X1 U11481 ( .A1(n12293), .A2(n16305), .ZN(n12288) );
  NOR2_X1 U11482 ( .A1(n13164), .A2(n12288), .ZN(n9755) );
  NAND2_X1 U11483 ( .A1(n13472), .A2(n16333), .ZN(n13167) );
  NAND2_X1 U11484 ( .A1(n11983), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U11485 ( .A1(n10048), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9760) );
  AND2_X1 U11486 ( .A1(n9756), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9757) );
  OR2_X1 U11487 ( .A1(n9757), .A2(n9769), .ZN(n12448) );
  NAND2_X1 U11488 ( .A1(n10035), .A2(n12448), .ZN(n9759) );
  NAND2_X1 U11489 ( .A1(n7367), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9758) );
  INV_X1 U11490 ( .A(SI_7_), .ZN(n13711) );
  NAND2_X1 U11491 ( .A1(n9777), .A2(n13711), .ZN(n9766) );
  XNOR2_X1 U11492 ( .A(n9763), .B(n9762), .ZN(n10963) );
  NAND2_X1 U11493 ( .A1(n10032), .A2(n10963), .ZN(n9765) );
  NAND2_X1 U11494 ( .A1(n9908), .A2(n15992), .ZN(n9764) );
  NAND2_X1 U11495 ( .A1(n12294), .A2(n12449), .ZN(n13171) );
  INV_X1 U11496 ( .A(n12294), .ZN(n13470) );
  INV_X1 U11497 ( .A(n12449), .ZN(n16345) );
  NAND2_X1 U11498 ( .A1(n13470), .A2(n16345), .ZN(n13170) );
  NAND2_X1 U11499 ( .A1(n13171), .A2(n13170), .ZN(n13305) );
  NAND2_X1 U11500 ( .A1(n12442), .A2(n13305), .ZN(n9768) );
  NAND2_X1 U11501 ( .A1(n13470), .A2(n12449), .ZN(n9767) );
  NAND2_X1 U11502 ( .A1(n11983), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9774) );
  NAND2_X1 U11503 ( .A1(n10048), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9773) );
  NOR2_X1 U11504 ( .A1(n9769), .A2(n13737), .ZN(n9770) );
  OR2_X1 U11505 ( .A1(n9783), .A2(n9770), .ZN(n12415) );
  NAND2_X1 U11506 ( .A1(n10035), .A2(n12415), .ZN(n9772) );
  NAND2_X1 U11507 ( .A1(n7367), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9771) );
  XNOR2_X1 U11508 ( .A(n9776), .B(n9775), .ZN(n10975) );
  NAND2_X1 U11509 ( .A1(n9777), .A2(SI_8_), .ZN(n9780) );
  NAND2_X1 U11510 ( .A1(n9908), .A2(n9778), .ZN(n9779) );
  OAI211_X1 U11511 ( .C1(n9781), .C2(n10975), .A(n9780), .B(n9779), .ZN(n12416) );
  NAND2_X1 U11512 ( .A1(n12588), .A2(n12416), .ZN(n13175) );
  INV_X1 U11513 ( .A(n12588), .ZN(n13469) );
  INV_X1 U11514 ( .A(n12416), .ZN(n16368) );
  NAND2_X1 U11515 ( .A1(n13469), .A2(n16368), .ZN(n13176) );
  NAND2_X1 U11516 ( .A1(n12588), .A2(n16368), .ZN(n9782) );
  NAND2_X1 U11517 ( .A1(n7367), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U11518 ( .A1(n11983), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9787) );
  OR2_X1 U11519 ( .A1(n9783), .A2(n13551), .ZN(n9784) );
  NAND2_X1 U11520 ( .A1(n9795), .A2(n9784), .ZN(n12593) );
  NAND2_X1 U11521 ( .A1(n10035), .A2(n12593), .ZN(n9786) );
  INV_X4 U11522 ( .A(n9964), .ZN(n10048) );
  NAND2_X1 U11523 ( .A1(n10048), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9785) );
  XNOR2_X1 U11524 ( .A(n9790), .B(n9789), .ZN(n10977) );
  NAND2_X1 U11525 ( .A1(n10032), .A2(n10977), .ZN(n9793) );
  NAND2_X1 U11526 ( .A1(n13279), .A2(n13506), .ZN(n9792) );
  NAND2_X1 U11527 ( .A1(n9908), .A2(n16032), .ZN(n9791) );
  NAND2_X1 U11528 ( .A1(n13468), .A2(n16381), .ZN(n9794) );
  INV_X1 U11529 ( .A(n16381), .ZN(n10071) );
  NAND2_X1 U11530 ( .A1(n7367), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U11531 ( .A1(n11983), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U11532 ( .A1(n9795), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9796) );
  NAND2_X1 U11533 ( .A1(n9807), .A2(n9796), .ZN(n12598) );
  NAND2_X1 U11534 ( .A1(n10035), .A2(n12598), .ZN(n9798) );
  NAND2_X1 U11535 ( .A1(n10048), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9797) );
  XNOR2_X1 U11536 ( .A(n9802), .B(n9801), .ZN(n10982) );
  NAND2_X1 U11537 ( .A1(n10032), .A2(n10982), .ZN(n9805) );
  INV_X1 U11538 ( .A(SI_10_), .ZN(n13702) );
  NAND2_X1 U11539 ( .A1(n13279), .A2(n13702), .ZN(n9804) );
  NAND2_X1 U11540 ( .A1(n9908), .A2(n12547), .ZN(n9803) );
  NAND2_X1 U11541 ( .A1(n12696), .A2(n16411), .ZN(n13184) );
  INV_X1 U11542 ( .A(n12696), .ZN(n13467) );
  INV_X1 U11543 ( .A(n16411), .ZN(n12763) );
  NAND2_X1 U11544 ( .A1(n13467), .A2(n12763), .ZN(n13192) );
  NAND2_X1 U11545 ( .A1(n12760), .A2(n12759), .ZN(n12758) );
  NAND2_X1 U11546 ( .A1(n13467), .A2(n16411), .ZN(n9806) );
  NAND2_X1 U11547 ( .A1(n12758), .A2(n9806), .ZN(n12992) );
  NAND2_X1 U11548 ( .A1(n7367), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9812) );
  NAND2_X1 U11549 ( .A1(n11983), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U11550 ( .A1(n9807), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9808) );
  NAND2_X1 U11551 ( .A1(n9819), .A2(n9808), .ZN(n12692) );
  NAND2_X1 U11552 ( .A1(n10035), .A2(n12692), .ZN(n9810) );
  NAND2_X1 U11553 ( .A1(n10048), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9809) );
  XNOR2_X1 U11554 ( .A(n9814), .B(n9813), .ZN(n10991) );
  NAND2_X1 U11555 ( .A1(n10032), .A2(n10991), .ZN(n9817) );
  NAND2_X1 U11556 ( .A1(n13279), .A2(n13698), .ZN(n9816) );
  NAND2_X1 U11557 ( .A1(n9908), .A2(n12238), .ZN(n9815) );
  NAND2_X1 U11558 ( .A1(n12780), .A2(n16441), .ZN(n10153) );
  NAND2_X1 U11559 ( .A1(n12992), .A2(n10153), .ZN(n9818) );
  OR2_X1 U11560 ( .A1(n12780), .A2(n16441), .ZN(n10155) );
  NAND2_X1 U11561 ( .A1(n11983), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U11562 ( .A1(n7367), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9823) );
  AND2_X1 U11563 ( .A1(n9819), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9820) );
  OR2_X1 U11564 ( .A1(n9820), .A2(n9833), .ZN(n12920) );
  NAND2_X1 U11565 ( .A1(n10035), .A2(n12920), .ZN(n9822) );
  NAND2_X1 U11566 ( .A1(n10048), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9821) );
  XNOR2_X1 U11567 ( .A(n9826), .B(n9825), .ZN(n11003) );
  NAND2_X1 U11568 ( .A1(n10032), .A2(n11003), .ZN(n9829) );
  NAND2_X1 U11569 ( .A1(n13279), .A2(n13699), .ZN(n9828) );
  NAND2_X1 U11570 ( .A1(n9908), .A2(n12524), .ZN(n9827) );
  NOR2_X1 U11571 ( .A1(n12928), .A2(n16468), .ZN(n10159) );
  NAND2_X1 U11572 ( .A1(n12928), .A2(n16468), .ZN(n10160) );
  XNOR2_X1 U11573 ( .A(n9830), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U11574 ( .A1(n11018), .A2(n10032), .ZN(n9832) );
  INV_X1 U11575 ( .A(SI_13_), .ZN(n13695) );
  AOI22_X1 U11576 ( .A1(n9995), .A2(n13695), .B1(n9908), .B2(n11019), .ZN(
        n9831) );
  NAND2_X1 U11577 ( .A1(n9832), .A2(n9831), .ZN(n14238) );
  NAND2_X1 U11578 ( .A1(n7367), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U11579 ( .A1(n11983), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9837) );
  OR2_X1 U11580 ( .A1(n9833), .A2(n13555), .ZN(n9834) );
  NAND2_X1 U11581 ( .A1(n9846), .A2(n9834), .ZN(n13020) );
  NAND2_X1 U11582 ( .A1(n10035), .A2(n13020), .ZN(n9836) );
  NAND2_X1 U11583 ( .A1(n10048), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9835) );
  NAND4_X1 U11584 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(n13026) );
  INV_X1 U11585 ( .A(n13026), .ZN(n9840) );
  AND2_X1 U11586 ( .A1(n14238), .A2(n9840), .ZN(n9839) );
  OR2_X1 U11587 ( .A1(n14238), .A2(n9840), .ZN(n10161) );
  XNOR2_X1 U11588 ( .A(n9843), .B(n9842), .ZN(n11033) );
  NAND2_X1 U11589 ( .A1(n11033), .A2(n10032), .ZN(n9845) );
  AOI22_X1 U11590 ( .A1(n9995), .A2(n11032), .B1(n9908), .B2(n11031), .ZN(
        n9844) );
  NAND2_X1 U11591 ( .A1(n7367), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U11592 ( .A1(n11983), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U11593 ( .A1(n9846), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9847) );
  NAND2_X1 U11594 ( .A1(n9859), .A2(n9847), .ZN(n13029) );
  NAND2_X1 U11595 ( .A1(n10035), .A2(n13029), .ZN(n9849) );
  NAND2_X1 U11596 ( .A1(n10048), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9848) );
  XNOR2_X1 U11597 ( .A(n14236), .B(n14160), .ZN(n13320) );
  INV_X1 U11598 ( .A(n13320), .ZN(n9852) );
  OR2_X1 U11599 ( .A1(n14236), .A2(n14160), .ZN(n9853) );
  INV_X1 U11600 ( .A(n9854), .ZN(n9855) );
  XNOR2_X1 U11601 ( .A(n9856), .B(n9855), .ZN(n11074) );
  NAND2_X1 U11602 ( .A1(n11074), .A2(n10032), .ZN(n9858) );
  AOI22_X1 U11603 ( .A1(n9995), .A2(SI_15_), .B1(n9908), .B2(n11075), .ZN(
        n9857) );
  NAND2_X1 U11604 ( .A1(n9858), .A2(n9857), .ZN(n14229) );
  NAND2_X1 U11605 ( .A1(n7367), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U11606 ( .A1(n11983), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9863) );
  AND2_X1 U11607 ( .A1(n9859), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9860) );
  OR2_X1 U11608 ( .A1(n9860), .A2(n9871), .ZN(n14162) );
  NAND2_X1 U11609 ( .A1(n10035), .A2(n14162), .ZN(n9862) );
  NAND2_X1 U11610 ( .A1(n10048), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9861) );
  OR2_X1 U11611 ( .A1(n14229), .A2(n14146), .ZN(n13211) );
  NAND2_X1 U11612 ( .A1(n14229), .A2(n14146), .ZN(n13210) );
  NAND2_X1 U11613 ( .A1(n13211), .A2(n13210), .ZN(n14154) );
  INV_X1 U11614 ( .A(n14143), .ZN(n9878) );
  INV_X1 U11615 ( .A(n9865), .ZN(n9866) );
  XNOR2_X1 U11616 ( .A(n9867), .B(n9866), .ZN(n11135) );
  NAND2_X1 U11617 ( .A1(n11135), .A2(n10032), .ZN(n9869) );
  AOI22_X1 U11618 ( .A1(n9995), .A2(SI_16_), .B1(n9908), .B2(n16042), .ZN(
        n9868) );
  NAND2_X1 U11619 ( .A1(n9869), .A2(n9868), .ZN(n13216) );
  NAND2_X1 U11620 ( .A1(n11983), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U11621 ( .A1(n7367), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9875) );
  NOR2_X1 U11622 ( .A1(n9871), .A2(n9870), .ZN(n9872) );
  OR2_X1 U11623 ( .A1(n9886), .A2(n9872), .ZN(n14148) );
  NAND2_X1 U11624 ( .A1(n10035), .A2(n14148), .ZN(n9874) );
  NAND2_X1 U11625 ( .A1(n10048), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9873) );
  NAND4_X1 U11626 ( .A1(n9876), .A2(n9875), .A3(n9874), .A4(n9873), .ZN(n14131) );
  XNOR2_X1 U11627 ( .A(n13216), .B(n14131), .ZN(n14144) );
  OR2_X1 U11628 ( .A1(n13216), .A2(n14131), .ZN(n9879) );
  INV_X1 U11629 ( .A(n9880), .ZN(n9881) );
  XNOR2_X1 U11630 ( .A(n9882), .B(n9881), .ZN(n11228) );
  NAND2_X1 U11631 ( .A1(n11228), .A2(n10032), .ZN(n9885) );
  AOI22_X1 U11632 ( .A1(n9995), .A2(SI_17_), .B1(n9908), .B2(n9883), .ZN(n9884) );
  NAND2_X1 U11633 ( .A1(n7367), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U11634 ( .A1(n11983), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9890) );
  OR2_X1 U11635 ( .A1(n9886), .A2(n13748), .ZN(n9887) );
  NAND2_X1 U11636 ( .A1(n9899), .A2(n9887), .ZN(n14135) );
  NAND2_X1 U11637 ( .A1(n10035), .A2(n14135), .ZN(n9889) );
  NAND2_X1 U11638 ( .A1(n10048), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9888) );
  NOR2_X1 U11639 ( .A1(n14220), .A2(n14147), .ZN(n13130) );
  INV_X1 U11640 ( .A(n13130), .ZN(n9892) );
  INV_X1 U11641 ( .A(n9893), .ZN(n9894) );
  XNOR2_X1 U11642 ( .A(n9895), .B(n9894), .ZN(n11373) );
  NAND2_X1 U11643 ( .A1(n11373), .A2(n10032), .ZN(n9898) );
  AOI22_X1 U11644 ( .A1(n9995), .A2(SI_18_), .B1(n9908), .B2(n9896), .ZN(n9897) );
  NAND2_X1 U11645 ( .A1(n9898), .A2(n9897), .ZN(n13436) );
  NAND2_X1 U11646 ( .A1(n7367), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U11647 ( .A1(n10036), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9903) );
  NAND2_X1 U11648 ( .A1(n9899), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U11649 ( .A1(n9911), .A2(n9900), .ZN(n14123) );
  NAND2_X1 U11650 ( .A1(n10035), .A2(n14123), .ZN(n9902) );
  NAND2_X1 U11651 ( .A1(n10048), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9901) );
  OR2_X1 U11652 ( .A1(n13436), .A2(n14108), .ZN(n13132) );
  INV_X1 U11653 ( .A(n14147), .ZN(n13397) );
  AND2_X1 U11654 ( .A1(n14220), .A2(n13397), .ZN(n14117) );
  NOR2_X1 U11655 ( .A1(n14116), .A2(n14117), .ZN(n9905) );
  OR2_X1 U11656 ( .A1(n13436), .A2(n14132), .ZN(n14104) );
  XNOR2_X1 U11657 ( .A(n9907), .B(n9906), .ZN(n11450) );
  NAND2_X1 U11658 ( .A1(n11450), .A2(n10032), .ZN(n9910) );
  AOI22_X1 U11659 ( .A1(n9995), .A2(n11451), .B1(n9908), .B2(n11452), .ZN(
        n9909) );
  NAND2_X1 U11660 ( .A1(n7367), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U11661 ( .A1(n10036), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9915) );
  AND2_X1 U11662 ( .A1(n9911), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9912) );
  OR2_X1 U11663 ( .A1(n9912), .A2(n9923), .ZN(n14110) );
  NAND2_X1 U11664 ( .A1(n10035), .A2(n14110), .ZN(n9914) );
  NAND2_X1 U11665 ( .A1(n10048), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U11666 ( .A1(n14287), .A2(n14122), .ZN(n9917) );
  AND2_X1 U11667 ( .A1(n14104), .A2(n9917), .ZN(n14083) );
  INV_X1 U11668 ( .A(n9918), .ZN(n9919) );
  XNOR2_X1 U11669 ( .A(n9920), .B(n9919), .ZN(n11772) );
  NAND2_X1 U11670 ( .A1(n11772), .A2(n10032), .ZN(n9922) );
  NAND2_X1 U11671 ( .A1(n9995), .A2(SI_20_), .ZN(n9921) );
  NAND2_X1 U11672 ( .A1(n7367), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9928) );
  NAND2_X1 U11673 ( .A1(n10036), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9927) );
  NOR2_X1 U11674 ( .A1(n9923), .A2(n13556), .ZN(n9924) );
  OR2_X1 U11675 ( .A1(n9937), .A2(n9924), .ZN(n14093) );
  NAND2_X1 U11676 ( .A1(n10035), .A2(n14093), .ZN(n9926) );
  NAND2_X1 U11677 ( .A1(n10048), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9925) );
  XNOR2_X1 U11678 ( .A(n14205), .B(n13464), .ZN(n14098) );
  INV_X1 U11679 ( .A(n14098), .ZN(n9929) );
  AND2_X1 U11680 ( .A1(n14083), .A2(n9929), .ZN(n9930) );
  NAND2_X1 U11681 ( .A1(n14119), .A2(n9930), .ZN(n14088) );
  NAND2_X1 U11682 ( .A1(n14205), .A2(n13464), .ZN(n9931) );
  NAND2_X1 U11683 ( .A1(n10175), .A2(n13442), .ZN(n14084) );
  OR2_X1 U11684 ( .A1(n14098), .A2(n14084), .ZN(n14087) );
  AND2_X1 U11685 ( .A1(n9931), .A2(n14087), .ZN(n9932) );
  NAND2_X1 U11686 ( .A1(n14088), .A2(n9932), .ZN(n14070) );
  AOI22_X1 U11687 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(
        P1_DATAO_REG_21__SCAN_IN), .B1(n12879), .B2(n12876), .ZN(n9933) );
  XNOR2_X1 U11688 ( .A(n7531), .B(n9933), .ZN(n11929) );
  NAND2_X1 U11689 ( .A1(n11929), .A2(n10032), .ZN(n9936) );
  NAND2_X1 U11690 ( .A1(n13279), .A2(SI_21_), .ZN(n9935) );
  OR2_X1 U11691 ( .A1(n9937), .A2(n13740), .ZN(n9938) );
  NAND2_X1 U11692 ( .A1(n9948), .A2(n9938), .ZN(n14079) );
  NAND2_X1 U11693 ( .A1(n14079), .A2(n10035), .ZN(n9942) );
  NAND2_X1 U11694 ( .A1(n7367), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9941) );
  NAND2_X1 U11695 ( .A1(n10036), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U11696 ( .A1(n10048), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9939) );
  OR2_X1 U11697 ( .A1(n14202), .A2(n14055), .ZN(n10186) );
  NAND2_X1 U11698 ( .A1(n14070), .A2(n10186), .ZN(n9943) );
  NAND2_X1 U11699 ( .A1(n14202), .A2(n14055), .ZN(n10183) );
  XNOR2_X1 U11700 ( .A(n9945), .B(n8026), .ZN(n11952) );
  NAND2_X1 U11701 ( .A1(n11952), .A2(n10032), .ZN(n9947) );
  NAND2_X1 U11702 ( .A1(n9995), .A2(SI_22_), .ZN(n9946) );
  NAND2_X1 U11703 ( .A1(n9948), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U11704 ( .A1(n9960), .A2(n9949), .ZN(n14063) );
  NAND2_X1 U11705 ( .A1(n14063), .A2(n10035), .ZN(n9954) );
  NAND2_X1 U11706 ( .A1(n7367), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U11707 ( .A1(n10036), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9950) );
  AND2_X1 U11708 ( .A1(n9951), .A2(n9950), .ZN(n9953) );
  NAND2_X1 U11709 ( .A1(n10048), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9952) );
  AND2_X1 U11710 ( .A1(n14199), .A2(n14041), .ZN(n9955) );
  XNOR2_X1 U11711 ( .A(n9957), .B(n9956), .ZN(n12147) );
  NAND2_X1 U11712 ( .A1(n12147), .A2(n10032), .ZN(n9959) );
  NAND2_X1 U11713 ( .A1(n9995), .A2(SI_23_), .ZN(n9958) );
  INV_X1 U11714 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14267) );
  NAND2_X1 U11715 ( .A1(n9960), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9961) );
  NAND2_X1 U11716 ( .A1(n9969), .A2(n9961), .ZN(n14045) );
  NAND2_X1 U11717 ( .A1(n14045), .A2(n10035), .ZN(n9963) );
  AOI22_X1 U11718 ( .A1(n7367), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n10036), 
        .B2(P3_REG1_REG_23__SCAN_IN), .ZN(n9962) );
  XNOR2_X1 U11719 ( .A(n13367), .B(n14056), .ZN(n14038) );
  NAND2_X1 U11720 ( .A1(n13367), .A2(n14056), .ZN(n9965) );
  XNOR2_X1 U11721 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9966), .ZN(n12535) );
  NAND2_X1 U11722 ( .A1(n12535), .A2(n10032), .ZN(n9968) );
  NAND2_X1 U11723 ( .A1(n13279), .A2(SI_24_), .ZN(n9967) );
  AND2_X1 U11724 ( .A1(n9969), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9970) );
  OR2_X1 U11725 ( .A1(n9970), .A2(n9984), .ZN(n14031) );
  NAND2_X1 U11726 ( .A1(n14031), .A2(n10035), .ZN(n9976) );
  INV_X1 U11727 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U11728 ( .A1(n10048), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9972) );
  NAND2_X1 U11729 ( .A1(n10036), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9971) );
  OAI211_X1 U11730 ( .C1(n11987), .C2(n9973), .A(n9972), .B(n9971), .ZN(n9974)
         );
  INV_X1 U11731 ( .A(n9974), .ZN(n9975) );
  NAND2_X1 U11732 ( .A1(n14265), .A2(n14042), .ZN(n13256) );
  INV_X1 U11733 ( .A(n14265), .ZN(n9977) );
  NAND2_X1 U11734 ( .A1(n9977), .A2(n14009), .ZN(n13253) );
  OR2_X2 U11735 ( .A1(n14025), .A2(n14030), .ZN(n14023) );
  NAND2_X1 U11736 ( .A1(n14265), .A2(n14009), .ZN(n9978) );
  XNOR2_X1 U11737 ( .A(n9981), .B(n9670), .ZN(n12634) );
  NAND2_X1 U11738 ( .A1(n12634), .A2(n10032), .ZN(n9983) );
  NAND2_X1 U11739 ( .A1(n13279), .A2(SI_25_), .ZN(n9982) );
  OR2_X1 U11740 ( .A1(n9984), .A2(n13541), .ZN(n9985) );
  NAND2_X1 U11741 ( .A1(n9998), .A2(n9985), .ZN(n14018) );
  NAND2_X1 U11742 ( .A1(n14018), .A2(n10035), .ZN(n9991) );
  INV_X1 U11743 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U11744 ( .A1(n10048), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U11745 ( .A1(n10036), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9986) );
  OAI211_X1 U11746 ( .C1(n11987), .C2(n9988), .A(n9987), .B(n9986), .ZN(n9989)
         );
  INV_X1 U11747 ( .A(n9989), .ZN(n9990) );
  XNOR2_X1 U11748 ( .A(n14260), .B(n13463), .ZN(n14014) );
  INV_X1 U11749 ( .A(n14014), .ZN(n14007) );
  NAND2_X1 U11750 ( .A1(n14260), .A2(n13463), .ZN(n13996) );
  INV_X1 U11751 ( .A(n9992), .ZN(n9993) );
  XNOR2_X1 U11752 ( .A(n9994), .B(n9993), .ZN(n12881) );
  NAND2_X1 U11753 ( .A1(n12881), .A2(n10032), .ZN(n9997) );
  NAND2_X1 U11754 ( .A1(n9995), .A2(SI_26_), .ZN(n9996) );
  NAND2_X2 U11755 ( .A1(n9997), .A2(n9996), .ZN(n14255) );
  NAND2_X1 U11756 ( .A1(n9998), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U11757 ( .A1(n10012), .A2(n9999), .ZN(n14003) );
  NAND2_X1 U11758 ( .A1(n14003), .A2(n10035), .ZN(n10004) );
  INV_X1 U11759 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U11760 ( .A1(n10036), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U11761 ( .A1(n10048), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n10000) );
  OAI211_X1 U11762 ( .C1(n14002), .C2(n11987), .A(n10001), .B(n10000), .ZN(
        n10002) );
  INV_X1 U11763 ( .A(n10002), .ZN(n10003) );
  NAND2_X1 U11764 ( .A1(n14255), .A2(n13462), .ZN(n10005) );
  AND2_X1 U11765 ( .A1(n13996), .A2(n10005), .ZN(n13108) );
  INV_X1 U11766 ( .A(n10006), .ZN(n10007) );
  XNOR2_X1 U11767 ( .A(n10008), .B(n10007), .ZN(n12981) );
  NAND2_X1 U11768 ( .A1(n12981), .A2(n10032), .ZN(n10010) );
  NAND2_X1 U11769 ( .A1(n13279), .A2(SI_27_), .ZN(n10009) );
  NAND2_X2 U11770 ( .A1(n10010), .A2(n10009), .ZN(n13987) );
  INV_X1 U11771 ( .A(n10011), .ZN(n10014) );
  NAND2_X1 U11772 ( .A1(n10012), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U11773 ( .A1(n10014), .A2(n10013), .ZN(n13986) );
  NAND2_X1 U11774 ( .A1(n13986), .A2(n10035), .ZN(n10020) );
  INV_X1 U11775 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U11776 ( .A1(n10036), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U11777 ( .A1(n10048), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n10015) );
  OAI211_X1 U11778 ( .C1(n11987), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        n10018) );
  INV_X1 U11779 ( .A(n10018), .ZN(n10019) );
  NAND2_X1 U11780 ( .A1(n13249), .A2(n13250), .ZN(n13124) );
  INV_X1 U11781 ( .A(n13124), .ZN(n13111) );
  AND2_X1 U11782 ( .A1(n13108), .A2(n13124), .ZN(n10021) );
  XNOR2_X2 U11783 ( .A(n10022), .B(n13116), .ZN(n13977) );
  INV_X1 U11784 ( .A(n13977), .ZN(n10024) );
  OR2_X1 U11785 ( .A1(n13987), .A2(n13461), .ZN(n10023) );
  OR2_X1 U11786 ( .A1(n14255), .A2(n13462), .ZN(n13109) );
  OR2_X1 U11787 ( .A1(n13111), .A2(n13109), .ZN(n13107) );
  AND2_X1 U11788 ( .A1(n10023), .A2(n13107), .ZN(n13968) );
  AND2_X1 U11789 ( .A1(n10024), .A2(n13968), .ZN(n10025) );
  AND2_X2 U11790 ( .A1(n13969), .A2(n10025), .ZN(n13973) );
  NAND2_X1 U11791 ( .A1(n13093), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10029) );
  INV_X1 U11792 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14800) );
  AOI22_X1 U11793 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(
        P1_DATAO_REG_29__SCAN_IN), .B1(n14800), .B2(n13089), .ZN(n13269) );
  INV_X1 U11794 ( .A(n13269), .ZN(n10031) );
  XNOR2_X1 U11795 ( .A(n13270), .B(n10031), .ZN(n14314) );
  NAND2_X1 U11796 ( .A1(n14314), .A2(n10032), .ZN(n10034) );
  NAND2_X1 U11797 ( .A1(n13279), .A2(SI_29_), .ZN(n10033) );
  NAND2_X1 U11798 ( .A1(n10034), .A2(n10033), .ZN(n10112) );
  NAND2_X1 U11799 ( .A1(n13961), .A2(n10035), .ZN(n11990) );
  INV_X1 U11800 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U11801 ( .A1(n10048), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U11802 ( .A1(n10036), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n10037) );
  OAI211_X1 U11803 ( .C1(n11987), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10040) );
  INV_X1 U11804 ( .A(n10040), .ZN(n10041) );
  NAND2_X1 U11805 ( .A1(n10112), .A2(n13974), .ZN(n13291) );
  XNOR2_X1 U11806 ( .A(n10042), .B(n8009), .ZN(n10058) );
  NAND2_X1 U11807 ( .A1(n13338), .A2(n13330), .ZN(n10106) );
  INV_X1 U11808 ( .A(n10043), .ZN(n10044) );
  NAND2_X1 U11809 ( .A1(n10044), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10046) );
  INV_X1 U11810 ( .A(n11774), .ZN(n10104) );
  AND2_X1 U11811 ( .A1(n10118), .A2(n10104), .ZN(n13333) );
  INV_X1 U11812 ( .A(n13333), .ZN(n10047) );
  INV_X1 U11813 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U11814 ( .A1(n10048), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10050) );
  NAND2_X1 U11815 ( .A1(n11983), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10049) );
  OAI211_X1 U11816 ( .C1(n11987), .C2(n10051), .A(n10050), .B(n10049), .ZN(
        n10052) );
  INV_X1 U11817 ( .A(n10052), .ZN(n10053) );
  AND2_X1 U11818 ( .A1(n11990), .A2(n10053), .ZN(n13282) );
  INV_X1 U11819 ( .A(n13282), .ZN(n13460) );
  NAND2_X1 U11820 ( .A1(n10055), .A2(n10054), .ZN(n10226) );
  AOI21_X1 U11821 ( .B1(n10056), .B2(P3_B_REG_SCAN_IN), .A(n14159), .ZN(n13954) );
  INV_X1 U11822 ( .A(n10226), .ZN(n10225) );
  AOI22_X1 U11823 ( .A1(n13460), .A2(n13954), .B1(n13116), .B2(n16180), .ZN(
        n10057) );
  OAI21_X2 U11824 ( .B1(n10058), .B2(n14156), .A(n10057), .ZN(n13960) );
  OR2_X1 U11825 ( .A1(n10118), .A2(n10104), .ZN(n10059) );
  XNOR2_X1 U11826 ( .A(n13338), .B(n10059), .ZN(n10061) );
  OR2_X1 U11827 ( .A1(n10118), .A2(n13330), .ZN(n10060) );
  NAND2_X1 U11828 ( .A1(n10061), .A2(n10060), .ZN(n10212) );
  NAND2_X1 U11829 ( .A1(n11774), .A2(n11452), .ZN(n13290) );
  INV_X1 U11830 ( .A(n13290), .ZN(n10215) );
  AND2_X1 U11831 ( .A1(n16467), .A2(n10215), .ZN(n10062) );
  NAND2_X1 U11832 ( .A1(n10212), .A2(n10062), .ZN(n10064) );
  AND2_X1 U11833 ( .A1(n13290), .A2(n11452), .ZN(n10063) );
  NAND2_X1 U11834 ( .A1(n13338), .A2(n10063), .ZN(n10238) );
  INV_X1 U11835 ( .A(n13289), .ZN(n10237) );
  OR2_X1 U11836 ( .A1(n13338), .A2(n10237), .ZN(n16413) );
  INV_X1 U11837 ( .A(n13893), .ZN(n11884) );
  NAND2_X1 U11838 ( .A1(n11884), .A2(n11883), .ZN(n13142) );
  NAND2_X1 U11839 ( .A1(n13143), .A2(n13142), .ZN(n10065) );
  NAND2_X1 U11840 ( .A1(n12117), .A2(n13308), .ZN(n12116) );
  NAND2_X1 U11841 ( .A1(n12116), .A2(n13153), .ZN(n12135) );
  AND2_X1 U11842 ( .A1(n13306), .A2(n10068), .ZN(n10067) );
  NAND2_X1 U11843 ( .A1(n12135), .A2(n10067), .ZN(n12281) );
  INV_X1 U11844 ( .A(n13472), .ZN(n12154) );
  NAND2_X1 U11845 ( .A1(n12154), .A2(n16333), .ZN(n10069) );
  INV_X1 U11846 ( .A(n13164), .ZN(n12289) );
  INV_X1 U11847 ( .A(n13305), .ZN(n12439) );
  NAND2_X1 U11848 ( .A1(n12440), .A2(n12439), .ZN(n12438) );
  NAND2_X1 U11849 ( .A1(n12438), .A2(n13171), .ZN(n12413) );
  NAND2_X1 U11850 ( .A1(n12413), .A2(n13173), .ZN(n12412) );
  NAND2_X1 U11851 ( .A1(n12602), .A2(n16381), .ZN(n13180) );
  INV_X1 U11852 ( .A(n13180), .ZN(n10070) );
  NAND2_X1 U11853 ( .A1(n13468), .A2(n10071), .ZN(n13181) );
  NAND2_X1 U11854 ( .A1(n12755), .A2(n13184), .ZN(n12989) );
  NAND2_X1 U11855 ( .A1(n12780), .A2(n12996), .ZN(n13190) );
  INV_X1 U11856 ( .A(n12780), .ZN(n13466) );
  NAND2_X1 U11857 ( .A1(n13466), .A2(n16441), .ZN(n13188) );
  NAND2_X1 U11858 ( .A1(n12989), .A2(n13312), .ZN(n10072) );
  NAND2_X1 U11859 ( .A1(n10072), .A2(n13190), .ZN(n12919) );
  NAND2_X1 U11860 ( .A1(n12928), .A2(n12782), .ZN(n13194) );
  INV_X1 U11861 ( .A(n12928), .ZN(n13018) );
  NAND2_X1 U11862 ( .A1(n13018), .A2(n16468), .ZN(n13187) );
  NAND2_X1 U11863 ( .A1(n13194), .A2(n13187), .ZN(n13318) );
  NAND2_X1 U11864 ( .A1(n14238), .A2(n13026), .ZN(n13200) );
  NAND2_X1 U11865 ( .A1(n13034), .A2(n13320), .ZN(n10074) );
  OR2_X1 U11866 ( .A1(n14236), .A2(n13465), .ZN(n10073) );
  NAND2_X1 U11867 ( .A1(n10074), .A2(n10073), .ZN(n14153) );
  INV_X1 U11868 ( .A(n14154), .ZN(n13209) );
  NAND2_X1 U11869 ( .A1(n14153), .A2(n13209), .ZN(n10075) );
  NAND2_X1 U11870 ( .A1(n10075), .A2(n13210), .ZN(n14140) );
  NAND2_X1 U11871 ( .A1(n14140), .A2(n14144), .ZN(n10076) );
  INV_X1 U11872 ( .A(n14131), .ZN(n14158) );
  NAND2_X1 U11873 ( .A1(n13216), .A2(n14158), .ZN(n13217) );
  NAND2_X1 U11874 ( .A1(n10076), .A2(n13217), .ZN(n14128) );
  NAND2_X1 U11875 ( .A1(n14128), .A2(n13321), .ZN(n10078) );
  NAND2_X1 U11876 ( .A1(n10078), .A2(n10077), .ZN(n14115) );
  NAND2_X1 U11877 ( .A1(n14115), .A2(n14116), .ZN(n10079) );
  NOR2_X1 U11878 ( .A1(n14205), .A2(n14109), .ZN(n13227) );
  INV_X1 U11879 ( .A(n13227), .ZN(n10080) );
  NAND2_X1 U11880 ( .A1(n14202), .A2(n14089), .ZN(n14050) );
  NAND2_X1 U11881 ( .A1(n10184), .A2(n14050), .ZN(n14069) );
  NAND2_X1 U11882 ( .A1(n14199), .A2(n14073), .ZN(n13127) );
  NAND2_X1 U11883 ( .A1(n13237), .A2(n13127), .ZN(n14051) );
  INV_X1 U11884 ( .A(n14050), .ZN(n13231) );
  NOR2_X1 U11885 ( .A1(n14051), .A2(n13231), .ZN(n10081) );
  NAND2_X1 U11886 ( .A1(n14269), .A2(n14056), .ZN(n13234) );
  NAND2_X1 U11887 ( .A1(n14255), .A2(n14010), .ZN(n13245) );
  NAND2_X1 U11888 ( .A1(n14260), .A2(n14027), .ZN(n13992) );
  INV_X1 U11889 ( .A(n13992), .ZN(n10082) );
  NOR2_X1 U11890 ( .A1(n13993), .A2(n10082), .ZN(n10083) );
  NAND2_X1 U11891 ( .A1(n13978), .A2(n13977), .ZN(n13980) );
  INV_X1 U11892 ( .A(n13116), .ZN(n13359) );
  NAND2_X1 U11893 ( .A1(n10022), .A2(n13359), .ZN(n13242) );
  XNOR2_X1 U11894 ( .A(n13294), .B(n8009), .ZN(n13965) );
  NOR2_X1 U11895 ( .A1(n13960), .A2(n10084), .ZN(n10243) );
  INV_X1 U11896 ( .A(P3_B_REG_SCAN_IN), .ZN(n10085) );
  XNOR2_X1 U11897 ( .A(n12537), .B(n10085), .ZN(n10086) );
  OR2_X1 U11898 ( .A1(n11024), .A2(P3_D_REG_0__SCAN_IN), .ZN(n10089) );
  OR2_X1 U11899 ( .A1(n12880), .A2(n10087), .ZN(n10088) );
  OR2_X1 U11900 ( .A1(n11024), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10091) );
  OR2_X1 U11901 ( .A1(n12633), .A2(n12880), .ZN(n10090) );
  NAND2_X1 U11902 ( .A1(n14307), .A2(n14305), .ZN(n10235) );
  INV_X1 U11903 ( .A(n10235), .ZN(n10103) );
  NOR2_X1 U11904 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n10095) );
  NOR4_X1 U11905 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n10094) );
  NOR4_X1 U11906 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n10093) );
  NOR4_X1 U11907 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n10092) );
  NAND4_X1 U11908 ( .A1(n10095), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n10101) );
  NOR4_X1 U11909 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n10099) );
  NOR4_X1 U11910 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n10098) );
  NOR4_X1 U11911 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n10097) );
  NOR4_X1 U11912 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n10096) );
  NAND4_X1 U11913 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n10100) );
  NOR2_X1 U11914 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  NAND2_X1 U11915 ( .A1(n10103), .A2(n10108), .ZN(n10213) );
  INV_X1 U11916 ( .A(n13332), .ZN(n10105) );
  OR2_X1 U11917 ( .A1(n10106), .A2(n10105), .ZN(n10214) );
  INV_X1 U11918 ( .A(n14307), .ZN(n10107) );
  NAND2_X1 U11919 ( .A1(n10107), .A2(n11917), .ZN(n10234) );
  NAND2_X1 U11920 ( .A1(n10224), .A2(n10212), .ZN(n10109) );
  OAI21_X1 U11921 ( .B1(n10213), .B2(n10110), .A(n10109), .ZN(n10111) );
  INV_X1 U11922 ( .A(n13337), .ZN(n10208) );
  OR2_X1 U11923 ( .A1(n10243), .A2(n16562), .ZN(n10117) );
  INV_X1 U11924 ( .A(n10112), .ZN(n13963) );
  NOR2_X1 U11925 ( .A1(n13963), .A2(n14296), .ZN(n10115) );
  INV_X1 U11926 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10113) );
  NOR2_X1 U11927 ( .A1(n16447), .A2(n10113), .ZN(n10114) );
  NAND2_X1 U11928 ( .A1(n10117), .A2(n10116), .ZN(P3_U3456) );
  NAND2_X1 U11929 ( .A1(n14307), .A2(n13332), .ZN(n10120) );
  OAI21_X1 U11930 ( .B1(n10118), .B2(n11452), .A(n11774), .ZN(n10119) );
  XNOR2_X1 U11931 ( .A(n10121), .B(n10129), .ZN(n10123) );
  INV_X1 U11932 ( .A(n10123), .ZN(n10124) );
  NAND2_X1 U11933 ( .A1(n10122), .A2(n10124), .ZN(n10125) );
  XNOR2_X1 U11934 ( .A(n11645), .B(n10129), .ZN(n10126) );
  XNOR2_X1 U11935 ( .A(n10126), .B(n12118), .ZN(n11644) );
  INV_X1 U11936 ( .A(n10126), .ZN(n10127) );
  AND2_X1 U11937 ( .A1(n12118), .A2(n10127), .ZN(n10128) );
  XNOR2_X1 U11938 ( .A(n12128), .B(n10191), .ZN(n10130) );
  XNOR2_X1 U11939 ( .A(n10130), .B(n12136), .ZN(n11660) );
  INV_X1 U11940 ( .A(n10130), .ZN(n10131) );
  OR2_X1 U11941 ( .A1(n12136), .A2(n10131), .ZN(n10132) );
  XNOR2_X1 U11942 ( .A(n12141), .B(n10199), .ZN(n10134) );
  XNOR2_X1 U11943 ( .A(n10134), .B(n12119), .ZN(n11731) );
  NAND2_X1 U11944 ( .A1(n12119), .A2(n10134), .ZN(n10135) );
  NAND2_X1 U11945 ( .A1(n11728), .A2(n10135), .ZN(n11846) );
  XNOR2_X1 U11946 ( .A(n12333), .B(n10191), .ZN(n10136) );
  XNOR2_X1 U11947 ( .A(n10136), .B(n12293), .ZN(n11845) );
  INV_X1 U11948 ( .A(n10136), .ZN(n10137) );
  NAND2_X1 U11949 ( .A1(n12293), .A2(n10137), .ZN(n10138) );
  XNOR2_X1 U11950 ( .A(n16333), .B(n10191), .ZN(n10140) );
  XNOR2_X1 U11951 ( .A(n10140), .B(n13472), .ZN(n11992) );
  INV_X1 U11952 ( .A(n11992), .ZN(n10139) );
  NAND2_X1 U11953 ( .A1(n10140), .A2(n13472), .ZN(n10141) );
  NAND2_X1 U11954 ( .A1(n11994), .A2(n10141), .ZN(n12152) );
  XNOR2_X1 U11955 ( .A(n12449), .B(n10191), .ZN(n10142) );
  XNOR2_X1 U11956 ( .A(n10142), .B(n12294), .ZN(n12151) );
  NAND2_X1 U11957 ( .A1(n12152), .A2(n12151), .ZN(n12150) );
  INV_X1 U11958 ( .A(n10142), .ZN(n10143) );
  OR2_X1 U11959 ( .A1(n12294), .A2(n10143), .ZN(n10144) );
  NAND2_X1 U11960 ( .A1(n12150), .A2(n10144), .ZN(n12224) );
  XNOR2_X1 U11961 ( .A(n12416), .B(n10191), .ZN(n10145) );
  XNOR2_X1 U11962 ( .A(n12588), .B(n10145), .ZN(n12223) );
  INV_X1 U11963 ( .A(n10145), .ZN(n10146) );
  OR2_X1 U11964 ( .A1(n12588), .A2(n10146), .ZN(n10147) );
  XNOR2_X1 U11965 ( .A(n16381), .B(n10199), .ZN(n10148) );
  XNOR2_X1 U11966 ( .A(n10148), .B(n12602), .ZN(n12512) );
  NAND2_X1 U11967 ( .A1(n12602), .A2(n10148), .ZN(n10149) );
  XNOR2_X1 U11968 ( .A(n16411), .B(n10191), .ZN(n10150) );
  XNOR2_X1 U11969 ( .A(n10150), .B(n12696), .ZN(n12600) );
  INV_X1 U11970 ( .A(n10150), .ZN(n10151) );
  OR2_X1 U11971 ( .A1(n12696), .A2(n10151), .ZN(n10152) );
  NAND2_X1 U11972 ( .A1(n12599), .A2(n10152), .ZN(n12695) );
  AND2_X1 U11973 ( .A1(n10155), .A2(n10153), .ZN(n10154) );
  MUX2_X1 U11974 ( .A(n10154), .B(n13312), .S(n10199), .Z(n12694) );
  NAND2_X1 U11975 ( .A1(n12695), .A2(n12694), .ZN(n12693) );
  MUX2_X1 U11976 ( .A(n10155), .B(n13188), .S(n10199), .Z(n10156) );
  INV_X1 U11977 ( .A(n13187), .ZN(n10158) );
  MUX2_X1 U11978 ( .A(n10159), .B(n10158), .S(n10199), .Z(n12773) );
  MUX2_X1 U11979 ( .A(n10160), .B(n13194), .S(n10199), .Z(n12772) );
  INV_X1 U11980 ( .A(n13197), .ZN(n13317) );
  MUX2_X1 U11981 ( .A(n13197), .B(n13317), .S(n10199), .Z(n12924) );
  MUX2_X1 U11982 ( .A(n10161), .B(n13200), .S(n10199), .Z(n10162) );
  XNOR2_X1 U11983 ( .A(n14236), .B(n10199), .ZN(n10163) );
  XNOR2_X1 U11984 ( .A(n10163), .B(n13465), .ZN(n13001) );
  INV_X1 U11985 ( .A(n10163), .ZN(n10164) );
  XNOR2_X1 U11986 ( .A(n14229), .B(n10199), .ZN(n10165) );
  XNOR2_X1 U11987 ( .A(n10165), .B(n13027), .ZN(n13038) );
  INV_X1 U11988 ( .A(n10165), .ZN(n10166) );
  NAND2_X1 U11989 ( .A1(n10166), .A2(n13027), .ZN(n10167) );
  XNOR2_X1 U11990 ( .A(n13216), .B(n10199), .ZN(n10168) );
  XNOR2_X1 U11991 ( .A(n10168), .B(n14131), .ZN(n13395) );
  INV_X1 U11992 ( .A(n10168), .ZN(n10169) );
  NAND2_X1 U11993 ( .A1(n10169), .A2(n14131), .ZN(n10170) );
  NAND2_X1 U11994 ( .A1(n10171), .A2(n10170), .ZN(n13405) );
  XNOR2_X1 U11995 ( .A(n14220), .B(n10191), .ZN(n13403) );
  INV_X1 U11996 ( .A(n13403), .ZN(n10172) );
  XNOR2_X1 U11997 ( .A(n13436), .B(n10199), .ZN(n10173) );
  XNOR2_X1 U11998 ( .A(n10173), .B(n14132), .ZN(n13439) );
  INV_X1 U11999 ( .A(n10173), .ZN(n10174) );
  XNOR2_X1 U12000 ( .A(n10175), .B(n10199), .ZN(n10176) );
  XNOR2_X1 U12001 ( .A(n10176), .B(n13442), .ZN(n13371) );
  NAND2_X1 U12002 ( .A1(n13372), .A2(n13371), .ZN(n13370) );
  INV_X1 U12003 ( .A(n10176), .ZN(n10177) );
  NAND2_X1 U12004 ( .A1(n10177), .A2(n13442), .ZN(n10178) );
  NAND2_X1 U12005 ( .A1(n13370), .A2(n10178), .ZN(n13424) );
  XNOR2_X1 U12006 ( .A(n14205), .B(n10199), .ZN(n13422) );
  NAND2_X1 U12007 ( .A1(n13422), .A2(n14109), .ZN(n10179) );
  NAND2_X1 U12008 ( .A1(n13424), .A2(n10179), .ZN(n10182) );
  INV_X1 U12009 ( .A(n13422), .ZN(n10180) );
  NAND2_X1 U12010 ( .A1(n10180), .A2(n13464), .ZN(n10181) );
  INV_X1 U12011 ( .A(n10183), .ZN(n10185) );
  INV_X1 U12012 ( .A(n10184), .ZN(n13230) );
  MUX2_X1 U12013 ( .A(n10185), .B(n13230), .S(n10199), .Z(n13380) );
  MUX2_X1 U12014 ( .A(n10186), .B(n14050), .S(n10199), .Z(n13378) );
  XNOR2_X1 U12015 ( .A(n14199), .B(n10191), .ZN(n10187) );
  INV_X1 U12016 ( .A(n10187), .ZN(n10188) );
  AND2_X1 U12017 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  XNOR2_X1 U12018 ( .A(n14265), .B(n10191), .ZN(n13414) );
  INV_X1 U12019 ( .A(n14056), .ZN(n14028) );
  XNOR2_X1 U12020 ( .A(n13367), .B(n10191), .ZN(n13411) );
  INV_X1 U12021 ( .A(n13411), .ZN(n10192) );
  OAI22_X1 U12022 ( .A1(n13414), .A2(n14009), .B1(n14028), .B2(n10192), .ZN(
        n10196) );
  OAI21_X1 U12023 ( .B1(n13411), .B2(n14056), .A(n14042), .ZN(n10194) );
  NOR2_X1 U12024 ( .A1(n14042), .A2(n14056), .ZN(n10193) );
  AOI22_X1 U12025 ( .A1(n13414), .A2(n10194), .B1(n10193), .B2(n10192), .ZN(
        n10195) );
  XNOR2_X1 U12026 ( .A(n14260), .B(n10199), .ZN(n10197) );
  XNOR2_X1 U12027 ( .A(n10197), .B(n13463), .ZN(n13389) );
  XNOR2_X1 U12028 ( .A(n14255), .B(n10199), .ZN(n10200) );
  XNOR2_X1 U12029 ( .A(n10200), .B(n14010), .ZN(n13449) );
  INV_X1 U12030 ( .A(n10200), .ZN(n10201) );
  XNOR2_X1 U12031 ( .A(n13987), .B(n10199), .ZN(n10202) );
  XNOR2_X1 U12032 ( .A(n10202), .B(n13461), .ZN(n13358) );
  XOR2_X1 U12033 ( .A(n10199), .B(n13977), .Z(n10203) );
  XNOR2_X1 U12034 ( .A(n10204), .B(n10203), .ZN(n10210) );
  NAND2_X1 U12035 ( .A1(n10212), .A2(n16467), .ZN(n10207) );
  INV_X1 U12036 ( .A(n10214), .ZN(n10205) );
  NAND2_X1 U12037 ( .A1(n10224), .A2(n10205), .ZN(n10206) );
  OAI21_X1 U12038 ( .B1(n10213), .B2(n10207), .A(n10206), .ZN(n10209) );
  NAND2_X1 U12039 ( .A1(n10210), .A2(n13437), .ZN(n10233) );
  NAND2_X1 U12040 ( .A1(n10213), .A2(n10237), .ZN(n10211) );
  NAND2_X1 U12041 ( .A1(n10213), .A2(n10212), .ZN(n10218) );
  OR2_X1 U12042 ( .A1(n10224), .A2(n10214), .ZN(n10216) );
  OR2_X1 U12043 ( .A1(n13266), .A2(n10215), .ZN(n10240) );
  NAND4_X1 U12044 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10240), .ZN(
        n10219) );
  NAND2_X1 U12045 ( .A1(n10219), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10222) );
  NOR2_X1 U12046 ( .A1(n13337), .A2(n13336), .ZN(n10223) );
  INV_X1 U12047 ( .A(n10223), .ZN(n10220) );
  OR2_X1 U12048 ( .A1(n10224), .A2(n10220), .ZN(n10221) );
  AND2_X1 U12049 ( .A1(n10222), .A2(n10221), .ZN(n11411) );
  NAND2_X1 U12050 ( .A1(n10224), .A2(n10223), .ZN(n10227) );
  NOR2_X1 U12051 ( .A1(n13974), .A2(n13451), .ZN(n10229) );
  OR2_X2 U12052 ( .A1(n10227), .A2(n10226), .ZN(n13450) );
  OAI22_X1 U12053 ( .A1(n13999), .A2(n13450), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13664), .ZN(n10228) );
  AOI211_X1 U12054 ( .C1(n13981), .C2(n13454), .A(n10229), .B(n10228), .ZN(
        n10230) );
  NAND2_X1 U12055 ( .A1(n10233), .A2(n10232), .ZN(P3_U3160) );
  INV_X1 U12056 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10244) );
  AND2_X1 U12057 ( .A1(n10235), .A2(n10234), .ZN(n11921) );
  NOR2_X1 U12058 ( .A1(n16467), .A2(n10237), .ZN(n10239) );
  NAND2_X1 U12059 ( .A1(n13266), .A2(n10238), .ZN(n11915) );
  OAI21_X1 U12060 ( .B1(n10239), .B2(n11915), .A(n11917), .ZN(n10242) );
  NAND2_X1 U12061 ( .A1(n10240), .A2(n11915), .ZN(n11916) );
  NAND2_X1 U12062 ( .A1(n11916), .A2(n14305), .ZN(n10241) );
  NAND2_X1 U12063 ( .A1(n10245), .A2(n8337), .ZN(P3_U3488) );
  NAND2_X1 U12064 ( .A1(n10309), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10326) );
  INV_X1 U12065 ( .A(n10326), .ZN(n10246) );
  NAND2_X1 U12066 ( .A1(n10246), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10334) );
  INV_X1 U12067 ( .A(n10334), .ZN(n10247) );
  NAND2_X1 U12068 ( .A1(n10247), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10343) );
  INV_X1 U12069 ( .A(n10352), .ZN(n10248) );
  NAND2_X1 U12070 ( .A1(n10248), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10361) );
  INV_X1 U12071 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10360) );
  INV_X1 U12072 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10382) );
  INV_X1 U12073 ( .A(n10394), .ZN(n10250) );
  NAND2_X1 U12074 ( .A1(n10250), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n10400) );
  INV_X1 U12075 ( .A(n10400), .ZN(n10251) );
  NAND2_X1 U12076 ( .A1(n10251), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10408) );
  INV_X1 U12077 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n12791) );
  INV_X1 U12078 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10421) );
  AND2_X1 U12079 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n10253) );
  INV_X1 U12080 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U12081 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n10255) );
  INV_X1 U12082 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14415) );
  INV_X1 U12083 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10256) );
  OAI21_X1 U12084 ( .B1(n10437), .B2(n14415), .A(n10256), .ZN(n10257) );
  AND2_X1 U12085 ( .A1(n10448), .A2(n10257), .ZN(n14574) );
  AND2_X4 U12086 ( .A1(n10258), .A2(n10259), .ZN(n10483) );
  NAND2_X1 U12087 ( .A1(n14574), .A2(n10483), .ZN(n10265) );
  INV_X1 U12088 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U12089 ( .A1(n10505), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U12090 ( .A1(n10507), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n10260) );
  OAI211_X1 U12091 ( .C1(n10262), .C2(n10499), .A(n10261), .B(n10260), .ZN(
        n10263) );
  INV_X1 U12092 ( .A(n10263), .ZN(n10264) );
  NAND2_X1 U12093 ( .A1(n10265), .A2(n10264), .ZN(n14558) );
  XNOR2_X1 U12094 ( .A(n10437), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n14586) );
  NAND2_X1 U12095 ( .A1(n14586), .A2(n10483), .ZN(n10271) );
  INV_X1 U12096 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U12097 ( .A1(n10505), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n10267) );
  NAND2_X1 U12098 ( .A1(n10507), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n10266) );
  OAI211_X1 U12099 ( .C1(n10268), .C2(n10499), .A(n10267), .B(n10266), .ZN(
        n10269) );
  INV_X1 U12100 ( .A(n10269), .ZN(n10270) );
  NAND2_X1 U12101 ( .A1(n10271), .A2(n10270), .ZN(n14455) );
  INV_X1 U12102 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10273) );
  INV_X1 U12103 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10272) );
  OAI21_X1 U12104 ( .B1(n10424), .B2(n10273), .A(n10272), .ZN(n10274) );
  NAND2_X1 U12105 ( .A1(n10274), .A2(n10435), .ZN(n14613) );
  OR2_X1 U12106 ( .A1(n14613), .A2(n10496), .ZN(n10279) );
  INV_X1 U12107 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n14614) );
  NAND2_X1 U12108 ( .A1(n10505), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n10276) );
  NAND2_X1 U12109 ( .A1(n10507), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n10275) );
  OAI211_X1 U12110 ( .C1(n14614), .C2(n10499), .A(n10276), .B(n10275), .ZN(
        n10277) );
  INV_X1 U12111 ( .A(n10277), .ZN(n10278) );
  NAND2_X1 U12112 ( .A1(n10279), .A2(n10278), .ZN(n14629) );
  INV_X1 U12113 ( .A(n14629), .ZN(n14596) );
  OR2_X1 U12114 ( .A1(n14739), .A2(n14596), .ZN(n10434) );
  NAND2_X1 U12115 ( .A1(n14739), .A2(n14596), .ZN(n10280) );
  NAND2_X1 U12116 ( .A1(n10434), .A2(n10280), .ZN(n14606) );
  INV_X1 U12117 ( .A(n14606), .ZN(n14609) );
  XNOR2_X1 U12118 ( .A(n10424), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n14634) );
  NAND2_X1 U12119 ( .A1(n14634), .A2(n10483), .ZN(n10286) );
  INV_X1 U12120 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U12121 ( .A1(n10507), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12122 ( .A1(n10505), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n10281) );
  OAI211_X1 U12123 ( .C1(n10283), .C2(n10499), .A(n10282), .B(n10281), .ZN(
        n10284) );
  INV_X1 U12124 ( .A(n10284), .ZN(n10285) );
  NAND2_X1 U12125 ( .A1(n10286), .A2(n10285), .ZN(n14457) );
  INV_X1 U12126 ( .A(n14457), .ZN(n14654) );
  NAND2_X1 U12127 ( .A1(n10296), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U12128 ( .A1(n10302), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U12129 ( .A1(n10483), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10287) );
  INV_X1 U12130 ( .A(n14475), .ZN(n11405) );
  NAND2_X1 U12131 ( .A1(n11405), .A2(n16106), .ZN(n10806) );
  INV_X1 U12132 ( .A(n10806), .ZN(n11740) );
  NAND2_X1 U12133 ( .A1(n10483), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n10294) );
  NAND2_X1 U12134 ( .A1(n10302), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U12135 ( .A1(n10296), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10292) );
  NAND2_X1 U12136 ( .A1(n10506), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10291) );
  INV_X1 U12137 ( .A(n14473), .ZN(n16109) );
  NAND2_X1 U12138 ( .A1(n16109), .A2(n11752), .ZN(n10295) );
  NAND2_X1 U12139 ( .A1(n10296), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U12140 ( .A1(n10483), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n10298) );
  NAND2_X2 U12141 ( .A1(n10506), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10297) );
  NAND4_X4 U12142 ( .A1(n10300), .A2(n10299), .A3(n10298), .A4(n10297), .ZN(
        n14472) );
  INV_X1 U12143 ( .A(n14472), .ZN(n10513) );
  AND2_X1 U12144 ( .A1(n16225), .A2(n10513), .ZN(n10301) );
  AOI21_X1 U12145 ( .B1(n16215), .B2(n10807), .A(n10301), .ZN(n16253) );
  INV_X1 U12146 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n16271) );
  NAND2_X1 U12147 ( .A1(n10483), .A2(n16271), .ZN(n10306) );
  NAND2_X1 U12148 ( .A1(n10302), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U12149 ( .A1(n10506), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U12150 ( .A1(n16270), .A2(n11695), .ZN(n10307) );
  NAND2_X1 U12151 ( .A1(n10296), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U12152 ( .A1(n10302), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n10313) );
  INV_X1 U12153 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10308) );
  NAND2_X1 U12154 ( .A1(n16271), .A2(n10308), .ZN(n10310) );
  INV_X1 U12155 ( .A(n10309), .ZN(n10318) );
  AND2_X1 U12156 ( .A1(n10310), .A2(n10318), .ZN(n11690) );
  NAND2_X1 U12157 ( .A1(n10483), .A2(n11690), .ZN(n10312) );
  NAND2_X1 U12158 ( .A1(n10506), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10311) );
  NAND4_X1 U12159 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n14470) );
  NAND2_X1 U12160 ( .A1(n11857), .A2(n11856), .ZN(n10316) );
  INV_X1 U12161 ( .A(n14470), .ZN(n11424) );
  NAND2_X1 U12162 ( .A1(n11853), .A2(n11424), .ZN(n10315) );
  NAND2_X1 U12163 ( .A1(n10296), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U12164 ( .A1(n10302), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n10322) );
  INV_X1 U12165 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10317) );
  NAND2_X1 U12166 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  AND2_X1 U12167 ( .A1(n10326), .A2(n10319), .ZN(n12100) );
  NAND2_X1 U12168 ( .A1(n10483), .A2(n12100), .ZN(n10321) );
  NAND2_X1 U12169 ( .A1(n10506), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10320) );
  INV_X1 U12170 ( .A(n14469), .ZN(n10324) );
  INV_X1 U12171 ( .A(n12101), .ZN(n16323) );
  NAND2_X1 U12172 ( .A1(n10507), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U12173 ( .A1(n10296), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10330) );
  INV_X1 U12174 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10325) );
  NAND2_X1 U12175 ( .A1(n10326), .A2(n10325), .ZN(n10327) );
  AND2_X1 U12176 ( .A1(n10334), .A2(n10327), .ZN(n11651) );
  NAND2_X1 U12177 ( .A1(n10483), .A2(n11651), .ZN(n10329) );
  NAND2_X1 U12178 ( .A1(n10506), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10328) );
  NAND4_X1 U12179 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n14468) );
  XNOR2_X1 U12180 ( .A(n11906), .B(n14468), .ZN(n11456) );
  INV_X1 U12181 ( .A(n14468), .ZN(n11635) );
  NAND2_X1 U12182 ( .A1(n11906), .A2(n11635), .ZN(n10332) );
  NAND2_X1 U12183 ( .A1(n11455), .A2(n10332), .ZN(n12090) );
  NAND2_X1 U12184 ( .A1(n10507), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10339) );
  NAND2_X1 U12185 ( .A1(n10296), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10338) );
  INV_X1 U12186 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10333) );
  NAND2_X1 U12187 ( .A1(n10334), .A2(n10333), .ZN(n10335) );
  AND2_X1 U12188 ( .A1(n10343), .A2(n10335), .ZN(n12085) );
  NAND2_X1 U12189 ( .A1(n10483), .A2(n12085), .ZN(n10337) );
  NAND2_X1 U12190 ( .A1(n10506), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10336) );
  NAND4_X1 U12191 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n14467) );
  NAND2_X1 U12192 ( .A1(n16360), .A2(n14467), .ZN(n10340) );
  NAND2_X1 U12193 ( .A1(n12090), .A2(n10340), .ZN(n10342) );
  NAND2_X1 U12194 ( .A1(n12086), .A2(n11505), .ZN(n10341) );
  NAND2_X1 U12195 ( .A1(n10342), .A2(n10341), .ZN(n11894) );
  NAND2_X1 U12196 ( .A1(n10505), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U12197 ( .A1(n10507), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U12198 ( .A1(n10343), .A2(n11509), .ZN(n10344) );
  AND2_X1 U12199 ( .A1(n10352), .A2(n10344), .ZN(n12057) );
  NAND2_X1 U12200 ( .A1(n10483), .A2(n12057), .ZN(n10346) );
  NAND2_X1 U12201 ( .A1(n10506), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10345) );
  NAND4_X1 U12202 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n14466) );
  XNOR2_X1 U12203 ( .A(n12058), .B(n14466), .ZN(n11895) );
  NAND2_X1 U12204 ( .A1(n11894), .A2(n11895), .ZN(n10350) );
  INV_X1 U12205 ( .A(n14466), .ZN(n11680) );
  NAND2_X1 U12206 ( .A1(n12058), .A2(n11680), .ZN(n10349) );
  NAND2_X1 U12207 ( .A1(n10505), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U12208 ( .A1(n10507), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10356) );
  INV_X1 U12209 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11685) );
  NAND2_X1 U12210 ( .A1(n10352), .A2(n11685), .ZN(n10353) );
  AND2_X1 U12211 ( .A1(n10361), .A2(n10353), .ZN(n16398) );
  NAND2_X1 U12212 ( .A1(n10483), .A2(n16398), .ZN(n10355) );
  NAND2_X1 U12213 ( .A1(n10506), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10354) );
  NAND4_X1 U12214 ( .A1(n10357), .A2(n10356), .A3(n10355), .A4(n10354), .ZN(
        n14465) );
  XNOR2_X1 U12215 ( .A(n16400), .B(n14465), .ZN(n12198) );
  NAND2_X1 U12216 ( .A1(n12199), .A2(n12198), .ZN(n10359) );
  INV_X1 U12217 ( .A(n14465), .ZN(n12026) );
  NAND2_X1 U12218 ( .A1(n16400), .A2(n12026), .ZN(n10358) );
  NAND2_X1 U12219 ( .A1(n10505), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U12220 ( .A1(n10507), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10365) );
  NAND2_X1 U12221 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  AND2_X1 U12222 ( .A1(n10369), .A2(n10362), .ZN(n12214) );
  NAND2_X1 U12223 ( .A1(n10483), .A2(n12214), .ZN(n10364) );
  NAND2_X1 U12224 ( .A1(n10506), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U12225 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n14464) );
  INV_X1 U12226 ( .A(n14464), .ZN(n12247) );
  AND2_X1 U12227 ( .A1(n12037), .A2(n12247), .ZN(n10368) );
  OR2_X1 U12228 ( .A1(n12037), .A2(n12247), .ZN(n10367) );
  NAND2_X1 U12229 ( .A1(n10505), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U12230 ( .A1(n10507), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10373) );
  INV_X1 U12231 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n15610) );
  NAND2_X1 U12232 ( .A1(n10369), .A2(n15610), .ZN(n10370) );
  AND2_X1 U12233 ( .A1(n10383), .A2(n10370), .ZN(n10948) );
  NAND2_X1 U12234 ( .A1(n10483), .A2(n10948), .ZN(n10372) );
  NAND2_X1 U12235 ( .A1(n10506), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10371) );
  NAND4_X1 U12236 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n14463) );
  XNOR2_X1 U12237 ( .A(n12254), .B(n12432), .ZN(n12255) );
  NAND2_X1 U12238 ( .A1(n12254), .A2(n12432), .ZN(n12426) );
  NAND2_X1 U12239 ( .A1(n10507), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U12240 ( .A1(n10505), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10377) );
  XNOR2_X1 U12241 ( .A(n10383), .B(P2_REG3_REG_12__SCAN_IN), .ZN(n12399) );
  NAND2_X1 U12242 ( .A1(n10483), .A2(n12399), .ZN(n10376) );
  NAND2_X1 U12243 ( .A1(n10506), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U12244 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n14462) );
  INV_X1 U12245 ( .A(n14462), .ZN(n12246) );
  NAND2_X1 U12246 ( .A1(n14677), .A2(n12246), .ZN(n12494) );
  OR2_X1 U12247 ( .A1(n14677), .A2(n12246), .ZN(n10379) );
  NAND2_X1 U12248 ( .A1(n12494), .A2(n10379), .ZN(n12427) );
  INV_X1 U12249 ( .A(n12427), .ZN(n12421) );
  NAND2_X1 U12250 ( .A1(n10380), .A2(n12421), .ZN(n12496) );
  NAND2_X1 U12251 ( .A1(n12496), .A2(n12494), .ZN(n10390) );
  NAND2_X1 U12252 ( .A1(n10505), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10388) );
  NAND2_X1 U12253 ( .A1(n10507), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10387) );
  OAI21_X1 U12254 ( .B1(n10383), .B2(n10382), .A(n10381), .ZN(n10384) );
  AND2_X1 U12255 ( .A1(n10384), .A2(n10394), .ZN(n12501) );
  NAND2_X1 U12256 ( .A1(n10483), .A2(n12501), .ZN(n10386) );
  NAND2_X1 U12257 ( .A1(n10506), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10385) );
  NAND4_X1 U12258 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n12400) );
  XNOR2_X1 U12259 ( .A(n12504), .B(n12431), .ZN(n12495) );
  INV_X1 U12260 ( .A(n12495), .ZN(n10389) );
  NAND2_X1 U12261 ( .A1(n10390), .A2(n10389), .ZN(n12493) );
  NAND2_X1 U12262 ( .A1(n12504), .A2(n12431), .ZN(n10391) );
  NAND2_X1 U12263 ( .A1(n10505), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U12264 ( .A1(n10507), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U12265 ( .A1(n10393), .A2(n10392), .ZN(n10397) );
  INV_X1 U12266 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n15624) );
  NAND2_X1 U12267 ( .A1(n10394), .A2(n15624), .ZN(n10395) );
  NAND2_X1 U12268 ( .A1(n10400), .A2(n10395), .ZN(n14663) );
  INV_X1 U12269 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n14664) );
  OAI22_X1 U12270 ( .A1(n14663), .A2(n10496), .B1(n10499), .B2(n14664), .ZN(
        n10396) );
  INV_X1 U12271 ( .A(n14461), .ZN(n10678) );
  OR2_X1 U12272 ( .A1(n14666), .A2(n10678), .ZN(n10398) );
  INV_X1 U12273 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10406) );
  INV_X1 U12274 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U12275 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  NAND2_X1 U12276 ( .A1(n10408), .A2(n10401), .ZN(n12896) );
  OR2_X1 U12277 ( .A1(n12896), .A2(n10496), .ZN(n10405) );
  NAND2_X1 U12278 ( .A1(n10507), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U12279 ( .A1(n10506), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n10402) );
  AND2_X1 U12280 ( .A1(n10403), .A2(n10402), .ZN(n10404) );
  OAI211_X1 U12281 ( .C1(n10407), .C2(n10406), .A(n10405), .B(n10404), .ZN(
        n14460) );
  XNOR2_X1 U12282 ( .A(n12902), .B(n14460), .ZN(n12627) );
  INV_X1 U12283 ( .A(n14460), .ZN(n12786) );
  OR2_X1 U12284 ( .A1(n12902), .A2(n12786), .ZN(n12743) );
  NAND2_X1 U12285 ( .A1(n10408), .A2(n12791), .ZN(n10409) );
  NAND2_X1 U12286 ( .A1(n10415), .A2(n10409), .ZN(n12790) );
  AOI22_X1 U12287 ( .A1(n10505), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n10507), 
        .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U12288 ( .A1(n10506), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n10410) );
  OAI211_X1 U12289 ( .C1(n12790), .C2(n10496), .A(n10411), .B(n10410), .ZN(
        n14459) );
  INV_X1 U12290 ( .A(n14459), .ZN(n10412) );
  NAND2_X1 U12291 ( .A1(n12795), .A2(n10412), .ZN(n10413) );
  NAND2_X1 U12292 ( .A1(n12943), .A2(n12941), .ZN(n10419) );
  INV_X1 U12293 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n15659) );
  INV_X1 U12294 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10414) );
  NAND2_X1 U12295 ( .A1(n10415), .A2(n10414), .ZN(n10416) );
  NAND2_X1 U12296 ( .A1(n10422), .A2(n10416), .ZN(n12938) );
  OR2_X1 U12297 ( .A1(n12938), .A2(n10496), .ZN(n10418) );
  AOI22_X1 U12298 ( .A1(n10505), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n10507), 
        .B2(P2_REG0_REG_17__SCAN_IN), .ZN(n10417) );
  OAI211_X1 U12299 ( .C1(n10499), .C2(n15659), .A(n10418), .B(n10417), .ZN(
        n14458) );
  INV_X1 U12300 ( .A(n14458), .ZN(n14653) );
  XNOR2_X1 U12301 ( .A(n14791), .B(n14653), .ZN(n12942) );
  INV_X1 U12302 ( .A(n12942), .ZN(n12933) );
  NAND2_X1 U12303 ( .A1(n10419), .A2(n12933), .ZN(n12945) );
  OR2_X1 U12304 ( .A1(n14791), .A2(n14653), .ZN(n10420) );
  NAND2_X1 U12305 ( .A1(n12945), .A2(n10420), .ZN(n14651) );
  NAND2_X1 U12306 ( .A1(n10422), .A2(n10421), .ZN(n10423) );
  AND2_X1 U12307 ( .A1(n10424), .A2(n10423), .ZN(n14646) );
  NAND2_X1 U12308 ( .A1(n14646), .A2(n10483), .ZN(n10430) );
  INV_X1 U12309 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U12310 ( .A1(n10505), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n10426) );
  NAND2_X1 U12311 ( .A1(n10507), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n10425) );
  OAI211_X1 U12312 ( .C1(n10427), .C2(n10499), .A(n10426), .B(n10425), .ZN(
        n10428) );
  INV_X1 U12313 ( .A(n10428), .ZN(n10429) );
  NAND2_X1 U12314 ( .A1(n10430), .A2(n10429), .ZN(n14626) );
  NAND2_X1 U12315 ( .A1(n7745), .A2(n14360), .ZN(n10431) );
  OAI21_X1 U12316 ( .B1(n14654), .B2(n14742), .A(n14621), .ZN(n10433) );
  NAND2_X1 U12317 ( .A1(n14742), .A2(n14654), .ZN(n10432) );
  AND2_X1 U12318 ( .A1(n10433), .A2(n10432), .ZN(n14608) );
  NAND2_X1 U12319 ( .A1(n10435), .A2(n10938), .ZN(n10436) );
  NAND2_X1 U12320 ( .A1(n10437), .A2(n10436), .ZN(n14599) );
  OR2_X1 U12321 ( .A1(n14599), .A2(n10496), .ZN(n10442) );
  INV_X1 U12322 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n14600) );
  NAND2_X1 U12323 ( .A1(n10507), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n10439) );
  NAND2_X1 U12324 ( .A1(n10505), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n10438) );
  OAI211_X1 U12325 ( .C1(n10499), .C2(n14600), .A(n10439), .B(n10438), .ZN(
        n10440) );
  INV_X1 U12326 ( .A(n10440), .ZN(n10441) );
  NAND2_X1 U12327 ( .A1(n10442), .A2(n10441), .ZN(n14456) );
  INV_X1 U12328 ( .A(n14456), .ZN(n14581) );
  NOR2_X1 U12329 ( .A1(n14732), .A2(n14581), .ZN(n10802) );
  INV_X1 U12330 ( .A(n10802), .ZN(n10443) );
  AND2_X1 U12331 ( .A1(n14732), .A2(n14581), .ZN(n10801) );
  INV_X1 U12332 ( .A(n14455), .ZN(n14597) );
  OR2_X1 U12333 ( .A1(n14569), .A2(n14566), .ZN(n10445) );
  OR2_X1 U12334 ( .A1(n14721), .A2(n14582), .ZN(n10444) );
  NAND2_X1 U12335 ( .A1(n10445), .A2(n10444), .ZN(n14556) );
  INV_X1 U12336 ( .A(n10448), .ZN(n10446) );
  NAND2_X1 U12337 ( .A1(n10446), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n10460) );
  INV_X1 U12338 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U12339 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  NAND2_X1 U12340 ( .A1(n10460), .A2(n10449), .ZN(n14551) );
  OR2_X1 U12341 ( .A1(n14551), .A2(n10496), .ZN(n10454) );
  INV_X1 U12342 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14550) );
  NAND2_X1 U12343 ( .A1(n10505), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n10451) );
  NAND2_X1 U12344 ( .A1(n10507), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n10450) );
  OAI211_X1 U12345 ( .C1(n14550), .C2(n10499), .A(n10451), .B(n10450), .ZN(
        n10452) );
  INV_X1 U12346 ( .A(n10452), .ZN(n10453) );
  NAND2_X1 U12347 ( .A1(n10454), .A2(n10453), .ZN(n14454) );
  INV_X1 U12348 ( .A(n14454), .ZN(n14567) );
  NAND2_X1 U12349 ( .A1(n10455), .A2(n14567), .ZN(n10457) );
  INV_X1 U12350 ( .A(n10460), .ZN(n10458) );
  NAND2_X1 U12351 ( .A1(n10458), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n10470) );
  INV_X1 U12352 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10459) );
  NAND2_X1 U12353 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  NAND2_X1 U12354 ( .A1(n10470), .A2(n10461), .ZN(n14384) );
  OR2_X1 U12355 ( .A1(n14384), .A2(n10496), .ZN(n10467) );
  INV_X1 U12356 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10464) );
  NAND2_X1 U12357 ( .A1(n10505), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n10463) );
  NAND2_X1 U12358 ( .A1(n10507), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n10462) );
  OAI211_X1 U12359 ( .C1(n10464), .C2(n10499), .A(n10463), .B(n10462), .ZN(
        n10465) );
  INV_X1 U12360 ( .A(n10465), .ZN(n10466) );
  OR2_X1 U12361 ( .A1(n14768), .A2(n14559), .ZN(n10468) );
  NAND2_X1 U12362 ( .A1(n10469), .A2(n10468), .ZN(n14518) );
  INV_X1 U12363 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n14441) );
  NAND2_X1 U12364 ( .A1(n10470), .A2(n14441), .ZN(n10471) );
  NAND2_X1 U12365 ( .A1(n14524), .A2(n10483), .ZN(n10476) );
  INV_X1 U12366 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U12367 ( .A1(n10507), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U12368 ( .A1(n10505), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n10472) );
  OAI211_X1 U12369 ( .C1(n10499), .C2(n14526), .A(n10473), .B(n10472), .ZN(
        n10474) );
  INV_X1 U12370 ( .A(n10474), .ZN(n10475) );
  NAND2_X1 U12371 ( .A1(n10476), .A2(n10475), .ZN(n14453) );
  INV_X1 U12372 ( .A(n14453), .ZN(n14340) );
  NAND2_X1 U12373 ( .A1(n14518), .A2(n14529), .ZN(n10478) );
  NAND2_X1 U12374 ( .A1(n14705), .A2(n14340), .ZN(n10477) );
  NAND2_X1 U12375 ( .A1(n10478), .A2(n10477), .ZN(n14504) );
  XNOR2_X1 U12376 ( .A(n10487), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14509) );
  INV_X1 U12377 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U12378 ( .A1(n10505), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n10480) );
  NAND2_X1 U12379 ( .A1(n10507), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n10479) );
  OAI211_X1 U12380 ( .C1(n10481), .C2(n10499), .A(n10480), .B(n10479), .ZN(
        n10482) );
  INV_X1 U12381 ( .A(n14440), .ZN(n14452) );
  OR2_X1 U12382 ( .A1(n14511), .A2(n14452), .ZN(n10484) );
  INV_X1 U12383 ( .A(n10487), .ZN(n10486) );
  AND2_X1 U12384 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n10485) );
  NAND2_X1 U12385 ( .A1(n10486), .A2(n10485), .ZN(n13096) );
  INV_X1 U12386 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n14341) );
  INV_X1 U12387 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n14374) );
  OAI21_X1 U12388 ( .B1(n10487), .B2(n14341), .A(n14374), .ZN(n10488) );
  NAND2_X1 U12389 ( .A1(n13096), .A2(n10488), .ZN(n14495) );
  INV_X1 U12390 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n14494) );
  NAND2_X1 U12391 ( .A1(n10507), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U12392 ( .A1(n10505), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n10489) );
  OAI211_X1 U12393 ( .C1(n10499), .C2(n14494), .A(n10490), .B(n10489), .ZN(
        n10491) );
  INV_X1 U12394 ( .A(n10491), .ZN(n10492) );
  NAND2_X1 U12395 ( .A1(n14695), .A2(n14369), .ZN(n10494) );
  NAND2_X1 U12396 ( .A1(n14488), .A2(n10495), .ZN(n10503) );
  OR2_X1 U12397 ( .A1(n13096), .A2(n10496), .ZN(n10502) );
  INV_X1 U12398 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13095) );
  NAND2_X1 U12399 ( .A1(n10505), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n10498) );
  NAND2_X1 U12400 ( .A1(n10507), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n10497) );
  OAI211_X1 U12401 ( .C1(n13095), .C2(n10499), .A(n10498), .B(n10497), .ZN(
        n10500) );
  INV_X1 U12402 ( .A(n10500), .ZN(n10501) );
  XNOR2_X1 U12403 ( .A(n13098), .B(n14450), .ZN(n10817) );
  OR2_X1 U12404 ( .A1(n12987), .A2(n10842), .ZN(n10795) );
  NAND2_X1 U12405 ( .A1(n10930), .A2(n10825), .ZN(n10504) );
  NAND2_X1 U12406 ( .A1(n10925), .A2(n11102), .ZN(n14652) );
  NAND2_X1 U12407 ( .A1(n10505), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n10510) );
  NAND2_X1 U12408 ( .A1(n10506), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n10509) );
  NAND2_X1 U12409 ( .A1(n10507), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n10508) );
  AND3_X1 U12410 ( .A1(n10510), .A2(n10509), .A3(n10508), .ZN(n10755) );
  OAI22_X1 U12411 ( .A1(n14369), .A2(n14652), .B1(n10755), .B2(n10511), .ZN(
        n10512) );
  AND2_X1 U12412 ( .A1(n14475), .A2(n16106), .ZN(n11756) );
  INV_X1 U12413 ( .A(n10807), .ZN(n16216) );
  NAND2_X1 U12414 ( .A1(n16212), .A2(n16216), .ZN(n10515) );
  NAND2_X1 U12415 ( .A1(n16214), .A2(n10513), .ZN(n10514) );
  NAND2_X1 U12416 ( .A1(n10515), .A2(n10514), .ZN(n16252) );
  NAND2_X1 U12417 ( .A1(n16252), .A2(n16254), .ZN(n10517) );
  OR2_X1 U12418 ( .A1(n16270), .A2(n14471), .ZN(n10516) );
  NAND2_X1 U12419 ( .A1(n10517), .A2(n10516), .ZN(n11851) );
  INV_X1 U12420 ( .A(n11856), .ZN(n10518) );
  NAND2_X1 U12421 ( .A1(n11851), .A2(n10518), .ZN(n10520) );
  OR2_X1 U12422 ( .A1(n11853), .A2(n14470), .ZN(n10519) );
  NAND2_X1 U12423 ( .A1(n12101), .A2(n14469), .ZN(n10521) );
  OR2_X1 U12424 ( .A1(n11906), .A2(n14468), .ZN(n10522) );
  XNOR2_X1 U12425 ( .A(n12086), .B(n11505), .ZN(n12088) );
  NAND2_X1 U12426 ( .A1(n16360), .A2(n11505), .ZN(n10523) );
  INV_X1 U12427 ( .A(n11895), .ZN(n10524) );
  NAND2_X1 U12428 ( .A1(n12058), .A2(n14466), .ZN(n10525) );
  INV_X1 U12429 ( .A(n16400), .ZN(n12206) );
  OR2_X1 U12430 ( .A1(n12037), .A2(n14464), .ZN(n10804) );
  NAND2_X1 U12431 ( .A1(n12216), .A2(n10804), .ZN(n10526) );
  NAND2_X1 U12432 ( .A1(n12037), .A2(n14464), .ZN(n10803) );
  NAND2_X1 U12433 ( .A1(n10526), .A2(n10803), .ZN(n12256) );
  NAND2_X1 U12434 ( .A1(n12256), .A2(n12255), .ZN(n12257) );
  NAND2_X1 U12435 ( .A1(n12254), .A2(n14463), .ZN(n10527) );
  OR2_X1 U12436 ( .A1(n14677), .A2(n14462), .ZN(n10528) );
  NAND2_X1 U12437 ( .A1(n12422), .A2(n10528), .ZN(n10530) );
  NAND2_X1 U12438 ( .A1(n14677), .A2(n14462), .ZN(n10529) );
  NAND2_X1 U12439 ( .A1(n10530), .A2(n10529), .ZN(n12492) );
  NAND2_X1 U12440 ( .A1(n12492), .A2(n12495), .ZN(n10532) );
  NAND2_X1 U12441 ( .A1(n12504), .A2(n12400), .ZN(n10531) );
  XNOR2_X1 U12442 ( .A(n14666), .B(n14461), .ZN(n12660) );
  INV_X1 U12443 ( .A(n12660), .ZN(n12666) );
  NAND2_X1 U12444 ( .A1(n14666), .A2(n14461), .ZN(n10533) );
  OR2_X1 U12445 ( .A1(n12902), .A2(n14460), .ZN(n10535) );
  OR2_X1 U12446 ( .A1(n14791), .A2(n14458), .ZN(n10536) );
  NAND2_X1 U12447 ( .A1(n14788), .A2(n14360), .ZN(n10537) );
  NAND2_X1 U12448 ( .A1(n14742), .A2(n14457), .ZN(n10539) );
  AND2_X1 U12449 ( .A1(n14739), .A2(n14629), .ZN(n10540) );
  NOR2_X1 U12450 ( .A1(n14732), .A2(n14456), .ZN(n10541) );
  NAND2_X1 U12451 ( .A1(n14585), .A2(n14455), .ZN(n10542) );
  NAND2_X1 U12452 ( .A1(n14721), .A2(n14558), .ZN(n10544) );
  NAND2_X1 U12453 ( .A1(n10545), .A2(n10544), .ZN(n14547) );
  NAND2_X1 U12454 ( .A1(n14547), .A2(n14557), .ZN(n10547) );
  NAND2_X1 U12455 ( .A1(n10455), .A2(n14454), .ZN(n10546) );
  NOR2_X1 U12456 ( .A1(n14768), .A2(n14439), .ZN(n10549) );
  NAND2_X1 U12457 ( .A1(n14768), .A2(n14439), .ZN(n10548) );
  NAND2_X1 U12458 ( .A1(n14705), .A2(n14453), .ZN(n10550) );
  OR2_X1 U12459 ( .A1(n14511), .A2(n14440), .ZN(n10551) );
  NAND2_X1 U12460 ( .A1(n10844), .A2(n12987), .ZN(n10554) );
  NAND3_X1 U12461 ( .A1(n10554), .A2(n12843), .A3(n10831), .ZN(n16431) );
  NAND2_X1 U12462 ( .A1(n8334), .A2(n12987), .ZN(n16430) );
  NAND2_X1 U12463 ( .A1(n16431), .A2(n16430), .ZN(n14751) );
  AOI21_X1 U12464 ( .B1(n14490), .B2(n13098), .A(n14491), .ZN(n10555) );
  NAND2_X1 U12465 ( .A1(n10555), .A2(n14480), .ZN(n13100) );
  INV_X1 U12466 ( .A(n15570), .ZN(n10924) );
  INV_X1 U12467 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10557) );
  NAND2_X1 U12468 ( .A1(n14686), .A2(n10557), .ZN(n10558) );
  NAND2_X1 U12469 ( .A1(n16512), .A2(n16265), .ZN(n14750) );
  NAND2_X1 U12470 ( .A1(n10560), .A2(n10559), .ZN(P2_U3528) );
  NAND2_X1 U12471 ( .A1(n10563), .A2(n10562), .ZN(n10565) );
  NAND2_X1 U12472 ( .A1(n13098), .A2(n14792), .ZN(n10564) );
  NAND2_X1 U12473 ( .A1(n10565), .A2(n10564), .ZN(P2_U3496) );
  AND2_X1 U12474 ( .A1(n10795), .A2(n10835), .ZN(n10566) );
  OAI21_X1 U12475 ( .B1(n16106), .B2(n10566), .A(n11753), .ZN(n10567) );
  NAND2_X1 U12476 ( .A1(n14475), .A2(n10567), .ZN(n10570) );
  OAI21_X1 U12477 ( .B1(n16106), .B2(n10844), .A(n10568), .ZN(n10569) );
  OAI211_X1 U12478 ( .C1(n14475), .C2(n10760), .A(n10570), .B(n10569), .ZN(
        n10579) );
  INV_X1 U12479 ( .A(n10641), .ZN(n10758) );
  AOI22_X1 U12480 ( .A1(n10571), .A2(n10641), .B1(n11752), .B2(n10758), .ZN(
        n10578) );
  NAND2_X1 U12481 ( .A1(n10571), .A2(n10758), .ZN(n10573) );
  INV_X4 U12482 ( .A(n10577), .ZN(n10747) );
  NAND2_X1 U12483 ( .A1(n11752), .A2(n10747), .ZN(n10572) );
  NAND2_X1 U12484 ( .A1(n10573), .A2(n10572), .ZN(n10574) );
  OAI21_X1 U12485 ( .B1(n10579), .B2(n10578), .A(n10574), .ZN(n10582) );
  NAND2_X1 U12486 ( .A1(n16225), .A2(n10747), .ZN(n10576) );
  NAND2_X1 U12487 ( .A1(n14472), .A2(n10760), .ZN(n10575) );
  NAND2_X1 U12488 ( .A1(n10576), .A2(n10575), .ZN(n10583) );
  NAND2_X1 U12489 ( .A1(n10583), .A2(n10584), .ZN(n10581) );
  NAND2_X1 U12490 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  NAND3_X1 U12491 ( .A1(n10582), .A2(n10581), .A3(n10580), .ZN(n10588) );
  INV_X1 U12492 ( .A(n10583), .ZN(n10586) );
  INV_X1 U12493 ( .A(n10584), .ZN(n10585) );
  NAND2_X1 U12494 ( .A1(n10586), .A2(n10585), .ZN(n10587) );
  NAND2_X1 U12495 ( .A1(n10588), .A2(n10587), .ZN(n10594) );
  NAND2_X1 U12496 ( .A1(n16270), .A2(n10789), .ZN(n10590) );
  NAND2_X1 U12497 ( .A1(n14471), .A2(n10747), .ZN(n10589) );
  NAND2_X1 U12498 ( .A1(n10590), .A2(n10589), .ZN(n10595) );
  NAND2_X1 U12499 ( .A1(n10594), .A2(n10595), .ZN(n10593) );
  CLKBUF_X3 U12500 ( .A(n10641), .Z(n10759) );
  AOI22_X1 U12501 ( .A1(n16270), .A2(n10759), .B1(n14471), .B2(n10758), .ZN(
        n10591) );
  INV_X1 U12502 ( .A(n10591), .ZN(n10592) );
  NAND2_X1 U12503 ( .A1(n10593), .A2(n10592), .ZN(n10599) );
  NAND2_X1 U12504 ( .A1(n10597), .A2(n10596), .ZN(n10598) );
  NAND2_X1 U12505 ( .A1(n11853), .A2(n10747), .ZN(n10601) );
  NAND2_X1 U12506 ( .A1(n14470), .A2(n10789), .ZN(n10600) );
  NAND2_X1 U12507 ( .A1(n10601), .A2(n10600), .ZN(n10606) );
  AND2_X1 U12508 ( .A1(n14469), .A2(n10767), .ZN(n10602) );
  NAND2_X1 U12509 ( .A1(n12101), .A2(n10789), .ZN(n10604) );
  NAND2_X1 U12510 ( .A1(n14469), .A2(n10747), .ZN(n10603) );
  NAND2_X1 U12511 ( .A1(n10604), .A2(n10603), .ZN(n10607) );
  AOI22_X1 U12512 ( .A1(n11853), .A2(n10767), .B1(n10759), .B2(n14470), .ZN(
        n10605) );
  INV_X1 U12513 ( .A(n10607), .ZN(n10610) );
  INV_X1 U12514 ( .A(n10608), .ZN(n10609) );
  NAND2_X1 U12515 ( .A1(n10610), .A2(n10609), .ZN(n10611) );
  NAND2_X1 U12516 ( .A1(n10612), .A2(n10611), .ZN(n10618) );
  NAND2_X1 U12517 ( .A1(n11906), .A2(n10759), .ZN(n10614) );
  NAND2_X1 U12518 ( .A1(n14468), .A2(n10789), .ZN(n10613) );
  NAND2_X1 U12519 ( .A1(n10614), .A2(n10613), .ZN(n10619) );
  NAND2_X1 U12520 ( .A1(n10618), .A2(n10619), .ZN(n10617) );
  AOI22_X1 U12521 ( .A1(n11906), .A2(n10767), .B1(n10759), .B2(n14468), .ZN(
        n10615) );
  INV_X1 U12522 ( .A(n10615), .ZN(n10616) );
  NAND2_X1 U12523 ( .A1(n10617), .A2(n10616), .ZN(n10623) );
  INV_X1 U12524 ( .A(n10618), .ZN(n10621) );
  INV_X1 U12525 ( .A(n10619), .ZN(n10620) );
  NAND2_X1 U12526 ( .A1(n10621), .A2(n10620), .ZN(n10622) );
  NAND2_X1 U12527 ( .A1(n12086), .A2(n10789), .ZN(n10625) );
  NAND2_X1 U12528 ( .A1(n14467), .A2(n10759), .ZN(n10624) );
  NAND2_X1 U12529 ( .A1(n12086), .A2(n10759), .ZN(n10626) );
  OAI21_X1 U12530 ( .B1(n11505), .B2(n10759), .A(n10626), .ZN(n10627) );
  NAND2_X1 U12531 ( .A1(n12058), .A2(n10759), .ZN(n10629) );
  NAND2_X1 U12532 ( .A1(n14466), .A2(n10789), .ZN(n10628) );
  NAND2_X1 U12533 ( .A1(n10629), .A2(n10628), .ZN(n10631) );
  AOI22_X1 U12534 ( .A1(n12058), .A2(n10767), .B1(n10759), .B2(n14466), .ZN(
        n10630) );
  NAND2_X1 U12535 ( .A1(n16400), .A2(n10789), .ZN(n10635) );
  NAND2_X1 U12536 ( .A1(n14465), .A2(n10759), .ZN(n10634) );
  NAND2_X1 U12537 ( .A1(n10635), .A2(n10634), .ZN(n10638) );
  AOI22_X1 U12538 ( .A1(n16400), .A2(n10759), .B1(n14465), .B2(n10758), .ZN(
        n10636) );
  INV_X1 U12539 ( .A(n10636), .ZN(n10637) );
  NAND2_X1 U12540 ( .A1(n12037), .A2(n10747), .ZN(n10640) );
  NAND2_X1 U12541 ( .A1(n14464), .A2(n10767), .ZN(n10639) );
  NAND2_X1 U12542 ( .A1(n10640), .A2(n10639), .ZN(n10646) );
  NAND2_X1 U12543 ( .A1(n10645), .A2(n10646), .ZN(n10644) );
  INV_X1 U12544 ( .A(n10641), .ZN(n10789) );
  NAND2_X1 U12545 ( .A1(n12037), .A2(n10767), .ZN(n10642) );
  NAND2_X1 U12546 ( .A1(n10644), .A2(n10643), .ZN(n10650) );
  INV_X1 U12547 ( .A(n10645), .ZN(n10648) );
  INV_X1 U12548 ( .A(n10646), .ZN(n10647) );
  NAND2_X1 U12549 ( .A1(n10648), .A2(n10647), .ZN(n10649) );
  NAND2_X1 U12550 ( .A1(n12254), .A2(n10767), .ZN(n10652) );
  NAND2_X1 U12551 ( .A1(n14463), .A2(n10759), .ZN(n10651) );
  NAND2_X1 U12552 ( .A1(n10652), .A2(n10651), .ZN(n10655) );
  AOI22_X1 U12553 ( .A1(n12254), .A2(n10759), .B1(n14463), .B2(n10789), .ZN(
        n10653) );
  AOI21_X1 U12554 ( .B1(n10656), .B2(n10655), .A(n10653), .ZN(n10654) );
  INV_X1 U12555 ( .A(n10654), .ZN(n10657) );
  NAND2_X1 U12556 ( .A1(n14677), .A2(n10747), .ZN(n10659) );
  NAND2_X1 U12557 ( .A1(n14462), .A2(n10767), .ZN(n10658) );
  NAND2_X1 U12558 ( .A1(n10659), .A2(n10658), .ZN(n10662) );
  NAND2_X1 U12559 ( .A1(n14677), .A2(n10767), .ZN(n10660) );
  OAI21_X1 U12560 ( .B1(n12246), .B2(n10789), .A(n10660), .ZN(n10661) );
  INV_X1 U12561 ( .A(n10662), .ZN(n10663) );
  NAND2_X1 U12562 ( .A1(n12504), .A2(n10767), .ZN(n10665) );
  NAND2_X1 U12563 ( .A1(n12400), .A2(n10759), .ZN(n10664) );
  NAND2_X1 U12564 ( .A1(n10665), .A2(n10664), .ZN(n10670) );
  NAND2_X1 U12565 ( .A1(n10669), .A2(n10670), .ZN(n10668) );
  AOI22_X1 U12566 ( .A1(n12504), .A2(n10759), .B1(n12400), .B2(n10758), .ZN(
        n10666) );
  INV_X1 U12567 ( .A(n10666), .ZN(n10667) );
  NAND2_X1 U12568 ( .A1(n10668), .A2(n10667), .ZN(n10674) );
  INV_X1 U12569 ( .A(n10669), .ZN(n10672) );
  NAND2_X1 U12570 ( .A1(n10672), .A2(n10671), .ZN(n10673) );
  NAND2_X1 U12571 ( .A1(n14666), .A2(n10759), .ZN(n10676) );
  NAND2_X1 U12572 ( .A1(n14461), .A2(n10767), .ZN(n10675) );
  NAND2_X1 U12573 ( .A1(n14666), .A2(n10767), .ZN(n10677) );
  OAI21_X1 U12574 ( .B1(n10678), .B2(n10789), .A(n10677), .ZN(n10679) );
  INV_X1 U12575 ( .A(n10685), .ZN(n10683) );
  NAND2_X1 U12576 ( .A1(n12902), .A2(n10767), .ZN(n10681) );
  NAND2_X1 U12577 ( .A1(n14460), .A2(n10759), .ZN(n10680) );
  NAND2_X1 U12578 ( .A1(n10681), .A2(n10680), .ZN(n10684) );
  INV_X1 U12579 ( .A(n10684), .ZN(n10682) );
  NAND2_X1 U12580 ( .A1(n10685), .A2(n10684), .ZN(n10688) );
  AOI22_X1 U12581 ( .A1(n12902), .A2(n10759), .B1(n14460), .B2(n10758), .ZN(
        n10686) );
  INV_X1 U12582 ( .A(n10686), .ZN(n10687) );
  NAND2_X1 U12583 ( .A1(n10688), .A2(n10687), .ZN(n10689) );
  NAND2_X1 U12584 ( .A1(n10690), .A2(n10689), .ZN(n10695) );
  NAND2_X1 U12585 ( .A1(n12795), .A2(n10759), .ZN(n10692) );
  NAND2_X1 U12586 ( .A1(n14459), .A2(n10767), .ZN(n10691) );
  NAND2_X1 U12587 ( .A1(n10692), .A2(n10691), .ZN(n10694) );
  AOI22_X1 U12588 ( .A1(n12795), .A2(n10767), .B1(n10759), .B2(n14459), .ZN(
        n10693) );
  NOR2_X1 U12589 ( .A1(n10695), .A2(n10694), .ZN(n10696) );
  NAND2_X1 U12590 ( .A1(n14791), .A2(n10767), .ZN(n10698) );
  NAND2_X1 U12591 ( .A1(n14458), .A2(n10759), .ZN(n10697) );
  NAND2_X1 U12592 ( .A1(n14791), .A2(n10759), .ZN(n10700) );
  NAND2_X1 U12593 ( .A1(n14458), .A2(n10789), .ZN(n10699) );
  NAND2_X1 U12594 ( .A1(n10700), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U12595 ( .A1(n14645), .A2(n10759), .ZN(n10703) );
  NAND2_X1 U12596 ( .A1(n14626), .A2(n10767), .ZN(n10702) );
  NAND2_X1 U12597 ( .A1(n10703), .A2(n10702), .ZN(n10705) );
  AOI22_X1 U12598 ( .A1(n7745), .A2(n10767), .B1(n10759), .B2(n14626), .ZN(
        n10704) );
  AOI21_X1 U12599 ( .B1(n10706), .B2(n10705), .A(n10704), .ZN(n10708) );
  NOR2_X1 U12600 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  NAND2_X1 U12601 ( .A1(n14742), .A2(n10789), .ZN(n10710) );
  NAND2_X1 U12602 ( .A1(n14457), .A2(n10747), .ZN(n10709) );
  NAND2_X1 U12603 ( .A1(n14742), .A2(n10759), .ZN(n10712) );
  NAND2_X1 U12604 ( .A1(n14457), .A2(n10789), .ZN(n10711) );
  NAND2_X1 U12605 ( .A1(n10712), .A2(n10711), .ZN(n10713) );
  NAND2_X1 U12606 ( .A1(n14739), .A2(n10759), .ZN(n10715) );
  NAND2_X1 U12607 ( .A1(n14629), .A2(n10767), .ZN(n10714) );
  NAND2_X1 U12608 ( .A1(n10715), .A2(n10714), .ZN(n10718) );
  AOI22_X1 U12609 ( .A1(n14739), .A2(n10767), .B1(n10747), .B2(n14629), .ZN(
        n10716) );
  AOI21_X1 U12610 ( .B1(n10719), .B2(n10718), .A(n10716), .ZN(n10717) );
  INV_X1 U12611 ( .A(n10717), .ZN(n10720) );
  NAND2_X1 U12612 ( .A1(n14732), .A2(n10767), .ZN(n10722) );
  NAND2_X1 U12613 ( .A1(n14456), .A2(n10759), .ZN(n10721) );
  NAND2_X1 U12614 ( .A1(n10722), .A2(n10721), .ZN(n10728) );
  NAND2_X1 U12615 ( .A1(n10727), .A2(n10728), .ZN(n10726) );
  NAND2_X1 U12616 ( .A1(n14732), .A2(n10759), .ZN(n10724) );
  NAND2_X1 U12617 ( .A1(n14456), .A2(n10767), .ZN(n10723) );
  NAND2_X1 U12618 ( .A1(n10724), .A2(n10723), .ZN(n10725) );
  INV_X1 U12619 ( .A(n10727), .ZN(n10730) );
  INV_X1 U12620 ( .A(n10728), .ZN(n10729) );
  NAND2_X1 U12621 ( .A1(n14585), .A2(n10759), .ZN(n10732) );
  NAND2_X1 U12622 ( .A1(n14455), .A2(n10767), .ZN(n10731) );
  NAND2_X1 U12623 ( .A1(n10732), .A2(n10731), .ZN(n10734) );
  AOI22_X1 U12624 ( .A1(n14585), .A2(n10767), .B1(n10759), .B2(n14455), .ZN(
        n10733) );
  NAND2_X1 U12625 ( .A1(n14721), .A2(n10767), .ZN(n10736) );
  NAND2_X1 U12626 ( .A1(n14558), .A2(n10759), .ZN(n10735) );
  NAND2_X1 U12627 ( .A1(n10736), .A2(n10735), .ZN(n10738) );
  NAND2_X1 U12628 ( .A1(n10739), .A2(n10738), .ZN(n10741) );
  AOI22_X1 U12629 ( .A1(n14721), .A2(n10747), .B1(n14558), .B2(n10758), .ZN(
        n10737) );
  INV_X1 U12630 ( .A(n10737), .ZN(n10740) );
  AOI22_X1 U12631 ( .A1(n10455), .A2(n10759), .B1(n14454), .B2(n10758), .ZN(
        n10742) );
  AOI22_X1 U12632 ( .A1(n10455), .A2(n10767), .B1(n10759), .B2(n14454), .ZN(
        n10743) );
  AOI22_X1 U12633 ( .A1(n7754), .A2(n10747), .B1(n14559), .B2(n10758), .ZN(
        n10744) );
  NOR2_X1 U12634 ( .A1(n10746), .A2(n10745), .ZN(n10753) );
  AOI22_X1 U12635 ( .A1(n14700), .A2(n10767), .B1(n10759), .B2(n14452), .ZN(
        n10768) );
  OAI22_X1 U12636 ( .A1(n14511), .A2(n10789), .B1(n14440), .B2(n10759), .ZN(
        n10770) );
  NAND2_X1 U12637 ( .A1(n14705), .A2(n10747), .ZN(n10749) );
  NAND2_X1 U12638 ( .A1(n14453), .A2(n10767), .ZN(n10748) );
  NAND2_X1 U12639 ( .A1(n10749), .A2(n10748), .ZN(n10763) );
  AND2_X1 U12640 ( .A1(n14453), .A2(n10759), .ZN(n10750) );
  AOI21_X1 U12641 ( .B1(n14705), .B2(n10767), .A(n10750), .ZN(n10764) );
  OAI21_X1 U12642 ( .B1(n10754), .B2(n10753), .A(n10752), .ZN(n10773) );
  OAI22_X1 U12643 ( .A1(n8926), .A2(n10759), .B1(n10755), .B2(n10789), .ZN(
        n10784) );
  INV_X1 U12644 ( .A(n10755), .ZN(n14449) );
  NAND2_X1 U12645 ( .A1(n11026), .A2(n10767), .ZN(n10790) );
  INV_X1 U12646 ( .A(n10795), .ZN(n10797) );
  NAND2_X1 U12647 ( .A1(n10797), .A2(n12739), .ZN(n10756) );
  NAND4_X1 U12648 ( .A1(n10790), .A2(n10825), .A3(n10835), .A4(n10756), .ZN(
        n10757) );
  AOI22_X1 U12649 ( .A1(n14691), .A2(n10759), .B1(n14449), .B2(n10757), .ZN(
        n10783) );
  AOI22_X1 U12650 ( .A1(n13098), .A2(n10759), .B1(n14450), .B2(n10758), .ZN(
        n10774) );
  OAI22_X1 U12651 ( .A1(n10761), .A2(n10759), .B1(n14373), .B2(n10760), .ZN(
        n10775) );
  OAI22_X1 U12652 ( .A1(n10784), .A2(n10783), .B1(n10774), .B2(n10775), .ZN(
        n10762) );
  XNOR2_X1 U12653 ( .A(n14687), .B(n11026), .ZN(n10822) );
  NAND2_X1 U12654 ( .A1(n10762), .A2(n10822), .ZN(n10780) );
  INV_X1 U12655 ( .A(n10763), .ZN(n10766) );
  INV_X1 U12656 ( .A(n10764), .ZN(n10765) );
  NOR2_X1 U12657 ( .A1(n10766), .A2(n10765), .ZN(n10769) );
  INV_X1 U12658 ( .A(n14369), .ZN(n14451) );
  AOI22_X1 U12659 ( .A1(n14695), .A2(n10767), .B1(n10759), .B2(n14451), .ZN(
        n10777) );
  OAI22_X1 U12660 ( .A1(n14493), .A2(n10789), .B1(n14369), .B2(n10759), .ZN(
        n10776) );
  AOI22_X1 U12661 ( .A1(n10770), .A2(n10769), .B1(n10777), .B2(n10776), .ZN(
        n10772) );
  OAI21_X1 U12662 ( .B1(n10770), .B2(n10769), .A(n10768), .ZN(n10771) );
  NAND2_X1 U12663 ( .A1(n10773), .A2(n8341), .ZN(n10788) );
  INV_X1 U12664 ( .A(n10822), .ZN(n10782) );
  INV_X1 U12665 ( .A(n10774), .ZN(n10779) );
  INV_X1 U12666 ( .A(n10775), .ZN(n10778) );
  OAI22_X1 U12667 ( .A1(n10779), .A2(n10778), .B1(n10777), .B2(n10776), .ZN(
        n10781) );
  OAI21_X1 U12668 ( .B1(n10782), .B2(n10781), .A(n10780), .ZN(n10786) );
  NAND2_X1 U12669 ( .A1(n10788), .A2(n10787), .ZN(n10794) );
  NAND2_X1 U12670 ( .A1(n11026), .A2(n10759), .ZN(n10792) );
  NAND2_X1 U12671 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  MUX2_X1 U12672 ( .A(n10792), .B(n10791), .S(n14687), .Z(n10793) );
  NAND2_X1 U12673 ( .A1(n10794), .A2(n10793), .ZN(n10828) );
  AOI22_X1 U12674 ( .A1(n12849), .A2(n10844), .B1(n10930), .B2(n12877), .ZN(
        n10796) );
  OAI211_X1 U12675 ( .C1(n10797), .C2(n10930), .A(n10825), .B(n12849), .ZN(
        n10798) );
  NAND2_X1 U12676 ( .A1(n10828), .A2(n10798), .ZN(n10800) );
  INV_X1 U12677 ( .A(n10935), .ZN(n10832) );
  NAND2_X1 U12678 ( .A1(n10832), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13010) );
  INV_X1 U12679 ( .A(n13010), .ZN(n10799) );
  OAI211_X1 U12680 ( .C1(n10828), .C2(n8332), .A(n10800), .B(n10799), .ZN(
        n10839) );
  XNOR2_X1 U12681 ( .A(n14691), .B(n14449), .ZN(n10819) );
  NOR2_X1 U12682 ( .A1(n10802), .A2(n10801), .ZN(n14593) );
  NAND2_X1 U12683 ( .A1(n10804), .A2(n10803), .ZN(n12217) );
  INV_X1 U12684 ( .A(n16106), .ZN(n11404) );
  NAND2_X1 U12685 ( .A1(n14475), .A2(n11404), .ZN(n10805) );
  AND2_X1 U12686 ( .A1(n10806), .A2(n10805), .ZN(n16111) );
  NAND4_X1 U12687 ( .A1(n10807), .A2(n16111), .A3(n10930), .A4(n11757), .ZN(
        n10808) );
  NOR2_X1 U12688 ( .A1(n16254), .A2(n10808), .ZN(n10809) );
  XNOR2_X1 U12689 ( .A(n12101), .B(n14469), .ZN(n12103) );
  NAND4_X1 U12690 ( .A1(n11856), .A2(n10809), .A3(n11456), .A4(n12103), .ZN(
        n10810) );
  NOR2_X1 U12691 ( .A1(n12088), .A2(n10810), .ZN(n10811) );
  NAND4_X1 U12692 ( .A1(n12217), .A2(n12198), .A3(n10811), .A4(n11895), .ZN(
        n10812) );
  NOR4_X1 U12693 ( .A1(n12495), .A2(n12255), .A3(n12427), .A4(n10812), .ZN(
        n10813) );
  NAND4_X1 U12694 ( .A1(n12742), .A2(n10813), .A3(n12660), .A4(n12627), .ZN(
        n10814) );
  NOR4_X1 U12695 ( .A1(n14606), .A2(n14650), .A3(n12942), .A4(n10814), .ZN(
        n10815) );
  NAND4_X1 U12696 ( .A1(n14583), .A2(n14593), .A3(n10815), .A4(n14623), .ZN(
        n10816) );
  NOR4_X1 U12697 ( .A1(n14499), .A2(n14557), .A3(n14569), .A4(n10816), .ZN(
        n10818) );
  NAND3_X1 U12698 ( .A1(n10819), .A2(n10818), .A3(n10817), .ZN(n10821) );
  XOR2_X1 U12699 ( .A(n14559), .B(n7754), .Z(n14538) );
  NAND2_X1 U12700 ( .A1(n10823), .A2(n10822), .ZN(n10824) );
  XOR2_X1 U12701 ( .A(n12849), .B(n10824), .Z(n10826) );
  OAI21_X1 U12702 ( .B1(n10828), .B2(n10930), .A(n10827), .ZN(n10838) );
  INV_X1 U12703 ( .A(n12987), .ZN(n10843) );
  AND2_X1 U12704 ( .A1(n10935), .A2(n10829), .ZN(n10840) );
  INV_X1 U12705 ( .A(n10840), .ZN(n10834) );
  OAI21_X1 U12706 ( .B1(n10832), .B2(n10831), .A(n10830), .ZN(n10833) );
  AND2_X1 U12707 ( .A1(n10834), .A2(n10833), .ZN(n11124) );
  AND2_X1 U12708 ( .A1(n11124), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15684) );
  INV_X1 U12709 ( .A(n10835), .ZN(n10939) );
  NAND4_X1 U12710 ( .A1(n15684), .A2(n11121), .A3(n11102), .A4(n10939), .ZN(
        n10836) );
  OAI211_X1 U12711 ( .C1(n10843), .C2(n13010), .A(n10836), .B(P2_B_REG_SCAN_IN), .ZN(n10837) );
  NAND3_X1 U12712 ( .A1(n10839), .A2(n10838), .A3(n10837), .ZN(P2_U3328) );
  INV_X1 U12713 ( .A(n10996), .ZN(n10841) );
  NAND2_X1 U12714 ( .A1(n10843), .A2(n10842), .ZN(n10845) );
  XNOR2_X1 U12715 ( .A(n14732), .B(n10854), .ZN(n14319) );
  NAND2_X1 U12716 ( .A1(n14456), .A2(n14491), .ZN(n14320) );
  XNOR2_X1 U12717 ( .A(n14319), .B(n14320), .ZN(n10929) );
  NAND2_X1 U12718 ( .A1(n14457), .A2(n14491), .ZN(n10918) );
  XNOR2_X1 U12719 ( .A(n14399), .B(n10918), .ZN(n14359) );
  AND2_X1 U12720 ( .A1(n14626), .A2(n14491), .ZN(n10846) );
  NAND2_X1 U12721 ( .A1(n14358), .A2(n10846), .ZN(n10848) );
  INV_X1 U12722 ( .A(n10848), .ZN(n10917) );
  XNOR2_X1 U12723 ( .A(n16400), .B(n10853), .ZN(n12031) );
  NAND2_X1 U12724 ( .A1(n14465), .A2(n14491), .ZN(n10885) );
  XNOR2_X1 U12725 ( .A(n12031), .B(n10885), .ZN(n11679) );
  XNOR2_X1 U12726 ( .A(n12058), .B(n10853), .ZN(n10881) );
  NAND2_X1 U12727 ( .A1(n14466), .A2(n14491), .ZN(n10882) );
  XNOR2_X1 U12728 ( .A(n10881), .B(n10882), .ZN(n11504) );
  XNOR2_X1 U12729 ( .A(n11853), .B(n10853), .ZN(n10864) );
  NAND2_X1 U12730 ( .A1(n14470), .A2(n14491), .ZN(n10865) );
  XNOR2_X1 U12731 ( .A(n10864), .B(n10865), .ZN(n11699) );
  XNOR2_X1 U12732 ( .A(n16270), .B(n10853), .ZN(n10849) );
  AND2_X1 U12733 ( .A1(n14471), .A2(n14491), .ZN(n10850) );
  NAND2_X1 U12734 ( .A1(n10849), .A2(n10850), .ZN(n10863) );
  INV_X1 U12735 ( .A(n10849), .ZN(n11696) );
  INV_X1 U12736 ( .A(n10850), .ZN(n10851) );
  NAND2_X1 U12737 ( .A1(n11696), .A2(n10851), .ZN(n10852) );
  NAND2_X1 U12738 ( .A1(n10863), .A2(n10852), .ZN(n10954) );
  XNOR2_X1 U12739 ( .A(n16225), .B(n10853), .ZN(n10859) );
  NAND2_X1 U12740 ( .A1(n14472), .A2(n14491), .ZN(n10860) );
  XNOR2_X1 U12741 ( .A(n10859), .B(n10860), .ZN(n11765) );
  XNOR2_X1 U12742 ( .A(n11752), .B(n10853), .ZN(n11763) );
  NAND2_X1 U12743 ( .A1(n14473), .A2(n14491), .ZN(n10856) );
  XNOR2_X1 U12744 ( .A(n11763), .B(n10856), .ZN(n11144) );
  NAND2_X1 U12745 ( .A1(n11756), .A2(n14491), .ZN(n11406) );
  NAND2_X1 U12746 ( .A1(n11404), .A2(n10854), .ZN(n10855) );
  AND2_X1 U12747 ( .A1(n11406), .A2(n10855), .ZN(n11145) );
  INV_X1 U12748 ( .A(n11763), .ZN(n10857) );
  NAND2_X1 U12749 ( .A1(n10857), .A2(n10856), .ZN(n10858) );
  INV_X1 U12750 ( .A(n10859), .ZN(n10861) );
  NAND2_X1 U12751 ( .A1(n10861), .A2(n10860), .ZN(n10862) );
  INV_X1 U12752 ( .A(n10864), .ZN(n11423) );
  NAND2_X1 U12753 ( .A1(n11423), .A2(n10865), .ZN(n10866) );
  NAND2_X1 U12754 ( .A1(n11704), .A2(n10866), .ZN(n10867) );
  XNOR2_X1 U12755 ( .A(n12101), .B(n10853), .ZN(n10868) );
  NAND2_X1 U12756 ( .A1(n14469), .A2(n14491), .ZN(n10869) );
  XNOR2_X1 U12757 ( .A(n10868), .B(n10869), .ZN(n11422) );
  INV_X1 U12758 ( .A(n10868), .ZN(n10870) );
  NAND2_X1 U12759 ( .A1(n10870), .A2(n10869), .ZN(n10871) );
  XNOR2_X1 U12760 ( .A(n11906), .B(n10853), .ZN(n10872) );
  AND2_X1 U12761 ( .A1(n14468), .A2(n14491), .ZN(n10873) );
  NAND2_X1 U12762 ( .A1(n10872), .A2(n10873), .ZN(n10876) );
  INV_X1 U12763 ( .A(n10872), .ZN(n11630) );
  INV_X1 U12764 ( .A(n10873), .ZN(n10874) );
  NAND2_X1 U12765 ( .A1(n11630), .A2(n10874), .ZN(n10875) );
  NAND2_X1 U12766 ( .A1(n10876), .A2(n10875), .ZN(n11654) );
  XNOR2_X1 U12767 ( .A(n12086), .B(n10853), .ZN(n10877) );
  NAND2_X1 U12768 ( .A1(n14467), .A2(n14491), .ZN(n10878) );
  XNOR2_X1 U12769 ( .A(n10877), .B(n10878), .ZN(n11641) );
  INV_X1 U12770 ( .A(n10877), .ZN(n11506) );
  NAND2_X1 U12771 ( .A1(n11506), .A2(n10878), .ZN(n10879) );
  NAND2_X1 U12772 ( .A1(n11504), .A2(n10880), .ZN(n11683) );
  INV_X1 U12773 ( .A(n10881), .ZN(n11681) );
  NAND2_X1 U12774 ( .A1(n11681), .A2(n10882), .ZN(n10883) );
  NAND2_X1 U12775 ( .A1(n11683), .A2(n10883), .ZN(n10884) );
  INV_X1 U12776 ( .A(n12031), .ZN(n10886) );
  NAND2_X1 U12777 ( .A1(n10886), .A2(n10885), .ZN(n10887) );
  XNOR2_X1 U12778 ( .A(n12037), .B(n10853), .ZN(n10888) );
  NAND2_X1 U12779 ( .A1(n14464), .A2(n14491), .ZN(n10889) );
  XNOR2_X1 U12780 ( .A(n10888), .B(n10889), .ZN(n12032) );
  INV_X1 U12781 ( .A(n10888), .ZN(n10890) );
  XNOR2_X1 U12782 ( .A(n12254), .B(n10853), .ZN(n10891) );
  AND2_X1 U12783 ( .A1(n14463), .A2(n14491), .ZN(n10892) );
  NAND2_X1 U12784 ( .A1(n10891), .A2(n10892), .ZN(n10895) );
  INV_X1 U12785 ( .A(n10891), .ZN(n12396) );
  INV_X1 U12786 ( .A(n10892), .ZN(n10893) );
  NAND2_X1 U12787 ( .A1(n12396), .A2(n10893), .ZN(n10894) );
  NAND2_X1 U12788 ( .A1(n10895), .A2(n10894), .ZN(n10946) );
  XNOR2_X1 U12789 ( .A(n14677), .B(n10853), .ZN(n12388) );
  NAND2_X1 U12790 ( .A1(n14462), .A2(n14491), .ZN(n10896) );
  XNOR2_X1 U12791 ( .A(n12388), .B(n10896), .ZN(n12407) );
  INV_X1 U12792 ( .A(n12388), .ZN(n10897) );
  NAND2_X1 U12793 ( .A1(n10897), .A2(n10896), .ZN(n10898) );
  XNOR2_X1 U12794 ( .A(n12504), .B(n10853), .ZN(n10899) );
  NAND2_X1 U12795 ( .A1(n12400), .A2(n14491), .ZN(n10900) );
  XNOR2_X1 U12796 ( .A(n10899), .B(n10900), .ZN(n12389) );
  INV_X1 U12797 ( .A(n10899), .ZN(n12379) );
  XNOR2_X1 U12798 ( .A(n14666), .B(n10853), .ZN(n10901) );
  NAND2_X1 U12799 ( .A1(n14461), .A2(n14491), .ZN(n10902) );
  XNOR2_X1 U12800 ( .A(n10901), .B(n10902), .ZN(n12378) );
  INV_X1 U12801 ( .A(n10901), .ZN(n10903) );
  XNOR2_X1 U12802 ( .A(n12902), .B(n10853), .ZN(n10904) );
  AND2_X1 U12803 ( .A1(n14460), .A2(n14491), .ZN(n10905) );
  NAND2_X1 U12804 ( .A1(n10904), .A2(n10905), .ZN(n10908) );
  INV_X1 U12805 ( .A(n10904), .ZN(n12787) );
  INV_X1 U12806 ( .A(n10905), .ZN(n10906) );
  NAND2_X1 U12807 ( .A1(n12787), .A2(n10906), .ZN(n10907) );
  NAND2_X1 U12808 ( .A1(n10908), .A2(n10907), .ZN(n12898) );
  XNOR2_X1 U12809 ( .A(n12795), .B(n10853), .ZN(n12907) );
  NAND2_X1 U12810 ( .A1(n14459), .A2(n14491), .ZN(n10909) );
  XNOR2_X1 U12811 ( .A(n12907), .B(n10909), .ZN(n12798) );
  NAND3_X1 U12812 ( .A1(n12785), .A2(n10908), .A3(n12798), .ZN(n12789) );
  INV_X1 U12813 ( .A(n12907), .ZN(n10910) );
  NAND2_X1 U12814 ( .A1(n10910), .A2(n10909), .ZN(n10911) );
  XNOR2_X1 U12815 ( .A(n14791), .B(n10853), .ZN(n10913) );
  NAND2_X1 U12816 ( .A1(n14458), .A2(n14491), .ZN(n10914) );
  XNOR2_X1 U12817 ( .A(n10913), .B(n10914), .ZN(n12909) );
  INV_X1 U12818 ( .A(n10913), .ZN(n10915) );
  NAND2_X1 U12819 ( .A1(n10915), .A2(n10914), .ZN(n10916) );
  XNOR2_X1 U12820 ( .A(n14739), .B(n10853), .ZN(n10919) );
  NAND2_X1 U12821 ( .A1(n14629), .A2(n14491), .ZN(n10920) );
  XNOR2_X1 U12822 ( .A(n10919), .B(n10920), .ZN(n14397) );
  INV_X1 U12823 ( .A(n10919), .ZN(n10921) );
  NAND2_X1 U12824 ( .A1(n10921), .A2(n10920), .ZN(n10922) );
  INV_X1 U12825 ( .A(n10923), .ZN(n11738) );
  NAND3_X1 U12826 ( .A1(n10924), .A2(n11739), .A3(n11738), .ZN(n10933) );
  NOR2_X1 U12827 ( .A1(n16265), .A2(n10925), .ZN(n10926) );
  INV_X1 U12828 ( .A(n14324), .ZN(n10927) );
  AOI211_X1 U12829 ( .C1(n10929), .C2(n10928), .A(n14427), .B(n10927), .ZN(
        n10944) );
  AND2_X1 U12830 ( .A1(n16105), .A2(n10930), .ZN(n11743) );
  NAND2_X1 U12831 ( .A1(n10940), .A2(n11743), .ZN(n10931) );
  INV_X1 U12832 ( .A(n14432), .ZN(n14448) );
  NOR2_X1 U12833 ( .A1(n7743), .A2(n14448), .ZN(n10943) );
  NAND2_X1 U12834 ( .A1(n10933), .A2(n10932), .ZN(n10937) );
  AND3_X1 U12835 ( .A1(n11736), .A2(n10935), .A3(n10934), .ZN(n10936) );
  NAND2_X1 U12836 ( .A1(n10937), .A2(n10936), .ZN(n11143) );
  OAI22_X1 U12837 ( .A1(n14442), .A2(n14599), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10938), .ZN(n10942) );
  NAND2_X1 U12838 ( .A1(n14445), .A2(n14627), .ZN(n14416) );
  NAND2_X1 U12839 ( .A1(n14445), .A2(n14628), .ZN(n14417) );
  OAI22_X1 U12840 ( .A1(n14596), .A2(n14416), .B1(n14417), .B2(n14597), .ZN(
        n10941) );
  OR4_X1 U12841 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        P2_U3195) );
  INV_X1 U12842 ( .A(n10945), .ZN(n12398) );
  AOI211_X1 U12843 ( .C1(n10947), .C2(n10946), .A(n14427), .B(n12398), .ZN(
        n10952) );
  INV_X1 U12844 ( .A(n12254), .ZN(n16459) );
  NOR2_X1 U12845 ( .A1(n16459), .A2(n14448), .ZN(n10951) );
  INV_X1 U12846 ( .A(n10948), .ZN(n12248) );
  OAI22_X1 U12847 ( .A1(n14442), .A2(n12248), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15610), .ZN(n10950) );
  OAI22_X1 U12848 ( .A1(n12246), .A2(n14417), .B1(n14416), .B2(n12247), .ZN(
        n10949) );
  OR4_X1 U12849 ( .A1(n10952), .A2(n10951), .A3(n10950), .A4(n10949), .ZN(
        P2_U3208) );
  MUX2_X1 U12850 ( .A(n14420), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n10959) );
  INV_X1 U12851 ( .A(n10953), .ZN(n11698) );
  AOI211_X1 U12852 ( .C1(n10955), .C2(n10954), .A(n14427), .B(n11698), .ZN(
        n10958) );
  INV_X1 U12853 ( .A(n16270), .ZN(n10956) );
  INV_X1 U12854 ( .A(n14445), .ZN(n14386) );
  AOI22_X1 U12855 ( .A1(n14627), .A2(n14472), .B1(n14470), .B2(n14628), .ZN(
        n16255) );
  OAI22_X1 U12856 ( .A1(n10956), .A2(n14448), .B1(n14386), .B2(n16255), .ZN(
        n10957) );
  OR3_X1 U12857 ( .A1(n10959), .A2(n10958), .A3(n10957), .ZN(P2_U3190) );
  MUX2_X1 U12858 ( .A(n10961), .B(n10960), .S(P3_STATE_REG_SCAN_IN), .Z(n10962) );
  INV_X1 U12859 ( .A(n10962), .ZN(P3_U3295) );
  AND2_X1 U12860 ( .A1(n10976), .A2(P3_U3151), .ZN(n12146) );
  INV_X2 U12861 ( .A(n12146), .ZN(n14312) );
  AND2_X1 U12862 ( .A1(n10984), .A2(P3_U3151), .ZN(n14310) );
  INV_X2 U12863 ( .A(n14310), .ZN(n14315) );
  OAI222_X1 U12864 ( .A1(n14312), .A2(n10963), .B1(n14315), .B2(n13711), .C1(
        n15992), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U12865 ( .A1(n10965), .A2(P3_U3151), .B1(n14312), .B2(n10964), 
        .C1(n13715), .C2(n14315), .ZN(P3_U3292) );
  INV_X1 U12866 ( .A(n10966), .ZN(n10967) );
  OAI222_X1 U12867 ( .A1(n7889), .A2(P3_U3151), .B1(n14312), .B2(n10967), .C1(
        n7839), .C2(n14315), .ZN(P3_U3294) );
  OAI222_X1 U12868 ( .A1(n15952), .A2(P3_U3151), .B1(n14312), .B2(n10968), 
        .C1(n13666), .C2(n14315), .ZN(P3_U3290) );
  INV_X1 U12869 ( .A(SI_2_), .ZN(n10969) );
  OAI222_X1 U12870 ( .A1(n7370), .A2(P3_U3151), .B1(n14312), .B2(n10970), .C1(
        n10969), .C2(n14315), .ZN(P3_U3293) );
  INV_X1 U12871 ( .A(SI_6_), .ZN(n10971) );
  OAI222_X1 U12872 ( .A1(n10973), .A2(P3_U3151), .B1(n14312), .B2(n10972), 
        .C1(n10971), .C2(n14315), .ZN(P3_U3289) );
  OAI222_X1 U12873 ( .A1(n15932), .A2(P3_U3151), .B1(n14312), .B2(n10974), 
        .C1(n7656), .C2(n14315), .ZN(P3_U3291) );
  OAI222_X1 U12874 ( .A1(n14315), .A2(n13705), .B1(n16011), .B2(P3_U3151), 
        .C1(n14312), .C2(n10975), .ZN(P3_U3287) );
  AND2_X1 U12875 ( .A1(n10976), .A2(P1_U3086), .ZN(n13012) );
  INV_X2 U12876 ( .A(n13012), .ZN(n15556) );
  OAI222_X1 U12877 ( .A1(n15556), .A2(n10988), .B1(n15558), .B2(n8585), .C1(
        P1_U3086), .C2(n11288), .ZN(P1_U3354) );
  OAI222_X1 U12878 ( .A1(n14312), .A2(n10977), .B1(n14315), .B2(n13506), .C1(
        n16032), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U12879 ( .A(n10978), .ZN(n10990) );
  INV_X1 U12880 ( .A(n11386), .ZN(n10979) );
  OAI222_X1 U12881 ( .A1(n15558), .A2(n10980), .B1(n15556), .B2(n10990), .C1(
        n10979), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U12882 ( .A(n15163), .ZN(n10981) );
  OAI222_X1 U12883 ( .A1(n15558), .A2(n7529), .B1(n15556), .B2(n10986), .C1(
        n10981), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U12884 ( .A1(n14312), .A2(n10982), .B1(n14315), .B2(n13702), .C1(
        n12547), .C2(P3_U3151), .ZN(P3_U3285) );
  AND2_X1 U12885 ( .A1(n10984), .A2(P2_U3088), .ZN(n14803) );
  INV_X2 U12886 ( .A(n14803), .ZN(n14819) );
  NOR2_X1 U12887 ( .A1(n10984), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14798) );
  AOI22_X1 U12888 ( .A1(n15572), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n14798), .ZN(n10985) );
  OAI21_X1 U12889 ( .B1(n10986), .B2(n14819), .A(n10985), .ZN(P2_U3324) );
  INV_X2 U12890 ( .A(n14798), .ZN(n14821) );
  OAI222_X1 U12891 ( .A1(P2_U3088), .A2(n11191), .B1(n14819), .B2(n10988), 
        .C1(n10987), .C2(n14821), .ZN(P2_U3326) );
  OAI222_X1 U12892 ( .A1(P2_U3088), .A2(n11220), .B1(n14819), .B2(n10990), 
        .C1(n10989), .C2(n14821), .ZN(P2_U3325) );
  OAI222_X1 U12893 ( .A1(n14312), .A2(n10991), .B1(n12238), .B2(P3_U3151), 
        .C1(n14315), .C2(n13698), .ZN(P3_U3284) );
  INV_X1 U12894 ( .A(n10992), .ZN(n15551) );
  NAND2_X1 U12895 ( .A1(n15551), .A2(P1_B_REG_SCAN_IN), .ZN(n10993) );
  MUX2_X1 U12896 ( .A(n10993), .B(P1_B_REG_SCAN_IN), .S(n11056), .Z(n10995) );
  INV_X1 U12897 ( .A(n15550), .ZN(n10994) );
  NAND2_X1 U12898 ( .A1(n11555), .A2(n11557), .ZN(n15563) );
  INV_X1 U12899 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U12900 ( .A1(n15550), .A2(n15551), .ZN(n11556) );
  INV_X1 U12901 ( .A(n11556), .ZN(n10997) );
  AOI22_X1 U12902 ( .A1(n15563), .A2(n11052), .B1(n10997), .B2(n10996), .ZN(
        P1_U3446) );
  INV_X1 U12903 ( .A(n10998), .ZN(n10999) );
  INV_X1 U12904 ( .A(n15172), .ZN(n15170) );
  OAI222_X1 U12905 ( .A1(n15558), .A2(n7696), .B1(n15556), .B2(n10999), .C1(
        P1_U3086), .C2(n15170), .ZN(P1_U3351) );
  OAI222_X1 U12906 ( .A1(n14821), .A2(n11016), .B1(n14819), .B2(n10999), .C1(
        P2_U3088), .C2(n11205), .ZN(P2_U3323) );
  INV_X1 U12907 ( .A(n11293), .ZN(n11339) );
  INV_X1 U12908 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n11000) );
  OAI222_X1 U12909 ( .A1(P1_U3086), .A2(n11339), .B1(n15556), .B2(n11001), 
        .C1(n11000), .C2(n15558), .ZN(P1_U3350) );
  OAI222_X1 U12910 ( .A1(n14821), .A2(n11002), .B1(n14819), .B2(n11001), .C1(
        n11162), .C2(P2_U3088), .ZN(P2_U3322) );
  OAI222_X1 U12911 ( .A1(n14312), .A2(n11003), .B1(n12524), .B2(P3_U3151), 
        .C1(n14315), .C2(n13699), .ZN(P3_U3283) );
  OR2_X1 U12912 ( .A1(n11005), .A2(n11004), .ZN(n11006) );
  AND2_X1 U12913 ( .A1(n11006), .A2(n9059), .ZN(n11279) );
  INV_X1 U12914 ( .A(n11279), .ZN(n11007) );
  INV_X1 U12915 ( .A(n11555), .ZN(n11071) );
  NAND2_X1 U12916 ( .A1(n11071), .A2(n13013), .ZN(n11280) );
  AND2_X1 U12917 ( .A1(n11007), .A2(n11280), .ZN(n15696) );
  NOR2_X1 U12918 ( .A1(n15696), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U12919 ( .A1(n11565), .A2(P1_U4016), .ZN(n11008) );
  OAI21_X1 U12920 ( .B1(P1_U4016), .B2(n9629), .A(n11008), .ZN(P1_U3560) );
  INV_X1 U12921 ( .A(n11009), .ZN(n11011) );
  OAI222_X1 U12922 ( .A1(n14821), .A2(n11010), .B1(n14819), .B2(n11011), .C1(
        n11117), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U12923 ( .A(n11434), .ZN(n11443) );
  OAI222_X1 U12924 ( .A1(n15558), .A2(n11012), .B1(n15556), .B2(n11011), .C1(
        n11443), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12925 ( .A(n11322), .ZN(n11315) );
  OAI222_X1 U12926 ( .A1(n15558), .A2(n11013), .B1(n15556), .B2(n11014), .C1(
        n11315), .C2(P1_U3086), .ZN(P1_U3348) );
  OAI222_X1 U12927 ( .A1(n14821), .A2(n11015), .B1(n14819), .B2(n11014), .C1(
        n11236), .C2(P2_U3088), .ZN(P2_U3320) );
  MUX2_X1 U12928 ( .A(n11016), .B(n12048), .S(P1_U4016), .Z(n11017) );
  INV_X1 U12929 ( .A(n11017), .ZN(P1_U3564) );
  OAI222_X1 U12930 ( .A1(n11019), .A2(P3_U3151), .B1(n14312), .B2(n11018), 
        .C1(n13695), .C2(n14315), .ZN(P3_U3282) );
  MUX2_X1 U12931 ( .A(n11134), .B(n12365), .S(P1_U4016), .Z(n11020) );
  INV_X1 U12932 ( .A(n11020), .ZN(P1_U3569) );
  NAND2_X1 U12933 ( .A1(n12400), .A2(P2_U3947), .ZN(n11021) );
  OAI21_X1 U12934 ( .B1(n11401), .B2(P2_U3947), .A(n11021), .ZN(P2_U3544) );
  INV_X1 U12935 ( .A(n11022), .ZN(n11029) );
  INV_X1 U12936 ( .A(n15558), .ZN(n15545) );
  AOI22_X1 U12937 ( .A1(n15196), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n15545), .ZN(n11023) );
  OAI21_X1 U12938 ( .B1(n11029), .B2(n15556), .A(n11023), .ZN(P1_U3347) );
  INV_X1 U12939 ( .A(n14306), .ZN(n11410) );
  AND2_X1 U12940 ( .A1(n11025), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12941 ( .A1(n11025), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12942 ( .A1(n11025), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12943 ( .A1(n11025), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12944 ( .A1(n11025), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12945 ( .A1(n11025), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12946 ( .A1(n11025), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12947 ( .A1(n11025), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12948 ( .A1(n11025), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12949 ( .A1(n11025), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12950 ( .A1(n11025), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12951 ( .A1(n11025), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12952 ( .A1(n11025), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12953 ( .A1(n11025), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12954 ( .A1(n11025), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12955 ( .A1(n11025), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12956 ( .A1(n11025), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12957 ( .A1(n11025), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12958 ( .A1(n11025), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12959 ( .A1(n11025), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12960 ( .A1(n11025), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12961 ( .A1(n11025), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12962 ( .A1(n11025), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12963 ( .A1(n11025), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12964 ( .A1(n11025), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12965 ( .A1(n11025), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12966 ( .A1(n11025), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12967 ( .A1(n11025), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12968 ( .A1(n11025), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12969 ( .A1(n11025), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  NAND2_X1 U12970 ( .A1(n11026), .A2(P2_U3947), .ZN(n11027) );
  OAI21_X1 U12971 ( .B1(n9470), .B2(P2_U3947), .A(n11027), .ZN(P2_U3562) );
  INV_X1 U12972 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n11030) );
  INV_X1 U12973 ( .A(n15594), .ZN(n11028) );
  OAI222_X1 U12974 ( .A1(n14821), .A2(n11030), .B1(n14819), .B2(n11029), .C1(
        P2_U3088), .C2(n11028), .ZN(P2_U3319) );
  OAI222_X1 U12975 ( .A1(n14312), .A2(n11033), .B1(n14315), .B2(n11032), .C1(
        n11031), .C2(P3_U3151), .ZN(P3_U3281) );
  NAND2_X1 U12976 ( .A1(n11068), .A2(n12559), .ZN(n15269) );
  INV_X1 U12977 ( .A(n11579), .ZN(n11034) );
  INV_X2 U12978 ( .A(n11037), .ZN(n15005) );
  OAI22_X1 U12979 ( .A1(n16142), .A2(n15005), .B1(n15691), .B2(n11496), .ZN(
        n11035) );
  INV_X1 U12980 ( .A(n11035), .ZN(n11036) );
  INV_X1 U12981 ( .A(n11041), .ZN(n11040) );
  INV_X1 U12982 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n11039) );
  NAND2_X1 U12983 ( .A1(n11040), .A2(n11082), .ZN(n11042) );
  AND2_X1 U12984 ( .A1(n11042), .A2(n11084), .ZN(n11376) );
  NOR4_X1 U12985 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n11051) );
  NOR4_X1 U12986 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n11050) );
  NOR4_X1 U12987 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n11046) );
  NOR4_X1 U12988 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n11045) );
  NOR4_X1 U12989 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n11044) );
  NOR4_X1 U12990 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n11043) );
  NAND4_X1 U12991 ( .A1(n11046), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(
        n11047) );
  NOR4_X1 U12992 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n11048), .A4(n11047), .ZN(n11049) );
  NAND3_X1 U12993 ( .A1(n11051), .A2(n11050), .A3(n11049), .ZN(n11558) );
  NOR2_X1 U12994 ( .A1(n11558), .A2(n11052), .ZN(n11053) );
  OAI21_X1 U12995 ( .B1(n11557), .B2(n11053), .A(n11556), .ZN(n11054) );
  INV_X1 U12996 ( .A(n11054), .ZN(n11791) );
  INV_X1 U12997 ( .A(n11557), .ZN(n11559) );
  INV_X1 U12998 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U12999 ( .A1(n11559), .A2(n11055), .ZN(n11057) );
  INV_X1 U13000 ( .A(n11056), .ZN(n15554) );
  NAND2_X1 U13001 ( .A1(n15550), .A2(n15554), .ZN(n15541) );
  NAND2_X1 U13002 ( .A1(n11791), .A2(n11599), .ZN(n11069) );
  INV_X1 U13003 ( .A(n11069), .ZN(n11058) );
  NAND2_X1 U13004 ( .A1(n11058), .A2(n11555), .ZN(n11065) );
  INV_X1 U13005 ( .A(n16086), .ZN(n11059) );
  OR2_X1 U13006 ( .A1(n11059), .A2(n12559), .ZN(n11060) );
  OR2_X1 U13007 ( .A1(n16528), .A2(n11063), .ZN(n11061) );
  INV_X1 U13008 ( .A(n11554), .ZN(n11062) );
  NOR2_X1 U13009 ( .A1(n11064), .A2(n15401), .ZN(n16092) );
  AOI22_X1 U13010 ( .A1(n11376), .A2(n16546), .B1(n16548), .B2(n16092), .ZN(
        n11073) );
  OR2_X1 U13011 ( .A1(n11065), .A2(n11798), .ZN(n11067) );
  AND2_X1 U13012 ( .A1(n11555), .A2(n7363), .ZN(n11066) );
  NAND2_X1 U13013 ( .A1(n15501), .A2(n7363), .ZN(n11562) );
  NAND2_X1 U13014 ( .A1(n11069), .A2(n11562), .ZN(n11070) );
  NAND2_X1 U13015 ( .A1(n11070), .A2(n11554), .ZN(n11498) );
  OR2_X1 U13016 ( .A1(n11498), .A2(n11071), .ZN(n11177) );
  AOI22_X1 U13017 ( .A1(n9047), .A2(n16551), .B1(n11177), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n11072) );
  NAND2_X1 U13018 ( .A1(n11073), .A2(n11072), .ZN(P1_U3232) );
  INV_X1 U13019 ( .A(n11074), .ZN(n11077) );
  OAI22_X1 U13020 ( .A1(n11075), .A2(P3_U3151), .B1(SI_15_), .B2(n14315), .ZN(
        n11076) );
  AOI21_X1 U13021 ( .B1(n11077), .B2(n12146), .A(n11076), .ZN(P3_U3280) );
  INV_X1 U13022 ( .A(n16551), .ZN(n15108) );
  NAND2_X1 U13023 ( .A1(n15143), .A2(n11037), .ZN(n11079) );
  NAND2_X1 U13024 ( .A1(n11079), .A2(n11078), .ZN(n11080) );
  NAND2_X2 U13025 ( .A1(n11580), .A2(n11579), .ZN(n15001) );
  XNOR2_X1 U13026 ( .A(n11080), .B(n15001), .ZN(n11163) );
  NOR2_X1 U13027 ( .A1(n16155), .A2(n15005), .ZN(n11081) );
  AOI21_X1 U13028 ( .B1(n14955), .B2(n15143), .A(n11081), .ZN(n11164) );
  XNOR2_X1 U13029 ( .A(n11163), .B(n11164), .ZN(n11086) );
  NAND2_X1 U13030 ( .A1(n11082), .A2(n14925), .ZN(n11083) );
  AND2_X1 U13031 ( .A1(n11084), .A2(n11083), .ZN(n11085) );
  NAND2_X1 U13032 ( .A1(n11086), .A2(n11085), .ZN(n11167) );
  OAI21_X1 U13033 ( .B1(n11086), .B2(n11085), .A(n11167), .ZN(n11087) );
  NAND2_X1 U13034 ( .A1(n11087), .A2(n16546), .ZN(n11090) );
  INV_X1 U13035 ( .A(n11565), .ZN(n11088) );
  INV_X1 U13036 ( .A(n15100), .ZN(n15399) );
  OAI22_X1 U13037 ( .A1(n11088), .A2(n15399), .B1(n11582), .B2(n15401), .ZN(
        n16147) );
  AOI22_X1 U13038 ( .A1(n16548), .A2(n16147), .B1(n11177), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n11089) );
  OAI211_X1 U13039 ( .C1(n16155), .C2(n15108), .A(n11090), .B(n11089), .ZN(
        P1_U3222) );
  INV_X1 U13040 ( .A(n11091), .ZN(n11140) );
  AOI22_X1 U13041 ( .A1(n15212), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n15545), .ZN(n11092) );
  OAI21_X1 U13042 ( .B1(n11140), .B2(n15556), .A(n11092), .ZN(P1_U3345) );
  INV_X1 U13043 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n16327) );
  INV_X1 U13044 ( .A(n11205), .ZN(n11096) );
  INV_X1 U13045 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n11094) );
  INV_X1 U13046 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n16171) );
  MUX2_X1 U13047 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n16171), .S(n11191), .Z(
        n11180) );
  NAND2_X1 U13048 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n11093) );
  NOR2_X1 U13049 ( .A1(n11180), .A2(n11093), .ZN(n11211) );
  NOR2_X1 U13050 ( .A1(n11191), .A2(n16171), .ZN(n11210) );
  MUX2_X1 U13051 ( .A(n11094), .B(P2_REG1_REG_2__SCAN_IN), .S(n11220), .Z(
        n11209) );
  OAI21_X1 U13052 ( .B1(n11211), .B2(n11210), .A(n11209), .ZN(n11208) );
  OAI21_X1 U13053 ( .B1(n11094), .B2(n11220), .A(n11208), .ZN(n15578) );
  INV_X1 U13054 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11095) );
  MUX2_X1 U13055 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n11095), .S(n15572), .Z(
        n15577) );
  NAND2_X1 U13056 ( .A1(n15578), .A2(n15577), .ZN(n15576) );
  NAND2_X1 U13057 ( .A1(n15572), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n11198) );
  INV_X1 U13058 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n16302) );
  MUX2_X1 U13059 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n16302), .S(n11205), .Z(
        n11197) );
  AOI21_X1 U13060 ( .B1(n15576), .B2(n11198), .A(n11197), .ZN(n11196) );
  AOI21_X1 U13061 ( .B1(n11096), .B2(P2_REG1_REG_4__SCAN_IN), .A(n11196), .ZN(
        n11150) );
  MUX2_X1 U13062 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n16327), .S(n11162), .Z(
        n11149) );
  OR2_X1 U13063 ( .A1(n11150), .A2(n11149), .ZN(n11151) );
  OAI21_X1 U13064 ( .B1(n16327), .B2(n11162), .A(n11151), .ZN(n15589) );
  INV_X1 U13065 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11097) );
  MUX2_X1 U13066 ( .A(n11097), .B(P2_REG1_REG_6__SCAN_IN), .S(n11117), .Z(
        n15588) );
  NAND2_X1 U13067 ( .A1(n15589), .A2(n15588), .ZN(n15587) );
  INV_X1 U13068 ( .A(n11117), .ZN(n15583) );
  NAND2_X1 U13069 ( .A1(n15583), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11099) );
  INV_X1 U13070 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n16364) );
  MUX2_X1 U13071 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n16364), .S(n11236), .Z(
        n11098) );
  AOI21_X1 U13072 ( .B1(n15587), .B2(n11099), .A(n11098), .ZN(n11230) );
  NAND3_X1 U13073 ( .A1(n15587), .A2(n11099), .A3(n11098), .ZN(n11101) );
  NAND2_X1 U13074 ( .A1(n11102), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14805) );
  INV_X1 U13075 ( .A(n14805), .ZN(n11122) );
  NAND2_X1 U13076 ( .A1(n11122), .A2(n14808), .ZN(n11100) );
  OR2_X1 U13077 ( .A1(n11124), .A2(n11100), .ZN(n15681) );
  NAND2_X1 U13078 ( .A1(n11101), .A2(n15668), .ZN(n11130) );
  INV_X1 U13079 ( .A(n11236), .ZN(n11231) );
  INV_X1 U13080 ( .A(n15684), .ZN(n11934) );
  INV_X1 U13081 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U13082 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11633) );
  OAI21_X1 U13083 ( .B1(n11934), .B2(n11103), .A(n11633), .ZN(n11104) );
  AOI21_X1 U13084 ( .B1(n11231), .B2(n15678), .A(n11104), .ZN(n11129) );
  INV_X1 U13085 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11105) );
  MUX2_X1 U13086 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11105), .S(n15572), .Z(
        n15574) );
  INV_X1 U13087 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11744) );
  MUX2_X1 U13088 ( .A(n11744), .B(P2_REG2_REG_1__SCAN_IN), .S(n11191), .Z(
        n11107) );
  AND2_X1 U13089 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n11106) );
  NAND2_X1 U13090 ( .A1(n11107), .A2(n11106), .ZN(n11187) );
  OAI21_X1 U13091 ( .B1(n11744), .B2(n11191), .A(n11187), .ZN(n11215) );
  XNOR2_X1 U13092 ( .A(n11220), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n11216) );
  NAND2_X1 U13093 ( .A1(n11215), .A2(n11216), .ZN(n11110) );
  INV_X1 U13094 ( .A(n11220), .ZN(n11108) );
  NAND2_X1 U13095 ( .A1(n11108), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U13096 ( .A1(n11110), .A2(n11109), .ZN(n15575) );
  NAND2_X1 U13097 ( .A1(n15574), .A2(n15575), .ZN(n15573) );
  NAND2_X1 U13098 ( .A1(n15572), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U13099 ( .A1(n15573), .A2(n11193), .ZN(n11112) );
  INV_X1 U13100 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11860) );
  MUX2_X1 U13101 ( .A(n11860), .B(P2_REG2_REG_4__SCAN_IN), .S(n11205), .Z(
        n11111) );
  NAND2_X1 U13102 ( .A1(n11112), .A2(n11111), .ZN(n11195) );
  OR2_X1 U13103 ( .A1(n11205), .A2(n11860), .ZN(n11157) );
  NAND2_X1 U13104 ( .A1(n11195), .A2(n11157), .ZN(n11114) );
  INV_X1 U13105 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11155) );
  MUX2_X1 U13106 ( .A(n11155), .B(P2_REG2_REG_5__SCAN_IN), .S(n11162), .Z(
        n11113) );
  NAND2_X1 U13107 ( .A1(n11114), .A2(n11113), .ZN(n11159) );
  INV_X1 U13108 ( .A(n11162), .ZN(n11115) );
  NAND2_X1 U13109 ( .A1(n11115), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n11116) );
  NAND2_X1 U13110 ( .A1(n11159), .A2(n11116), .ZN(n15586) );
  INV_X1 U13111 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11903) );
  MUX2_X1 U13112 ( .A(n11903), .B(P2_REG2_REG_6__SCAN_IN), .S(n11117), .Z(
        n15585) );
  NAND2_X1 U13113 ( .A1(n15586), .A2(n15585), .ZN(n15584) );
  OR2_X1 U13114 ( .A1(n11117), .A2(n11903), .ZN(n11126) );
  NAND2_X1 U13115 ( .A1(n15584), .A2(n11126), .ZN(n11120) );
  INV_X1 U13116 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11118) );
  MUX2_X1 U13117 ( .A(n11118), .B(P2_REG2_REG_7__SCAN_IN), .S(n11236), .Z(
        n11119) );
  NAND2_X1 U13118 ( .A1(n11120), .A2(n11119), .ZN(n11238) );
  NAND2_X1 U13119 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  INV_X1 U13120 ( .A(n15686), .ZN(n15661) );
  MUX2_X1 U13121 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11118), .S(n11236), .Z(
        n11125) );
  NAND3_X1 U13122 ( .A1(n15584), .A2(n11126), .A3(n11125), .ZN(n11127) );
  NAND3_X1 U13123 ( .A1(n11238), .A2(n15661), .A3(n11127), .ZN(n11128) );
  OAI211_X1 U13124 ( .C1(n11230), .C2(n11130), .A(n11129), .B(n11128), .ZN(
        P2_U3221) );
  INV_X1 U13125 ( .A(n11356), .ZN(n11350) );
  INV_X1 U13126 ( .A(n11131), .ZN(n11133) );
  OAI222_X1 U13127 ( .A1(P1_U3086), .A2(n11350), .B1(n15558), .B2(n11132), 
        .C1(n15556), .C2(n11133), .ZN(P1_U3346) );
  INV_X1 U13128 ( .A(n11258), .ZN(n11264) );
  OAI222_X1 U13129 ( .A1(P2_U3088), .A2(n11264), .B1(n14821), .B2(n11134), 
        .C1(n14819), .C2(n11133), .ZN(P2_U3318) );
  INV_X1 U13130 ( .A(n11135), .ZN(n11138) );
  INV_X1 U13131 ( .A(SI_16_), .ZN(n11137) );
  OAI222_X1 U13132 ( .A1(n14312), .A2(n11138), .B1(n14315), .B2(n11137), .C1(
        n11136), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U13133 ( .A(n11538), .ZN(n11249) );
  INV_X1 U13134 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n11139) );
  OAI222_X1 U13135 ( .A1(P2_U3088), .A2(n11249), .B1(n14819), .B2(n11140), 
        .C1(n11139), .C2(n14821), .ZN(P2_U3317) );
  INV_X1 U13136 ( .A(n11752), .ZN(n16168) );
  NAND2_X1 U13137 ( .A1(n14472), .A2(n14628), .ZN(n11142) );
  NAND2_X1 U13138 ( .A1(n14475), .A2(n14627), .ZN(n11141) );
  NAND2_X1 U13139 ( .A1(n11142), .A2(n11141), .ZN(n11741) );
  OR2_X1 U13140 ( .A1(n11143), .A2(P2_U3088), .ZN(n11760) );
  AOI22_X1 U13141 ( .A1(n14445), .A2(n11741), .B1(n11760), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n11148) );
  OAI21_X1 U13142 ( .B1(n11145), .B2(n11144), .A(n11764), .ZN(n11146) );
  NAND2_X1 U13143 ( .A1(n14437), .A2(n11146), .ZN(n11147) );
  OAI211_X1 U13144 ( .C1(n14448), .C2(n16168), .A(n11148), .B(n11147), .ZN(
        P2_U3194) );
  NAND2_X1 U13145 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n11418) );
  AOI21_X1 U13146 ( .B1(n11150), .B2(n11149), .A(n15681), .ZN(n11152) );
  NAND2_X1 U13147 ( .A1(n11152), .A2(n11151), .ZN(n11153) );
  NAND2_X1 U13148 ( .A1(n11418), .A2(n11153), .ZN(n11154) );
  AOI21_X1 U13149 ( .B1(n15684), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n11154), .ZN(
        n11161) );
  MUX2_X1 U13150 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11155), .S(n11162), .Z(
        n11156) );
  NAND3_X1 U13151 ( .A1(n11195), .A2(n11157), .A3(n11156), .ZN(n11158) );
  NAND3_X1 U13152 ( .A1(n15661), .A2(n11159), .A3(n11158), .ZN(n11160) );
  OAI211_X1 U13153 ( .C1(n15626), .C2(n11162), .A(n11161), .B(n11160), .ZN(
        P2_U3219) );
  INV_X1 U13154 ( .A(n11163), .ZN(n11165) );
  NAND2_X1 U13155 ( .A1(n11165), .A2(n11164), .ZN(n11166) );
  NAND2_X1 U13156 ( .A1(n11171), .A2(n14900), .ZN(n11169) );
  INV_X2 U13157 ( .A(n15000), .ZN(n14950) );
  NAND2_X1 U13158 ( .A1(n11802), .A2(n14950), .ZN(n11168) );
  NAND2_X1 U13159 ( .A1(n11169), .A2(n11168), .ZN(n11170) );
  XNOR2_X1 U13160 ( .A(n11170), .B(n14925), .ZN(n11474) );
  NAND2_X1 U13161 ( .A1(n14955), .A2(n11171), .ZN(n11173) );
  INV_X2 U13162 ( .A(n15005), .ZN(n14900) );
  NAND2_X1 U13163 ( .A1(n11802), .A2(n14900), .ZN(n11172) );
  NAND2_X1 U13164 ( .A1(n11173), .A2(n11172), .ZN(n11472) );
  XNOR2_X1 U13165 ( .A(n11471), .B(n11470), .ZN(n11174) );
  NAND2_X1 U13166 ( .A1(n11174), .A2(n16546), .ZN(n11179) );
  NAND2_X1 U13167 ( .A1(n15141), .A2(n15099), .ZN(n11176) );
  NAND2_X1 U13168 ( .A1(n15143), .A2(n15100), .ZN(n11175) );
  NAND2_X1 U13169 ( .A1(n11176), .A2(n11175), .ZN(n11795) );
  AOI22_X1 U13170 ( .A1(n16548), .A2(n11795), .B1(n11177), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n11178) );
  OAI211_X1 U13171 ( .C1(n16204), .C2(n15108), .A(n11179), .B(n11178), .ZN(
        P1_U3237) );
  INV_X1 U13172 ( .A(n11211), .ZN(n11182) );
  INV_X1 U13173 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n16113) );
  OAI21_X1 U13174 ( .B1(n16113), .B2(n11185), .A(n11180), .ZN(n11181) );
  NAND2_X1 U13175 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  INV_X1 U13176 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11749) );
  OAI22_X1 U13177 ( .A1(n15681), .A2(n11183), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11749), .ZN(n11189) );
  INV_X1 U13178 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n16124) );
  MUX2_X1 U13179 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11744), .S(n11191), .Z(
        n11184) );
  OAI21_X1 U13180 ( .B1(n16124), .B2(n11185), .A(n11184), .ZN(n11186) );
  AND3_X1 U13181 ( .A1(n15661), .A2(n11187), .A3(n11186), .ZN(n11188) );
  AOI211_X1 U13182 ( .C1(n15684), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n11189), .B(
        n11188), .ZN(n11190) );
  OAI21_X1 U13183 ( .B1(n11191), .B2(n15626), .A(n11190), .ZN(P2_U3215) );
  MUX2_X1 U13184 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11860), .S(n11205), .Z(
        n11192) );
  NAND3_X1 U13185 ( .A1(n15573), .A2(n11193), .A3(n11192), .ZN(n11194) );
  NAND3_X1 U13186 ( .A1(n15661), .A2(n11195), .A3(n11194), .ZN(n11203) );
  INV_X1 U13187 ( .A(n11196), .ZN(n11200) );
  NAND3_X1 U13188 ( .A1(n15576), .A2(n11198), .A3(n11197), .ZN(n11199) );
  NAND3_X1 U13189 ( .A1(n15668), .A2(n11200), .A3(n11199), .ZN(n11202) );
  NAND2_X1 U13190 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n11693) );
  NAND2_X1 U13191 ( .A1(n15684), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n11201) );
  AND4_X1 U13192 ( .A1(n11203), .A2(n11202), .A3(n11693), .A4(n11201), .ZN(
        n11204) );
  OAI21_X1 U13193 ( .B1(n11205), .B2(n15626), .A(n11204), .ZN(P2_U3218) );
  INV_X1 U13194 ( .A(n11206), .ZN(n11226) );
  AOI22_X1 U13195 ( .A1(n11614), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n15545), .ZN(n11207) );
  OAI21_X1 U13196 ( .B1(n11226), .B2(n15556), .A(n11207), .ZN(P1_U3344) );
  INV_X1 U13197 ( .A(n11208), .ZN(n11213) );
  NOR3_X1 U13198 ( .A1(n11211), .A2(n11210), .A3(n11209), .ZN(n11212) );
  NOR3_X1 U13199 ( .A1(n15681), .A2(n11213), .A3(n11212), .ZN(n11214) );
  AOI21_X1 U13200 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .A(n11214), 
        .ZN(n11219) );
  XOR2_X1 U13201 ( .A(n11216), .B(n11215), .Z(n11217) );
  AOI22_X1 U13202 ( .A1(n15661), .A2(n11217), .B1(n15684), .B2(
        P2_ADDR_REG_2__SCAN_IN), .ZN(n11218) );
  OAI211_X1 U13203 ( .C1(n11220), .C2(n15626), .A(n11219), .B(n11218), .ZN(
        P2_U3216) );
  AOI22_X1 U13204 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15661), .B1(n15668), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n11223) );
  OAI22_X1 U13205 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15686), .B1(n15681), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n11221) );
  NOR2_X1 U13206 ( .A1(n11221), .A2(n15678), .ZN(n11222) );
  MUX2_X1 U13207 ( .A(n11223), .B(n11222), .S(P2_IR_REG_0__SCAN_IN), .Z(n11225) );
  AOI22_X1 U13208 ( .A1(n15684), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n11224) );
  NAND2_X1 U13209 ( .A1(n11225), .A2(n11224), .ZN(P2_U3214) );
  INV_X1 U13210 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n11227) );
  INV_X1 U13211 ( .A(n11541), .ZN(n15611) );
  OAI222_X1 U13212 ( .A1(n14821), .A2(n11227), .B1(n14819), .B2(n11226), .C1(
        P2_U3088), .C2(n15611), .ZN(P2_U3316) );
  INV_X1 U13213 ( .A(n11228), .ZN(n11229) );
  INV_X1 U13214 ( .A(SI_17_), .ZN(n13690) );
  OAI222_X1 U13215 ( .A1(n14312), .A2(n11229), .B1(n16075), .B2(P3_U3151), 
        .C1(n13690), .C2(n14315), .ZN(P3_U3278) );
  AOI21_X1 U13216 ( .B1(n11231), .B2(P2_REG1_REG_7__SCAN_IN), .A(n11230), .ZN(
        n15597) );
  INV_X1 U13217 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11232) );
  MUX2_X1 U13218 ( .A(n11232), .B(P2_REG1_REG_8__SCAN_IN), .S(n15594), .Z(
        n15596) );
  NOR2_X1 U13219 ( .A1(n15597), .A2(n15596), .ZN(n15595) );
  AOI21_X1 U13220 ( .B1(n15594), .B2(P2_REG1_REG_8__SCAN_IN), .A(n15595), .ZN(
        n11255) );
  INV_X1 U13221 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11233) );
  MUX2_X1 U13222 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11233), .S(n11258), .Z(
        n11254) );
  NAND2_X1 U13223 ( .A1(n11255), .A2(n11254), .ZN(n11253) );
  OAI21_X1 U13224 ( .B1(n11258), .B2(P2_REG1_REG_9__SCAN_IN), .A(n11253), .ZN(
        n11235) );
  INV_X1 U13225 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n16437) );
  MUX2_X1 U13226 ( .A(n16437), .B(P2_REG1_REG_10__SCAN_IN), .S(n11538), .Z(
        n11234) );
  NOR2_X1 U13227 ( .A1(n11235), .A2(n11234), .ZN(n11534) );
  AOI211_X1 U13228 ( .C1(n11235), .C2(n11234), .A(n15681), .B(n11534), .ZN(
        n11252) );
  OR2_X1 U13229 ( .A1(n11236), .A2(n11118), .ZN(n11237) );
  NAND2_X1 U13230 ( .A1(n11238), .A2(n11237), .ZN(n15601) );
  INV_X1 U13231 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11239) );
  MUX2_X1 U13232 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11239), .S(n15594), .Z(
        n15600) );
  NAND2_X1 U13233 ( .A1(n15601), .A2(n15600), .ZN(n15599) );
  NAND2_X1 U13234 ( .A1(n15594), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U13235 ( .A1(n15599), .A2(n11240), .ZN(n11257) );
  INV_X1 U13236 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11241) );
  MUX2_X1 U13237 ( .A(n11241), .B(P2_REG2_REG_9__SCAN_IN), .S(n11258), .Z(
        n11242) );
  OR2_X1 U13238 ( .A1(n11257), .A2(n11242), .ZN(n11259) );
  OR2_X1 U13239 ( .A1(n11258), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U13240 ( .A1(n11259), .A2(n11243), .ZN(n11247) );
  INV_X1 U13241 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11244) );
  MUX2_X1 U13242 ( .A(n11244), .B(P2_REG2_REG_10__SCAN_IN), .S(n11538), .Z(
        n11246) );
  INV_X1 U13243 ( .A(n11540), .ZN(n11245) );
  AOI211_X1 U13244 ( .C1(n11247), .C2(n11246), .A(n15686), .B(n11245), .ZN(
        n11251) );
  NAND2_X1 U13245 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n12027)
         );
  NAND2_X1 U13246 ( .A1(n15684), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n11248) );
  OAI211_X1 U13247 ( .C1(n15626), .C2(n11249), .A(n12027), .B(n11248), .ZN(
        n11250) );
  OR3_X1 U13248 ( .A1(n11252), .A2(n11251), .A3(n11250), .ZN(P2_U3224) );
  OAI21_X1 U13249 ( .B1(n11255), .B2(n11254), .A(n11253), .ZN(n11256) );
  NAND2_X1 U13250 ( .A1(n11256), .A2(n15668), .ZN(n11268) );
  INV_X1 U13251 ( .A(n11257), .ZN(n11261) );
  MUX2_X1 U13252 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11241), .S(n11258), .Z(
        n11260) );
  OAI21_X1 U13253 ( .B1(n11261), .B2(n11260), .A(n11259), .ZN(n11266) );
  NAND2_X1 U13254 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11263) );
  NAND2_X1 U13255 ( .A1(n15684), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11262) );
  OAI211_X1 U13256 ( .C1(n15626), .C2(n11264), .A(n11263), .B(n11262), .ZN(
        n11265) );
  AOI21_X1 U13257 ( .B1(n11266), .B2(n15661), .A(n11265), .ZN(n11267) );
  NAND2_X1 U13258 ( .A1(n11268), .A2(n11267), .ZN(P2_U3223) );
  INV_X1 U13259 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11269) );
  MUX2_X1 U13260 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n11269), .S(n11386), .Z(
        n11270) );
  MUX2_X1 U13261 ( .A(n9048), .B(P1_REG2_REG_1__SCAN_IN), .S(n11288), .Z(
        n15145) );
  AND2_X1 U13262 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15146) );
  NAND2_X1 U13263 ( .A1(n15145), .A2(n15146), .ZN(n15144) );
  OAI21_X1 U13264 ( .B1(n9048), .B2(n11288), .A(n15144), .ZN(n11379) );
  NAND2_X1 U13265 ( .A1(n11270), .A2(n11379), .ZN(n15157) );
  NAND2_X1 U13266 ( .A1(n11386), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n15156) );
  NAND2_X1 U13267 ( .A1(n15157), .A2(n15156), .ZN(n11272) );
  INV_X1 U13268 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n12051) );
  MUX2_X1 U13269 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n12051), .S(n15163), .Z(
        n11271) );
  NAND2_X1 U13270 ( .A1(n11272), .A2(n11271), .ZN(n15175) );
  NAND2_X1 U13271 ( .A1(n15163), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U13272 ( .A1(n15175), .A2(n15174), .ZN(n11275) );
  INV_X1 U13273 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11273) );
  MUX2_X1 U13274 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11273), .S(n15172), .Z(
        n11274) );
  NAND2_X1 U13275 ( .A1(n11275), .A2(n11274), .ZN(n15177) );
  NAND2_X1 U13276 ( .A1(n15172), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n11343) );
  INV_X1 U13277 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11276) );
  MUX2_X1 U13278 ( .A(n11276), .B(P1_REG2_REG_5__SCAN_IN), .S(n11293), .Z(
        n11342) );
  AOI21_X1 U13279 ( .B1(n15177), .B2(n11343), .A(n11342), .ZN(n11439) );
  NOR2_X1 U13280 ( .A1(n11339), .A2(n11276), .ZN(n11433) );
  INV_X1 U13281 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11277) );
  MUX2_X1 U13282 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11277), .S(n11434), .Z(
        n11278) );
  OAI21_X1 U13283 ( .B1(n11439), .B2(n11433), .A(n11278), .ZN(n11437) );
  NAND2_X1 U13284 ( .A1(n11434), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11283) );
  INV_X1 U13285 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11314) );
  MUX2_X1 U13286 ( .A(n11314), .B(P1_REG2_REG_7__SCAN_IN), .S(n11322), .Z(
        n11282) );
  AOI21_X1 U13287 ( .B1(n11437), .B2(n11283), .A(n11282), .ZN(n15195) );
  NAND2_X1 U13288 ( .A1(n11280), .A2(n11279), .ZN(n15699) );
  NOR2_X1 U13289 ( .A1(n15699), .A2(n15689), .ZN(n15231) );
  INV_X1 U13290 ( .A(n15231), .ZN(n11281) );
  NAND3_X1 U13291 ( .A1(n11437), .A2(n11283), .A3(n11282), .ZN(n11284) );
  NAND2_X1 U13292 ( .A1(n7362), .A2(n11284), .ZN(n11301) );
  OR2_X1 U13293 ( .A1(n15699), .A2(n11285), .ZN(n15704) );
  INV_X1 U13294 ( .A(n15704), .ZN(n15722) );
  INV_X1 U13295 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n11286) );
  NAND2_X1 U13296 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11879) );
  OAI21_X1 U13297 ( .B1(n15728), .B2(n11286), .A(n11879), .ZN(n11287) );
  AOI21_X1 U13298 ( .B1(n11322), .B2(n15722), .A(n11287), .ZN(n11300) );
  INV_X1 U13299 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n16356) );
  MUX2_X1 U13300 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n16356), .S(n11322), .Z(
        n11298) );
  INV_X1 U13301 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n16209) );
  MUX2_X1 U13302 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n16209), .S(n11386), .Z(
        n11385) );
  INV_X1 U13303 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n16150) );
  MUX2_X1 U13304 ( .A(n16150), .B(P1_REG1_REG_1__SCAN_IN), .S(n11288), .Z(
        n15149) );
  AND2_X1 U13305 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n15148) );
  NAND2_X1 U13306 ( .A1(n15149), .A2(n15148), .ZN(n15147) );
  INV_X1 U13307 ( .A(n11288), .ZN(n15150) );
  NAND2_X1 U13308 ( .A1(n15150), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U13309 ( .A1(n15147), .A2(n11289), .ZN(n11384) );
  NAND2_X1 U13310 ( .A1(n11385), .A2(n11384), .ZN(n11383) );
  NAND2_X1 U13311 ( .A1(n11386), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n11290) );
  NAND2_X1 U13312 ( .A1(n11383), .A2(n11290), .ZN(n15161) );
  INV_X1 U13313 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n16249) );
  MUX2_X1 U13314 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n16249), .S(n15163), .Z(
        n15162) );
  NAND2_X1 U13315 ( .A1(n15161), .A2(n15162), .ZN(n15160) );
  NAND2_X1 U13316 ( .A1(n15163), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U13317 ( .A1(n15160), .A2(n11291), .ZN(n15179) );
  INV_X1 U13318 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n16292) );
  MUX2_X1 U13319 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n16292), .S(n15172), .Z(
        n15180) );
  NAND2_X1 U13320 ( .A1(n15179), .A2(n15180), .ZN(n15178) );
  NAND2_X1 U13321 ( .A1(n15172), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n11292) );
  NAND2_X1 U13322 ( .A1(n15178), .A2(n11292), .ZN(n11337) );
  XNOR2_X1 U13323 ( .A(n11293), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n11338) );
  OR2_X1 U13324 ( .A1(n11337), .A2(n11338), .ZN(n11335) );
  OR2_X1 U13325 ( .A1(n11293), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n11294) );
  NAND2_X1 U13326 ( .A1(n11335), .A2(n11294), .ZN(n11446) );
  XNOR2_X1 U13327 ( .A(n11434), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n11447) );
  NAND2_X1 U13328 ( .A1(n11434), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11295) );
  NAND2_X1 U13329 ( .A1(n11444), .A2(n11295), .ZN(n11297) );
  NAND2_X1 U13330 ( .A1(n11297), .A2(n11298), .ZN(n11324) );
  OAI211_X1 U13331 ( .C1(n11298), .C2(n11297), .A(n15720), .B(n11324), .ZN(
        n11299) );
  OAI211_X1 U13332 ( .C1(n15195), .C2(n11301), .A(n11300), .B(n11299), .ZN(
        P1_U3250) );
  INV_X1 U13333 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U13334 ( .A1(n13397), .A2(P3_U3897), .ZN(n11302) );
  OAI21_X1 U13335 ( .B1(P3_U3897), .B2(n11303), .A(n11302), .ZN(P3_U3508) );
  INV_X1 U13336 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n13812) );
  NAND2_X1 U13337 ( .A1(n13026), .A2(P3_U3897), .ZN(n11304) );
  OAI21_X1 U13338 ( .B1(P3_U3897), .B2(n13812), .A(n11304), .ZN(P3_U3504) );
  INV_X1 U13339 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U13340 ( .A1(n13027), .A2(P3_U3897), .ZN(n11305) );
  OAI21_X1 U13341 ( .B1(P3_U3897), .B2(n11306), .A(n11305), .ZN(P3_U3506) );
  INV_X1 U13342 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n13805) );
  NAND2_X1 U13343 ( .A1(n14131), .A2(P3_U3897), .ZN(n11307) );
  OAI21_X1 U13344 ( .B1(P3_U3897), .B2(n13805), .A(n11307), .ZN(P3_U3507) );
  INV_X1 U13345 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n13830) );
  NAND2_X1 U13346 ( .A1(n11308), .A2(P3_U3897), .ZN(n11309) );
  OAI21_X1 U13347 ( .B1(P3_U3897), .B2(n13830), .A(n11309), .ZN(P3_U3492) );
  INV_X1 U13348 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n13831) );
  NAND2_X1 U13349 ( .A1(n11310), .A2(P3_U3897), .ZN(n11311) );
  OAI21_X1 U13350 ( .B1(P3_U3897), .B2(n13831), .A(n11311), .ZN(P3_U3493) );
  INV_X1 U13351 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U13352 ( .A1(n13018), .A2(P3_U3897), .ZN(n11312) );
  OAI21_X1 U13353 ( .B1(P3_U3897), .B2(n11313), .A(n11312), .ZN(P3_U3503) );
  NOR2_X1 U13354 ( .A1(n11315), .A2(n11314), .ZN(n15190) );
  INV_X1 U13355 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11316) );
  MUX2_X1 U13356 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11316), .S(n15196), .Z(
        n11317) );
  OAI21_X1 U13357 ( .B1(n15195), .B2(n15190), .A(n11317), .ZN(n15193) );
  NAND2_X1 U13358 ( .A1(n15196), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11319) );
  INV_X1 U13359 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11349) );
  MUX2_X1 U13360 ( .A(n11349), .B(P1_REG2_REG_9__SCAN_IN), .S(n11356), .Z(
        n11318) );
  AOI21_X1 U13361 ( .B1(n15193), .B2(n11319), .A(n11318), .ZN(n15206) );
  NAND3_X1 U13362 ( .A1(n15193), .A2(n11319), .A3(n11318), .ZN(n11320) );
  NAND2_X1 U13363 ( .A1(n11320), .A2(n7362), .ZN(n11334) );
  INV_X1 U13364 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11321) );
  MUX2_X1 U13365 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n11321), .S(n11356), .Z(
        n11328) );
  NAND2_X1 U13366 ( .A1(n11322), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11323) );
  AND2_X1 U13367 ( .A1(n11324), .A2(n11323), .ZN(n15187) );
  INV_X1 U13368 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11325) );
  MUX2_X1 U13369 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n11325), .S(n15196), .Z(
        n15186) );
  OR2_X1 U13370 ( .A1(n15196), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11326) );
  NAND2_X1 U13371 ( .A1(n15185), .A2(n11326), .ZN(n11327) );
  NAND2_X1 U13372 ( .A1(n11327), .A2(n11328), .ZN(n11358) );
  OAI21_X1 U13373 ( .B1(n11328), .B2(n11327), .A(n11358), .ZN(n11329) );
  NAND2_X1 U13374 ( .A1(n11329), .A2(n15720), .ZN(n11333) );
  INV_X1 U13375 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U13376 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n12370) );
  OAI21_X1 U13377 ( .B1(n15728), .B2(n11330), .A(n12370), .ZN(n11331) );
  AOI21_X1 U13378 ( .B1(n11356), .B2(n15722), .A(n11331), .ZN(n11332) );
  OAI211_X1 U13379 ( .C1(n15206), .C2(n11334), .A(n11333), .B(n11332), .ZN(
        P1_U3252) );
  INV_X1 U13380 ( .A(n11335), .ZN(n11336) );
  AOI21_X1 U13381 ( .B1(n11338), .B2(n11337), .A(n11336), .ZN(n11348) );
  NAND2_X1 U13382 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11529) );
  INV_X1 U13383 ( .A(n11529), .ZN(n11341) );
  NOR2_X1 U13384 ( .A1(n15704), .A2(n11339), .ZN(n11340) );
  AOI211_X1 U13385 ( .C1(n15696), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n11341), .B(
        n11340), .ZN(n11347) );
  INV_X1 U13386 ( .A(n11439), .ZN(n11345) );
  NAND3_X1 U13387 ( .A1(n15177), .A2(n11343), .A3(n11342), .ZN(n11344) );
  NAND3_X1 U13388 ( .A1(n7362), .A2(n11345), .A3(n11344), .ZN(n11346) );
  OAI211_X1 U13389 ( .C1(n11348), .C2(n15227), .A(n11347), .B(n11346), .ZN(
        P1_U3248) );
  NOR2_X1 U13390 ( .A1(n11350), .A2(n11349), .ZN(n15201) );
  INV_X1 U13391 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12266) );
  MUX2_X1 U13392 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12266), .S(n15212), .Z(
        n11351) );
  OAI21_X1 U13393 ( .B1(n15206), .B2(n15201), .A(n11351), .ZN(n15204) );
  NAND2_X1 U13394 ( .A1(n15212), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11354) );
  INV_X1 U13395 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11352) );
  MUX2_X1 U13396 ( .A(n11352), .B(P1_REG2_REG_11__SCAN_IN), .S(n11614), .Z(
        n11353) );
  AOI21_X1 U13397 ( .B1(n15204), .B2(n11354), .A(n11353), .ZN(n11613) );
  NAND3_X1 U13398 ( .A1(n15204), .A2(n11354), .A3(n11353), .ZN(n11355) );
  NAND2_X1 U13399 ( .A1(n11355), .A2(n7362), .ZN(n11370) );
  OR2_X1 U13400 ( .A1(n11356), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11357) );
  NAND2_X1 U13401 ( .A1(n11358), .A2(n11357), .ZN(n15208) );
  INV_X1 U13402 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11359) );
  MUX2_X1 U13403 ( .A(n11359), .B(P1_REG1_REG_10__SCAN_IN), .S(n15212), .Z(
        n15207) );
  NAND2_X1 U13404 ( .A1(n15212), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11360) );
  INV_X1 U13405 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11361) );
  MUX2_X1 U13406 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11361), .S(n11614), .Z(
        n11362) );
  OAI21_X1 U13407 ( .B1(n11363), .B2(n11362), .A(n15717), .ZN(n11364) );
  NAND2_X1 U13408 ( .A1(n11364), .A2(n15720), .ZN(n11369) );
  NAND2_X1 U13409 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12654)
         );
  INV_X1 U13410 ( .A(n12654), .ZN(n11367) );
  INV_X1 U13411 ( .A(n11614), .ZN(n11365) );
  NOR2_X1 U13412 ( .A1(n15704), .A2(n11365), .ZN(n11366) );
  AOI211_X1 U13413 ( .C1(n15696), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11367), 
        .B(n11366), .ZN(n11368) );
  OAI211_X1 U13414 ( .C1(n11613), .C2(n11370), .A(n11369), .B(n11368), .ZN(
        P1_U3254) );
  INV_X1 U13415 ( .A(n11371), .ZN(n11402) );
  AOI22_X1 U13416 ( .A1(n15723), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15545), .ZN(n11372) );
  OAI21_X1 U13417 ( .B1(n11402), .B2(n15556), .A(n11372), .ZN(P1_U3343) );
  INV_X1 U13418 ( .A(n11373), .ZN(n11375) );
  OAI222_X1 U13419 ( .A1(n14312), .A2(n11375), .B1(n14315), .B2(n11374), .C1(
        n13943), .C2(P3_U3151), .ZN(P3_U3277) );
  MUX2_X1 U13420 ( .A(n15691), .B(n11376), .S(n15689), .Z(n11378) );
  NOR2_X1 U13421 ( .A1(n15689), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n11377) );
  OR2_X1 U13422 ( .A1(n9598), .A2(n11377), .ZN(n15688) );
  NAND2_X1 U13423 ( .A1(n15688), .A2(n15691), .ZN(n15694) );
  OAI211_X1 U13424 ( .C1(n11378), .C2(n15688), .A(P1_U4016), .B(n15694), .ZN(
        n15184) );
  INV_X1 U13425 ( .A(n15184), .ZN(n11392) );
  INV_X1 U13426 ( .A(n11379), .ZN(n11381) );
  MUX2_X1 U13427 ( .A(n11269), .B(P1_REG2_REG_2__SCAN_IN), .S(n11386), .Z(
        n11380) );
  NAND2_X1 U13428 ( .A1(n11381), .A2(n11380), .ZN(n11382) );
  NAND3_X1 U13429 ( .A1(n7362), .A2(n15157), .A3(n11382), .ZN(n11390) );
  AOI22_X1 U13430 ( .A1(n15696), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n11389) );
  OAI211_X1 U13431 ( .C1(n11385), .C2(n11384), .A(n15720), .B(n11383), .ZN(
        n11388) );
  NAND2_X1 U13432 ( .A1(n15722), .A2(n11386), .ZN(n11387) );
  NAND4_X1 U13433 ( .A1(n11390), .A2(n11389), .A3(n11388), .A4(n11387), .ZN(
        n11391) );
  OR2_X1 U13434 ( .A1(n11392), .A2(n11391), .ZN(P1_U3245) );
  INV_X1 U13435 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11393) );
  INV_X1 U13436 ( .A(n11950), .ZN(n12833) );
  OAI222_X1 U13437 ( .A1(n14821), .A2(n11393), .B1(n14819), .B2(n11400), .C1(
        n12833), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13438 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n11395) );
  NAND2_X1 U13439 ( .A1(n16179), .A2(P3_U3897), .ZN(n11394) );
  OAI21_X1 U13440 ( .B1(P3_U3897), .B2(n11395), .A(n11394), .ZN(P3_U3494) );
  INV_X1 U13441 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U13442 ( .A1(n14132), .A2(P3_U3897), .ZN(n11396) );
  OAI21_X1 U13443 ( .B1(P3_U3897), .B2(n11397), .A(n11396), .ZN(P3_U3509) );
  INV_X1 U13444 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n11399) );
  NAND2_X1 U13445 ( .A1(n13442), .A2(P3_U3897), .ZN(n11398) );
  OAI21_X1 U13446 ( .B1(P3_U3897), .B2(n11399), .A(n11398), .ZN(P3_U3510) );
  INV_X1 U13447 ( .A(n11617), .ZN(n11675) );
  OAI222_X1 U13448 ( .A1(P1_U3086), .A2(n11675), .B1(n15558), .B2(n11401), 
        .C1(n11400), .C2(n15556), .ZN(P1_U3342) );
  OAI222_X1 U13449 ( .A1(n14821), .A2(n11403), .B1(n14819), .B2(n11402), .C1(
        n11943), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI22_X1 U13450 ( .A1(n14398), .A2(n11405), .B1(n11404), .B2(n14408), .ZN(
        n11407) );
  NAND2_X1 U13451 ( .A1(n11407), .A2(n11406), .ZN(n11409) );
  AOI22_X1 U13452 ( .A1(n14432), .A2(n16106), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n11760), .ZN(n11408) );
  OAI211_X1 U13453 ( .C1(n16109), .C2(n14417), .A(n11409), .B(n11408), .ZN(
        P2_U3204) );
  NAND2_X1 U13454 ( .A1(n11411), .A2(n11410), .ZN(n11648) );
  INV_X1 U13455 ( .A(n11648), .ZN(n11432) );
  INV_X1 U13456 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n16131) );
  NAND2_X1 U13457 ( .A1(n11414), .A2(n13437), .ZN(n11417) );
  INV_X1 U13458 ( .A(n13450), .ZN(n13003) );
  OAI22_X1 U13459 ( .A1(n12118), .A2(n13451), .B1(n16130), .B2(n13447), .ZN(
        n11415) );
  AOI21_X1 U13460 ( .B1(n13003), .B2(n13893), .A(n11415), .ZN(n11416) );
  OAI211_X1 U13461 ( .C1(n11432), .C2(n16131), .A(n11417), .B(n11416), .ZN(
        P3_U3162) );
  INV_X1 U13462 ( .A(n14417), .ZN(n14423) );
  INV_X1 U13463 ( .A(n12100), .ZN(n11419) );
  OAI21_X1 U13464 ( .B1(n14442), .B2(n11419), .A(n11418), .ZN(n11421) );
  OAI22_X1 U13465 ( .A1(n16323), .A2(n14448), .B1(n14416), .B2(n11424), .ZN(
        n11420) );
  AOI211_X1 U13466 ( .C1(n14423), .C2(n14468), .A(n11421), .B(n11420), .ZN(
        n11428) );
  INV_X1 U13467 ( .A(n11422), .ZN(n11426) );
  OAI22_X1 U13468 ( .A1(n14398), .A2(n11424), .B1(n11423), .B2(n14408), .ZN(
        n11425) );
  NAND3_X1 U13469 ( .A1(n11426), .A2(n11704), .A3(n11425), .ZN(n11427) );
  OAI211_X1 U13470 ( .C1(n14427), .C2(n11429), .A(n11428), .B(n11427), .ZN(
        P2_U3199) );
  INV_X1 U13471 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15904) );
  NAND2_X1 U13472 ( .A1(n13893), .A2(n11928), .ZN(n13140) );
  NAND2_X1 U13473 ( .A1(n13142), .A2(n13140), .ZN(n13309) );
  OAI22_X1 U13474 ( .A1(n10122), .A2(n13451), .B1(n11928), .B2(n13447), .ZN(
        n11430) );
  AOI21_X1 U13475 ( .B1(n13437), .B2(n13309), .A(n11430), .ZN(n11431) );
  OAI21_X1 U13476 ( .B1(n11432), .B2(n15904), .A(n11431), .ZN(P3_U3172) );
  INV_X1 U13477 ( .A(n11433), .ZN(n11436) );
  MUX2_X1 U13478 ( .A(n11277), .B(P1_REG2_REG_6__SCAN_IN), .S(n11434), .Z(
        n11435) );
  NAND2_X1 U13479 ( .A1(n11436), .A2(n11435), .ZN(n11438) );
  OAI211_X1 U13480 ( .C1(n11439), .C2(n11438), .A(n7362), .B(n11437), .ZN(
        n11442) );
  NAND2_X1 U13481 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11723) );
  INV_X1 U13482 ( .A(n11723), .ZN(n11440) );
  AOI21_X1 U13483 ( .B1(n15696), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n11440), .ZN(
        n11441) );
  OAI211_X1 U13484 ( .C1(n15704), .C2(n11443), .A(n11442), .B(n11441), .ZN(
        n11449) );
  INV_X1 U13485 ( .A(n11444), .ZN(n11445) );
  AOI211_X1 U13486 ( .C1(n11447), .C2(n11446), .A(n11445), .B(n15227), .ZN(
        n11448) );
  OR2_X1 U13487 ( .A1(n11449), .A2(n11448), .ZN(P1_U3249) );
  OAI222_X1 U13488 ( .A1(P3_U3151), .A2(n11452), .B1(n14315), .B2(n11451), 
        .C1(n14312), .C2(n11450), .ZN(P3_U3276) );
  INV_X1 U13489 ( .A(n14751), .ZN(n16456) );
  INV_X1 U13490 ( .A(n11456), .ZN(n11454) );
  XNOR2_X1 U13491 ( .A(n11454), .B(n11453), .ZN(n11913) );
  OAI21_X1 U13492 ( .B1(n11457), .B2(n11456), .A(n11455), .ZN(n11458) );
  NAND2_X1 U13493 ( .A1(n11458), .A2(n16107), .ZN(n11460) );
  AOI22_X1 U13494 ( .A1(n14628), .A2(n14467), .B1(n14469), .B2(n14627), .ZN(
        n11459) );
  AND2_X1 U13495 ( .A1(n11460), .A2(n11459), .ZN(n11904) );
  NAND2_X1 U13496 ( .A1(n11906), .A2(n12099), .ZN(n11461) );
  NAND2_X1 U13497 ( .A1(n11461), .A2(n16261), .ZN(n11462) );
  OR2_X1 U13498 ( .A1(n11462), .A2(n12084), .ZN(n11905) );
  OAI211_X1 U13499 ( .C1(n16456), .C2(n11913), .A(n11904), .B(n11905), .ZN(
        n11465) );
  NAND2_X1 U13500 ( .A1(n11465), .A2(n16512), .ZN(n11464) );
  AOI22_X1 U13501 ( .A1(n14757), .A2(n11906), .B1(n16510), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11463) );
  NAND2_X1 U13502 ( .A1(n11464), .A2(n11463), .ZN(P2_U3505) );
  NAND2_X1 U13503 ( .A1(n11465), .A2(n16516), .ZN(n11469) );
  INV_X1 U13504 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11466) );
  NOR2_X1 U13505 ( .A1(n16516), .A2(n11466), .ZN(n11467) );
  AOI21_X1 U13506 ( .B1(n14792), .B2(n11906), .A(n11467), .ZN(n11468) );
  NAND2_X1 U13507 ( .A1(n11469), .A2(n11468), .ZN(P2_U3448) );
  INV_X1 U13508 ( .A(n11472), .ZN(n11473) );
  NAND2_X1 U13509 ( .A1(n11474), .A2(n11473), .ZN(n11475) );
  NAND2_X1 U13510 ( .A1(n14985), .A2(n14950), .ZN(n11478) );
  NAND2_X1 U13511 ( .A1(n15141), .A2(n14900), .ZN(n11477) );
  NAND2_X1 U13512 ( .A1(n11478), .A2(n11477), .ZN(n11479) );
  XNOR2_X1 U13513 ( .A(n11479), .B(n15001), .ZN(n11482) );
  INV_X2 U13514 ( .A(n15005), .ZN(n14954) );
  NAND2_X1 U13515 ( .A1(n14985), .A2(n14954), .ZN(n11481) );
  NAND2_X1 U13516 ( .A1(n14955), .A2(n15141), .ZN(n11480) );
  NAND2_X1 U13517 ( .A1(n11481), .A2(n11480), .ZN(n11483) );
  NAND2_X1 U13518 ( .A1(n11482), .A2(n11483), .ZN(n11487) );
  INV_X1 U13519 ( .A(n11482), .ZN(n11485) );
  INV_X1 U13520 ( .A(n11483), .ZN(n11484) );
  NAND2_X1 U13521 ( .A1(n11485), .A2(n11484), .ZN(n11486) );
  NAND2_X1 U13522 ( .A1(n11487), .A2(n11486), .ZN(n14981) );
  NAND2_X1 U13523 ( .A1(n11816), .A2(n14900), .ZN(n11489) );
  OR2_X1 U13524 ( .A1(n12048), .A2(n15003), .ZN(n11488) );
  NAND2_X1 U13525 ( .A1(n11489), .A2(n11488), .ZN(n11490) );
  OR2_X1 U13526 ( .A1(n11491), .A2(n11490), .ZN(n11519) );
  NAND2_X1 U13527 ( .A1(n11491), .A2(n11490), .ZN(n11518) );
  NAND2_X1 U13528 ( .A1(n11519), .A2(n11518), .ZN(n11495) );
  NAND2_X1 U13529 ( .A1(n11816), .A2(n14950), .ZN(n11493) );
  OR2_X1 U13530 ( .A1(n12048), .A2(n15005), .ZN(n11492) );
  NAND2_X1 U13531 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  XNOR2_X1 U13532 ( .A(n11494), .B(n14925), .ZN(n11517) );
  XNOR2_X1 U13533 ( .A(n11495), .B(n11517), .ZN(n11503) );
  AOI22_X1 U13534 ( .A1(n15140), .A2(n15099), .B1(n15100), .B2(n15141), .ZN(
        n16286) );
  INV_X1 U13535 ( .A(n11496), .ZN(n11497) );
  OAI21_X1 U13536 ( .B1(n11498), .B2(n11497), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U13537 ( .A1(n15104), .A2(n11811), .ZN(n11500) );
  NAND2_X1 U13538 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n15169) );
  OAI211_X1 U13539 ( .C1(n16286), .C2(n15102), .A(n11500), .B(n15169), .ZN(
        n11501) );
  AOI21_X1 U13540 ( .B1(n11816), .B2(n16551), .A(n11501), .ZN(n11502) );
  OAI21_X1 U13541 ( .B1(n11503), .B2(n15115), .A(n11502), .ZN(P1_U3230) );
  INV_X1 U13542 ( .A(n11504), .ZN(n11508) );
  OAI22_X1 U13543 ( .A1(n11506), .A2(n14408), .B1(n11505), .B2(n14398), .ZN(
        n11507) );
  NAND3_X1 U13544 ( .A1(n11508), .A2(n11632), .A3(n11507), .ZN(n11514) );
  AOI22_X1 U13545 ( .A1(n14628), .A2(n14465), .B1(n14467), .B2(n14627), .ZN(
        n11896) );
  OAI22_X1 U13546 ( .A1(n14386), .A2(n11896), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11509), .ZN(n11512) );
  INV_X1 U13547 ( .A(n12058), .ZN(n11510) );
  NOR2_X1 U13548 ( .A1(n11510), .A2(n14448), .ZN(n11511) );
  AOI211_X1 U13549 ( .C1(n14420), .C2(n12057), .A(n11512), .B(n11511), .ZN(
        n11513) );
  OAI211_X1 U13550 ( .C1(n11683), .C2(n14408), .A(n11514), .B(n11513), .ZN(
        P2_U3193) );
  INV_X1 U13551 ( .A(n11515), .ZN(n11604) );
  AOI22_X1 U13552 ( .A1(n12311), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n15545), .ZN(n11516) );
  OAI21_X1 U13553 ( .B1(n11604), .B2(n15556), .A(n11516), .ZN(P1_U3341) );
  NAND2_X1 U13554 ( .A1(n11518), .A2(n11517), .ZN(n11520) );
  NAND2_X1 U13555 ( .A1(n16314), .A2(n14950), .ZN(n11522) );
  NAND2_X1 U13556 ( .A1(n15140), .A2(n14900), .ZN(n11521) );
  NAND2_X1 U13557 ( .A1(n11522), .A2(n11521), .ZN(n11523) );
  XNOR2_X1 U13558 ( .A(n11523), .B(n14925), .ZN(n11705) );
  NOR2_X1 U13559 ( .A1(n11823), .A2(n15003), .ZN(n11524) );
  AOI21_X1 U13560 ( .B1(n16314), .B2(n14900), .A(n11524), .ZN(n11706) );
  XNOR2_X1 U13561 ( .A(n11705), .B(n11706), .ZN(n11525) );
  XNOR2_X1 U13562 ( .A(n11711), .B(n11525), .ZN(n11533) );
  INV_X1 U13563 ( .A(n11526), .ZN(n16311) );
  OR2_X1 U13564 ( .A1(n12048), .A2(n15399), .ZN(n11528) );
  NAND2_X1 U13565 ( .A1(n15139), .A2(n15099), .ZN(n11527) );
  AND2_X1 U13566 ( .A1(n11528), .A2(n11527), .ZN(n11591) );
  NAND2_X1 U13567 ( .A1(n16314), .A2(n16551), .ZN(n11530) );
  OAI211_X1 U13568 ( .C1(n11591), .C2(n15102), .A(n11530), .B(n11529), .ZN(
        n11531) );
  AOI21_X1 U13569 ( .B1(n15104), .B2(n16311), .A(n11531), .ZN(n11532) );
  OAI21_X1 U13570 ( .B1(n11533), .B2(n15115), .A(n11532), .ZN(P1_U3227) );
  AOI21_X1 U13571 ( .B1(n11538), .B2(P2_REG1_REG_10__SCAN_IN), .A(n11534), 
        .ZN(n15616) );
  INV_X1 U13572 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n16463) );
  MUX2_X1 U13573 ( .A(n16463), .B(P2_REG1_REG_11__SCAN_IN), .S(n11541), .Z(
        n15615) );
  NOR2_X1 U13574 ( .A1(n15616), .A2(n15615), .ZN(n15614) );
  AOI21_X1 U13575 ( .B1(n11541), .B2(P2_REG1_REG_11__SCAN_IN), .A(n15614), 
        .ZN(n11537) );
  INV_X1 U13576 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11535) );
  MUX2_X1 U13577 ( .A(n11535), .B(P2_REG1_REG_12__SCAN_IN), .S(n11943), .Z(
        n11536) );
  NAND2_X1 U13578 ( .A1(n11537), .A2(n11536), .ZN(n11935) );
  OAI21_X1 U13579 ( .B1(n11537), .B2(n11536), .A(n11935), .ZN(n11552) );
  NAND2_X1 U13580 ( .A1(n11538), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11539) );
  NAND2_X1 U13581 ( .A1(n11540), .A2(n11539), .ZN(n15607) );
  INV_X1 U13582 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12249) );
  MUX2_X1 U13583 ( .A(n12249), .B(P2_REG2_REG_11__SCAN_IN), .S(n11541), .Z(
        n15606) );
  NOR2_X1 U13584 ( .A1(n15607), .A2(n15606), .ZN(n15609) );
  AND2_X1 U13585 ( .A1(n15611), .A2(n12249), .ZN(n11544) );
  INV_X1 U13586 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11542) );
  MUX2_X1 U13587 ( .A(n11542), .B(P2_REG2_REG_12__SCAN_IN), .S(n11943), .Z(
        n11543) );
  OAI21_X1 U13588 ( .B1(n15609), .B2(n11544), .A(n11543), .ZN(n11941) );
  INV_X1 U13589 ( .A(n15609), .ZN(n11547) );
  INV_X1 U13590 ( .A(n11543), .ZN(n11546) );
  INV_X1 U13591 ( .A(n11544), .ZN(n11545) );
  NAND3_X1 U13592 ( .A1(n11547), .A2(n11546), .A3(n11545), .ZN(n11548) );
  AOI21_X1 U13593 ( .B1(n11941), .B2(n11548), .A(n15686), .ZN(n11551) );
  NAND2_X1 U13594 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n12401)
         );
  NAND2_X1 U13595 ( .A1(n15684), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n11549) );
  OAI211_X1 U13596 ( .C1(n15626), .C2(n11943), .A(n12401), .B(n11549), .ZN(
        n11550) );
  AOI211_X1 U13597 ( .C1(n11552), .C2(n15668), .A(n11551), .B(n11550), .ZN(
        n11553) );
  INV_X1 U13598 ( .A(n11553), .ZN(P2_U3226) );
  AND2_X1 U13599 ( .A1(n11555), .A2(n11554), .ZN(n11790) );
  OAI21_X1 U13600 ( .B1(n11557), .B2(P1_D_REG_1__SCAN_IN), .A(n11556), .ZN(
        n11561) );
  NAND2_X1 U13601 ( .A1(n11559), .A2(n11558), .ZN(n11560) );
  NAND4_X1 U13602 ( .A1(n11790), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n11600) );
  INV_X1 U13603 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n11598) );
  AND2_X1 U13604 ( .A1(n12770), .A2(n7363), .ZN(n11563) );
  NAND2_X1 U13605 ( .A1(n11564), .A2(n11563), .ZN(n16485) );
  INV_X1 U13606 ( .A(n11793), .ZN(n11569) );
  NAND2_X1 U13607 ( .A1(n11565), .A2(n9047), .ZN(n16138) );
  NAND2_X1 U13608 ( .A1(n16139), .A2(n16138), .ZN(n11568) );
  OR2_X1 U13609 ( .A1(n15143), .A2(n11566), .ZN(n11567) );
  NAND2_X1 U13610 ( .A1(n11569), .A2(n11788), .ZN(n11571) );
  INV_X1 U13611 ( .A(n12042), .ZN(n11572) );
  NAND2_X1 U13612 ( .A1(n12040), .A2(n11572), .ZN(n11575) );
  NAND2_X1 U13613 ( .A1(n16242), .A2(n11573), .ZN(n11574) );
  NAND2_X1 U13614 ( .A1(n11575), .A2(n11574), .ZN(n11806) );
  NAND2_X1 U13615 ( .A1(n11806), .A2(n11807), .ZN(n11578) );
  OR2_X1 U13616 ( .A1(n11816), .A2(n11576), .ZN(n11577) );
  XNOR2_X1 U13617 ( .A(n11822), .B(n11587), .ZN(n16316) );
  INV_X1 U13618 ( .A(n16316), .ZN(n11596) );
  OR2_X1 U13619 ( .A1(n11580), .A2(n11579), .ZN(n11581) );
  NAND2_X1 U13620 ( .A1(n11805), .A2(n12559), .ZN(n16085) );
  INV_X1 U13621 ( .A(n16085), .ZN(n16488) );
  NAND2_X1 U13622 ( .A1(n11794), .A2(n11793), .ZN(n11792) );
  NAND2_X1 U13623 ( .A1(n11582), .A2(n11802), .ZN(n11583) );
  NAND2_X1 U13624 ( .A1(n11792), .A2(n11583), .ZN(n12043) );
  NAND2_X1 U13625 ( .A1(n12043), .A2(n12042), .ZN(n12041) );
  NAND2_X1 U13626 ( .A1(n12041), .A2(n11584), .ZN(n11808) );
  OR2_X1 U13627 ( .A1(n11816), .A2(n12048), .ZN(n11585) );
  NAND2_X1 U13628 ( .A1(n11816), .A2(n12048), .ZN(n11586) );
  XNOR2_X1 U13629 ( .A(n11827), .B(n11587), .ZN(n11592) );
  NAND2_X1 U13630 ( .A1(n15559), .A2(n7363), .ZN(n11590) );
  NAND2_X1 U13631 ( .A1(n11588), .A2(n7690), .ZN(n11589) );
  OAI21_X1 U13632 ( .B1(n11592), .B2(n16532), .A(n11591), .ZN(n11593) );
  AOI21_X1 U13633 ( .B1(n16488), .B2(n16316), .A(n11593), .ZN(n16321) );
  INV_X1 U13634 ( .A(n11816), .ZN(n16288) );
  AND2_X1 U13635 ( .A1(n16155), .A2(n16142), .ZN(n16140) );
  NAND2_X1 U13636 ( .A1(n16140), .A2(n16204), .ZN(n12045) );
  INV_X1 U13637 ( .A(n11594), .ZN(n11813) );
  INV_X1 U13638 ( .A(n16314), .ZN(n11824) );
  NAND2_X1 U13639 ( .A1(n11824), .A2(n11594), .ZN(n11833) );
  INV_X1 U13640 ( .A(n11833), .ZN(n11835) );
  AOI211_X1 U13641 ( .C1(n16314), .C2(n11813), .A(n16495), .B(n11835), .ZN(
        n16318) );
  AOI21_X1 U13642 ( .B1(n16314), .B2(n16528), .A(n16318), .ZN(n11595) );
  OAI211_X1 U13643 ( .C1(n16485), .C2(n11596), .A(n16321), .B(n11595), .ZN(
        n11601) );
  NAND2_X1 U13644 ( .A1(n11601), .A2(n16539), .ZN(n11597) );
  OAI21_X1 U13645 ( .B1(n16539), .B2(n11598), .A(n11597), .ZN(P1_U3533) );
  INV_X1 U13646 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U13647 ( .A1(n11601), .A2(n16543), .ZN(n11602) );
  OAI21_X1 U13648 ( .B1(n16543), .B2(n11603), .A(n11602), .ZN(P1_U3474) );
  OAI222_X1 U13649 ( .A1(n14821), .A2(n11605), .B1(n14819), .B2(n11604), .C1(
        P2_U3088), .C2(n15625), .ZN(P2_U3313) );
  OR2_X1 U13650 ( .A1(n11614), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n15716) );
  NAND2_X1 U13651 ( .A1(n15717), .A2(n15716), .ZN(n11608) );
  INV_X1 U13652 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11606) );
  MUX2_X1 U13653 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n11606), .S(n15723), .Z(
        n11607) );
  NAND2_X1 U13654 ( .A1(n11608), .A2(n11607), .ZN(n15719) );
  OR2_X1 U13655 ( .A1(n15723), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11609) );
  NAND2_X1 U13656 ( .A1(n15719), .A2(n11609), .ZN(n11671) );
  INV_X1 U13657 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11610) );
  MUX2_X1 U13658 ( .A(n11610), .B(P1_REG1_REG_13__SCAN_IN), .S(n11617), .Z(
        n11672) );
  NAND2_X1 U13659 ( .A1(n11617), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11611) );
  XNOR2_X1 U13660 ( .A(n12304), .B(n12311), .ZN(n12305) );
  INV_X1 U13661 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11612) );
  XNOR2_X1 U13662 ( .A(n12305), .B(n11612), .ZN(n11628) );
  AOI21_X1 U13663 ( .B1(n11614), .B2(P1_REG2_REG_11__SCAN_IN), .A(n11613), 
        .ZN(n15713) );
  INV_X1 U13664 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11615) );
  MUX2_X1 U13665 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11615), .S(n15723), .Z(
        n15714) );
  NAND2_X1 U13666 ( .A1(n15713), .A2(n15714), .ZN(n15712) );
  OAI21_X1 U13667 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n15723), .A(n15712), 
        .ZN(n11668) );
  INV_X1 U13668 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11616) );
  MUX2_X1 U13669 ( .A(n11616), .B(P1_REG2_REG_13__SCAN_IN), .S(n11617), .Z(
        n11667) );
  NAND2_X1 U13670 ( .A1(n11617), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11620) );
  INV_X1 U13671 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11618) );
  MUX2_X1 U13672 ( .A(n11618), .B(P1_REG2_REG_14__SCAN_IN), .S(n12311), .Z(
        n11619) );
  AOI21_X1 U13673 ( .B1(n11665), .B2(n11620), .A(n11619), .ZN(n12310) );
  INV_X1 U13674 ( .A(n12310), .ZN(n11622) );
  NAND3_X1 U13675 ( .A1(n11665), .A2(n11620), .A3(n11619), .ZN(n11621) );
  NAND3_X1 U13676 ( .A1(n11622), .A2(n7362), .A3(n11621), .ZN(n11627) );
  NAND2_X1 U13677 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n16524)
         );
  INV_X1 U13678 ( .A(n16524), .ZN(n11625) );
  INV_X1 U13679 ( .A(n12311), .ZN(n11623) );
  NOR2_X1 U13680 ( .A1(n15704), .A2(n11623), .ZN(n11624) );
  AOI211_X1 U13681 ( .C1(n15696), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11625), 
        .B(n11624), .ZN(n11626) );
  OAI211_X1 U13682 ( .C1(n11628), .C2(n15227), .A(n11627), .B(n11626), .ZN(
        P1_U3257) );
  INV_X1 U13683 ( .A(n11629), .ZN(n11653) );
  NOR3_X1 U13684 ( .A1(n11630), .A2(n11635), .A3(n14398), .ZN(n11631) );
  AOI21_X1 U13685 ( .B1(n11653), .B2(n14437), .A(n11631), .ZN(n11642) );
  NOR2_X1 U13686 ( .A1(n11632), .A2(n14408), .ZN(n11639) );
  AND2_X1 U13687 ( .A1(n12086), .A2(n14432), .ZN(n11638) );
  INV_X1 U13688 ( .A(n12085), .ZN(n11634) );
  OAI21_X1 U13689 ( .B1(n14442), .B2(n11634), .A(n11633), .ZN(n11637) );
  OAI22_X1 U13690 ( .A1(n11680), .A2(n14417), .B1(n14416), .B2(n11635), .ZN(
        n11636) );
  NOR4_X1 U13691 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n11640) );
  OAI21_X1 U13692 ( .B1(n11642), .B2(n11641), .A(n11640), .ZN(P2_U3185) );
  XOR2_X1 U13693 ( .A(n11644), .B(n11643), .Z(n11650) );
  INV_X1 U13694 ( .A(n13437), .ZN(n13458) );
  INV_X1 U13695 ( .A(n13451), .ZN(n13441) );
  AOI22_X1 U13696 ( .A1(n16179), .A2(n13441), .B1(n13455), .B2(n11645), .ZN(
        n11646) );
  OAI21_X1 U13697 ( .B1(n10122), .B2(n13450), .A(n11646), .ZN(n11647) );
  AOI21_X1 U13698 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n11648), .A(n11647), .ZN(
        n11649) );
  OAI21_X1 U13699 ( .B1(n11650), .B2(n13458), .A(n11649), .ZN(P3_U3177) );
  INV_X1 U13700 ( .A(n11651), .ZN(n11907) );
  INV_X1 U13701 ( .A(n14416), .ZN(n14424) );
  AOI22_X1 U13702 ( .A1(n14423), .A2(n14467), .B1(n14424), .B2(n14469), .ZN(
        n11652) );
  NAND2_X1 U13703 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15592) );
  OAI211_X1 U13704 ( .C1(n11907), .C2(n14442), .A(n11652), .B(n15592), .ZN(
        n11657) );
  AOI211_X1 U13705 ( .C1(n11655), .C2(n11654), .A(n14427), .B(n11653), .ZN(
        n11656) );
  AOI211_X1 U13706 ( .C1(n11906), .C2(n14432), .A(n11657), .B(n11656), .ZN(
        n11658) );
  INV_X1 U13707 ( .A(n11658), .ZN(P2_U3211) );
  OAI211_X1 U13708 ( .C1(n11661), .C2(n11660), .A(n11659), .B(n13437), .ZN(
        n11664) );
  NOR2_X1 U13709 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13734), .ZN(n15908) );
  OAI22_X1 U13710 ( .A1(n12119), .A2(n13451), .B1(n12118), .B2(n13450), .ZN(
        n11662) );
  AOI211_X1 U13711 ( .C1(n13455), .C2(n12128), .A(n15908), .B(n11662), .ZN(
        n11663) );
  OAI211_X1 U13712 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12702), .A(n11664), .B(
        n11663), .ZN(P3_U3158) );
  INV_X1 U13714 ( .A(n11665), .ZN(n11666) );
  AOI211_X1 U13715 ( .C1(n11668), .C2(n11667), .A(n16567), .B(n11666), .ZN(
        n11678) );
  INV_X1 U13716 ( .A(n11669), .ZN(n11670) );
  AOI211_X1 U13717 ( .C1(n11672), .C2(n11671), .A(n15227), .B(n11670), .ZN(
        n11677) );
  NAND2_X1 U13718 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n12869)
         );
  INV_X1 U13719 ( .A(n12869), .ZN(n11673) );
  AOI21_X1 U13720 ( .B1(n15696), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11673), 
        .ZN(n11674) );
  OAI21_X1 U13721 ( .B1(n11675), .B2(n15704), .A(n11674), .ZN(n11676) );
  OR3_X1 U13722 ( .A1(n11678), .A2(n11677), .A3(n11676), .ZN(P1_U3256) );
  INV_X1 U13723 ( .A(n11679), .ZN(n11684) );
  OAI22_X1 U13724 ( .A1(n11681), .A2(n14408), .B1(n11680), .B2(n14398), .ZN(
        n11682) );
  NAND3_X1 U13725 ( .A1(n11684), .A2(n11683), .A3(n11682), .ZN(n11689) );
  AOI22_X1 U13726 ( .A1(n14627), .A2(n14466), .B1(n14464), .B2(n14628), .ZN(
        n12200) );
  OAI22_X1 U13727 ( .A1(n14386), .A2(n12200), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11685), .ZN(n11687) );
  NOR2_X1 U13728 ( .A1(n12206), .A2(n14448), .ZN(n11686) );
  AOI211_X1 U13729 ( .C1(n14420), .C2(n16398), .A(n11687), .B(n11686), .ZN(
        n11688) );
  OAI211_X1 U13730 ( .C1(n12030), .C2(n14408), .A(n11689), .B(n11688), .ZN(
        P2_U3203) );
  INV_X1 U13731 ( .A(n11690), .ZN(n11854) );
  NAND2_X1 U13732 ( .A1(n14469), .A2(n14628), .ZN(n11692) );
  NAND2_X1 U13733 ( .A1(n14471), .A2(n14627), .ZN(n11691) );
  NAND2_X1 U13734 ( .A1(n11692), .A2(n11691), .ZN(n11858) );
  NAND2_X1 U13735 ( .A1(n14445), .A2(n11858), .ZN(n11694) );
  OAI211_X1 U13736 ( .C1(n14442), .C2(n11854), .A(n11694), .B(n11693), .ZN(
        n11702) );
  NOR3_X1 U13737 ( .A1(n14398), .A2(n11696), .A3(n11695), .ZN(n11697) );
  AOI21_X1 U13738 ( .B1(n14437), .B2(n11698), .A(n11697), .ZN(n11700) );
  NOR2_X1 U13739 ( .A1(n11700), .A2(n11699), .ZN(n11701) );
  AOI211_X1 U13740 ( .C1(n11853), .C2(n14432), .A(n11702), .B(n11701), .ZN(
        n11703) );
  OAI21_X1 U13741 ( .B1(n11704), .B2(n14408), .A(n11703), .ZN(P2_U3202) );
  AND2_X1 U13742 ( .A1(n11705), .A2(n11706), .ZN(n11710) );
  INV_X1 U13743 ( .A(n11705), .ZN(n11708) );
  INV_X1 U13744 ( .A(n11706), .ZN(n11707) );
  NAND2_X1 U13745 ( .A1(n11708), .A2(n11707), .ZN(n11709) );
  NAND2_X1 U13746 ( .A1(n11838), .A2(n14950), .ZN(n11713) );
  NAND2_X1 U13747 ( .A1(n15139), .A2(n14954), .ZN(n11712) );
  NAND2_X1 U13748 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  XNOR2_X1 U13749 ( .A(n11714), .B(n15001), .ZN(n11720) );
  INV_X1 U13750 ( .A(n11720), .ZN(n11718) );
  NAND2_X1 U13751 ( .A1(n11838), .A2(n14954), .ZN(n11716) );
  NAND2_X1 U13752 ( .A1(n14955), .A2(n15139), .ZN(n11715) );
  NAND2_X1 U13753 ( .A1(n11716), .A2(n11715), .ZN(n11719) );
  INV_X1 U13754 ( .A(n11719), .ZN(n11717) );
  NAND2_X1 U13755 ( .A1(n11718), .A2(n11717), .ZN(n11867) );
  INV_X1 U13756 ( .A(n11867), .ZN(n11721) );
  AND2_X1 U13757 ( .A1(n11720), .A2(n11719), .ZN(n11868) );
  NOR2_X1 U13758 ( .A1(n11721), .A2(n11868), .ZN(n11722) );
  XNOR2_X1 U13759 ( .A(n11869), .B(n11722), .ZN(n11727) );
  AOI22_X1 U13760 ( .A1(n15140), .A2(n15100), .B1(n15099), .B2(n15138), .ZN(
        n11829) );
  NAND2_X1 U13761 ( .A1(n15104), .A2(n11831), .ZN(n11724) );
  OAI211_X1 U13762 ( .C1(n11829), .C2(n15102), .A(n11724), .B(n11723), .ZN(
        n11725) );
  AOI21_X1 U13763 ( .B1(n11838), .B2(n16551), .A(n11725), .ZN(n11726) );
  OAI21_X1 U13764 ( .B1(n11727), .B2(n15115), .A(n11726), .ZN(P1_U3239) );
  INV_X1 U13765 ( .A(n11728), .ZN(n11729) );
  AOI21_X1 U13766 ( .B1(n11731), .B2(n11730), .A(n11729), .ZN(n11735) );
  INV_X1 U13767 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n13756) );
  NOR2_X1 U13768 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13756), .ZN(n15935) );
  OAI22_X1 U13769 ( .A1(n12293), .A2(n13451), .B1(n12136), .B2(n13450), .ZN(
        n11732) );
  AOI211_X1 U13770 ( .C1(n13455), .C2(n12141), .A(n15935), .B(n11732), .ZN(
        n11734) );
  NAND2_X1 U13771 ( .A1(n13454), .A2(n12140), .ZN(n11733) );
  OAI211_X1 U13772 ( .C1(n11735), .C2(n13458), .A(n11734), .B(n11733), .ZN(
        P3_U3170) );
  AND2_X1 U13773 ( .A1(n11736), .A2(n15571), .ZN(n11737) );
  NAND4_X1 U13774 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n15570), .ZN(
        n11745) );
  INV_X2 U13775 ( .A(n14675), .ZN(n16408) );
  XNOR2_X1 U13776 ( .A(n11740), .B(n11757), .ZN(n11742) );
  AOI21_X1 U13777 ( .B1(n11742), .B2(n16107), .A(n11741), .ZN(n16167) );
  NOR2_X1 U13778 ( .A1(n14675), .A2(n11744), .ZN(n11751) );
  INV_X1 U13779 ( .A(n11745), .ZN(n11746) );
  INV_X1 U13780 ( .A(n16213), .ZN(n11748) );
  AOI21_X1 U13781 ( .B1(n11752), .B2(n16106), .A(n14491), .ZN(n11747) );
  NAND2_X1 U13782 ( .A1(n11748), .A2(n11747), .ZN(n16166) );
  OAI22_X1 U13783 ( .A1(n16228), .A2(n16166), .B1(n11749), .B2(n16117), .ZN(
        n11750) );
  AOI211_X1 U13784 ( .C1(n16399), .C2(n11752), .A(n11751), .B(n11750), .ZN(
        n11759) );
  AND2_X1 U13785 ( .A1(n11753), .A2(n12849), .ZN(n16122) );
  INV_X1 U13786 ( .A(n16122), .ZN(n11754) );
  NAND2_X1 U13787 ( .A1(n16431), .A2(n11754), .ZN(n11755) );
  XNOR2_X1 U13788 ( .A(n11757), .B(n11756), .ZN(n16164) );
  NAND2_X1 U13789 ( .A1(n14678), .A2(n16164), .ZN(n11758) );
  OAI211_X1 U13790 ( .C1(n16408), .C2(n16167), .A(n11759), .B(n11758), .ZN(
        P2_U3264) );
  AOI22_X1 U13791 ( .A1(n14627), .A2(n14473), .B1(n14471), .B2(n14628), .ZN(
        n16217) );
  INV_X1 U13792 ( .A(n11760), .ZN(n11762) );
  INV_X1 U13793 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11761) );
  OAI22_X1 U13794 ( .A1(n14386), .A2(n16217), .B1(n11762), .B2(n11761), .ZN(
        n11769) );
  INV_X1 U13795 ( .A(n14398), .ZN(n14411) );
  AOI22_X1 U13796 ( .A1(n14411), .A2(n14473), .B1(n14437), .B2(n11763), .ZN(
        n11767) );
  INV_X1 U13797 ( .A(n11764), .ZN(n11766) );
  NOR3_X1 U13798 ( .A1(n11767), .A2(n11766), .A3(n11765), .ZN(n11768) );
  AOI211_X1 U13799 ( .C1(n16225), .C2(n14432), .A(n11769), .B(n11768), .ZN(
        n11770) );
  OAI21_X1 U13800 ( .B1(n11771), .B2(n14408), .A(n11770), .ZN(P2_U3209) );
  INV_X1 U13801 ( .A(n11772), .ZN(n11773) );
  OAI222_X1 U13802 ( .A1(P3_U3151), .A2(n11774), .B1(n14315), .B2(n13668), 
        .C1(n14312), .C2(n11773), .ZN(P3_U3275) );
  INV_X1 U13803 ( .A(n11775), .ZN(n12016) );
  AOI21_X1 U13804 ( .B1(n11776), .B2(n15898), .A(n12016), .ZN(n11787) );
  XNOR2_X1 U13805 ( .A(n11777), .B(P3_REG1_REG_1__SCAN_IN), .ZN(n11783) );
  OAI22_X1 U13806 ( .A1(n15981), .A2(n15733), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n16131), .ZN(n11782) );
  NAND2_X1 U13807 ( .A1(n11778), .A2(n16137), .ZN(n11779) );
  AOI21_X1 U13808 ( .B1(n11780), .B2(n11779), .A(n16082), .ZN(n11781) );
  AOI211_X1 U13809 ( .C1(n16079), .C2(n11783), .A(n11782), .B(n11781), .ZN(
        n11786) );
  NAND2_X1 U13810 ( .A1(n16043), .A2(n11784), .ZN(n11785) );
  OAI211_X1 U13811 ( .C1(n11787), .C2(n16069), .A(n11786), .B(n11785), .ZN(
        P3_U3183) );
  XNOR2_X1 U13812 ( .A(n11788), .B(n11793), .ZN(n16203) );
  NAND3_X1 U13813 ( .A1(n11791), .A2(n11790), .A3(n11789), .ZN(n13079) );
  OAI21_X1 U13814 ( .B1(n11794), .B2(n11793), .A(n11792), .ZN(n11796) );
  AOI21_X1 U13815 ( .B1(n11796), .B2(n16248), .A(n11795), .ZN(n11797) );
  OAI21_X1 U13816 ( .B1(n16085), .B2(n16203), .A(n11797), .ZN(n16206) );
  NAND2_X1 U13817 ( .A1(n16206), .A2(n15352), .ZN(n11804) );
  OR2_X1 U13818 ( .A1(n13079), .A2(n15269), .ZN(n16099) );
  OAI21_X1 U13819 ( .B1(n16140), .B2(n16204), .A(n12045), .ZN(n16205) );
  INV_X1 U13820 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11799) );
  OAI22_X1 U13821 ( .A1(n16099), .A2(n16205), .B1(n11799), .B2(n16104), .ZN(
        n11801) );
  NOR2_X1 U13822 ( .A1(n15352), .A2(n11269), .ZN(n11800) );
  AOI211_X1 U13823 ( .C1(n16313), .C2(n11802), .A(n11801), .B(n11800), .ZN(
        n11803) );
  OAI211_X1 U13824 ( .C1(n16203), .C2(n13351), .A(n11804), .B(n11803), .ZN(
        P1_U3291) );
  INV_X1 U13825 ( .A(n11805), .ZN(n12276) );
  XNOR2_X1 U13826 ( .A(n11806), .B(n9106), .ZN(n16285) );
  XNOR2_X1 U13827 ( .A(n11808), .B(n11807), .ZN(n11809) );
  NOR2_X1 U13828 ( .A1(n11809), .A2(n16532), .ZN(n16289) );
  INV_X1 U13829 ( .A(n16286), .ZN(n11810) );
  OAI21_X1 U13830 ( .B1(n16289), .B2(n11810), .A(n15352), .ZN(n11818) );
  INV_X1 U13831 ( .A(n11811), .ZN(n11812) );
  OAI22_X1 U13832 ( .A1(n15352), .A2(n11273), .B1(n11812), .B2(n16104), .ZN(
        n11815) );
  OAI211_X1 U13833 ( .C1(n16288), .C2(n12044), .A(n11813), .B(n15501), .ZN(
        n16287) );
  OR2_X1 U13834 ( .A1(n13079), .A2(n7363), .ZN(n15372) );
  NOR2_X1 U13835 ( .A1(n16287), .A2(n15372), .ZN(n11814) );
  AOI211_X1 U13836 ( .C1(n16313), .C2(n11816), .A(n11815), .B(n11814), .ZN(
        n11817) );
  OAI211_X1 U13837 ( .C1(n15412), .C2(n16285), .A(n11818), .B(n11817), .ZN(
        P1_U3289) );
  INV_X1 U13838 ( .A(n13336), .ZN(n11819) );
  NOR2_X1 U13839 ( .A1(n11819), .A2(n16410), .ZN(n11820) );
  AOI22_X1 U13840 ( .A1(n13309), .A2(n11820), .B1(n16178), .B2(n11308), .ZN(
        n11925) );
  INV_X1 U13841 ( .A(n14227), .ZN(n14189) );
  AOI22_X1 U13842 ( .A1(n14189), .A2(n11883), .B1(n16470), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n11821) );
  OAI21_X1 U13843 ( .B1(n11925), .B2(n16470), .A(n11821), .ZN(P3_U3459) );
  INV_X1 U13844 ( .A(n11955), .ZN(n11967) );
  XNOR2_X1 U13845 ( .A(n11968), .B(n11967), .ZN(n16341) );
  INV_X1 U13846 ( .A(n16341), .ZN(n11841) );
  AND2_X1 U13847 ( .A1(n16314), .A2(n11823), .ZN(n11826) );
  NAND2_X1 U13848 ( .A1(n11824), .A2(n15140), .ZN(n11825) );
  XNOR2_X1 U13849 ( .A(n11956), .B(n11955), .ZN(n11830) );
  NAND2_X1 U13850 ( .A1(n16341), .A2(n16488), .ZN(n11828) );
  OAI211_X1 U13851 ( .C1(n11830), .C2(n16532), .A(n11829), .B(n11828), .ZN(
        n16339) );
  NAND2_X1 U13852 ( .A1(n16339), .A2(n15352), .ZN(n11840) );
  INV_X1 U13853 ( .A(n11831), .ZN(n11832) );
  OAI22_X1 U13854 ( .A1(n15352), .A2(n11277), .B1(n11832), .B2(n16104), .ZN(
        n11837) );
  INV_X1 U13855 ( .A(n11838), .ZN(n16338) );
  INV_X1 U13856 ( .A(n12069), .ZN(n11834) );
  OAI211_X1 U13857 ( .C1(n16338), .C2(n11835), .A(n11834), .B(n15501), .ZN(
        n16337) );
  NOR2_X1 U13858 ( .A1(n16337), .A2(n15372), .ZN(n11836) );
  AOI211_X1 U13859 ( .C1(n16313), .C2(n11838), .A(n11837), .B(n11836), .ZN(
        n11839) );
  OAI211_X1 U13860 ( .C1(n11841), .C2(n13351), .A(n11840), .B(n11839), .ZN(
        P1_U3287) );
  INV_X1 U13861 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11842) );
  OAI22_X1 U13862 ( .A1(n14296), .A2(n11928), .B1(n16447), .B2(n11842), .ZN(
        n11843) );
  INV_X1 U13863 ( .A(n11843), .ZN(n11844) );
  OAI21_X1 U13864 ( .B1(n11925), .B2(n16562), .A(n11844), .ZN(P3_U3390) );
  XOR2_X1 U13865 ( .A(n11846), .B(n11845), .Z(n11850) );
  NOR2_X1 U13866 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13745), .ZN(n15955) );
  OAI22_X1 U13867 ( .A1(n12154), .A2(n13451), .B1(n12119), .B2(n13450), .ZN(
        n11847) );
  AOI211_X1 U13868 ( .C1(n13455), .C2(n12333), .A(n15955), .B(n11847), .ZN(
        n11849) );
  NAND2_X1 U13869 ( .A1(n13454), .A2(n12332), .ZN(n11848) );
  OAI211_X1 U13870 ( .C1(n11850), .C2(n13458), .A(n11849), .B(n11848), .ZN(
        P3_U3167) );
  XNOR2_X1 U13871 ( .A(n11851), .B(n11856), .ZN(n16299) );
  INV_X1 U13872 ( .A(n16264), .ZN(n11852) );
  AOI211_X1 U13873 ( .C1(n11853), .C2(n11852), .A(n14491), .B(n7510), .ZN(
        n16295) );
  OAI22_X1 U13874 ( .A1(n14648), .A2(n16298), .B1(n11854), .B2(n16117), .ZN(
        n11855) );
  AOI21_X1 U13875 ( .B1(n16295), .B2(n16403), .A(n11855), .ZN(n11862) );
  XNOR2_X1 U13876 ( .A(n11857), .B(n11856), .ZN(n11859) );
  AOI21_X1 U13877 ( .B1(n11859), .B2(n16107), .A(n11858), .ZN(n16296) );
  MUX2_X1 U13878 ( .A(n11860), .B(n16296), .S(n14675), .Z(n11861) );
  OAI211_X1 U13879 ( .C1(n14620), .C2(n16299), .A(n11862), .B(n11861), .ZN(
        P2_U3261) );
  INV_X1 U13880 ( .A(n11863), .ZN(n11865) );
  INV_X1 U13881 ( .A(n15637), .ZN(n12818) );
  OAI222_X1 U13882 ( .A1(n14821), .A2(n11864), .B1(n14819), .B2(n11865), .C1(
        n12818), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U13883 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11866) );
  OAI222_X1 U13884 ( .A1(n15558), .A2(n11866), .B1(n15556), .B2(n11865), .C1(
        n15705), .C2(P1_U3086), .ZN(P1_U3340) );
  NAND2_X1 U13885 ( .A1(n12071), .A2(n14950), .ZN(n11871) );
  NAND2_X1 U13886 ( .A1(n15138), .A2(n14900), .ZN(n11870) );
  NAND2_X1 U13887 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  XNOR2_X1 U13888 ( .A(n11872), .B(n14925), .ZN(n12163) );
  AND2_X1 U13889 ( .A1(n14955), .A2(n15138), .ZN(n11873) );
  AOI21_X1 U13890 ( .B1(n12071), .B2(n14900), .A(n11873), .ZN(n12164) );
  XNOR2_X1 U13891 ( .A(n12163), .B(n12164), .ZN(n11874) );
  AOI21_X1 U13892 ( .B1(n11875), .B2(n11874), .A(n15115), .ZN(n11876) );
  NAND2_X1 U13893 ( .A1(n11876), .A2(n12168), .ZN(n11882) );
  NAND2_X1 U13894 ( .A1(n15137), .A2(n15099), .ZN(n11878) );
  NAND2_X1 U13895 ( .A1(n15139), .A2(n15100), .ZN(n11877) );
  AND2_X1 U13896 ( .A1(n11878), .A2(n11877), .ZN(n12076) );
  OAI21_X1 U13897 ( .B1(n15102), .B2(n12076), .A(n11879), .ZN(n11880) );
  AOI21_X1 U13898 ( .B1(n15104), .B2(n12070), .A(n11880), .ZN(n11881) );
  OAI211_X1 U13899 ( .C1(n16351), .C2(n15108), .A(n11882), .B(n11881), .ZN(
        P1_U3213) );
  XOR2_X1 U13900 ( .A(n13142), .B(n13307), .Z(n16135) );
  NAND3_X1 U13901 ( .A1(n13307), .A2(n11883), .A3(n16183), .ZN(n11885) );
  AOI21_X1 U13902 ( .B1(n11885), .B2(n14161), .A(n11884), .ZN(n11887) );
  OAI22_X1 U13903 ( .A1(n16182), .A2(n14156), .B1(n12118), .B2(n14159), .ZN(
        n11886) );
  AOI211_X1 U13904 ( .C1(n16135), .C2(n16475), .A(n11887), .B(n11886), .ZN(
        n16132) );
  OAI21_X1 U13905 ( .B1(n16130), .B2(n16467), .A(n16132), .ZN(n16127) );
  INV_X1 U13906 ( .A(n16127), .ZN(n11889) );
  NAND2_X1 U13907 ( .A1(n16447), .A2(n16382), .ZN(n14303) );
  INV_X1 U13908 ( .A(n14303), .ZN(n16476) );
  AOI22_X1 U13909 ( .A1(n16135), .A2(n16476), .B1(P3_REG0_REG_1__SCAN_IN), 
        .B2(n16562), .ZN(n11888) );
  OAI21_X1 U13910 ( .B1(n11889), .B2(n16562), .A(n11888), .ZN(P3_U3393) );
  INV_X1 U13911 ( .A(n11890), .ZN(n11891) );
  AOI21_X1 U13912 ( .B1(n11895), .B2(n11892), .A(n11891), .ZN(n12064) );
  INV_X1 U13913 ( .A(n12197), .ZN(n11893) );
  AOI211_X1 U13914 ( .C1(n12058), .C2(n12083), .A(n14491), .B(n11893), .ZN(
        n12056) );
  XOR2_X1 U13915 ( .A(n11895), .B(n11894), .Z(n11897) );
  OAI21_X1 U13916 ( .B1(n11897), .B2(n16256), .A(n11896), .ZN(n12061) );
  AOI211_X1 U13917 ( .C1(n12064), .C2(n14751), .A(n12056), .B(n12061), .ZN(
        n11902) );
  INV_X1 U13918 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11898) );
  NOR2_X1 U13919 ( .A1(n16516), .A2(n11898), .ZN(n11899) );
  AOI21_X1 U13920 ( .B1(n12058), .B2(n14792), .A(n11899), .ZN(n11900) );
  OAI21_X1 U13921 ( .B1(n11902), .B2(n16513), .A(n11900), .ZN(P2_U3454) );
  AOI22_X1 U13922 ( .A1(n12058), .A2(n14757), .B1(n16510), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n11901) );
  OAI21_X1 U13923 ( .B1(n11902), .B2(n16510), .A(n11901), .ZN(P2_U3507) );
  MUX2_X1 U13924 ( .A(n11904), .B(n11903), .S(n16408), .Z(n11912) );
  INV_X1 U13925 ( .A(n11905), .ZN(n11910) );
  INV_X1 U13926 ( .A(n11906), .ZN(n11908) );
  OAI22_X1 U13927 ( .A1(n11908), .A2(n14648), .B1(n16117), .B2(n11907), .ZN(
        n11909) );
  AOI21_X1 U13928 ( .B1(n11910), .B2(n16403), .A(n11909), .ZN(n11911) );
  OAI211_X1 U13929 ( .C1(n11913), .C2(n14620), .A(n11912), .B(n11911), .ZN(
        P2_U3259) );
  NAND2_X1 U13930 ( .A1(n13471), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11914) );
  OAI21_X1 U13931 ( .B1(n13974), .B2(n13471), .A(n11914), .ZN(P3_U3520) );
  NAND2_X1 U13932 ( .A1(n14305), .A2(n11915), .ZN(n11919) );
  NAND2_X1 U13933 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  NAND4_X1 U13934 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n11924) );
  INV_X1 U13935 ( .A(n11924), .ZN(n11922) );
  NOR2_X1 U13936 ( .A1(n16467), .A2(n13289), .ZN(n16129) );
  MUX2_X1 U13937 ( .A(n7881), .B(n11925), .S(n14169), .Z(n11927) );
  NAND2_X1 U13938 ( .A1(n14163), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n11926) );
  OAI211_X1 U13939 ( .C1(n11928), .C2(n14166), .A(n11927), .B(n11926), .ZN(
        P3_U3233) );
  INV_X1 U13940 ( .A(n11929), .ZN(n11931) );
  INV_X1 U13941 ( .A(SI_21_), .ZN(n11930) );
  OAI222_X1 U13942 ( .A1(n11932), .A2(P3_U3151), .B1(n14312), .B2(n11931), 
        .C1(n11930), .C2(n14315), .ZN(P3_U3274) );
  INV_X1 U13943 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n11933) );
  NAND2_X1 U13944 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n12385)
         );
  OAI21_X1 U13945 ( .B1(n11934), .B2(n11933), .A(n12385), .ZN(n11949) );
  INV_X1 U13946 ( .A(n11943), .ZN(n11936) );
  OAI21_X1 U13947 ( .B1(n11936), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11935), 
        .ZN(n11939) );
  NAND2_X1 U13948 ( .A1(n11950), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11937) );
  OAI21_X1 U13949 ( .B1(n11950), .B2(P2_REG1_REG_13__SCAN_IN), .A(n11937), 
        .ZN(n11938) );
  AOI21_X1 U13950 ( .B1(n11939), .B2(n11938), .A(n15681), .ZN(n11940) );
  NAND2_X1 U13951 ( .A1(n11940), .A2(n12815), .ZN(n11947) );
  INV_X1 U13952 ( .A(n11941), .ZN(n11942) );
  AOI21_X1 U13953 ( .B1(n11542), .B2(n11943), .A(n11942), .ZN(n11945) );
  INV_X1 U13954 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U13955 ( .A1(n11950), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12834), 
        .B2(n12833), .ZN(n11944) );
  NAND2_X1 U13956 ( .A1(n11945), .A2(n11944), .ZN(n12832) );
  OAI211_X1 U13957 ( .C1(n11945), .C2(n11944), .A(n15661), .B(n12832), .ZN(
        n11946) );
  NAND2_X1 U13958 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  AOI211_X1 U13959 ( .C1(n15678), .C2(n11950), .A(n11949), .B(n11948), .ZN(
        n11951) );
  INV_X1 U13960 ( .A(n11951), .ZN(P2_U3227) );
  INV_X1 U13961 ( .A(n11952), .ZN(n11954) );
  OAI22_X1 U13962 ( .A1(n13338), .A2(P3_U3151), .B1(SI_22_), .B2(n14315), .ZN(
        n11953) );
  AOI21_X1 U13963 ( .B1(n11954), .B2(n12146), .A(n11953), .ZN(P3_U3273) );
  NAND2_X1 U13964 ( .A1(n16338), .A2(n15139), .ZN(n11957) );
  NAND2_X1 U13965 ( .A1(n11958), .A2(n11957), .ZN(n12073) );
  NAND2_X1 U13966 ( .A1(n12073), .A2(n12074), .ZN(n11960) );
  NAND2_X1 U13967 ( .A1(n16351), .A2(n15138), .ZN(n11959) );
  NAND2_X1 U13968 ( .A1(n11960), .A2(n11959), .ZN(n12188) );
  NAND2_X1 U13969 ( .A1(n12188), .A2(n12189), .ZN(n11963) );
  INV_X1 U13970 ( .A(n15137), .ZN(n11961) );
  OR2_X1 U13971 ( .A1(n12186), .A2(n11961), .ZN(n11962) );
  XNOR2_X1 U13972 ( .A(n12267), .B(n12262), .ZN(n11966) );
  AND2_X1 U13973 ( .A1(n15137), .A2(n15100), .ZN(n11964) );
  AOI21_X1 U13974 ( .B1(n15136), .B2(n15099), .A(n11964), .ZN(n12372) );
  INV_X1 U13975 ( .A(n12372), .ZN(n11965) );
  AOI21_X1 U13976 ( .B1(n11966), .B2(n16248), .A(n11965), .ZN(n11977) );
  INV_X1 U13977 ( .A(n15139), .ZN(n11969) );
  NAND2_X1 U13978 ( .A1(n16338), .A2(n11969), .ZN(n11970) );
  INV_X1 U13979 ( .A(n12074), .ZN(n12066) );
  NAND2_X1 U13980 ( .A1(n12067), .A2(n12066), .ZN(n11973) );
  INV_X1 U13981 ( .A(n15138), .ZN(n11971) );
  NAND2_X1 U13982 ( .A1(n16351), .A2(n11971), .ZN(n11972) );
  NAND2_X1 U13983 ( .A1(n11973), .A2(n11972), .ZN(n12181) );
  NAND2_X1 U13984 ( .A1(n12181), .A2(n12182), .ZN(n11975) );
  OR2_X1 U13985 ( .A1(n12186), .A2(n15137), .ZN(n11974) );
  XNOR2_X1 U13986 ( .A(n12263), .B(n12262), .ZN(n16392) );
  NAND2_X1 U13987 ( .A1(n16392), .A2(n16488), .ZN(n11976) );
  AND2_X1 U13988 ( .A1(n11977), .A2(n11976), .ZN(n16394) );
  INV_X1 U13989 ( .A(n13351), .ZN(n16315) );
  INV_X1 U13990 ( .A(n12186), .ZN(n16374) );
  NAND2_X1 U13991 ( .A1(n16388), .A2(n12183), .ZN(n11978) );
  NAND2_X1 U13992 ( .A1(n12273), .A2(n11978), .ZN(n16389) );
  INV_X1 U13993 ( .A(n16104), .ZN(n16312) );
  AOI22_X1 U13994 ( .A1(n16153), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n12369), 
        .B2(n16312), .ZN(n11980) );
  NAND2_X1 U13995 ( .A1(n16388), .A2(n16313), .ZN(n11979) );
  OAI211_X1 U13996 ( .C1(n16389), .C2(n16099), .A(n11980), .B(n11979), .ZN(
        n11981) );
  AOI21_X1 U13997 ( .B1(n16392), .B2(n16315), .A(n11981), .ZN(n11982) );
  OAI21_X1 U13998 ( .B1(n16394), .B2(n16153), .A(n11982), .ZN(P1_U3284) );
  INV_X1 U13999 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n13773) );
  INV_X1 U14000 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n11986) );
  NAND2_X1 U14001 ( .A1(n11983), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11985) );
  NAND2_X1 U14002 ( .A1(n9746), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11984) );
  OAI211_X1 U14003 ( .C1(n11987), .C2(n11986), .A(n11985), .B(n11984), .ZN(
        n11988) );
  INV_X1 U14004 ( .A(n11988), .ZN(n11989) );
  NAND2_X1 U14005 ( .A1(n11990), .A2(n11989), .ZN(n13955) );
  NAND2_X1 U14006 ( .A1(n13955), .A2(P3_U3897), .ZN(n11991) );
  OAI21_X1 U14007 ( .B1(P3_U3897), .B2(n13773), .A(n11991), .ZN(P3_U3522) );
  INV_X1 U14008 ( .A(n12301), .ZN(n12000) );
  AOI21_X1 U14009 ( .B1(n11993), .B2(n11992), .A(n13458), .ZN(n11995) );
  NAND2_X1 U14010 ( .A1(n11995), .A2(n11994), .ZN(n11999) );
  NAND2_X1 U14011 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15979) );
  INV_X1 U14012 ( .A(n15979), .ZN(n11997) );
  OAI22_X1 U14013 ( .A1(n12294), .A2(n13451), .B1(n12293), .B2(n13450), .ZN(
        n11996) );
  AOI211_X1 U14014 ( .C1(n13455), .C2(n16333), .A(n11997), .B(n11996), .ZN(
        n11998) );
  OAI211_X1 U14015 ( .C1(n12000), .C2(n12702), .A(n11999), .B(n11998), .ZN(
        P3_U3179) );
  OAI21_X1 U14016 ( .B1(n12003), .B2(n12002), .A(n12001), .ZN(n12012) );
  INV_X1 U14017 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n13617) );
  INV_X1 U14018 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n16193) );
  OAI22_X1 U14019 ( .A1(n15981), .A2(n13617), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n16193), .ZN(n12011) );
  INV_X1 U14020 ( .A(n12004), .ZN(n12007) );
  INV_X1 U14021 ( .A(n12005), .ZN(n12006) );
  NAND2_X1 U14022 ( .A1(n12007), .A2(n12006), .ZN(n12008) );
  INV_X1 U14023 ( .A(n16079), .ZN(n15969) );
  AOI21_X1 U14024 ( .B1(n12009), .B2(n12008), .A(n15969), .ZN(n12010) );
  AOI211_X1 U14025 ( .C1(n16054), .C2(n12012), .A(n12011), .B(n12010), .ZN(
        n12020) );
  INV_X1 U14026 ( .A(n12013), .ZN(n12015) );
  NOR3_X1 U14027 ( .A1(n12016), .A2(n12015), .A3(n12014), .ZN(n12018) );
  INV_X1 U14028 ( .A(n15913), .ZN(n12017) );
  INV_X1 U14029 ( .A(n16069), .ZN(n16052) );
  OAI21_X1 U14030 ( .B1(n12018), .B2(n12017), .A(n16052), .ZN(n12019) );
  OAI211_X1 U14031 ( .C1(n16076), .C2(n7370), .A(n12020), .B(n12019), .ZN(
        P3_U3184) );
  INV_X1 U14032 ( .A(n12022), .ZN(n12025) );
  INV_X1 U14033 ( .A(n12609), .ZN(n12617) );
  OAI222_X1 U14034 ( .A1(n15558), .A2(n12023), .B1(n15556), .B2(n12025), .C1(
        n12617), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U14035 ( .A1(P2_U3088), .A2(n15644), .B1(n14819), .B2(n12025), 
        .C1(n12024), .C2(n14821), .ZN(P2_U3311) );
  INV_X1 U14036 ( .A(n12214), .ZN(n12029) );
  OAI22_X1 U14037 ( .A1(n12432), .A2(n16108), .B1(n12026), .B2(n14652), .ZN(
        n12211) );
  NAND2_X1 U14038 ( .A1(n14445), .A2(n12211), .ZN(n12028) );
  OAI211_X1 U14039 ( .C1(n14442), .C2(n12029), .A(n12028), .B(n12027), .ZN(
        n12036) );
  INV_X1 U14040 ( .A(n12030), .ZN(n12034) );
  AOI22_X1 U14041 ( .A1(n12031), .A2(n14437), .B1(n14411), .B2(n14465), .ZN(
        n12033) );
  NOR3_X1 U14042 ( .A1(n12034), .A2(n12033), .A3(n12032), .ZN(n12035) );
  AOI211_X1 U14043 ( .C1(n12037), .C2(n14432), .A(n12036), .B(n12035), .ZN(
        n12038) );
  OAI21_X1 U14044 ( .B1(n12039), .B2(n14408), .A(n12038), .ZN(P2_U3189) );
  XNOR2_X1 U14045 ( .A(n12042), .B(n12040), .ZN(n16244) );
  OAI21_X1 U14046 ( .B1(n12043), .B2(n12042), .A(n12041), .ZN(n16247) );
  INV_X1 U14047 ( .A(n12044), .ZN(n12047) );
  AOI21_X1 U14048 ( .B1(n12045), .B2(n14985), .A(n16495), .ZN(n12046) );
  NAND2_X1 U14049 ( .A1(n12047), .A2(n12046), .ZN(n16241) );
  AOI22_X1 U14050 ( .A1(n16313), .A2(n14985), .B1(n14987), .B2(n16312), .ZN(
        n12053) );
  OR2_X1 U14051 ( .A1(n12048), .A2(n15401), .ZN(n12050) );
  NAND2_X1 U14052 ( .A1(n11171), .A2(n15100), .ZN(n12049) );
  NAND2_X1 U14053 ( .A1(n12050), .A2(n12049), .ZN(n14986) );
  INV_X1 U14054 ( .A(n14986), .ZN(n16240) );
  MUX2_X1 U14055 ( .A(n16240), .B(n12051), .S(n16153), .Z(n12052) );
  OAI211_X1 U14056 ( .C1(n16241), .C2(n15372), .A(n12053), .B(n12052), .ZN(
        n12054) );
  AOI21_X1 U14057 ( .B1(n16247), .B2(n15374), .A(n12054), .ZN(n12055) );
  OAI21_X1 U14058 ( .B1(n16244), .B2(n15412), .A(n12055), .ZN(P1_U3290) );
  INV_X1 U14059 ( .A(n12056), .ZN(n12060) );
  AOI22_X1 U14060 ( .A1(n12058), .A2(n16399), .B1(n12057), .B2(n16397), .ZN(
        n12059) );
  OAI21_X1 U14061 ( .B1(n12060), .B2(n16228), .A(n12059), .ZN(n12063) );
  MUX2_X1 U14062 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n12061), .S(n14675), .Z(
        n12062) );
  AOI211_X1 U14063 ( .C1(n14678), .C2(n12064), .A(n12063), .B(n12062), .ZN(
        n12065) );
  INV_X1 U14064 ( .A(n12065), .ZN(P2_U3257) );
  XNOR2_X1 U14065 ( .A(n12067), .B(n12066), .ZN(n16355) );
  INV_X1 U14066 ( .A(n12184), .ZN(n12068) );
  OAI21_X1 U14067 ( .B1(n16351), .B2(n12069), .A(n12068), .ZN(n16352) );
  AOI22_X1 U14068 ( .A1(n12071), .A2(n16313), .B1(n16312), .B2(n12070), .ZN(
        n12072) );
  OAI21_X1 U14069 ( .B1(n16352), .B2(n16099), .A(n12072), .ZN(n12079) );
  XNOR2_X1 U14070 ( .A(n12073), .B(n12074), .ZN(n12077) );
  NAND2_X1 U14071 ( .A1(n16355), .A2(n16488), .ZN(n12075) );
  OAI211_X1 U14072 ( .C1(n12077), .C2(n16532), .A(n12076), .B(n12075), .ZN(
        n16353) );
  MUX2_X1 U14073 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n16353), .S(n15356), .Z(
        n12078) );
  AOI211_X1 U14074 ( .C1(n16355), .C2(n16315), .A(n12079), .B(n12078), .ZN(
        n12080) );
  INV_X1 U14075 ( .A(n12080), .ZN(P1_U3286) );
  AND2_X1 U14076 ( .A1(n14675), .A2(n16122), .ZN(n16401) );
  OAI21_X1 U14077 ( .B1(n12082), .B2(n12088), .A(n12081), .ZN(n16363) );
  OAI211_X1 U14078 ( .C1(n16360), .C2(n12084), .A(n16261), .B(n12083), .ZN(
        n16359) );
  AOI22_X1 U14079 ( .A1(n12086), .A2(n16399), .B1(n12085), .B2(n16397), .ZN(
        n12087) );
  OAI21_X1 U14080 ( .B1(n16359), .B2(n16228), .A(n12087), .ZN(n12096) );
  INV_X1 U14081 ( .A(n16431), .ZN(n16259) );
  NAND2_X1 U14082 ( .A1(n16363), .A2(n16259), .ZN(n12094) );
  INV_X1 U14083 ( .A(n12088), .ZN(n12089) );
  XNOR2_X1 U14084 ( .A(n12090), .B(n12089), .ZN(n12091) );
  NAND2_X1 U14085 ( .A1(n12091), .A2(n16107), .ZN(n12093) );
  AOI22_X1 U14086 ( .A1(n14628), .A2(n14466), .B1(n14468), .B2(n14627), .ZN(
        n12092) );
  NAND3_X1 U14087 ( .A1(n12094), .A2(n12093), .A3(n12092), .ZN(n16361) );
  MUX2_X1 U14088 ( .A(n16361), .B(P2_REG2_REG_7__SCAN_IN), .S(n16408), .Z(
        n12095) );
  AOI211_X1 U14089 ( .C1(n16401), .C2(n16363), .A(n12096), .B(n12095), .ZN(
        n12097) );
  INV_X1 U14090 ( .A(n12097), .ZN(P2_U3258) );
  XNOR2_X1 U14091 ( .A(n12098), .B(n12103), .ZN(n12109) );
  INV_X1 U14092 ( .A(n12109), .ZN(n16326) );
  OAI211_X1 U14093 ( .C1(n7510), .C2(n16323), .A(n16261), .B(n12099), .ZN(
        n16322) );
  AOI22_X1 U14094 ( .A1(n16399), .A2(n12101), .B1(n16397), .B2(n12100), .ZN(
        n12102) );
  OAI21_X1 U14095 ( .B1(n16322), .B2(n16228), .A(n12102), .ZN(n12113) );
  XNOR2_X1 U14096 ( .A(n12104), .B(n12103), .ZN(n12108) );
  NAND2_X1 U14097 ( .A1(n14470), .A2(n14627), .ZN(n12106) );
  NAND2_X1 U14098 ( .A1(n14468), .A2(n14628), .ZN(n12105) );
  NAND2_X1 U14099 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  AOI21_X1 U14100 ( .B1(n12108), .B2(n16107), .A(n12107), .ZN(n12111) );
  OR2_X1 U14101 ( .A1(n12109), .A2(n16431), .ZN(n12110) );
  NAND2_X1 U14102 ( .A1(n12111), .A2(n12110), .ZN(n16324) );
  MUX2_X1 U14103 ( .A(n16324), .B(P2_REG2_REG_5__SCAN_IN), .S(n16408), .Z(
        n12112) );
  AOI211_X1 U14104 ( .C1(n16326), .C2(n16401), .A(n12113), .B(n12112), .ZN(
        n12114) );
  INV_X1 U14105 ( .A(n12114), .ZN(P2_U3260) );
  INV_X1 U14106 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n13780) );
  NAND2_X1 U14107 ( .A1(n13116), .A2(P3_U3897), .ZN(n12115) );
  OAI21_X1 U14108 ( .B1(P3_U3897), .B2(n13780), .A(n12115), .ZN(P3_U3519) );
  OAI21_X1 U14109 ( .B1(n12117), .B2(n13308), .A(n12116), .ZN(n16237) );
  INV_X1 U14110 ( .A(n16237), .ZN(n12127) );
  INV_X1 U14111 ( .A(n16475), .ZN(n16188) );
  OAI22_X1 U14112 ( .A1(n12119), .A2(n14159), .B1(n12118), .B2(n14161), .ZN(
        n12120) );
  INV_X1 U14113 ( .A(n12120), .ZN(n12126) );
  INV_X1 U14114 ( .A(n12121), .ZN(n16185) );
  OAI21_X1 U14115 ( .B1(n16185), .B2(n12122), .A(n13308), .ZN(n12124) );
  NAND3_X1 U14116 ( .A1(n12124), .A2(n16183), .A3(n12123), .ZN(n12125) );
  OAI211_X1 U14117 ( .C1(n12127), .C2(n16188), .A(n12126), .B(n12125), .ZN(
        n16235) );
  INV_X1 U14118 ( .A(n16235), .ZN(n12132) );
  AND2_X1 U14119 ( .A1(n13289), .A2(n10118), .ZN(n16200) );
  NAND2_X1 U14120 ( .A1(n14169), .A2(n16200), .ZN(n14082) );
  INV_X1 U14121 ( .A(n14082), .ZN(n12596) );
  AOI22_X1 U14122 ( .A1(n14097), .A2(n12128), .B1(n14163), .B2(n13734), .ZN(
        n12129) );
  OAI21_X1 U14123 ( .B1(n8506), .B2(n14169), .A(n12129), .ZN(n12130) );
  AOI21_X1 U14124 ( .B1(n16237), .B2(n12596), .A(n12130), .ZN(n12131) );
  OAI21_X1 U14125 ( .B1(n12132), .B2(n14164), .A(n12131), .ZN(P3_U3230) );
  XNOR2_X1 U14126 ( .A(n12134), .B(n12133), .ZN(n12139) );
  NAND2_X1 U14127 ( .A1(n12135), .A2(n13306), .ZN(n12284) );
  OAI21_X1 U14128 ( .B1(n12135), .B2(n13306), .A(n12284), .ZN(n16281) );
  OAI22_X1 U14129 ( .A1(n12293), .A2(n14159), .B1(n12136), .B2(n14161), .ZN(
        n12137) );
  AOI21_X1 U14130 ( .B1(n16281), .B2(n16475), .A(n12137), .ZN(n12138) );
  OAI21_X1 U14131 ( .B1(n14156), .B2(n12139), .A(n12138), .ZN(n16279) );
  INV_X1 U14132 ( .A(n16279), .ZN(n12145) );
  AOI22_X1 U14133 ( .A1(n14097), .A2(n12141), .B1(n14163), .B2(n12140), .ZN(
        n12142) );
  OAI21_X1 U14134 ( .B1(n8511), .B2(n14169), .A(n12142), .ZN(n12143) );
  AOI21_X1 U14135 ( .B1(n16281), .B2(n12596), .A(n12143), .ZN(n12144) );
  OAI21_X1 U14136 ( .B1(n12145), .B2(n14164), .A(n12144), .ZN(P3_U3229) );
  NAND2_X1 U14137 ( .A1(n12147), .A2(n12146), .ZN(n12148) );
  OAI211_X1 U14138 ( .C1(n12149), .C2(n14315), .A(n12148), .B(n13341), .ZN(
        P3_U3272) );
  INV_X1 U14139 ( .A(n12448), .ZN(n12158) );
  OAI211_X1 U14140 ( .C1(n12152), .C2(n12151), .A(n12150), .B(n13437), .ZN(
        n12157) );
  INV_X1 U14141 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n12153) );
  NOR2_X1 U14142 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12153), .ZN(n15995) );
  OAI22_X1 U14143 ( .A1(n12154), .A2(n13450), .B1(n12588), .B2(n13451), .ZN(
        n12155) );
  AOI211_X1 U14144 ( .C1(n13455), .C2(n12449), .A(n15995), .B(n12155), .ZN(
        n12156) );
  OAI211_X1 U14145 ( .C1(n12158), .C2(n12702), .A(n12157), .B(n12156), .ZN(
        P3_U3153) );
  NAND2_X1 U14146 ( .A1(n12186), .A2(n14950), .ZN(n12160) );
  NAND2_X1 U14147 ( .A1(n15137), .A2(n14954), .ZN(n12159) );
  NAND2_X1 U14148 ( .A1(n12160), .A2(n12159), .ZN(n12161) );
  XNOR2_X1 U14149 ( .A(n12161), .B(n15001), .ZN(n12358) );
  AND2_X1 U14150 ( .A1(n14955), .A2(n15137), .ZN(n12162) );
  AOI21_X1 U14151 ( .B1(n12186), .B2(n14900), .A(n12162), .ZN(n12359) );
  XNOR2_X1 U14152 ( .A(n12358), .B(n12359), .ZN(n12170) );
  INV_X1 U14153 ( .A(n12163), .ZN(n12166) );
  INV_X1 U14154 ( .A(n12164), .ZN(n12165) );
  NAND2_X1 U14155 ( .A1(n12166), .A2(n12165), .ZN(n12167) );
  OAI21_X1 U14156 ( .B1(n12170), .B2(n12169), .A(n12362), .ZN(n12171) );
  NAND2_X1 U14157 ( .A1(n12171), .A2(n16546), .ZN(n12177) );
  OR2_X1 U14158 ( .A1(n12365), .A2(n15401), .ZN(n12173) );
  NAND2_X1 U14159 ( .A1(n15138), .A2(n15100), .ZN(n12172) );
  AND2_X1 U14160 ( .A1(n12173), .A2(n12172), .ZN(n12191) );
  OAI22_X1 U14161 ( .A1(n12191), .A2(n15102), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12174), .ZN(n12175) );
  AOI21_X1 U14162 ( .B1(n15104), .B2(n12185), .A(n12175), .ZN(n12176) );
  OAI211_X1 U14163 ( .C1(n16374), .C2(n15108), .A(n12177), .B(n12176), .ZN(
        P1_U3221) );
  INV_X1 U14164 ( .A(n12178), .ZN(n12179) );
  INV_X1 U14165 ( .A(n12970), .ZN(n12977) );
  OAI222_X1 U14166 ( .A1(n15558), .A2(n9656), .B1(n15556), .B2(n12179), .C1(
        P1_U3086), .C2(n12977), .ZN(P1_U3338) );
  OAI222_X1 U14167 ( .A1(n14821), .A2(n12180), .B1(n14819), .B2(n12179), .C1(
        P2_U3088), .C2(n15658), .ZN(P2_U3310) );
  XNOR2_X1 U14168 ( .A(n12181), .B(n12182), .ZN(n16378) );
  OAI21_X1 U14169 ( .B1(n16374), .B2(n12184), .A(n12183), .ZN(n16375) );
  AOI22_X1 U14170 ( .A1(n12186), .A2(n16313), .B1(n12185), .B2(n16312), .ZN(
        n12187) );
  OAI21_X1 U14171 ( .B1(n16375), .B2(n16099), .A(n12187), .ZN(n12194) );
  XNOR2_X1 U14172 ( .A(n12188), .B(n12189), .ZN(n12192) );
  NAND2_X1 U14173 ( .A1(n16378), .A2(n16488), .ZN(n12190) );
  OAI211_X1 U14174 ( .C1(n12192), .C2(n16532), .A(n12191), .B(n12190), .ZN(
        n16376) );
  MUX2_X1 U14175 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n16376), .S(n15356), .Z(
        n12193) );
  AOI211_X1 U14176 ( .C1(n16378), .C2(n16315), .A(n12194), .B(n12193), .ZN(
        n12195) );
  INV_X1 U14177 ( .A(n12195), .ZN(P1_U3285) );
  XOR2_X1 U14178 ( .A(n12196), .B(n12198), .Z(n16402) );
  AOI211_X1 U14179 ( .C1(n16400), .C2(n12197), .A(n14491), .B(n12213), .ZN(
        n16404) );
  XOR2_X1 U14180 ( .A(n12199), .B(n12198), .Z(n12201) );
  OAI21_X1 U14181 ( .B1(n12201), .B2(n16256), .A(n12200), .ZN(n12202) );
  AOI21_X1 U14182 ( .B1(n16259), .B2(n16402), .A(n12202), .ZN(n16407) );
  INV_X1 U14183 ( .A(n16407), .ZN(n12203) );
  AOI211_X1 U14184 ( .C1(n16509), .C2(n16402), .A(n16404), .B(n12203), .ZN(
        n12209) );
  AOI22_X1 U14185 ( .A1(n16400), .A2(n14757), .B1(n16510), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n12204) );
  OAI21_X1 U14186 ( .B1(n12209), .B2(n16510), .A(n12204), .ZN(P2_U3508) );
  INV_X1 U14187 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n12205) );
  OAI22_X1 U14188 ( .A1(n12206), .A2(n14787), .B1(n16516), .B2(n12205), .ZN(
        n12207) );
  INV_X1 U14189 ( .A(n12207), .ZN(n12208) );
  OAI21_X1 U14190 ( .B1(n12209), .B2(n16513), .A(n12208), .ZN(P2_U3457) );
  XNOR2_X1 U14191 ( .A(n12210), .B(n12217), .ZN(n12212) );
  AOI21_X1 U14192 ( .B1(n12212), .B2(n16107), .A(n12211), .ZN(n16433) );
  OAI211_X1 U14193 ( .C1(n12213), .C2(n16434), .A(n12250), .B(n16261), .ZN(
        n16432) );
  INV_X1 U14194 ( .A(n16432), .ZN(n12220) );
  AOI22_X1 U14195 ( .A1(n16408), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12214), 
        .B2(n16397), .ZN(n12215) );
  OAI21_X1 U14196 ( .B1(n16434), .B2(n14648), .A(n12215), .ZN(n12219) );
  XOR2_X1 U14197 ( .A(n12216), .B(n12217), .Z(n16429) );
  NOR2_X1 U14198 ( .A1(n16429), .A2(n14620), .ZN(n12218) );
  AOI211_X1 U14199 ( .C1(n12220), .C2(n16403), .A(n12219), .B(n12218), .ZN(
        n12221) );
  OAI21_X1 U14200 ( .B1(n16408), .B2(n16433), .A(n12221), .ZN(P2_U3255) );
  INV_X1 U14201 ( .A(n12415), .ZN(n12228) );
  OAI211_X1 U14202 ( .C1(n12224), .C2(n12223), .A(n12222), .B(n13437), .ZN(
        n12227) );
  NOR2_X1 U14203 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13737), .ZN(n16014) );
  OAI22_X1 U14204 ( .A1(n12602), .A2(n13451), .B1(n12294), .B2(n13450), .ZN(
        n12225) );
  AOI211_X1 U14205 ( .C1(n13455), .C2(n12416), .A(n16014), .B(n12225), .ZN(
        n12226) );
  OAI211_X1 U14206 ( .C1(n12228), .C2(n12702), .A(n12227), .B(n12226), .ZN(
        P3_U3161) );
  AOI21_X1 U14207 ( .B1(n12991), .B2(n12230), .A(n12229), .ZN(n12242) );
  OAI21_X1 U14208 ( .B1(n12232), .B2(n12231), .A(n12528), .ZN(n12240) );
  OAI21_X1 U14209 ( .B1(n12234), .B2(P3_REG1_REG_11__SCAN_IN), .A(n12233), 
        .ZN(n12236) );
  INV_X1 U14210 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15822) );
  NAND2_X1 U14211 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(P3_U3151), .ZN(n12697)
         );
  OAI21_X1 U14212 ( .B1(n15981), .B2(n15822), .A(n12697), .ZN(n12235) );
  AOI21_X1 U14213 ( .B1(n16079), .B2(n12236), .A(n12235), .ZN(n12237) );
  OAI21_X1 U14214 ( .B1(n12238), .B2(n16076), .A(n12237), .ZN(n12239) );
  AOI21_X1 U14215 ( .B1(n12240), .B2(n16052), .A(n12239), .ZN(n12241) );
  OAI21_X1 U14216 ( .B1(n12242), .B2(n16082), .A(n12241), .ZN(P3_U3193) );
  INV_X1 U14217 ( .A(n12428), .ZN(n12243) );
  AOI21_X1 U14218 ( .B1(n12255), .B2(n12244), .A(n12243), .ZN(n12245) );
  OAI222_X1 U14219 ( .A1(n14652), .A2(n12247), .B1(n16108), .B2(n12246), .C1(
        n16256), .C2(n12245), .ZN(n16460) );
  INV_X1 U14220 ( .A(n16460), .ZN(n12261) );
  OAI22_X1 U14221 ( .A1(n14675), .A2(n12249), .B1(n12248), .B2(n16117), .ZN(
        n12253) );
  INV_X1 U14222 ( .A(n12250), .ZN(n12251) );
  OAI211_X1 U14223 ( .C1(n12251), .C2(n16459), .A(n16261), .B(n12423), .ZN(
        n16458) );
  NOR2_X1 U14224 ( .A1(n16458), .A2(n16228), .ZN(n12252) );
  AOI211_X1 U14225 ( .C1(n16399), .C2(n12254), .A(n12253), .B(n12252), .ZN(
        n12260) );
  NOR2_X1 U14226 ( .A1(n12256), .A2(n12255), .ZN(n16457) );
  INV_X1 U14227 ( .A(n16457), .ZN(n12258) );
  NAND3_X1 U14228 ( .A1(n12258), .A2(n14678), .A3(n12257), .ZN(n12259) );
  OAI211_X1 U14229 ( .C1(n12261), .C2(n16408), .A(n12260), .B(n12259), .ZN(
        P2_U3254) );
  NAND2_X1 U14230 ( .A1(n12263), .A2(n12262), .ZN(n12265) );
  OR2_X1 U14231 ( .A1(n16388), .A2(n12270), .ZN(n12264) );
  NAND2_X1 U14232 ( .A1(n12265), .A2(n12264), .ZN(n12340) );
  XNOR2_X1 U14233 ( .A(n12340), .B(n12268), .ZN(n16419) );
  OAI22_X1 U14234 ( .A1(n15352), .A2(n12266), .B1(n12488), .B2(n16104), .ZN(
        n12272) );
  OAI211_X1 U14235 ( .C1(n12269), .C2(n12268), .A(n16248), .B(n12345), .ZN(
        n16424) );
  NAND2_X1 U14236 ( .A1(n12270), .A2(n15100), .ZN(n12486) );
  AOI21_X1 U14237 ( .B1(n16424), .B2(n12486), .A(n16153), .ZN(n12271) );
  AOI211_X1 U14238 ( .C1(n16313), .C2(n16421), .A(n12272), .B(n12271), .ZN(
        n12279) );
  NAND2_X1 U14239 ( .A1(n15135), .A2(n15099), .ZN(n12485) );
  INV_X1 U14240 ( .A(n12273), .ZN(n12275) );
  INV_X1 U14241 ( .A(n16421), .ZN(n12274) );
  OAI211_X1 U14242 ( .C1(n12275), .C2(n12274), .A(n15501), .B(n12350), .ZN(
        n16422) );
  OAI211_X1 U14243 ( .C1(n16419), .C2(n12276), .A(n12485), .B(n16422), .ZN(
        n12277) );
  INV_X1 U14244 ( .A(n15372), .ZN(n16317) );
  NAND2_X1 U14245 ( .A1(n12277), .A2(n16317), .ZN(n12278) );
  OAI211_X1 U14246 ( .C1(n16419), .C2(n13351), .A(n12279), .B(n12278), .ZN(
        P1_U3283) );
  AND2_X1 U14247 ( .A1(n12281), .A2(n12280), .ZN(n12283) );
  AND2_X1 U14248 ( .A1(n12283), .A2(n12282), .ZN(n12287) );
  NAND2_X1 U14249 ( .A1(n12284), .A2(n13157), .ZN(n12320) );
  NAND2_X1 U14250 ( .A1(n12320), .A2(n13302), .ZN(n12322) );
  NAND2_X1 U14251 ( .A1(n12322), .A2(n13162), .ZN(n12285) );
  OR2_X1 U14252 ( .A1(n12285), .A2(n13164), .ZN(n12286) );
  NAND2_X1 U14253 ( .A1(n12287), .A2(n12286), .ZN(n12292) );
  INV_X1 U14254 ( .A(n12292), .ZN(n16330) );
  INV_X1 U14255 ( .A(n12288), .ZN(n12290) );
  AOI21_X1 U14256 ( .B1(n12325), .B2(n12290), .A(n12289), .ZN(n12299) );
  NAND2_X1 U14257 ( .A1(n12291), .A2(n16183), .ZN(n12298) );
  NAND2_X1 U14258 ( .A1(n12292), .A2(n16475), .ZN(n12297) );
  OAI22_X1 U14259 ( .A1(n12294), .A2(n14159), .B1(n12293), .B2(n14161), .ZN(
        n12295) );
  INV_X1 U14260 ( .A(n12295), .ZN(n12296) );
  OAI211_X1 U14261 ( .C1(n12299), .C2(n12298), .A(n12297), .B(n12296), .ZN(
        n16332) );
  MUX2_X1 U14262 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n16332), .S(n14169), .Z(
        n12300) );
  INV_X1 U14263 ( .A(n12300), .ZN(n12303) );
  AOI22_X1 U14264 ( .A1(n14097), .A2(n16333), .B1(n14163), .B2(n12301), .ZN(
        n12302) );
  OAI211_X1 U14265 ( .C1(n16330), .C2(n14082), .A(n12303), .B(n12302), .ZN(
        P3_U3227) );
  OAI22_X1 U14266 ( .A1(n12305), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n12311), 
        .B2(n12304), .ZN(n12306) );
  NAND2_X1 U14267 ( .A1(n15705), .A2(n12306), .ZN(n12307) );
  INV_X1 U14268 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n16538) );
  NAND2_X1 U14269 ( .A1(n12307), .A2(n15700), .ZN(n12309) );
  XNOR2_X1 U14270 ( .A(n12609), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12308) );
  NOR2_X1 U14271 ( .A1(n12308), .A2(n12309), .ZN(n12608) );
  AOI211_X1 U14272 ( .C1(n12309), .C2(n12308), .A(n12608), .B(n15227), .ZN(
        n12319) );
  AOI21_X1 U14273 ( .B1(n12311), .B2(P1_REG2_REG_14__SCAN_IN), .A(n12310), 
        .ZN(n12312) );
  XNOR2_X1 U14274 ( .A(n12312), .B(n15705), .ZN(n15703) );
  NOR2_X1 U14275 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15703), .ZN(n15702) );
  AOI21_X1 U14276 ( .B1(n12312), .B2(n15705), .A(n15702), .ZN(n12314) );
  INV_X1 U14277 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15396) );
  XNOR2_X1 U14278 ( .A(n12609), .B(n15396), .ZN(n12313) );
  NAND2_X1 U14279 ( .A1(n12314), .A2(n12313), .ZN(n12616) );
  OAI211_X1 U14280 ( .C1(n12314), .C2(n12313), .A(n7362), .B(n12616), .ZN(
        n12317) );
  NAND2_X1 U14281 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n16552)
         );
  INV_X1 U14282 ( .A(n16552), .ZN(n12315) );
  AOI21_X1 U14283 ( .B1(n15696), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12315), 
        .ZN(n12316) );
  OAI211_X1 U14284 ( .C1(n15704), .C2(n12617), .A(n12317), .B(n12316), .ZN(
        n12318) );
  OR2_X1 U14285 ( .A1(n12319), .A2(n12318), .ZN(P1_U3259) );
  OR2_X1 U14286 ( .A1(n12320), .A2(n13302), .ZN(n12321) );
  NAND2_X1 U14287 ( .A1(n12322), .A2(n12321), .ZN(n12327) );
  INV_X1 U14288 ( .A(n12327), .ZN(n16306) );
  NAND2_X1 U14289 ( .A1(n12323), .A2(n13302), .ZN(n12324) );
  NAND2_X1 U14290 ( .A1(n12325), .A2(n12324), .ZN(n12326) );
  NAND2_X1 U14291 ( .A1(n12326), .A2(n16183), .ZN(n12330) );
  NAND2_X1 U14292 ( .A1(n12327), .A2(n16475), .ZN(n12329) );
  AOI22_X1 U14293 ( .A1(n13475), .A2(n16180), .B1(n16178), .B2(n13472), .ZN(
        n12328) );
  NAND3_X1 U14294 ( .A1(n12330), .A2(n12329), .A3(n12328), .ZN(n16307) );
  MUX2_X1 U14295 ( .A(n16307), .B(P3_REG2_REG_5__SCAN_IN), .S(n14164), .Z(
        n12331) );
  INV_X1 U14296 ( .A(n12331), .ZN(n12335) );
  AOI22_X1 U14297 ( .A1(n14097), .A2(n12333), .B1(n14163), .B2(n12332), .ZN(
        n12334) );
  OAI211_X1 U14298 ( .C1(n16306), .C2(n14082), .A(n12335), .B(n12334), .ZN(
        P3_U3228) );
  OAI222_X1 U14299 ( .A1(n15558), .A2(n12336), .B1(n15556), .B2(n12337), .C1(
        n7542), .C2(P1_U3086), .ZN(P1_U3337) );
  OAI222_X1 U14300 ( .A1(n14821), .A2(n12338), .B1(n14819), .B2(n12337), .C1(
        n12841), .C2(P2_U3088), .ZN(P2_U3309) );
  NAND2_X1 U14301 ( .A1(n12340), .A2(n12339), .ZN(n12342) );
  OR2_X1 U14302 ( .A1(n16421), .A2(n15136), .ZN(n12341) );
  XNOR2_X1 U14303 ( .A(n12453), .B(n12452), .ZN(n16453) );
  INV_X1 U14304 ( .A(n16453), .ZN(n12357) );
  OR2_X1 U14305 ( .A1(n16421), .A2(n12343), .ZN(n12344) );
  INV_X1 U14306 ( .A(n12457), .ZN(n12347) );
  AOI21_X1 U14307 ( .B1(n12452), .B2(n12348), .A(n12347), .ZN(n12349) );
  AOI22_X1 U14308 ( .A1(n15136), .A2(n15100), .B1(n15099), .B2(n15134), .ZN(
        n12655) );
  OAI21_X1 U14309 ( .B1(n12349), .B2(n16532), .A(n12655), .ZN(n16451) );
  INV_X1 U14310 ( .A(n16153), .ZN(n15352) );
  AND2_X1 U14311 ( .A1(n12350), .A2(n12642), .ZN(n12351) );
  OR2_X1 U14312 ( .A1(n12351), .A2(n12461), .ZN(n16450) );
  INV_X1 U14313 ( .A(n12352), .ZN(n12657) );
  AOI22_X1 U14314 ( .A1(n16153), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12657), 
        .B2(n16312), .ZN(n12354) );
  NAND2_X1 U14315 ( .A1(n12642), .A2(n16313), .ZN(n12353) );
  OAI211_X1 U14316 ( .C1(n16450), .C2(n16099), .A(n12354), .B(n12353), .ZN(
        n12355) );
  AOI21_X1 U14317 ( .B1(n16451), .B2(n15352), .A(n12355), .ZN(n12356) );
  OAI21_X1 U14318 ( .B1(n15412), .B2(n12357), .A(n12356), .ZN(P1_U3282) );
  INV_X1 U14319 ( .A(n12358), .ZN(n12360) );
  NAND2_X1 U14320 ( .A1(n12360), .A2(n12359), .ZN(n12361) );
  NAND2_X1 U14321 ( .A1(n12362), .A2(n12361), .ZN(n12472) );
  NAND2_X1 U14322 ( .A1(n16388), .A2(n14954), .ZN(n12364) );
  OR2_X1 U14323 ( .A1(n12365), .A2(n15003), .ZN(n12363) );
  NAND2_X1 U14324 ( .A1(n12364), .A2(n12363), .ZN(n12470) );
  XNOR2_X1 U14325 ( .A(n12472), .B(n12470), .ZN(n12469) );
  NAND2_X1 U14326 ( .A1(n16388), .A2(n14950), .ZN(n12367) );
  OR2_X1 U14327 ( .A1(n12365), .A2(n15005), .ZN(n12366) );
  NAND2_X1 U14328 ( .A1(n12367), .A2(n12366), .ZN(n12368) );
  XNOR2_X1 U14329 ( .A(n12368), .B(n14925), .ZN(n12468) );
  XOR2_X1 U14330 ( .A(n12469), .B(n12468), .Z(n12375) );
  NAND2_X1 U14331 ( .A1(n15104), .A2(n12369), .ZN(n12371) );
  OAI211_X1 U14332 ( .C1(n12372), .C2(n15102), .A(n12371), .B(n12370), .ZN(
        n12373) );
  AOI21_X1 U14333 ( .B1(n16388), .B2(n16551), .A(n12373), .ZN(n12374) );
  OAI21_X1 U14334 ( .B1(n12375), .B2(n15115), .A(n12374), .ZN(P1_U3231) );
  NOR2_X1 U14335 ( .A1(n14442), .A2(n14663), .ZN(n12377) );
  AOI22_X1 U14336 ( .A1(n14460), .A2(n14628), .B1(n14627), .B2(n12400), .ZN(
        n12667) );
  OAI22_X1 U14337 ( .A1(n14386), .A2(n12667), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15624), .ZN(n12376) );
  AOI211_X1 U14338 ( .C1(n14666), .C2(n14432), .A(n12377), .B(n12376), .ZN(
        n12383) );
  INV_X1 U14339 ( .A(n12378), .ZN(n12381) );
  OAI22_X1 U14340 ( .A1(n12379), .A2(n14408), .B1(n12431), .B2(n14398), .ZN(
        n12380) );
  NAND3_X1 U14341 ( .A1(n12381), .A2(n12395), .A3(n12380), .ZN(n12382) );
  OAI211_X1 U14342 ( .C1(n12384), .C2(n14427), .A(n12383), .B(n12382), .ZN(
        P2_U3187) );
  INV_X1 U14343 ( .A(n12501), .ZN(n12387) );
  AOI22_X1 U14344 ( .A1(n14424), .A2(n14462), .B1(n14423), .B2(n14461), .ZN(
        n12386) );
  OAI211_X1 U14345 ( .C1(n12387), .C2(n14442), .A(n12386), .B(n12385), .ZN(
        n12393) );
  INV_X1 U14346 ( .A(n12403), .ZN(n12391) );
  AOI22_X1 U14347 ( .A1(n12388), .A2(n14437), .B1(n14411), .B2(n14462), .ZN(
        n12390) );
  NOR3_X1 U14348 ( .A1(n12391), .A2(n12390), .A3(n12389), .ZN(n12392) );
  AOI211_X1 U14349 ( .C1(n12504), .C2(n14432), .A(n12393), .B(n12392), .ZN(
        n12394) );
  OAI21_X1 U14350 ( .B1(n12395), .B2(n14408), .A(n12394), .ZN(P2_U3206) );
  NOR3_X1 U14351 ( .A1(n12396), .A2(n12432), .A3(n14398), .ZN(n12397) );
  AOI21_X1 U14352 ( .B1(n12398), .B2(n14437), .A(n12397), .ZN(n12408) );
  INV_X1 U14353 ( .A(n12399), .ZN(n14674) );
  AOI22_X1 U14354 ( .A1(n14423), .A2(n12400), .B1(n14424), .B2(n14463), .ZN(
        n12402) );
  OAI211_X1 U14355 ( .C1(n14674), .C2(n14442), .A(n12402), .B(n12401), .ZN(
        n12405) );
  NOR2_X1 U14356 ( .A1(n12403), .A2(n14408), .ZN(n12404) );
  AOI211_X1 U14357 ( .C1(n14677), .C2(n14432), .A(n12405), .B(n12404), .ZN(
        n12406) );
  OAI21_X1 U14358 ( .B1(n12408), .B2(n12407), .A(n12406), .ZN(P2_U3196) );
  INV_X1 U14359 ( .A(n13173), .ZN(n13304) );
  OAI21_X1 U14360 ( .B1(n12410), .B2(n13304), .A(n12409), .ZN(n12411) );
  AOI222_X1 U14361 ( .A1(n16183), .A2(n12411), .B1(n13470), .B2(n16180), .C1(
        n13468), .C2(n16178), .ZN(n16367) );
  OAI21_X1 U14362 ( .B1(n12413), .B2(n13173), .A(n12412), .ZN(n16370) );
  OR2_X1 U14363 ( .A1(n16475), .A2(n16200), .ZN(n12414) );
  AOI22_X1 U14364 ( .A1(n14097), .A2(n12416), .B1(n14163), .B2(n12415), .ZN(
        n12417) );
  OAI21_X1 U14365 ( .B1(n12418), .B2(n14169), .A(n12417), .ZN(n12419) );
  AOI21_X1 U14366 ( .B1(n16370), .B2(n14100), .A(n12419), .ZN(n12420) );
  OAI21_X1 U14367 ( .B1(n16367), .B2(n14164), .A(n12420), .ZN(P3_U3225) );
  XNOR2_X1 U14368 ( .A(n12422), .B(n12421), .ZN(n14679) );
  NAND2_X1 U14369 ( .A1(n12423), .A2(n14677), .ZN(n12424) );
  NAND2_X1 U14370 ( .A1(n12424), .A2(n16261), .ZN(n12425) );
  NOR2_X1 U14371 ( .A1(n12503), .A2(n12425), .ZN(n14680) );
  NAND3_X1 U14372 ( .A1(n12428), .A2(n12427), .A3(n12426), .ZN(n12429) );
  AND2_X1 U14373 ( .A1(n12496), .A2(n12429), .ZN(n12430) );
  OAI222_X1 U14374 ( .A1(n14652), .A2(n12432), .B1(n16108), .B2(n12431), .C1(
        n16256), .C2(n12430), .ZN(n14673) );
  AOI211_X1 U14375 ( .C1(n14679), .C2(n14751), .A(n14680), .B(n14673), .ZN(
        n12437) );
  AOI22_X1 U14376 ( .A1(n14677), .A2(n14757), .B1(n16510), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n12433) );
  OAI21_X1 U14377 ( .B1(n12437), .B2(n16510), .A(n12433), .ZN(P2_U3511) );
  INV_X1 U14378 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n12434) );
  NOR2_X1 U14379 ( .A1(n16516), .A2(n12434), .ZN(n12435) );
  AOI21_X1 U14380 ( .B1(n14677), .B2(n14792), .A(n12435), .ZN(n12436) );
  OAI21_X1 U14381 ( .B1(n12437), .B2(n16513), .A(n12436), .ZN(P2_U3466) );
  OR2_X1 U14382 ( .A1(n12440), .A2(n12439), .ZN(n12441) );
  NAND2_X1 U14383 ( .A1(n12438), .A2(n12441), .ZN(n12443) );
  INV_X1 U14384 ( .A(n12443), .ZN(n16346) );
  XNOR2_X1 U14385 ( .A(n12442), .B(n13305), .ZN(n12446) );
  NAND2_X1 U14386 ( .A1(n12443), .A2(n16475), .ZN(n12445) );
  AOI22_X1 U14387 ( .A1(n13469), .A2(n16178), .B1(n16180), .B2(n13472), .ZN(
        n12444) );
  OAI211_X1 U14388 ( .C1(n14156), .C2(n12446), .A(n12445), .B(n12444), .ZN(
        n16347) );
  MUX2_X1 U14389 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n16347), .S(n14169), .Z(
        n12447) );
  INV_X1 U14390 ( .A(n12447), .ZN(n12451) );
  AOI22_X1 U14391 ( .A1(n14097), .A2(n12449), .B1(n14163), .B2(n12448), .ZN(
        n12450) );
  OAI211_X1 U14392 ( .C1(n16346), .C2(n14082), .A(n12451), .B(n12450), .ZN(
        P3_U3226) );
  NAND2_X1 U14393 ( .A1(n12453), .A2(n12452), .ZN(n12455) );
  OR2_X1 U14394 ( .A1(n12642), .A2(n15135), .ZN(n12454) );
  NAND2_X1 U14395 ( .A1(n12455), .A2(n12454), .ZN(n12577) );
  XNOR2_X1 U14396 ( .A(n12577), .B(n12575), .ZN(n16484) );
  NAND2_X1 U14397 ( .A1(n12642), .A2(n12640), .ZN(n12456) );
  OAI211_X1 U14398 ( .C1(n12458), .C2(n12575), .A(n12564), .B(n16248), .ZN(
        n12460) );
  AND2_X1 U14399 ( .A1(n15133), .A2(n15099), .ZN(n12459) );
  AOI21_X1 U14400 ( .B1(n15135), .B2(n15100), .A(n12459), .ZN(n12734) );
  NAND2_X1 U14401 ( .A1(n12460), .A2(n12734), .ZN(n16480) );
  INV_X1 U14402 ( .A(n16482), .ZN(n12465) );
  OAI21_X1 U14403 ( .B1(n12465), .B2(n12461), .A(n15501), .ZN(n12462) );
  AND2_X1 U14404 ( .A1(n12465), .A2(n12461), .ZN(n12676) );
  NOR2_X1 U14405 ( .A1(n12462), .A2(n12676), .ZN(n16481) );
  NAND2_X1 U14406 ( .A1(n16481), .A2(n16317), .ZN(n12464) );
  AOI22_X1 U14407 ( .A1(n16153), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12732), 
        .B2(n16312), .ZN(n12463) );
  OAI211_X1 U14408 ( .C1(n12465), .C2(n16156), .A(n12464), .B(n12463), .ZN(
        n12466) );
  AOI21_X1 U14409 ( .B1(n16480), .B2(n15352), .A(n12466), .ZN(n12467) );
  OAI21_X1 U14410 ( .B1(n15412), .B2(n16484), .A(n12467), .ZN(P1_U3281) );
  NAND2_X1 U14411 ( .A1(n12469), .A2(n12468), .ZN(n12474) );
  INV_X1 U14412 ( .A(n12470), .ZN(n12471) );
  NAND2_X1 U14413 ( .A1(n12472), .A2(n12471), .ZN(n12473) );
  NAND2_X1 U14414 ( .A1(n12474), .A2(n12473), .ZN(n12649) );
  NAND2_X1 U14415 ( .A1(n16421), .A2(n14950), .ZN(n12476) );
  NAND2_X1 U14416 ( .A1(n15136), .A2(n14954), .ZN(n12475) );
  NAND2_X1 U14417 ( .A1(n12476), .A2(n12475), .ZN(n12477) );
  XNOR2_X1 U14418 ( .A(n12477), .B(n15001), .ZN(n12483) );
  INV_X1 U14419 ( .A(n12483), .ZN(n12481) );
  NAND2_X1 U14420 ( .A1(n16421), .A2(n14954), .ZN(n12479) );
  NAND2_X1 U14421 ( .A1(n15136), .A2(n14955), .ZN(n12478) );
  NAND2_X1 U14422 ( .A1(n12479), .A2(n12478), .ZN(n12482) );
  INV_X1 U14423 ( .A(n12482), .ZN(n12480) );
  NAND2_X1 U14424 ( .A1(n12481), .A2(n12480), .ZN(n12650) );
  NAND2_X1 U14425 ( .A1(n12483), .A2(n12482), .ZN(n12648) );
  NAND2_X1 U14426 ( .A1(n12650), .A2(n12648), .ZN(n12484) );
  XNOR2_X1 U14427 ( .A(n12649), .B(n12484), .ZN(n12491) );
  NAND2_X1 U14428 ( .A1(n12486), .A2(n12485), .ZN(n16420) );
  AOI22_X1 U14429 ( .A1(n16548), .A2(n16420), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12487) );
  OAI21_X1 U14430 ( .B1(n16555), .B2(n12488), .A(n12487), .ZN(n12489) );
  AOI21_X1 U14431 ( .B1(n16421), .B2(n16551), .A(n12489), .ZN(n12490) );
  OAI21_X1 U14432 ( .B1(n12491), .B2(n15115), .A(n12490), .ZN(P1_U3217) );
  XNOR2_X1 U14433 ( .A(n12492), .B(n12495), .ZN(n12502) );
  AOI22_X1 U14434 ( .A1(n14461), .A2(n14628), .B1(n14462), .B2(n14627), .ZN(
        n12500) );
  INV_X1 U14435 ( .A(n12493), .ZN(n12498) );
  AND3_X1 U14436 ( .A1(n12496), .A2(n12495), .A3(n12494), .ZN(n12497) );
  OAI21_X1 U14437 ( .B1(n12498), .B2(n12497), .A(n16107), .ZN(n12499) );
  OAI211_X1 U14438 ( .C1(n12502), .C2(n16431), .A(n12500), .B(n12499), .ZN(
        n16506) );
  AOI21_X1 U14439 ( .B1(n12501), .B2(n16397), .A(n16506), .ZN(n12508) );
  INV_X1 U14440 ( .A(n12502), .ZN(n16508) );
  OAI211_X1 U14441 ( .C1(n16505), .C2(n12503), .A(n16261), .B(n12662), .ZN(
        n16503) );
  AOI22_X1 U14442 ( .A1(n12504), .A2(n16399), .B1(P2_REG2_REG_13__SCAN_IN), 
        .B2(n16408), .ZN(n12505) );
  OAI21_X1 U14443 ( .B1(n16503), .B2(n16228), .A(n12505), .ZN(n12506) );
  AOI21_X1 U14444 ( .B1(n16508), .B2(n16401), .A(n12506), .ZN(n12507) );
  OAI21_X1 U14445 ( .B1(n12508), .B2(n16408), .A(n12507), .ZN(P2_U3252) );
  INV_X1 U14446 ( .A(n12509), .ZN(n12510) );
  AOI21_X1 U14447 ( .B1(n12512), .B2(n12511), .A(n12510), .ZN(n12516) );
  AND2_X1 U14448 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n16035) );
  OAI22_X1 U14449 ( .A1(n12588), .A2(n13450), .B1(n12696), .B2(n13451), .ZN(
        n12513) );
  AOI211_X1 U14450 ( .C1(n13455), .C2(n16381), .A(n16035), .B(n12513), .ZN(
        n12515) );
  NAND2_X1 U14451 ( .A1(n13454), .A2(n12593), .ZN(n12514) );
  OAI211_X1 U14452 ( .C1(n12516), .C2(n13458), .A(n12515), .B(n12514), .ZN(
        P3_U3171) );
  AOI21_X1 U14453 ( .B1(n12519), .B2(n12518), .A(n12517), .ZN(n12534) );
  OAI21_X1 U14454 ( .B1(n12522), .B2(n12521), .A(n12520), .ZN(n12526) );
  INV_X1 U14455 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13738) );
  NOR2_X1 U14456 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13738), .ZN(n12777) );
  AOI21_X1 U14457 ( .B1(n16073), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12777), 
        .ZN(n12523) );
  OAI21_X1 U14458 ( .B1(n16076), .B2(n12524), .A(n12523), .ZN(n12525) );
  AOI21_X1 U14459 ( .B1(n12526), .B2(n16079), .A(n12525), .ZN(n12533) );
  AND2_X1 U14460 ( .A1(n12528), .A2(n12527), .ZN(n12531) );
  OAI211_X1 U14461 ( .C1(n12531), .C2(n12530), .A(n16052), .B(n12529), .ZN(
        n12532) );
  OAI211_X1 U14462 ( .C1(n12534), .C2(n16082), .A(n12533), .B(n12532), .ZN(
        P3_U3194) );
  INV_X1 U14463 ( .A(n12535), .ZN(n12536) );
  OAI222_X1 U14464 ( .A1(n12537), .A2(P3_U3151), .B1(n14315), .B2(n13681), 
        .C1(n14312), .C2(n12536), .ZN(P3_U3271) );
  OAI21_X1 U14465 ( .B1(n12540), .B2(n12539), .A(n12538), .ZN(n12555) );
  INV_X1 U14466 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n12541) );
  NOR2_X1 U14467 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12541), .ZN(n12604) );
  AOI21_X1 U14468 ( .B1(n12543), .B2(n12542), .A(n7390), .ZN(n12544) );
  NOR2_X1 U14469 ( .A1(n16082), .A2(n12544), .ZN(n12545) );
  AOI211_X1 U14470 ( .C1(n16073), .C2(P3_ADDR_REG_10__SCAN_IN), .A(n12604), 
        .B(n12545), .ZN(n12546) );
  OAI21_X1 U14471 ( .B1(n12547), .B2(n16076), .A(n12546), .ZN(n12554) );
  INV_X1 U14472 ( .A(n12548), .ZN(n12549) );
  NAND3_X1 U14473 ( .A1(n16028), .A2(n12550), .A3(n12549), .ZN(n12551) );
  AOI21_X1 U14474 ( .B1(n12552), .B2(n12551), .A(n16069), .ZN(n12553) );
  AOI211_X1 U14475 ( .C1(n16079), .C2(n12555), .A(n12554), .B(n12553), .ZN(
        n12556) );
  INV_X1 U14476 ( .A(n12556), .ZN(P3_U3192) );
  INV_X1 U14477 ( .A(n12557), .ZN(n12560) );
  OAI222_X1 U14478 ( .A1(n14821), .A2(n12558), .B1(n14819), .B2(n12560), .C1(
        P2_U3088), .C2(n12843), .ZN(P2_U3308) );
  OAI222_X1 U14479 ( .A1(n15558), .A2(n12561), .B1(n15556), .B2(n12560), .C1(
        n12559), .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U14480 ( .A(n15134), .ZN(n12562) );
  OR2_X1 U14481 ( .A1(n16482), .A2(n12562), .ZN(n12563) );
  NAND2_X1 U14482 ( .A1(n12677), .A2(n15133), .ZN(n12565) );
  NAND2_X1 U14483 ( .A1(n12686), .A2(n12565), .ZN(n12566) );
  NAND2_X1 U14484 ( .A1(n12566), .A2(n12582), .ZN(n12704) );
  OAI21_X1 U14485 ( .B1(n12566), .B2(n12582), .A(n12704), .ZN(n15524) );
  NAND2_X1 U14486 ( .A1(n16523), .A2(n12678), .ZN(n12567) );
  NAND2_X1 U14487 ( .A1(n12567), .A2(n15501), .ZN(n12568) );
  NOR2_X1 U14488 ( .A1(n7487), .A2(n12568), .ZN(n15520) );
  NAND2_X1 U14489 ( .A1(n16523), .A2(n16313), .ZN(n12573) );
  NAND2_X1 U14490 ( .A1(n15131), .A2(n15099), .ZN(n12570) );
  NAND2_X1 U14491 ( .A1(n15133), .A2(n15100), .ZN(n12569) );
  NAND2_X1 U14492 ( .A1(n12570), .A2(n12569), .ZN(n16522) );
  NOR2_X1 U14493 ( .A1(n16104), .A2(n16526), .ZN(n12571) );
  AOI21_X1 U14494 ( .B1(n15352), .B2(n16522), .A(n12571), .ZN(n12572) );
  OAI211_X1 U14495 ( .C1(n15356), .C2(n11618), .A(n12573), .B(n12572), .ZN(
        n12574) );
  AOI21_X1 U14496 ( .B1(n15520), .B2(n16317), .A(n12574), .ZN(n12585) );
  INV_X1 U14497 ( .A(n12575), .ZN(n12576) );
  NAND2_X1 U14498 ( .A1(n12577), .A2(n12576), .ZN(n12579) );
  OR2_X1 U14499 ( .A1(n16482), .A2(n15134), .ZN(n12578) );
  INV_X1 U14500 ( .A(n15133), .ZN(n12580) );
  NAND2_X1 U14501 ( .A1(n12677), .A2(n12580), .ZN(n12581) );
  NAND2_X1 U14502 ( .A1(n12583), .A2(n12582), .ZN(n15521) );
  NAND3_X1 U14503 ( .A1(n12714), .A2(n15521), .A3(n15393), .ZN(n12584) );
  OAI211_X1 U14504 ( .C1(n15524), .C2(n15345), .A(n12585), .B(n12584), .ZN(
        P1_U3279) );
  AND2_X1 U14505 ( .A1(n13180), .A2(n13181), .ZN(n13178) );
  XNOR2_X1 U14506 ( .A(n12586), .B(n13178), .ZN(n16383) );
  NAND2_X1 U14507 ( .A1(n16383), .A2(n16475), .ZN(n12592) );
  INV_X1 U14508 ( .A(n13178), .ZN(n13303) );
  XNOR2_X1 U14509 ( .A(n12587), .B(n13303), .ZN(n12590) );
  OAI22_X1 U14510 ( .A1(n12588), .A2(n14161), .B1(n12696), .B2(n14159), .ZN(
        n12589) );
  AOI21_X1 U14511 ( .B1(n12590), .B2(n16183), .A(n12589), .ZN(n12591) );
  AND2_X1 U14512 ( .A1(n12592), .A2(n12591), .ZN(n16385) );
  AOI22_X1 U14513 ( .A1(n14097), .A2(n16381), .B1(n14163), .B2(n12593), .ZN(
        n12594) );
  OAI21_X1 U14514 ( .B1(n16024), .B2(n14169), .A(n12594), .ZN(n12595) );
  AOI21_X1 U14515 ( .B1(n16383), .B2(n12596), .A(n12595), .ZN(n12597) );
  OAI21_X1 U14516 ( .B1(n16385), .B2(n14164), .A(n12597), .ZN(P3_U3224) );
  INV_X1 U14517 ( .A(n12598), .ZN(n12764) );
  OAI211_X1 U14518 ( .C1(n12601), .C2(n12600), .A(n12599), .B(n13437), .ZN(
        n12606) );
  OAI22_X1 U14519 ( .A1(n12602), .A2(n13450), .B1(n12763), .B2(n13447), .ZN(
        n12603) );
  AOI211_X1 U14520 ( .C1(n13441), .C2(n13466), .A(n12604), .B(n12603), .ZN(
        n12605) );
  OAI211_X1 U14521 ( .C1(n12764), .C2(n12702), .A(n12606), .B(n12605), .ZN(
        P3_U3157) );
  INV_X1 U14522 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n12607) );
  NAND2_X1 U14523 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15045)
         );
  OAI21_X1 U14524 ( .B1(n15728), .B2(n12607), .A(n15045), .ZN(n12613) );
  XNOR2_X1 U14525 ( .A(n12970), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n12610) );
  NOR2_X1 U14526 ( .A1(n12611), .A2(n12610), .ZN(n12969) );
  AOI211_X1 U14527 ( .C1(n12611), .C2(n12610), .A(n12969), .B(n15227), .ZN(
        n12612) );
  AOI211_X1 U14528 ( .C1(n15722), .C2(n12970), .A(n12613), .B(n12612), .ZN(
        n12621) );
  OR2_X1 U14529 ( .A1(n12970), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n12615) );
  NAND2_X1 U14530 ( .A1(n12970), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n12614) );
  AND2_X1 U14531 ( .A1(n12615), .A2(n12614), .ZN(n12619) );
  OAI21_X1 U14532 ( .B1(n12617), .B2(n15396), .A(n12616), .ZN(n12618) );
  NAND2_X1 U14533 ( .A1(n12619), .A2(n12618), .ZN(n12975) );
  OAI211_X1 U14534 ( .C1(n12619), .C2(n12618), .A(n7362), .B(n12975), .ZN(
        n12620) );
  NAND2_X1 U14535 ( .A1(n12621), .A2(n12620), .ZN(P1_U3260) );
  OAI21_X1 U14536 ( .B1(n7490), .B2(n7870), .A(n12622), .ZN(n12855) );
  INV_X1 U14537 ( .A(n12855), .ZN(n12632) );
  AOI211_X1 U14538 ( .C1(n12902), .C2(n12663), .A(n14491), .B(n12748), .ZN(
        n12853) );
  INV_X1 U14539 ( .A(n12902), .ZN(n12623) );
  NOR2_X1 U14540 ( .A1(n12623), .A2(n14648), .ZN(n12626) );
  INV_X1 U14541 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12624) );
  OAI22_X1 U14542 ( .A1(n14675), .A2(n12624), .B1(n12896), .B2(n16117), .ZN(
        n12625) );
  AOI211_X1 U14543 ( .C1(n12853), .C2(n16403), .A(n12626), .B(n12625), .ZN(
        n12631) );
  OAI211_X1 U14544 ( .C1(n12628), .C2(n12627), .A(n12744), .B(n16107), .ZN(
        n12629) );
  AOI22_X1 U14545 ( .A1(n14459), .A2(n14628), .B1(n14627), .B2(n14461), .ZN(
        n12893) );
  NAND2_X1 U14546 ( .A1(n12629), .A2(n12893), .ZN(n12854) );
  NAND2_X1 U14547 ( .A1(n12854), .A2(n14675), .ZN(n12630) );
  OAI211_X1 U14548 ( .C1(n14620), .C2(n12632), .A(n12631), .B(n12630), .ZN(
        P2_U3250) );
  INV_X1 U14549 ( .A(n12633), .ZN(n12636) );
  INV_X1 U14550 ( .A(n12634), .ZN(n12635) );
  OAI222_X1 U14551 ( .A1(n12636), .A2(P3_U3151), .B1(n14315), .B2(n13680), 
        .C1(n14312), .C2(n12635), .ZN(P3_U3270) );
  INV_X1 U14552 ( .A(n12642), .ZN(n16449) );
  NAND2_X1 U14553 ( .A1(n12642), .A2(n14950), .ZN(n12638) );
  NAND2_X1 U14554 ( .A1(n15135), .A2(n14954), .ZN(n12637) );
  NAND2_X1 U14555 ( .A1(n12638), .A2(n12637), .ZN(n12639) );
  XNOR2_X1 U14556 ( .A(n12639), .B(n14925), .ZN(n12643) );
  NOR2_X1 U14557 ( .A1(n12640), .A2(n15003), .ZN(n12641) );
  AOI21_X1 U14558 ( .B1(n12642), .B2(n14900), .A(n12641), .ZN(n12644) );
  NAND2_X1 U14559 ( .A1(n12643), .A2(n12644), .ZN(n12720) );
  INV_X1 U14560 ( .A(n12643), .ZN(n12646) );
  INV_X1 U14561 ( .A(n12644), .ZN(n12645) );
  NAND2_X1 U14562 ( .A1(n12646), .A2(n12645), .ZN(n12647) );
  AND2_X1 U14563 ( .A1(n12720), .A2(n12647), .ZN(n12652) );
  OAI21_X1 U14564 ( .B1(n12652), .B2(n12651), .A(n12721), .ZN(n12653) );
  NAND2_X1 U14565 ( .A1(n12653), .A2(n16546), .ZN(n12659) );
  OAI21_X1 U14566 ( .B1(n12655), .B2(n15102), .A(n12654), .ZN(n12656) );
  AOI21_X1 U14567 ( .B1(n15104), .B2(n12657), .A(n12656), .ZN(n12658) );
  OAI211_X1 U14568 ( .C1(n16449), .C2(n15108), .A(n12659), .B(n12658), .ZN(
        P1_U3236) );
  XNOR2_X1 U14569 ( .A(n12661), .B(n12660), .ZN(n14667) );
  AOI21_X1 U14570 ( .B1(n14666), .B2(n12662), .A(n14491), .ZN(n12664) );
  AND2_X1 U14571 ( .A1(n12664), .A2(n12663), .ZN(n14668) );
  XNOR2_X1 U14572 ( .A(n12666), .B(n12665), .ZN(n12668) );
  OAI21_X1 U14573 ( .B1(n12668), .B2(n16256), .A(n12667), .ZN(n14662) );
  AOI211_X1 U14574 ( .C1(n14751), .C2(n14667), .A(n14668), .B(n14662), .ZN(
        n12673) );
  AOI22_X1 U14575 ( .A1(n14666), .A2(n14757), .B1(n16510), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n12669) );
  OAI21_X1 U14576 ( .B1(n12673), .B2(n16510), .A(n12669), .ZN(P2_U3513) );
  INV_X1 U14577 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n12670) );
  NOR2_X1 U14578 ( .A1(n16516), .A2(n12670), .ZN(n12671) );
  AOI21_X1 U14579 ( .B1(n14666), .B2(n14792), .A(n12671), .ZN(n12672) );
  OAI21_X1 U14580 ( .B1(n12673), .B2(n16513), .A(n12672), .ZN(P2_U3472) );
  XNOR2_X1 U14581 ( .A(n12675), .B(n12674), .ZN(n16500) );
  OR2_X1 U14582 ( .A1(n12677), .A2(n12676), .ZN(n12679) );
  NAND2_X1 U14583 ( .A1(n12679), .A2(n12678), .ZN(n16496) );
  NAND2_X1 U14584 ( .A1(n15132), .A2(n15099), .ZN(n12681) );
  NAND2_X1 U14585 ( .A1(n15134), .A2(n15100), .ZN(n12680) );
  AND2_X1 U14586 ( .A1(n12681), .A2(n12680), .ZN(n16491) );
  NAND2_X1 U14587 ( .A1(n16153), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U14588 ( .A1(n16312), .A2(n12868), .ZN(n12682) );
  OAI211_X1 U14589 ( .C1(n16153), .C2(n16491), .A(n12683), .B(n12682), .ZN(
        n12684) );
  AOI21_X1 U14590 ( .B1(n16493), .B2(n16313), .A(n12684), .ZN(n12685) );
  OAI21_X1 U14591 ( .B1(n16496), .B2(n16099), .A(n12685), .ZN(n12690) );
  OAI21_X1 U14592 ( .B1(n12688), .B2(n12687), .A(n12686), .ZN(n16497) );
  NOR2_X1 U14593 ( .A1(n16497), .A2(n15345), .ZN(n12689) );
  AOI211_X1 U14594 ( .C1(n16500), .C2(n15393), .A(n12690), .B(n12689), .ZN(
        n12691) );
  INV_X1 U14595 ( .A(n12691), .ZN(P1_U3280) );
  INV_X1 U14596 ( .A(n12692), .ZN(n12990) );
  OAI211_X1 U14597 ( .C1(n12695), .C2(n12694), .A(n12693), .B(n13437), .ZN(
        n12701) );
  NOR2_X1 U14598 ( .A1(n12696), .A2(n13450), .ZN(n12699) );
  OAI21_X1 U14599 ( .B1(n12928), .B2(n13451), .A(n12697), .ZN(n12698) );
  AOI211_X1 U14600 ( .C1(n13455), .C2(n12996), .A(n12699), .B(n12698), .ZN(
        n12700) );
  OAI211_X1 U14601 ( .C1(n12990), .C2(n12702), .A(n12701), .B(n12700), .ZN(
        P3_U3176) );
  INV_X1 U14602 ( .A(n15132), .ZN(n12706) );
  OR2_X1 U14603 ( .A1(n16523), .A2(n12706), .ZN(n12703) );
  NAND2_X1 U14604 ( .A1(n12704), .A2(n12703), .ZN(n12705) );
  NAND2_X1 U14605 ( .A1(n12705), .A2(n12715), .ZN(n12955) );
  OAI21_X1 U14606 ( .B1(n12705), .B2(n12715), .A(n12955), .ZN(n16533) );
  OAI22_X1 U14607 ( .A1(n12957), .A2(n15401), .B1(n12706), .B2(n15399), .ZN(
        n16527) );
  INV_X1 U14608 ( .A(n15112), .ZN(n12707) );
  AOI22_X1 U14609 ( .A1(n16527), .A2(n15352), .B1(n12707), .B2(n16312), .ZN(
        n12708) );
  OAI21_X1 U14610 ( .B1(n12709), .B2(n15352), .A(n12708), .ZN(n12712) );
  INV_X1 U14611 ( .A(n16529), .ZN(n12710) );
  OAI211_X1 U14612 ( .C1(n12710), .C2(n7487), .A(n15501), .B(n15406), .ZN(
        n16530) );
  NOR2_X1 U14613 ( .A1(n16530), .A2(n15372), .ZN(n12711) );
  AOI211_X1 U14614 ( .C1(n16313), .C2(n16529), .A(n12712), .B(n12711), .ZN(
        n12719) );
  NAND2_X1 U14615 ( .A1(n16523), .A2(n15132), .ZN(n12713) );
  OAI21_X1 U14616 ( .B1(n12717), .B2(n12716), .A(n12952), .ZN(n16535) );
  NAND2_X1 U14617 ( .A1(n16535), .A2(n15393), .ZN(n12718) );
  OAI211_X1 U14618 ( .C1(n16533), .C2(n15345), .A(n12719), .B(n12718), .ZN(
        P1_U3278) );
  NAND2_X1 U14619 ( .A1(n16482), .A2(n14950), .ZN(n12723) );
  NAND2_X1 U14620 ( .A1(n15134), .A2(n14954), .ZN(n12722) );
  NAND2_X1 U14621 ( .A1(n12723), .A2(n12722), .ZN(n12724) );
  XNOR2_X1 U14622 ( .A(n12724), .B(n15001), .ZN(n12727) );
  NAND2_X1 U14623 ( .A1(n16482), .A2(n14954), .ZN(n12726) );
  NAND2_X1 U14624 ( .A1(n14955), .A2(n15134), .ZN(n12725) );
  NAND2_X1 U14625 ( .A1(n12726), .A2(n12725), .ZN(n12728) );
  NAND2_X1 U14626 ( .A1(n12727), .A2(n12728), .ZN(n12859) );
  INV_X1 U14627 ( .A(n12727), .ZN(n12730) );
  INV_X1 U14628 ( .A(n12728), .ZN(n12729) );
  NAND2_X1 U14629 ( .A1(n12730), .A2(n12729), .ZN(n12861) );
  NAND2_X1 U14630 ( .A1(n12859), .A2(n12861), .ZN(n12731) );
  XNOR2_X1 U14631 ( .A(n12860), .B(n12731), .ZN(n12737) );
  NAND2_X1 U14632 ( .A1(n15104), .A2(n12732), .ZN(n12733) );
  NAND2_X1 U14633 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n15726)
         );
  OAI211_X1 U14634 ( .C1(n12734), .C2(n15102), .A(n12733), .B(n15726), .ZN(
        n12735) );
  AOI21_X1 U14635 ( .B1(n16482), .B2(n16551), .A(n12735), .ZN(n12736) );
  OAI21_X1 U14636 ( .B1(n12737), .B2(n15115), .A(n12736), .ZN(P1_U3224) );
  INV_X1 U14637 ( .A(n12738), .ZN(n12769) );
  OAI222_X1 U14638 ( .A1(n14821), .A2(n12740), .B1(P2_U3088), .B2(n12739), 
        .C1(n12769), .C2(n14819), .ZN(P2_U3307) );
  XOR2_X1 U14639 ( .A(n12742), .B(n12741), .Z(n12889) );
  INV_X1 U14640 ( .A(n12889), .ZN(n12754) );
  NAND3_X1 U14641 ( .A1(n7934), .A2(n12744), .A3(n12743), .ZN(n12745) );
  NAND3_X1 U14642 ( .A1(n12943), .A2(n12745), .A3(n16107), .ZN(n12747) );
  AND2_X1 U14643 ( .A1(n14460), .A2(n14627), .ZN(n12746) );
  AOI21_X1 U14644 ( .B1(n14458), .B2(n14628), .A(n12746), .ZN(n12792) );
  NAND2_X1 U14645 ( .A1(n12747), .A2(n12792), .ZN(n12887) );
  OAI211_X1 U14646 ( .C1(n12886), .C2(n12748), .A(n16261), .B(n12936), .ZN(
        n12885) );
  INV_X1 U14647 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12749) );
  OAI22_X1 U14648 ( .A1(n14675), .A2(n12749), .B1(n12790), .B2(n16117), .ZN(
        n12750) );
  AOI21_X1 U14649 ( .B1(n12795), .B2(n16399), .A(n12750), .ZN(n12751) );
  OAI21_X1 U14650 ( .B1(n12885), .B2(n16228), .A(n12751), .ZN(n12752) );
  AOI21_X1 U14651 ( .B1(n12887), .B2(n14675), .A(n12752), .ZN(n12753) );
  OAI21_X1 U14652 ( .B1(n12754), .B2(n14620), .A(n12753), .ZN(P2_U3249) );
  INV_X1 U14653 ( .A(n12755), .ZN(n12756) );
  AOI21_X1 U14654 ( .B1(n12759), .B2(n12757), .A(n12756), .ZN(n16414) );
  OAI211_X1 U14655 ( .C1(n12760), .C2(n12759), .A(n12758), .B(n16183), .ZN(
        n12762) );
  NAND2_X1 U14656 ( .A1(n13468), .A2(n16180), .ZN(n12761) );
  OAI211_X1 U14657 ( .C1(n12780), .C2(n14159), .A(n12762), .B(n12761), .ZN(
        n16409) );
  NOR2_X1 U14658 ( .A1(n14166), .A2(n12763), .ZN(n12767) );
  OAI22_X1 U14659 ( .A1(n14169), .A2(n12765), .B1(n12764), .B2(n16194), .ZN(
        n12766) );
  AOI211_X1 U14660 ( .C1(n16409), .C2(n14169), .A(n12767), .B(n12766), .ZN(
        n12768) );
  OAI21_X1 U14661 ( .B1(n16414), .B2(n14171), .A(n12768), .ZN(P3_U3223) );
  OAI222_X1 U14662 ( .A1(n15558), .A2(n12771), .B1(P1_U3086), .B2(n12770), 
        .C1(n15556), .C2(n12769), .ZN(P1_U3335) );
  INV_X1 U14663 ( .A(n12772), .ZN(n12774) );
  NOR2_X1 U14664 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  XNOR2_X1 U14665 ( .A(n12776), .B(n12775), .ZN(n12784) );
  NAND2_X1 U14666 ( .A1(n13454), .A2(n12920), .ZN(n12779) );
  AOI21_X1 U14667 ( .B1(n13441), .B2(n13026), .A(n12777), .ZN(n12778) );
  OAI211_X1 U14668 ( .C1(n12780), .C2(n13450), .A(n12779), .B(n12778), .ZN(
        n12781) );
  AOI21_X1 U14669 ( .B1(n12782), .B2(n13455), .A(n12781), .ZN(n12783) );
  OAI21_X1 U14670 ( .B1(n12784), .B2(n13458), .A(n12783), .ZN(P3_U3164) );
  INV_X1 U14671 ( .A(n12785), .ZN(n12897) );
  NOR3_X1 U14672 ( .A1(n12787), .A2(n12786), .A3(n14398), .ZN(n12788) );
  AOI21_X1 U14673 ( .B1(n12897), .B2(n14437), .A(n12788), .ZN(n12799) );
  INV_X1 U14674 ( .A(n12789), .ZN(n12910) );
  NAND2_X1 U14675 ( .A1(n12910), .A2(n14437), .ZN(n12797) );
  NOR2_X1 U14676 ( .A1(n14442), .A2(n12790), .ZN(n12794) );
  OAI22_X1 U14677 ( .A1(n14386), .A2(n12792), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12791), .ZN(n12793) );
  AOI211_X1 U14678 ( .C1(n12795), .C2(n14432), .A(n12794), .B(n12793), .ZN(
        n12796) );
  OAI211_X1 U14679 ( .C1(n12799), .C2(n12798), .A(n12797), .B(n12796), .ZN(
        P2_U3198) );
  AOI21_X1 U14680 ( .B1(n12802), .B2(n12801), .A(n12800), .ZN(n12814) );
  OAI21_X1 U14681 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12804), .A(n12803), 
        .ZN(n12812) );
  INV_X1 U14682 ( .A(n13905), .ZN(n12805) );
  AOI21_X1 U14683 ( .B1(n12807), .B2(n12806), .A(n12805), .ZN(n12810) );
  NOR2_X1 U14684 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13555), .ZN(n12926) );
  INV_X1 U14685 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15836) );
  NOR2_X1 U14686 ( .A1(n15981), .A2(n15836), .ZN(n12808) );
  AOI211_X1 U14687 ( .C1(n16043), .C2(n7734), .A(n12926), .B(n12808), .ZN(
        n12809) );
  OAI21_X1 U14688 ( .B1(n12810), .B2(n16069), .A(n12809), .ZN(n12811) );
  AOI21_X1 U14689 ( .B1(n16079), .B2(n12812), .A(n12811), .ZN(n12813) );
  OAI21_X1 U14690 ( .B1(n12814), .B2(n16082), .A(n12813), .ZN(P3_U3195) );
  NAND2_X1 U14691 ( .A1(n12829), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n12821) );
  XNOR2_X1 U14692 ( .A(n15644), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15651) );
  INV_X1 U14693 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12817) );
  INV_X1 U14694 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n16511) );
  OAI21_X1 U14695 ( .B1(n16511), .B2(n12833), .A(n12815), .ZN(n15631) );
  INV_X1 U14696 ( .A(n15625), .ZN(n12830) );
  NOR2_X1 U14697 ( .A1(n12830), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n12816) );
  AOI21_X1 U14698 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n12830), .A(n12816), 
        .ZN(n15630) );
  NAND2_X1 U14699 ( .A1(n15631), .A2(n15630), .ZN(n15629) );
  OAI21_X1 U14700 ( .B1(n12817), .B2(n15625), .A(n15629), .ZN(n12819) );
  NAND2_X1 U14701 ( .A1(n15637), .A2(n12819), .ZN(n12820) );
  XNOR2_X1 U14702 ( .A(n12819), .B(n12818), .ZN(n15639) );
  NAND2_X1 U14703 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15639), .ZN(n15638) );
  NAND2_X1 U14704 ( .A1(n12820), .A2(n15638), .ZN(n15652) );
  NAND2_X1 U14705 ( .A1(n15651), .A2(n15652), .ZN(n15650) );
  NAND2_X1 U14706 ( .A1(n12821), .A2(n15650), .ZN(n15665) );
  XNOR2_X1 U14707 ( .A(n15658), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15666) );
  NAND2_X1 U14708 ( .A1(n15665), .A2(n15666), .ZN(n12824) );
  INV_X1 U14709 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n12822) );
  OR2_X1 U14710 ( .A1(n15658), .A2(n12822), .ZN(n12823) );
  NAND2_X1 U14711 ( .A1(n12824), .A2(n12823), .ZN(n12825) );
  INV_X1 U14712 ( .A(n12841), .ZN(n15677) );
  XNOR2_X1 U14713 ( .A(n12825), .B(n15677), .ZN(n15676) );
  INV_X1 U14714 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15675) );
  INV_X1 U14715 ( .A(n12825), .ZN(n12826) );
  OAI22_X1 U14716 ( .A1(n15676), .A2(n15675), .B1(n12826), .B2(n12841), .ZN(
        n12828) );
  XNOR2_X1 U14717 ( .A(n12843), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12827) );
  XNOR2_X1 U14718 ( .A(n12828), .B(n12827), .ZN(n12852) );
  NAND2_X1 U14719 ( .A1(n12829), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U14720 ( .A1(n12829), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12749), 
        .B2(n15644), .ZN(n15649) );
  NOR2_X1 U14721 ( .A1(n12830), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12835) );
  INV_X1 U14722 ( .A(n12835), .ZN(n12831) );
  OAI21_X1 U14723 ( .B1(n14664), .B2(n15625), .A(n12831), .ZN(n15623) );
  OAI21_X1 U14724 ( .B1(n12834), .B2(n12833), .A(n12832), .ZN(n15622) );
  NOR2_X1 U14725 ( .A1(n15623), .A2(n15622), .ZN(n15621) );
  NOR2_X1 U14726 ( .A1(n12835), .A2(n15621), .ZN(n12836) );
  NAND2_X1 U14727 ( .A1(n15637), .A2(n12836), .ZN(n12837) );
  XOR2_X1 U14728 ( .A(n15637), .B(n12836), .Z(n15636) );
  NAND2_X1 U14729 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15636), .ZN(n15635) );
  NAND2_X1 U14730 ( .A1(n12837), .A2(n15635), .ZN(n15648) );
  NAND2_X1 U14731 ( .A1(n15649), .A2(n15648), .ZN(n15647) );
  NAND2_X1 U14732 ( .A1(n12838), .A2(n15647), .ZN(n15662) );
  INV_X1 U14733 ( .A(n15662), .ZN(n12839) );
  NAND2_X1 U14734 ( .A1(n15659), .A2(n12839), .ZN(n12840) );
  INV_X1 U14735 ( .A(n15658), .ZN(n15664) );
  AOI22_X1 U14736 ( .A1(n12840), .A2(n15664), .B1(n15662), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n12842) );
  XNOR2_X1 U14737 ( .A(n12842), .B(n12841), .ZN(n15674) );
  NOR2_X1 U14738 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n15674), .ZN(n15673) );
  AOI21_X1 U14739 ( .B1(n12842), .B2(n12841), .A(n15673), .ZN(n12845) );
  MUX2_X1 U14740 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n10283), .S(n12843), .Z(
        n12844) );
  XNOR2_X1 U14741 ( .A(n12845), .B(n12844), .ZN(n12846) );
  NAND2_X1 U14742 ( .A1(n12846), .A2(n15661), .ZN(n12851) );
  NAND2_X1 U14743 ( .A1(n15684), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n12847) );
  NAND2_X1 U14744 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n14357)
         );
  NAND2_X1 U14745 ( .A1(n12847), .A2(n14357), .ZN(n12848) );
  AOI21_X1 U14746 ( .B1(n12849), .B2(n15678), .A(n12848), .ZN(n12850) );
  OAI211_X1 U14747 ( .C1(n12852), .C2(n15681), .A(n12851), .B(n12850), .ZN(
        P2_U3233) );
  AOI211_X1 U14748 ( .C1(n14751), .C2(n12855), .A(n12854), .B(n12853), .ZN(
        n12858) );
  AOI22_X1 U14749 ( .A1(n12902), .A2(n14792), .B1(P2_REG0_REG_15__SCAN_IN), 
        .B2(n16513), .ZN(n12856) );
  OAI21_X1 U14750 ( .B1(n12858), .B2(n16513), .A(n12856), .ZN(P2_U3475) );
  AOI22_X1 U14751 ( .A1(n12902), .A2(n14757), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n16510), .ZN(n12857) );
  OAI21_X1 U14752 ( .B1(n12858), .B2(n16510), .A(n12857), .ZN(P2_U3514) );
  NAND2_X1 U14753 ( .A1(n12860), .A2(n12859), .ZN(n12862) );
  NAND2_X1 U14754 ( .A1(n16493), .A2(n14950), .ZN(n12864) );
  NAND2_X1 U14755 ( .A1(n15133), .A2(n14954), .ZN(n12863) );
  NAND2_X1 U14756 ( .A1(n12864), .A2(n12863), .ZN(n12865) );
  XNOR2_X1 U14757 ( .A(n12865), .B(n14925), .ZN(n14837) );
  AND2_X1 U14758 ( .A1(n14955), .A2(n15133), .ZN(n12866) );
  AOI21_X1 U14759 ( .B1(n16493), .B2(n14900), .A(n12866), .ZN(n14838) );
  XNOR2_X1 U14760 ( .A(n14837), .B(n14838), .ZN(n12867) );
  XNOR2_X1 U14761 ( .A(n14836), .B(n12867), .ZN(n12873) );
  NAND2_X1 U14762 ( .A1(n15104), .A2(n12868), .ZN(n12870) );
  OAI211_X1 U14763 ( .C1(n16491), .C2(n15102), .A(n12870), .B(n12869), .ZN(
        n12871) );
  AOI21_X1 U14764 ( .B1(n16493), .B2(n16551), .A(n12871), .ZN(n12872) );
  OAI21_X1 U14765 ( .B1(n12873), .B2(n15115), .A(n12872), .ZN(P1_U3234) );
  INV_X1 U14766 ( .A(n12874), .ZN(n12878) );
  OAI222_X1 U14767 ( .A1(n15558), .A2(n12876), .B1(n15556), .B2(n12878), .C1(
        n12875), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U14768 ( .A1(n14821), .A2(n12879), .B1(n14819), .B2(n12878), .C1(
        P2_U3088), .C2(n12877), .ZN(P2_U3306) );
  INV_X1 U14769 ( .A(n12880), .ZN(n12884) );
  INV_X1 U14770 ( .A(n12881), .ZN(n12882) );
  OAI222_X1 U14771 ( .A1(n12884), .A2(P3_U3151), .B1(n14315), .B2(n13677), 
        .C1(n14312), .C2(n12882), .ZN(P3_U3269) );
  INV_X1 U14772 ( .A(n16265), .ZN(n16504) );
  OAI21_X1 U14773 ( .B1(n12886), .B2(n16504), .A(n12885), .ZN(n12888) );
  AOI211_X1 U14774 ( .C1(n12889), .C2(n14751), .A(n12888), .B(n12887), .ZN(
        n12892) );
  NAND2_X1 U14775 ( .A1(n16510), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n12890) );
  OAI21_X1 U14776 ( .B1(n12892), .B2(n16510), .A(n12890), .ZN(P2_U3515) );
  NAND2_X1 U14777 ( .A1(n16513), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n12891) );
  OAI21_X1 U14778 ( .B1(n12892), .B2(n16513), .A(n12891), .ZN(P2_U3478) );
  INV_X1 U14779 ( .A(n12893), .ZN(n12894) );
  AOI22_X1 U14780 ( .A1(n14445), .A2(n12894), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12895) );
  OAI21_X1 U14781 ( .B1(n12896), .B2(n14442), .A(n12895), .ZN(n12901) );
  AOI211_X1 U14782 ( .C1(n12899), .C2(n12898), .A(n14427), .B(n12897), .ZN(
        n12900) );
  AOI211_X1 U14783 ( .C1(n12902), .C2(n14432), .A(n12901), .B(n12900), .ZN(
        n12903) );
  INV_X1 U14784 ( .A(n12903), .ZN(P2_U3213) );
  AND2_X1 U14785 ( .A1(n14459), .A2(n14627), .ZN(n12904) );
  AOI21_X1 U14786 ( .B1(n14626), .B2(n14628), .A(n12904), .ZN(n12946) );
  INV_X1 U14787 ( .A(n12946), .ZN(n12905) );
  AOI22_X1 U14788 ( .A1(n14445), .A2(n12905), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12906) );
  OAI21_X1 U14789 ( .B1(n12938), .B2(n14442), .A(n12906), .ZN(n12912) );
  AOI22_X1 U14790 ( .A1(n12907), .A2(n14437), .B1(n14411), .B2(n14459), .ZN(
        n12908) );
  NOR3_X1 U14791 ( .A1(n12910), .A2(n12909), .A3(n12908), .ZN(n12911) );
  AOI211_X1 U14792 ( .C1(n14791), .C2(n14432), .A(n12912), .B(n12911), .ZN(
        n12913) );
  OAI21_X1 U14793 ( .B1(n12914), .B2(n14427), .A(n12913), .ZN(P2_U3200) );
  XNOR2_X1 U14794 ( .A(n12915), .B(n12918), .ZN(n12916) );
  AOI222_X1 U14795 ( .A1(n16183), .A2(n12916), .B1(n13026), .B2(n16178), .C1(
        n13466), .C2(n16180), .ZN(n16466) );
  OAI21_X1 U14796 ( .B1(n12919), .B2(n12918), .A(n12917), .ZN(n16477) );
  AOI22_X1 U14797 ( .A1(n14164), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n14163), 
        .B2(n12920), .ZN(n12921) );
  OAI21_X1 U14798 ( .B1(n16468), .B2(n14166), .A(n12921), .ZN(n12922) );
  AOI21_X1 U14799 ( .B1(n16477), .B2(n14100), .A(n12922), .ZN(n12923) );
  OAI21_X1 U14800 ( .B1(n16466), .B2(n14164), .A(n12923), .ZN(P3_U3221) );
  XNOR2_X1 U14801 ( .A(n12925), .B(n12924), .ZN(n12932) );
  AOI21_X1 U14802 ( .B1(n13465), .B2(n13441), .A(n12926), .ZN(n12927) );
  OAI21_X1 U14803 ( .B1(n12928), .B2(n13450), .A(n12927), .ZN(n12930) );
  NOR2_X1 U14804 ( .A1(n14238), .A2(n13447), .ZN(n12929) );
  AOI211_X1 U14805 ( .C1(n13020), .C2(n13454), .A(n12930), .B(n12929), .ZN(
        n12931) );
  OAI21_X1 U14806 ( .B1(n12932), .B2(n13458), .A(n12931), .ZN(P3_U3174) );
  XNOR2_X1 U14807 ( .A(n12934), .B(n12933), .ZN(n14752) );
  NAND2_X1 U14808 ( .A1(n12936), .A2(n14791), .ZN(n12937) );
  NAND3_X1 U14809 ( .A1(n14644), .A2(n16261), .A3(n12937), .ZN(n14753) );
  OAI22_X1 U14810 ( .A1(n14675), .A2(n15659), .B1(n12938), .B2(n16117), .ZN(
        n12939) );
  AOI21_X1 U14811 ( .B1(n14791), .B2(n16399), .A(n12939), .ZN(n12940) );
  OAI21_X1 U14812 ( .B1(n14753), .B2(n16228), .A(n12940), .ZN(n12949) );
  NAND3_X1 U14813 ( .A1(n12943), .A2(n12942), .A3(n12941), .ZN(n12944) );
  NAND3_X1 U14814 ( .A1(n12945), .A2(n16107), .A3(n12944), .ZN(n12947) );
  AND2_X1 U14815 ( .A1(n12947), .A2(n12946), .ZN(n14754) );
  NOR2_X1 U14816 ( .A1(n14754), .A2(n16408), .ZN(n12948) );
  AOI211_X1 U14817 ( .C1(n14678), .C2(n14752), .A(n12949), .B(n12948), .ZN(
        n12950) );
  INV_X1 U14818 ( .A(n12950), .ZN(P2_U3248) );
  OR2_X1 U14819 ( .A1(n16529), .A2(n15131), .ZN(n12951) );
  OAI21_X1 U14820 ( .B1(n12959), .B2(n12953), .A(n13045), .ZN(n15515) );
  INV_X1 U14821 ( .A(n15131), .ZN(n15400) );
  OR2_X1 U14822 ( .A1(n16529), .A2(n15400), .ZN(n12954) );
  NAND2_X1 U14823 ( .A1(n16550), .A2(n12957), .ZN(n12958) );
  NAND2_X1 U14824 ( .A1(n12960), .A2(n12959), .ZN(n15506) );
  NAND3_X1 U14825 ( .A1(n15507), .A2(n15506), .A3(n15374), .ZN(n12967) );
  NAND2_X1 U14826 ( .A1(n15508), .A2(n15404), .ZN(n12961) );
  AND2_X1 U14827 ( .A1(n15384), .A2(n12961), .ZN(n15512) );
  AND2_X1 U14828 ( .A1(n15130), .A2(n15100), .ZN(n12962) );
  AOI21_X1 U14829 ( .B1(n15128), .B2(n15099), .A(n12962), .ZN(n15509) );
  OAI21_X1 U14830 ( .B1(n15044), .B2(n16104), .A(n15509), .ZN(n12963) );
  MUX2_X1 U14831 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n12963), .S(n15352), .Z(
        n12965) );
  INV_X1 U14832 ( .A(n15508), .ZN(n15050) );
  NOR2_X1 U14833 ( .A1(n15050), .A2(n16156), .ZN(n12964) );
  AOI211_X1 U14834 ( .C1(n15512), .C2(n15387), .A(n12965), .B(n12964), .ZN(
        n12966) );
  OAI211_X1 U14835 ( .C1(n15515), .C2(n15412), .A(n12967), .B(n12966), .ZN(
        P1_U3276) );
  INV_X1 U14836 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n12968) );
  NAND2_X1 U14837 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15091)
         );
  OAI21_X1 U14838 ( .B1(n15728), .B2(n12968), .A(n15091), .ZN(n12974) );
  NOR2_X1 U14839 ( .A1(n12971), .A2(n12972), .ZN(n15219) );
  AOI211_X1 U14840 ( .C1(n12972), .C2(n12971), .A(n15219), .B(n15227), .ZN(
        n12973) );
  AOI211_X1 U14841 ( .C1(n15722), .C2(n15222), .A(n12974), .B(n12973), .ZN(
        n12980) );
  INV_X1 U14842 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12976) );
  OAI21_X1 U14843 ( .B1(n12977), .B2(n12976), .A(n12975), .ZN(n15221) );
  XNOR2_X1 U14844 ( .A(n7542), .B(n15221), .ZN(n12978) );
  NAND2_X1 U14845 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n12978), .ZN(n15223) );
  OAI211_X1 U14846 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n12978), .A(n7362), .B(
        n15223), .ZN(n12979) );
  NAND2_X1 U14847 ( .A1(n12980), .A2(n12979), .ZN(P1_U3261) );
  INV_X1 U14848 ( .A(n12981), .ZN(n12982) );
  OAI222_X1 U14849 ( .A1(P3_U3151), .A2(n12984), .B1(n14315), .B2(n12983), 
        .C1(n14312), .C2(n12982), .ZN(P3_U3268) );
  INV_X1 U14850 ( .A(n12985), .ZN(n12986) );
  OAI222_X1 U14851 ( .A1(n14821), .A2(n12988), .B1(P2_U3088), .B2(n12987), 
        .C1(n14819), .C2(n12986), .ZN(P2_U3305) );
  XNOR2_X1 U14852 ( .A(n12989), .B(n13312), .ZN(n16443) );
  INV_X1 U14853 ( .A(n16443), .ZN(n12998) );
  OAI22_X1 U14854 ( .A1(n14169), .A2(n12991), .B1(n12990), .B2(n16194), .ZN(
        n12995) );
  XNOR2_X1 U14855 ( .A(n12992), .B(n13312), .ZN(n12993) );
  AOI222_X1 U14856 ( .A1(n16183), .A2(n12993), .B1(n13018), .B2(n16178), .C1(
        n13467), .C2(n16180), .ZN(n16440) );
  NOR2_X1 U14857 ( .A1(n16440), .A2(n14164), .ZN(n12994) );
  AOI211_X1 U14858 ( .C1(n14097), .C2(n12996), .A(n12995), .B(n12994), .ZN(
        n12997) );
  OAI21_X1 U14859 ( .B1(n14171), .B2(n12998), .A(n12997), .ZN(P3_U3222) );
  AOI21_X1 U14860 ( .B1(n13001), .B2(n13000), .A(n12999), .ZN(n13008) );
  INV_X1 U14861 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13002) );
  NOR2_X1 U14862 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13002), .ZN(n13908) );
  AOI21_X1 U14863 ( .B1(n13003), .B2(n13026), .A(n13908), .ZN(n13004) );
  OAI21_X1 U14864 ( .B1(n14146), .B2(n13451), .A(n13004), .ZN(n13006) );
  NOR2_X1 U14865 ( .A1(n14236), .A2(n13447), .ZN(n13005) );
  AOI211_X1 U14866 ( .C1(n13029), .C2(n13454), .A(n13006), .B(n13005), .ZN(
        n13007) );
  OAI21_X1 U14867 ( .B1(n13008), .B2(n13458), .A(n13007), .ZN(P3_U3155) );
  NAND2_X1 U14868 ( .A1(n13009), .A2(n14803), .ZN(n13011) );
  OAI211_X1 U14869 ( .C1(n9665), .C2(n14821), .A(n13011), .B(n13010), .ZN(
        P2_U3304) );
  NAND2_X1 U14870 ( .A1(n13009), .A2(n13012), .ZN(n13014) );
  OAI211_X1 U14871 ( .C1(n13015), .C2(n15558), .A(n13014), .B(n13013), .ZN(
        P1_U3332) );
  XNOR2_X1 U14872 ( .A(n13016), .B(n13197), .ZN(n14240) );
  INV_X1 U14873 ( .A(n14240), .ZN(n14304) );
  XNOR2_X1 U14874 ( .A(n13017), .B(n13317), .ZN(n13019) );
  AOI222_X1 U14875 ( .A1(n16183), .A2(n13019), .B1(n13465), .B2(n16178), .C1(
        n13018), .C2(n16180), .ZN(n14237) );
  INV_X1 U14876 ( .A(n14237), .ZN(n13023) );
  AOI22_X1 U14877 ( .A1(n14164), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n14163), 
        .B2(n13020), .ZN(n13021) );
  OAI21_X1 U14878 ( .B1(n14238), .B2(n14166), .A(n13021), .ZN(n13022) );
  AOI21_X1 U14879 ( .B1(n13023), .B2(n14169), .A(n13022), .ZN(n13024) );
  OAI21_X1 U14880 ( .B1(n14171), .B2(n14304), .A(n13024), .ZN(P3_U3220) );
  XNOR2_X1 U14881 ( .A(n13025), .B(n13320), .ZN(n13028) );
  AOI222_X1 U14882 ( .A1(n16183), .A2(n13028), .B1(n13027), .B2(n16178), .C1(
        n13026), .C2(n16180), .ZN(n14235) );
  INV_X1 U14883 ( .A(n14236), .ZN(n13033) );
  INV_X1 U14884 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13031) );
  INV_X1 U14885 ( .A(n13029), .ZN(n13030) );
  OAI22_X1 U14886 ( .A1(n14169), .A2(n13031), .B1(n13030), .B2(n16194), .ZN(
        n13032) );
  AOI21_X1 U14887 ( .B1(n13033), .B2(n14097), .A(n13032), .ZN(n13036) );
  XNOR2_X1 U14888 ( .A(n13034), .B(n13320), .ZN(n14233) );
  NAND2_X1 U14889 ( .A1(n14233), .A2(n14100), .ZN(n13035) );
  OAI211_X1 U14890 ( .C1(n14235), .C2(n14164), .A(n13036), .B(n13035), .ZN(
        P3_U3219) );
  INV_X1 U14891 ( .A(n14229), .ZN(n14167) );
  OAI211_X1 U14892 ( .C1(n13039), .C2(n13038), .A(n13037), .B(n13437), .ZN(
        n13043) );
  INV_X1 U14893 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13775) );
  NOR2_X1 U14894 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13775), .ZN(n13926) );
  AOI21_X1 U14895 ( .B1(n13441), .B2(n14131), .A(n13926), .ZN(n13040) );
  OAI21_X1 U14896 ( .B1(n14160), .B2(n13450), .A(n13040), .ZN(n13041) );
  AOI21_X1 U14897 ( .B1(n14162), .B2(n13454), .A(n13041), .ZN(n13042) );
  OAI211_X1 U14898 ( .C1(n14167), .C2(n13447), .A(n13043), .B(n13042), .ZN(
        P3_U3181) );
  INV_X1 U14899 ( .A(n15378), .ZN(n15383) );
  NAND2_X1 U14900 ( .A1(n15508), .A2(n15129), .ZN(n13044) );
  INV_X1 U14901 ( .A(n15128), .ZN(n13046) );
  NAND2_X1 U14902 ( .A1(n15391), .A2(n13046), .ZN(n13047) );
  NAND2_X1 U14903 ( .A1(n15363), .A2(n13067), .ZN(n13049) );
  OR2_X1 U14904 ( .A1(n15370), .A2(n15127), .ZN(n13048) );
  NAND2_X1 U14905 ( .A1(n13049), .A2(n13048), .ZN(n15358) );
  INV_X1 U14906 ( .A(n15358), .ZN(n13051) );
  NAND2_X1 U14907 ( .A1(n15484), .A2(n15126), .ZN(n13052) );
  INV_X1 U14908 ( .A(n15330), .ZN(n15333) );
  OR2_X1 U14909 ( .A1(n15334), .A2(n15125), .ZN(n13053) );
  INV_X1 U14910 ( .A(n15124), .ZN(n14919) );
  NAND2_X1 U14911 ( .A1(n15326), .A2(n14919), .ZN(n13054) );
  OR2_X1 U14912 ( .A1(n15457), .A2(n15122), .ZN(n13057) );
  NAND2_X1 U14913 ( .A1(n9544), .A2(n15121), .ZN(n13058) );
  NAND2_X1 U14914 ( .A1(n15274), .A2(n15120), .ZN(n13059) );
  OR2_X1 U14915 ( .A1(n15436), .A2(n8086), .ZN(n13061) );
  OR2_X1 U14916 ( .A1(n15508), .A2(n15402), .ZN(n13065) );
  NAND2_X1 U14917 ( .A1(n15391), .A2(n15128), .ZN(n13066) );
  NAND2_X1 U14918 ( .A1(n15346), .A2(n15359), .ZN(n15347) );
  INV_X1 U14919 ( .A(n15126), .ZN(n13068) );
  NAND2_X1 U14920 ( .A1(n15347), .A2(n13069), .ZN(n15331) );
  INV_X1 U14921 ( .A(n15125), .ZN(n13070) );
  INV_X1 U14922 ( .A(n15457), .ZN(n15299) );
  INV_X1 U14923 ( .A(n15120), .ZN(n14965) );
  INV_X1 U14924 ( .A(n15370), .ZN(n15494) );
  NOR2_X2 U14925 ( .A1(n15500), .A2(n15384), .ZN(n15386) );
  NAND2_X1 U14926 ( .A1(n15494), .A2(n15386), .ZN(n15365) );
  AOI21_X1 U14927 ( .B1(n13075), .B2(n7396), .A(n15242), .ZN(n15424) );
  NAND2_X1 U14928 ( .A1(n15424), .A2(n15387), .ZN(n13083) );
  INV_X1 U14929 ( .A(P1_B_REG_SCAN_IN), .ZN(n13076) );
  OR2_X1 U14930 ( .A1(n15689), .A2(n13076), .ZN(n13077) );
  AND2_X1 U14931 ( .A1(n15099), .A2(n13077), .ZN(n15237) );
  NAND2_X1 U14932 ( .A1(n15117), .A2(n15237), .ZN(n15420) );
  OAI22_X1 U14933 ( .A1(n13079), .A2(n15420), .B1(n13078), .B2(n16104), .ZN(
        n13081) );
  NAND2_X1 U14934 ( .A1(n15119), .A2(n15100), .ZN(n15421) );
  NOR2_X1 U14935 ( .A1(n16153), .A2(n15421), .ZN(n13080) );
  AOI211_X1 U14936 ( .C1(n16153), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13081), 
        .B(n13080), .ZN(n13082) );
  OAI211_X1 U14937 ( .C1(n15422), .C2(n16156), .A(n13083), .B(n13082), .ZN(
        n13084) );
  AOI21_X1 U14938 ( .B1(n15419), .B2(n15374), .A(n13084), .ZN(n13085) );
  OAI21_X1 U14939 ( .B1(n15426), .B2(n15412), .A(n13085), .ZN(P1_U3356) );
  INV_X1 U14940 ( .A(n13086), .ZN(n14809) );
  OAI222_X1 U14941 ( .A1(n15558), .A2(n13087), .B1(n15556), .B2(n14809), .C1(
        n15689), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U14942 ( .A(n13088), .ZN(n14801) );
  OAI222_X1 U14943 ( .A1(P1_U3086), .A2(n13090), .B1(n15556), .B2(n14801), 
        .C1(n13089), .C2(n15558), .ZN(P1_U3326) );
  INV_X1 U14944 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13272) );
  OAI222_X1 U14945 ( .A1(n14819), .A2(n13122), .B1(P2_U3088), .B2(n13091), 
        .C1(n13272), .C2(n14821), .ZN(P2_U3297) );
  INV_X1 U14946 ( .A(n14804), .ZN(n13092) );
  OAI222_X1 U14947 ( .A1(n15558), .A2(n13093), .B1(n15556), .B2(n13092), .C1(
        n9598), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI22_X1 U14948 ( .A1(n13096), .A2(n16117), .B1(n13095), .B2(n14675), .ZN(
        n13097) );
  AOI21_X1 U14949 ( .B1(n13098), .B2(n16399), .A(n13097), .ZN(n13099) );
  OAI21_X1 U14950 ( .B1(n13100), .B2(n16228), .A(n13099), .ZN(n13101) );
  AOI21_X1 U14951 ( .B1(n13102), .B2(n14678), .A(n13101), .ZN(n13103) );
  OAI21_X1 U14952 ( .B1(n13094), .B2(n16408), .A(n13103), .ZN(P2_U3236) );
  NAND2_X1 U14953 ( .A1(n13104), .A2(n13124), .ZN(n13105) );
  AND2_X2 U14954 ( .A1(n13106), .A2(n13105), .ZN(n14250) );
  AND2_X1 U14955 ( .A1(n13969), .A2(n13107), .ZN(n13114) );
  AND2_X1 U14956 ( .A1(n13110), .A2(n13109), .ZN(n13112) );
  NAND2_X1 U14957 ( .A1(n13112), .A2(n13111), .ZN(n13113) );
  NAND2_X1 U14958 ( .A1(n13114), .A2(n13113), .ZN(n13115) );
  AOI22_X1 U14959 ( .A1(n13116), .A2(n16178), .B1(n16180), .B2(n13462), .ZN(
        n13117) );
  NAND2_X1 U14960 ( .A1(n16473), .A2(n16382), .ZN(n14243) );
  INV_X1 U14961 ( .A(n13987), .ZN(n14249) );
  OAI22_X1 U14962 ( .A1(n14250), .A2(n14243), .B1(n14249), .B2(n14227), .ZN(
        n13118) );
  INV_X1 U14963 ( .A(n13119), .ZN(n13121) );
  OAI222_X1 U14964 ( .A1(n14312), .A2(n13121), .B1(n13335), .B2(P3_U3151), 
        .C1(n13120), .C2(n14315), .ZN(P3_U3267) );
  NAND2_X1 U14965 ( .A1(n13997), .A2(n14014), .ZN(n13123) );
  INV_X1 U14966 ( .A(n13132), .ZN(n13128) );
  AOI211_X1 U14967 ( .C1(n13130), .C2(n13129), .A(n13128), .B(n13222), .ZN(
        n13135) );
  AOI211_X1 U14968 ( .C1(n13133), .C2(n13132), .A(n13131), .B(n13299), .ZN(
        n13134) );
  MUX2_X1 U14969 ( .A(n13135), .B(n13134), .S(n13266), .Z(n13225) );
  NAND2_X1 U14970 ( .A1(n13137), .A2(n13140), .ZN(n13136) );
  NAND2_X1 U14971 ( .A1(n13143), .A2(n13136), .ZN(n13139) );
  INV_X1 U14972 ( .A(n13137), .ZN(n13138) );
  MUX2_X1 U14973 ( .A(n13139), .B(n13138), .S(n13266), .Z(n13152) );
  NAND2_X1 U14974 ( .A1(n13140), .A2(n10118), .ZN(n13141) );
  NAND4_X1 U14975 ( .A1(n13143), .A2(n13142), .A3(n13266), .A4(n13141), .ZN(
        n13144) );
  NAND2_X1 U14976 ( .A1(n10066), .A2(n13144), .ZN(n13151) );
  NAND2_X1 U14977 ( .A1(n13154), .A2(n13145), .ZN(n13148) );
  NAND2_X1 U14978 ( .A1(n13153), .A2(n13146), .ZN(n13147) );
  MUX2_X1 U14979 ( .A(n13148), .B(n13147), .S(n13266), .Z(n13149) );
  INV_X1 U14980 ( .A(n13149), .ZN(n13150) );
  OAI21_X1 U14981 ( .B1(n13152), .B2(n13151), .A(n13150), .ZN(n13156) );
  MUX2_X1 U14982 ( .A(n13154), .B(n13153), .S(n13207), .Z(n13155) );
  NAND3_X1 U14983 ( .A1(n13156), .A2(n13306), .A3(n13155), .ZN(n13160) );
  MUX2_X1 U14984 ( .A(n13158), .B(n13157), .S(n13266), .Z(n13159) );
  NAND3_X1 U14985 ( .A1(n13160), .A2(n13302), .A3(n13159), .ZN(n13165) );
  MUX2_X1 U14986 ( .A(n13162), .B(n13161), .S(n13266), .Z(n13163) );
  NAND3_X1 U14987 ( .A1(n13165), .A2(n13164), .A3(n13163), .ZN(n13169) );
  MUX2_X1 U14988 ( .A(n13472), .B(n16333), .S(n13266), .Z(n13166) );
  AOI21_X1 U14989 ( .B1(n13167), .B2(n13166), .A(n13305), .ZN(n13168) );
  NAND2_X1 U14990 ( .A1(n13169), .A2(n13168), .ZN(n13174) );
  MUX2_X1 U14991 ( .A(n13171), .B(n13170), .S(n13266), .Z(n13172) );
  NAND3_X1 U14992 ( .A1(n13174), .A2(n13173), .A3(n13172), .ZN(n13179) );
  MUX2_X1 U14993 ( .A(n13176), .B(n13175), .S(n13266), .Z(n13177) );
  NAND3_X1 U14994 ( .A1(n13179), .A2(n13178), .A3(n13177), .ZN(n13183) );
  MUX2_X1 U14995 ( .A(n13181), .B(n13180), .S(n13207), .Z(n13182) );
  NAND2_X1 U14996 ( .A1(n13183), .A2(n13182), .ZN(n13186) );
  OAI21_X1 U14997 ( .B1(n13266), .B2(n13184), .A(n13312), .ZN(n13185) );
  AOI21_X1 U14998 ( .B1(n13186), .B2(n13313), .A(n13185), .ZN(n13193) );
  INV_X1 U14999 ( .A(n13193), .ZN(n13189) );
  NAND4_X1 U15000 ( .A1(n13189), .A2(n13207), .A3(n13188), .A4(n13187), .ZN(
        n13199) );
  INV_X1 U15001 ( .A(n13190), .ZN(n13191) );
  AOI21_X1 U15002 ( .B1(n13193), .B2(n13192), .A(n13191), .ZN(n13196) );
  XNOR2_X1 U15003 ( .A(n13194), .B(n13266), .ZN(n13195) );
  OAI21_X1 U15004 ( .B1(n13196), .B2(n13318), .A(n13195), .ZN(n13198) );
  NAND3_X1 U15005 ( .A1(n13199), .A2(n13198), .A3(n13197), .ZN(n13205) );
  INV_X1 U15006 ( .A(n13200), .ZN(n13202) );
  MUX2_X1 U15007 ( .A(n13202), .B(n7892), .S(n13266), .Z(n13203) );
  NOR2_X1 U15008 ( .A1(n14154), .A2(n13203), .ZN(n13204) );
  NAND3_X1 U15009 ( .A1(n13205), .A2(n13320), .A3(n13204), .ZN(n13215) );
  MUX2_X1 U15010 ( .A(n14160), .B(n13266), .S(n14236), .Z(n13206) );
  OAI21_X1 U15011 ( .B1(n13207), .B2(n13465), .A(n13206), .ZN(n13208) );
  NAND2_X1 U15012 ( .A1(n13209), .A2(n13208), .ZN(n13213) );
  MUX2_X1 U15013 ( .A(n13211), .B(n13210), .S(n13266), .Z(n13212) );
  NAND2_X1 U15014 ( .A1(n13213), .A2(n13212), .ZN(n13214) );
  NAND3_X1 U15015 ( .A1(n13215), .A2(n13214), .A3(n14144), .ZN(n13220) );
  INV_X1 U15016 ( .A(n13216), .ZN(n14297) );
  NAND2_X1 U15017 ( .A1(n14297), .A2(n14131), .ZN(n13218) );
  MUX2_X1 U15018 ( .A(n13218), .B(n13217), .S(n13266), .Z(n13219) );
  NAND2_X1 U15019 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  NAND3_X1 U15020 ( .A1(n14116), .A2(n13321), .A3(n13221), .ZN(n13224) );
  MUX2_X1 U15021 ( .A(n13299), .B(n13222), .S(n13266), .Z(n13223) );
  AOI21_X1 U15022 ( .B1(n13225), .B2(n13224), .A(n13223), .ZN(n13229) );
  AND2_X1 U15023 ( .A1(n14205), .A2(n14109), .ZN(n13226) );
  MUX2_X1 U15024 ( .A(n13227), .B(n13226), .S(n13266), .Z(n13228) );
  AOI211_X1 U15025 ( .C1(n13229), .C2(n14098), .A(n13228), .B(n14069), .ZN(
        n13233) );
  MUX2_X1 U15026 ( .A(n13231), .B(n13230), .S(n13266), .Z(n13232) );
  NOR3_X1 U15027 ( .A1(n13233), .A2(n13232), .A3(n14051), .ZN(n13238) );
  NOR3_X1 U15028 ( .A1(n13126), .A2(n13359), .A3(n10022), .ZN(n13235) );
  INV_X1 U15029 ( .A(n13237), .ZN(n13239) );
  NAND3_X1 U15030 ( .A1(n13240), .A2(n14028), .A3(n13367), .ZN(n13241) );
  OAI211_X1 U15031 ( .C1(n13126), .C2(n13242), .A(n13241), .B(n13291), .ZN(
        n13243) );
  NOR2_X1 U15032 ( .A1(n13244), .A2(n13243), .ZN(n13262) );
  INV_X1 U15033 ( .A(n13257), .ZN(n13254) );
  NAND2_X1 U15034 ( .A1(n13245), .A2(n13992), .ZN(n13247) );
  AND2_X1 U15035 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  NAND2_X1 U15036 ( .A1(n13249), .A2(n13248), .ZN(n13251) );
  NAND2_X1 U15037 ( .A1(n13251), .A2(n13250), .ZN(n13255) );
  INV_X1 U15038 ( .A(n13255), .ZN(n13252) );
  OAI21_X1 U15039 ( .B1(n13254), .B2(n13253), .A(n13252), .ZN(n13259) );
  AOI21_X1 U15040 ( .B1(n13257), .B2(n13256), .A(n13255), .ZN(n13258) );
  MUX2_X1 U15041 ( .A(n13259), .B(n13258), .S(n13266), .Z(n13260) );
  NAND3_X1 U15042 ( .A1(n8009), .A2(n13977), .A3(n13260), .ZN(n13261) );
  INV_X1 U15043 ( .A(n13263), .ZN(n13264) );
  NAND2_X1 U15044 ( .A1(n13265), .A2(n13264), .ZN(n13267) );
  AOI22_X1 U15045 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13272), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n13268), .ZN(n13277) );
  NAND2_X1 U15046 ( .A1(n13277), .A2(n13276), .ZN(n13271) );
  OAI21_X1 U15047 ( .B1(n13272), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n13271), 
        .ZN(n13275) );
  INV_X1 U15048 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13273) );
  AOI22_X1 U15049 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n13273), .B2(n9470), .ZN(n13274) );
  XNOR2_X1 U15050 ( .A(n13275), .B(n13274), .ZN(n14308) );
  INV_X1 U15051 ( .A(n13276), .ZN(n13278) );
  XNOR2_X1 U15052 ( .A(n13278), .B(n13277), .ZN(n13355) );
  NAND2_X1 U15053 ( .A1(n10032), .A2(n13355), .ZN(n13281) );
  NAND2_X1 U15054 ( .A1(n13279), .A2(SI_30_), .ZN(n13280) );
  NAND2_X1 U15055 ( .A1(n13281), .A2(n13280), .ZN(n16556) );
  AOI22_X1 U15056 ( .A1(n14173), .A2(n13955), .B1(n13282), .B2(n16556), .ZN(
        n13292) );
  INV_X1 U15057 ( .A(n13955), .ZN(n13283) );
  NAND2_X1 U15058 ( .A1(n16559), .A2(n13283), .ZN(n13285) );
  NAND2_X1 U15059 ( .A1(n13460), .A2(n14176), .ZN(n13284) );
  NAND2_X1 U15060 ( .A1(n13285), .A2(n13284), .ZN(n13286) );
  INV_X1 U15061 ( .A(n13286), .ZN(n13325) );
  NAND2_X1 U15062 ( .A1(n13286), .A2(n16559), .ZN(n13296) );
  OAI21_X1 U15063 ( .B1(n14176), .B2(n13955), .A(n13291), .ZN(n13293) );
  INV_X1 U15064 ( .A(n13292), .ZN(n13326) );
  AOI211_X1 U15065 ( .C1(n13295), .C2(n13294), .A(n13293), .B(n13326), .ZN(
        n13298) );
  INV_X1 U15066 ( .A(n13296), .ZN(n13297) );
  INV_X1 U15067 ( .A(n14051), .ZN(n14057) );
  INV_X1 U15068 ( .A(n14116), .ZN(n13323) );
  INV_X1 U15069 ( .A(n13299), .ZN(n13301) );
  NAND2_X1 U15070 ( .A1(n13301), .A2(n13300), .ZN(n14106) );
  NOR4_X1 U15071 ( .A1(n9743), .A2(n13305), .A3(n13304), .A4(n13303), .ZN(
        n13315) );
  NAND3_X1 U15072 ( .A1(n10066), .A2(n13307), .A3(n13306), .ZN(n13311) );
  INV_X1 U15073 ( .A(n13308), .ZN(n13310) );
  NOR4_X1 U15074 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n12289), .ZN(
        n13314) );
  NAND4_X1 U15075 ( .A1(n13315), .A2(n13314), .A3(n13313), .A4(n13312), .ZN(
        n13316) );
  NOR4_X1 U15076 ( .A1(n14154), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13319) );
  NAND4_X1 U15077 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n14144), .ZN(
        n13322) );
  NOR4_X1 U15078 ( .A1(n14069), .A2(n13323), .A3(n14106), .A4(n13322), .ZN(
        n13324) );
  NAND4_X1 U15079 ( .A1(n13325), .A2(n14057), .A3(n13324), .A4(n14098), .ZN(
        n13327) );
  NOR3_X1 U15080 ( .A1(n13328), .A2(n13327), .A3(n13326), .ZN(n13329) );
  XOR2_X1 U15081 ( .A(n13330), .B(n13329), .Z(n13331) );
  NOR4_X1 U15082 ( .A1(n13337), .A2(n13336), .A3(n13335), .A4(n13334), .ZN(
        n13340) );
  OAI21_X1 U15083 ( .B1(n13341), .B2(n13338), .A(P3_B_REG_SCAN_IN), .ZN(n13339) );
  OAI22_X1 U15084 ( .A1(n13342), .A2(n13341), .B1(n13340), .B2(n13339), .ZN(
        P3_U3296) );
  NAND2_X1 U15085 ( .A1(n13345), .A2(n13344), .ZN(n13346) );
  AOI22_X1 U15086 ( .A1(n15100), .A2(n8086), .B1(n15118), .B2(n15099), .ZN(
        n15011) );
  NAND2_X1 U15087 ( .A1(n15251), .A2(n15428), .ZN(n13349) );
  AOI22_X1 U15088 ( .A1(n16153), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n15013), 
        .B2(n16312), .ZN(n13350) );
  OAI21_X1 U15089 ( .B1(n15006), .B2(n16156), .A(n13350), .ZN(n13353) );
  NOR2_X1 U15090 ( .A1(n15431), .A2(n13351), .ZN(n13352) );
  AOI211_X1 U15091 ( .C1(n15387), .C2(n15429), .A(n13353), .B(n13352), .ZN(
        n13354) );
  OAI21_X1 U15092 ( .B1(n15434), .B2(n16153), .A(n13354), .ZN(P1_U3265) );
  INV_X1 U15093 ( .A(n13355), .ZN(n13357) );
  INV_X1 U15094 ( .A(SI_30_), .ZN(n13673) );
  OAI222_X1 U15095 ( .A1(n14312), .A2(n13357), .B1(n13356), .B2(P3_U3151), 
        .C1(n13673), .C2(n14315), .ZN(P3_U3265) );
  INV_X1 U15096 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n13723) );
  OAI22_X1 U15097 ( .A1(n14010), .A2(n13450), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13723), .ZN(n13361) );
  NOR2_X1 U15098 ( .A1(n13359), .A2(n13451), .ZN(n13360) );
  AOI211_X1 U15099 ( .C1(n13986), .C2(n13454), .A(n13361), .B(n13360), .ZN(
        n13362) );
  OAI211_X1 U15100 ( .C1(n14249), .C2(n13447), .A(n13363), .B(n13362), .ZN(
        P3_U3154) );
  XNOR2_X1 U15101 ( .A(n13412), .B(n13411), .ZN(n13413) );
  XNOR2_X1 U15102 ( .A(n13413), .B(n14028), .ZN(n13369) );
  AOI22_X1 U15103 ( .A1(n14042), .A2(n13441), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13365) );
  NAND2_X1 U15104 ( .A1(n13454), .A2(n14045), .ZN(n13364) );
  OAI211_X1 U15105 ( .C1(n14073), .C2(n13450), .A(n13365), .B(n13364), .ZN(
        n13366) );
  AOI21_X1 U15106 ( .B1(n13367), .B2(n13455), .A(n13366), .ZN(n13368) );
  OAI21_X1 U15107 ( .B1(n13369), .B2(n13458), .A(n13368), .ZN(P3_U3156) );
  OAI211_X1 U15108 ( .C1(n13372), .C2(n13371), .A(n13370), .B(n13437), .ZN(
        n13377) );
  AOI21_X1 U15109 ( .B1(n13464), .B2(n13441), .A(n13373), .ZN(n13374) );
  OAI21_X1 U15110 ( .B1(n14108), .B2(n13450), .A(n13374), .ZN(n13375) );
  AOI21_X1 U15111 ( .B1(n14110), .B2(n13454), .A(n13375), .ZN(n13376) );
  OAI211_X1 U15112 ( .C1(n13447), .C2(n14287), .A(n13377), .B(n13376), .ZN(
        P3_U3159) );
  INV_X1 U15113 ( .A(n13378), .ZN(n13379) );
  NOR2_X1 U15114 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  XNOR2_X1 U15115 ( .A(n13382), .B(n13381), .ZN(n13387) );
  OAI22_X1 U15116 ( .A1(n14109), .A2(n13450), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13740), .ZN(n13384) );
  NOR2_X1 U15117 ( .A1(n14073), .A2(n13451), .ZN(n13383) );
  AOI211_X1 U15118 ( .C1(n14079), .C2(n13454), .A(n13384), .B(n13383), .ZN(
        n13386) );
  NAND2_X1 U15119 ( .A1(n14202), .A2(n13455), .ZN(n13385) );
  OAI211_X1 U15120 ( .C1(n13387), .C2(n13458), .A(n13386), .B(n13385), .ZN(
        P3_U3163) );
  XOR2_X1 U15121 ( .A(n13389), .B(n13388), .Z(n13394) );
  OAI22_X1 U15122 ( .A1(n14009), .A2(n13450), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13541), .ZN(n13391) );
  NOR2_X1 U15123 ( .A1(n14010), .A2(n13451), .ZN(n13390) );
  AOI211_X1 U15124 ( .C1(n14018), .C2(n13454), .A(n13391), .B(n13390), .ZN(
        n13393) );
  NAND2_X1 U15125 ( .A1(n14260), .A2(n13455), .ZN(n13392) );
  OAI211_X1 U15126 ( .C1(n13394), .C2(n13458), .A(n13393), .B(n13392), .ZN(
        P3_U3165) );
  XNOR2_X1 U15127 ( .A(n13396), .B(n13395), .ZN(n13402) );
  NAND2_X1 U15128 ( .A1(n13397), .A2(n13441), .ZN(n13398) );
  NAND2_X1 U15129 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n16058)
         );
  OAI211_X1 U15130 ( .C1(n14146), .C2(n13450), .A(n13398), .B(n16058), .ZN(
        n13400) );
  NOR2_X1 U15131 ( .A1(n14297), .A2(n13447), .ZN(n13399) );
  AOI211_X1 U15132 ( .C1(n14148), .C2(n13454), .A(n13400), .B(n13399), .ZN(
        n13401) );
  OAI21_X1 U15133 ( .B1(n13402), .B2(n13458), .A(n13401), .ZN(P3_U3166) );
  XNOR2_X1 U15134 ( .A(n13403), .B(n14147), .ZN(n13404) );
  XNOR2_X1 U15135 ( .A(n13405), .B(n13404), .ZN(n13410) );
  NOR2_X1 U15136 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13748), .ZN(n16072) );
  AOI21_X1 U15137 ( .B1(n14132), .B2(n13441), .A(n16072), .ZN(n13407) );
  NAND2_X1 U15138 ( .A1(n13454), .A2(n14135), .ZN(n13406) );
  OAI211_X1 U15139 ( .C1(n14158), .C2(n13450), .A(n13407), .B(n13406), .ZN(
        n13408) );
  AOI21_X1 U15140 ( .B1(n14220), .B2(n13455), .A(n13408), .ZN(n13409) );
  OAI21_X1 U15141 ( .B1(n13410), .B2(n13458), .A(n13409), .ZN(P3_U3168) );
  OAI22_X1 U15142 ( .A1(n13413), .A2(n14056), .B1(n13412), .B2(n13411), .ZN(
        n13416) );
  XNOR2_X1 U15143 ( .A(n13414), .B(n14042), .ZN(n13415) );
  XNOR2_X1 U15144 ( .A(n13416), .B(n13415), .ZN(n13417) );
  NAND2_X1 U15145 ( .A1(n13417), .A2(n13437), .ZN(n13421) );
  INV_X1 U15146 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n13751) );
  OAI22_X1 U15147 ( .A1(n14028), .A2(n13450), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13751), .ZN(n13419) );
  NOR2_X1 U15148 ( .A1(n14027), .A2(n13451), .ZN(n13418) );
  AOI211_X1 U15149 ( .C1(n14031), .C2(n13454), .A(n13419), .B(n13418), .ZN(
        n13420) );
  OAI211_X1 U15150 ( .C1(n14265), .C2(n13447), .A(n13421), .B(n13420), .ZN(
        P3_U3169) );
  XNOR2_X1 U15151 ( .A(n13422), .B(n13464), .ZN(n13423) );
  XNOR2_X1 U15152 ( .A(n13424), .B(n13423), .ZN(n13429) );
  AOI22_X1 U15153 ( .A1(n14055), .A2(n13441), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13426) );
  NAND2_X1 U15154 ( .A1(n13454), .A2(n14093), .ZN(n13425) );
  OAI211_X1 U15155 ( .C1(n14122), .C2(n13450), .A(n13426), .B(n13425), .ZN(
        n13427) );
  AOI21_X1 U15156 ( .B1(n14205), .B2(n13455), .A(n13427), .ZN(n13428) );
  OAI21_X1 U15157 ( .B1(n13429), .B2(n13458), .A(n13428), .ZN(P3_U3173) );
  XNOR2_X1 U15158 ( .A(n13430), .B(n14041), .ZN(n13435) );
  INV_X1 U15159 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13761) );
  OAI22_X1 U15160 ( .A1(n14089), .A2(n13450), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13761), .ZN(n13432) );
  NOR2_X1 U15161 ( .A1(n14028), .A2(n13451), .ZN(n13431) );
  AOI211_X1 U15162 ( .C1(n14063), .C2(n13454), .A(n13432), .B(n13431), .ZN(
        n13434) );
  NAND2_X1 U15163 ( .A1(n14199), .A2(n13455), .ZN(n13433) );
  OAI211_X1 U15164 ( .C1(n13435), .C2(n13458), .A(n13434), .B(n13433), .ZN(
        P3_U3175) );
  INV_X1 U15165 ( .A(n13436), .ZN(n14291) );
  OAI211_X1 U15166 ( .C1(n13440), .C2(n13439), .A(n13438), .B(n13437), .ZN(
        n13446) );
  NAND2_X1 U15167 ( .A1(n13442), .A2(n13441), .ZN(n13443) );
  NAND2_X1 U15168 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13942)
         );
  OAI211_X1 U15169 ( .C1(n14147), .C2(n13450), .A(n13443), .B(n13942), .ZN(
        n13444) );
  AOI21_X1 U15170 ( .B1(n14123), .B2(n13454), .A(n13444), .ZN(n13445) );
  OAI211_X1 U15171 ( .C1(n14291), .C2(n13447), .A(n13446), .B(n13445), .ZN(
        P3_U3178) );
  XOR2_X1 U15172 ( .A(n13449), .B(n13448), .Z(n13459) );
  INV_X1 U15173 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n13772) );
  OAI22_X1 U15174 ( .A1(n14027), .A2(n13450), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13772), .ZN(n13453) );
  NOR2_X1 U15175 ( .A1(n13999), .A2(n13451), .ZN(n13452) );
  AOI211_X1 U15176 ( .C1(n14003), .C2(n13454), .A(n13453), .B(n13452), .ZN(
        n13457) );
  NAND2_X1 U15177 ( .A1(n14255), .A2(n13455), .ZN(n13456) );
  OAI211_X1 U15178 ( .C1(n13459), .C2(n13458), .A(n13457), .B(n13456), .ZN(
        P3_U3180) );
  MUX2_X1 U15179 ( .A(n13460), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13471), .Z(
        P3_U3521) );
  MUX2_X1 U15180 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13461), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15181 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13462), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15182 ( .A(n13463), .B(P3_DATAO_REG_25__SCAN_IN), .S(n13471), .Z(
        P3_U3516) );
  MUX2_X1 U15183 ( .A(n14042), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13471), .Z(
        P3_U3515) );
  MUX2_X1 U15184 ( .A(n14056), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13471), .Z(
        P3_U3514) );
  MUX2_X1 U15185 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n14041), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15186 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n14055), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15187 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13464), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15188 ( .A(n13465), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13471), .Z(
        P3_U3505) );
  MUX2_X1 U15189 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13466), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15190 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13467), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15191 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13468), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15192 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13469), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15193 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13470), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15194 ( .A(n13472), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13471), .Z(
        P3_U3497) );
  MUX2_X1 U15195 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13474), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15196 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13475), .S(P3_U3897), .Z(
        P3_U3495) );
  XNOR2_X1 U15197 ( .A(SI_31_), .B(keyinput_129), .ZN(n13478) );
  XNOR2_X1 U15198 ( .A(SI_30_), .B(keyinput_130), .ZN(n13477) );
  XNOR2_X1 U15199 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n13476) );
  NOR3_X1 U15200 ( .A1(n13478), .A2(n13477), .A3(n13476), .ZN(n13481) );
  XOR2_X1 U15201 ( .A(SI_28_), .B(keyinput_132), .Z(n13480) );
  XNOR2_X1 U15202 ( .A(SI_29_), .B(keyinput_131), .ZN(n13479) );
  NOR3_X1 U15203 ( .A1(n13481), .A2(n13480), .A3(n13479), .ZN(n13484) );
  XNOR2_X1 U15204 ( .A(SI_27_), .B(keyinput_133), .ZN(n13483) );
  XNOR2_X1 U15205 ( .A(SI_26_), .B(keyinput_134), .ZN(n13482) );
  OAI21_X1 U15206 ( .B1(n13484), .B2(n13483), .A(n13482), .ZN(n13488) );
  XOR2_X1 U15207 ( .A(SI_25_), .B(keyinput_135), .Z(n13487) );
  XNOR2_X1 U15208 ( .A(SI_24_), .B(keyinput_136), .ZN(n13486) );
  XNOR2_X1 U15209 ( .A(SI_23_), .B(keyinput_137), .ZN(n13485) );
  NAND4_X1 U15210 ( .A1(n13488), .A2(n13487), .A3(n13486), .A4(n13485), .ZN(
        n13491) );
  XNOR2_X1 U15211 ( .A(SI_22_), .B(keyinput_138), .ZN(n13490) );
  XNOR2_X1 U15212 ( .A(SI_21_), .B(keyinput_139), .ZN(n13489) );
  NAND3_X1 U15213 ( .A1(n13491), .A2(n13490), .A3(n13489), .ZN(n13495) );
  XOR2_X1 U15214 ( .A(SI_18_), .B(keyinput_142), .Z(n13494) );
  XNOR2_X1 U15215 ( .A(SI_19_), .B(keyinput_141), .ZN(n13493) );
  XNOR2_X1 U15216 ( .A(SI_20_), .B(keyinput_140), .ZN(n13492) );
  NAND4_X1 U15217 ( .A1(n13495), .A2(n13494), .A3(n13493), .A4(n13492), .ZN(
        n13501) );
  XNOR2_X1 U15218 ( .A(SI_17_), .B(keyinput_143), .ZN(n13500) );
  XOR2_X1 U15219 ( .A(SI_16_), .B(keyinput_144), .Z(n13498) );
  XNOR2_X1 U15220 ( .A(SI_14_), .B(keyinput_146), .ZN(n13497) );
  XNOR2_X1 U15221 ( .A(SI_15_), .B(keyinput_145), .ZN(n13496) );
  NAND3_X1 U15222 ( .A1(n13498), .A2(n13497), .A3(n13496), .ZN(n13499) );
  AOI21_X1 U15223 ( .B1(n13501), .B2(n13500), .A(n13499), .ZN(n13505) );
  XNOR2_X1 U15224 ( .A(n13695), .B(keyinput_147), .ZN(n13504) );
  XNOR2_X1 U15225 ( .A(n13698), .B(keyinput_149), .ZN(n13503) );
  XNOR2_X1 U15226 ( .A(n13699), .B(keyinput_148), .ZN(n13502) );
  OAI211_X1 U15227 ( .C1(n13505), .C2(n13504), .A(n13503), .B(n13502), .ZN(
        n13509) );
  XNOR2_X1 U15228 ( .A(n13506), .B(keyinput_151), .ZN(n13508) );
  XNOR2_X1 U15229 ( .A(SI_10_), .B(keyinput_150), .ZN(n13507) );
  NAND3_X1 U15230 ( .A1(n13509), .A2(n13508), .A3(n13507), .ZN(n13513) );
  XOR2_X1 U15231 ( .A(SI_6_), .B(keyinput_154), .Z(n13512) );
  XOR2_X1 U15232 ( .A(SI_8_), .B(keyinput_152), .Z(n13511) );
  XNOR2_X1 U15233 ( .A(SI_7_), .B(keyinput_153), .ZN(n13510) );
  NAND4_X1 U15234 ( .A1(n13513), .A2(n13512), .A3(n13511), .A4(n13510), .ZN(
        n13516) );
  XNOR2_X1 U15235 ( .A(n7656), .B(keyinput_156), .ZN(n13515) );
  XNOR2_X1 U15236 ( .A(n13666), .B(keyinput_155), .ZN(n13514) );
  NAND3_X1 U15237 ( .A1(n13516), .A2(n13515), .A3(n13514), .ZN(n13520) );
  XNOR2_X1 U15238 ( .A(n13715), .B(keyinput_157), .ZN(n13519) );
  XOR2_X1 U15239 ( .A(SI_1_), .B(keyinput_159), .Z(n13518) );
  XNOR2_X1 U15240 ( .A(SI_2_), .B(keyinput_158), .ZN(n13517) );
  NAND4_X1 U15241 ( .A1(n13520), .A2(n13519), .A3(n13518), .A4(n13517), .ZN(
        n13527) );
  XOR2_X1 U15242 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_162), .Z(n13524) );
  XOR2_X1 U15243 ( .A(SI_0_), .B(keyinput_160), .Z(n13523) );
  XOR2_X1 U15244 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_163), .Z(n13522) );
  XNOR2_X1 U15245 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n13521) );
  NOR4_X1 U15246 ( .A1(n13524), .A2(n13523), .A3(n13522), .A4(n13521), .ZN(
        n13526) );
  XOR2_X1 U15247 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_164), .Z(n13525)
         );
  AOI21_X1 U15248 ( .B1(n13527), .B2(n13526), .A(n13525), .ZN(n13530) );
  XOR2_X1 U15249 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_165), .Z(n13529)
         );
  XNOR2_X1 U15250 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n13528)
         );
  NOR3_X1 U15251 ( .A1(n13530), .A2(n13529), .A3(n13528), .ZN(n13533) );
  XOR2_X1 U15252 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_167), .Z(n13532)
         );
  XNOR2_X1 U15253 ( .A(n13734), .B(keyinput_168), .ZN(n13531) );
  OAI21_X1 U15254 ( .B1(n13533), .B2(n13532), .A(n13531), .ZN(n13536) );
  XOR2_X1 U15255 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_169), .Z(n13535)
         );
  XNOR2_X1 U15256 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n13534)
         );
  NAND3_X1 U15257 ( .A1(n13536), .A2(n13535), .A3(n13534), .ZN(n13547) );
  XNOR2_X1 U15258 ( .A(n13740), .B(keyinput_173), .ZN(n13540) );
  XNOR2_X1 U15259 ( .A(n13737), .B(keyinput_171), .ZN(n13539) );
  XNOR2_X1 U15260 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n13538)
         );
  XNOR2_X1 U15261 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n13537)
         );
  NOR4_X1 U15262 ( .A1(n13540), .A2(n13539), .A3(n13538), .A4(n13537), .ZN(
        n13546) );
  XNOR2_X1 U15263 ( .A(n13541), .B(keyinput_175), .ZN(n13544) );
  XNOR2_X1 U15264 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput_177), .ZN(n13543)
         );
  XNOR2_X1 U15265 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n13542)
         );
  NAND3_X1 U15266 ( .A1(n13544), .A2(n13543), .A3(n13542), .ZN(n13545) );
  AOI21_X1 U15267 ( .B1(n13547), .B2(n13546), .A(n13545), .ZN(n13550) );
  XNOR2_X1 U15268 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n13549)
         );
  XNOR2_X1 U15269 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_179), .ZN(n13548)
         );
  OAI21_X1 U15270 ( .B1(n13550), .B2(n13549), .A(n13548), .ZN(n13554) );
  XOR2_X1 U15271 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_180), .Z(n13553) );
  XNOR2_X1 U15272 ( .A(n13551), .B(keyinput_181), .ZN(n13552) );
  AOI21_X1 U15273 ( .B1(n13554), .B2(n13553), .A(n13552), .ZN(n13564) );
  XNOR2_X1 U15274 ( .A(n13555), .B(keyinput_184), .ZN(n13560) );
  XNOR2_X1 U15275 ( .A(n13556), .B(keyinput_183), .ZN(n13559) );
  XNOR2_X1 U15276 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n13558)
         );
  XNOR2_X1 U15277 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n13557)
         );
  NAND4_X1 U15278 ( .A1(n13560), .A2(n13559), .A3(n13558), .A4(n13557), .ZN(
        n13563) );
  XNOR2_X1 U15279 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n13562)
         );
  XNOR2_X1 U15280 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n13561)
         );
  OAI211_X1 U15281 ( .C1(n13564), .C2(n13563), .A(n13562), .B(n13561), .ZN(
        n13566) );
  XOR2_X1 U15282 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_188), .Z(n13565)
         );
  NAND2_X1 U15283 ( .A1(n13566), .A2(n13565), .ZN(n13572) );
  OAI22_X1 U15284 ( .A1(n13775), .A2(keyinput_191), .B1(keyinput_192), .B2(
        P3_B_REG_SCAN_IN), .ZN(n13567) );
  AOI221_X1 U15285 ( .B1(n13775), .B2(keyinput_191), .C1(P3_B_REG_SCAN_IN), 
        .C2(keyinput_192), .A(n13567), .ZN(n13571) );
  XOR2_X1 U15286 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_189), .Z(n13570) );
  OAI22_X1 U15287 ( .A1(n13773), .A2(keyinput_193), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_190), .ZN(n13568) );
  AOI221_X1 U15288 ( .B1(n13773), .B2(keyinput_193), .C1(keyinput_190), .C2(
        P3_REG3_REG_26__SCAN_IN), .A(n13568), .ZN(n13569) );
  NAND4_X1 U15289 ( .A1(n13572), .A2(n13571), .A3(n13570), .A4(n13569), .ZN(
        n13579) );
  XOR2_X1 U15290 ( .A(keyinput_195), .B(P3_DATAO_REG_29__SCAN_IN), .Z(n13576)
         );
  XOR2_X1 U15291 ( .A(keyinput_194), .B(P3_DATAO_REG_30__SCAN_IN), .Z(n13575)
         );
  XOR2_X1 U15292 ( .A(keyinput_197), .B(P3_DATAO_REG_27__SCAN_IN), .Z(n13574)
         );
  XNOR2_X1 U15293 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n13573) );
  NOR4_X1 U15294 ( .A1(n13576), .A2(n13575), .A3(n13574), .A4(n13573), .ZN(
        n13578) );
  XNOR2_X1 U15295 ( .A(keyinput_198), .B(P3_DATAO_REG_26__SCAN_IN), .ZN(n13577) );
  AOI21_X1 U15296 ( .B1(n13579), .B2(n13578), .A(n13577), .ZN(n13583) );
  XOR2_X1 U15297 ( .A(keyinput_199), .B(P3_DATAO_REG_25__SCAN_IN), .Z(n13582)
         );
  XNOR2_X1 U15298 ( .A(keyinput_201), .B(P3_DATAO_REG_23__SCAN_IN), .ZN(n13581) );
  XNOR2_X1 U15299 ( .A(keyinput_200), .B(P3_DATAO_REG_24__SCAN_IN), .ZN(n13580) );
  OAI211_X1 U15300 ( .C1(n13583), .C2(n13582), .A(n13581), .B(n13580), .ZN(
        n13586) );
  XOR2_X1 U15301 ( .A(keyinput_203), .B(P3_DATAO_REG_21__SCAN_IN), .Z(n13585)
         );
  XNOR2_X1 U15302 ( .A(keyinput_202), .B(P3_DATAO_REG_22__SCAN_IN), .ZN(n13584) );
  NAND3_X1 U15303 ( .A1(n13586), .A2(n13585), .A3(n13584), .ZN(n13589) );
  XNOR2_X1 U15304 ( .A(keyinput_204), .B(P3_DATAO_REG_20__SCAN_IN), .ZN(n13588) );
  XOR2_X1 U15305 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .Z(n13587)
         );
  AOI21_X1 U15306 ( .B1(n13589), .B2(n13588), .A(n13587), .ZN(n13593) );
  XOR2_X1 U15307 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .Z(n13592)
         );
  XNOR2_X1 U15308 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n13591) );
  XNOR2_X1 U15309 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n13590) );
  NOR4_X1 U15310 ( .A1(n13593), .A2(n13592), .A3(n13591), .A4(n13590), .ZN(
        n13597) );
  XOR2_X1 U15311 ( .A(keyinput_210), .B(P3_DATAO_REG_14__SCAN_IN), .Z(n13596)
         );
  XNOR2_X1 U15312 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n13595) );
  XNOR2_X1 U15313 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n13594) );
  NOR4_X1 U15314 ( .A1(n13597), .A2(n13596), .A3(n13595), .A4(n13594), .ZN(
        n13600) );
  XOR2_X1 U15315 ( .A(keyinput_213), .B(P3_DATAO_REG_11__SCAN_IN), .Z(n13599)
         );
  XNOR2_X1 U15316 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n13598) );
  NOR3_X1 U15317 ( .A1(n13600), .A2(n13599), .A3(n13598), .ZN(n13603) );
  XOR2_X1 U15318 ( .A(keyinput_214), .B(P3_DATAO_REG_10__SCAN_IN), .Z(n13602)
         );
  XOR2_X1 U15319 ( .A(keyinput_215), .B(P3_DATAO_REG_9__SCAN_IN), .Z(n13601)
         );
  NOR3_X1 U15320 ( .A1(n13603), .A2(n13602), .A3(n13601), .ZN(n13606) );
  INV_X1 U15321 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n13822) );
  XNOR2_X1 U15322 ( .A(n13822), .B(keyinput_216), .ZN(n13605) );
  INV_X1 U15323 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n13825) );
  XNOR2_X1 U15324 ( .A(n13825), .B(keyinput_217), .ZN(n13604) );
  OAI21_X1 U15325 ( .B1(n13606), .B2(n13605), .A(n13604), .ZN(n13610) );
  INV_X1 U15326 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n13827) );
  XNOR2_X1 U15327 ( .A(n13827), .B(keyinput_218), .ZN(n13609) );
  XOR2_X1 U15328 ( .A(keyinput_219), .B(P3_DATAO_REG_5__SCAN_IN), .Z(n13608)
         );
  XOR2_X1 U15329 ( .A(keyinput_220), .B(P3_DATAO_REG_4__SCAN_IN), .Z(n13607)
         );
  AOI211_X1 U15330 ( .C1(n13610), .C2(n13609), .A(n13608), .B(n13607), .ZN(
        n13614) );
  XNOR2_X1 U15331 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_221), .ZN(n13613)
         );
  XNOR2_X1 U15332 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_223), .ZN(n13612)
         );
  XNOR2_X1 U15333 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_222), .ZN(n13611)
         );
  NOR4_X1 U15334 ( .A1(n13614), .A2(n13613), .A3(n13612), .A4(n13611), .ZN(
        n13623) );
  XOR2_X1 U15335 ( .A(keyinput_224), .B(P3_DATAO_REG_0__SCAN_IN), .Z(n13622)
         );
  AOI22_X1 U15336 ( .A1(n8038), .A2(keyinput_228), .B1(keyinput_225), .B2(
        n15730), .ZN(n13615) );
  OAI221_X1 U15337 ( .B1(n8038), .B2(keyinput_228), .C1(n15730), .C2(
        keyinput_225), .A(n13615), .ZN(n13620) );
  AOI22_X1 U15338 ( .A1(n15733), .A2(keyinput_226), .B1(n13617), .B2(
        keyinput_227), .ZN(n13616) );
  OAI221_X1 U15339 ( .B1(n15733), .B2(keyinput_226), .C1(n13617), .C2(
        keyinput_227), .A(n13616), .ZN(n13619) );
  XNOR2_X1 U15340 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_229), .ZN(n13618)
         );
  NOR3_X1 U15341 ( .A1(n13620), .A2(n13619), .A3(n13618), .ZN(n13621) );
  OAI21_X1 U15342 ( .B1(n13623), .B2(n13622), .A(n13621), .ZN(n13630) );
  XOR2_X1 U15343 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_231), .Z(n13629) );
  XOR2_X1 U15344 ( .A(keyinput_230), .B(P3_ADDR_REG_5__SCAN_IN), .Z(n13626) );
  XOR2_X1 U15345 ( .A(keyinput_234), .B(P3_ADDR_REG_9__SCAN_IN), .Z(n13625) );
  XNOR2_X1 U15346 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_233), .ZN(n13624)
         );
  NOR3_X1 U15347 ( .A1(n13626), .A2(n13625), .A3(n13624), .ZN(n13628) );
  XNOR2_X1 U15348 ( .A(keyinput_232), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n13627)
         );
  NAND4_X1 U15349 ( .A1(n13630), .A2(n13629), .A3(n13628), .A4(n13627), .ZN(
        n13634) );
  XOR2_X1 U15350 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_235), .Z(n13633) );
  XOR2_X1 U15351 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_236), .Z(n13632) );
  XOR2_X1 U15352 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_237), .Z(n13631) );
  NAND4_X1 U15353 ( .A1(n13634), .A2(n13633), .A3(n13632), .A4(n13631), .ZN(
        n13637) );
  XOR2_X1 U15354 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_238), .Z(n13636) );
  XNOR2_X1 U15355 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .ZN(n13635) );
  AOI21_X1 U15356 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n13640) );
  XOR2_X1 U15357 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_240), .Z(n13639) );
  XNOR2_X1 U15358 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_241), .ZN(n13638) );
  NOR3_X1 U15359 ( .A1(n13640), .A2(n13639), .A3(n13638), .ZN(n13643) );
  XOR2_X1 U15360 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_243), .Z(n13642) );
  XOR2_X1 U15361 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_242), .Z(n13641) );
  NOR3_X1 U15362 ( .A1(n13643), .A2(n13642), .A3(n13641), .ZN(n13652) );
  INV_X1 U15363 ( .A(keyinput_247), .ZN(n13644) );
  XNOR2_X1 U15364 ( .A(n13644), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13648) );
  XNOR2_X1 U15365 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_246), .ZN(n13647)
         );
  XNOR2_X1 U15366 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_244), .ZN(n13646) );
  XNOR2_X1 U15367 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_245), .ZN(n13645)
         );
  NAND4_X1 U15368 ( .A1(n13648), .A2(n13647), .A3(n13646), .A4(n13645), .ZN(
        n13651) );
  XNOR2_X1 U15369 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_249), .ZN(n13650)
         );
  XNOR2_X1 U15370 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_248), .ZN(n13649)
         );
  OAI211_X1 U15371 ( .C1(n13652), .C2(n13651), .A(n13650), .B(n13649), .ZN(
        n13654) );
  XNOR2_X1 U15372 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_250), .ZN(n13653)
         );
  AND2_X1 U15373 ( .A1(n13654), .A2(n13653), .ZN(n13892) );
  XOR2_X1 U15374 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_251), .Z(n13891) );
  OAI22_X1 U15375 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(keyinput_100), .B1(
        P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_98), .ZN(n13655) );
  AOI221_X1 U15376 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_100), .C1(
        keyinput_98), .C2(P3_ADDR_REG_1__SCAN_IN), .A(n13655), .ZN(n13658) );
  OAI22_X1 U15377 ( .A1(n8036), .A2(keyinput_101), .B1(P3_ADDR_REG_2__SCAN_IN), 
        .B2(keyinput_99), .ZN(n13656) );
  AOI221_X1 U15378 ( .B1(n8036), .B2(keyinput_101), .C1(keyinput_99), .C2(
        P3_ADDR_REG_2__SCAN_IN), .A(n13656), .ZN(n13657) );
  OAI211_X1 U15379 ( .C1(P3_ADDR_REG_0__SCAN_IN), .C2(keyinput_97), .A(n13658), 
        .B(n13657), .ZN(n13659) );
  AOI21_X1 U15380 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(keyinput_97), .A(n13659), 
        .ZN(n13845) );
  INV_X1 U15381 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n13838) );
  INV_X1 U15382 ( .A(keyinput_96), .ZN(n13837) );
  INV_X1 U15383 ( .A(keyinput_90), .ZN(n13826) );
  INV_X1 U15384 ( .A(keyinput_89), .ZN(n13824) );
  INV_X1 U15385 ( .A(keyinput_88), .ZN(n13823) );
  INV_X1 U15386 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n13661) );
  OAI22_X1 U15387 ( .A1(n13661), .A2(keyinput_85), .B1(
        P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_84), .ZN(n13660) );
  AOI221_X1 U15388 ( .B1(n13661), .B2(keyinput_85), .C1(keyinput_84), .C2(
        P3_DATAO_REG_12__SCAN_IN), .A(n13660), .ZN(n13821) );
  XNOR2_X1 U15389 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n13809)
         );
  XOR2_X1 U15390 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .Z(n13787)
         );
  XNOR2_X1 U15391 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n13766)
         );
  INV_X1 U15392 ( .A(keyinput_50), .ZN(n13749) );
  INV_X1 U15393 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n13663) );
  OAI22_X1 U15394 ( .A1(n13664), .A2(keyinput_42), .B1(n13663), .B2(
        keyinput_41), .ZN(n13662) );
  AOI221_X1 U15395 ( .B1(n13664), .B2(keyinput_42), .C1(keyinput_41), .C2(
        n13663), .A(n13662), .ZN(n13743) );
  INV_X1 U15396 ( .A(keyinput_40), .ZN(n13735) );
  AOI22_X1 U15397 ( .A1(n7656), .A2(keyinput_28), .B1(n13666), .B2(keyinput_27), .ZN(n13665) );
  OAI221_X1 U15398 ( .B1(n7656), .B2(keyinput_28), .C1(n13666), .C2(
        keyinput_27), .A(n13665), .ZN(n13713) );
  INV_X1 U15399 ( .A(keyinput_19), .ZN(n13696) );
  AOI22_X1 U15400 ( .A1(SI_18_), .A2(keyinput_14), .B1(n13668), .B2(
        keyinput_12), .ZN(n13667) );
  OAI221_X1 U15401 ( .B1(SI_18_), .B2(keyinput_14), .C1(n13668), .C2(
        keyinput_12), .A(n13667), .ZN(n13689) );
  INV_X1 U15402 ( .A(keyinput_6), .ZN(n13678) );
  AOI22_X1 U15403 ( .A1(SI_28_), .A2(keyinput_4), .B1(SI_29_), .B2(keyinput_3), 
        .ZN(n13669) );
  OAI221_X1 U15404 ( .B1(SI_28_), .B2(keyinput_4), .C1(SI_29_), .C2(keyinput_3), .A(n13669), .ZN(n13675) );
  INV_X1 U15405 ( .A(keyinput_2), .ZN(n13672) );
  OAI221_X1 U15406 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n13670), .ZN(n13671) );
  AOI221_X1 U15407 ( .B1(SI_30_), .B2(keyinput_2), .C1(n13673), .C2(n13672), 
        .A(n13671), .ZN(n13674) );
  OAI22_X1 U15408 ( .A1(n13675), .A2(n13674), .B1(keyinput_5), .B2(SI_27_), 
        .ZN(n13676) );
  AOI22_X1 U15409 ( .A1(n13681), .A2(keyinput_8), .B1(n13680), .B2(keyinput_7), 
        .ZN(n13679) );
  OAI221_X1 U15410 ( .B1(n13681), .B2(keyinput_8), .C1(n13680), .C2(keyinput_7), .A(n13679), .ZN(n13682) );
  OAI22_X1 U15411 ( .A1(SI_22_), .A2(keyinput_10), .B1(keyinput_11), .B2(
        SI_21_), .ZN(n13683) );
  AOI221_X1 U15412 ( .B1(SI_22_), .B2(keyinput_10), .C1(SI_21_), .C2(
        keyinput_11), .A(n13683), .ZN(n13685) );
  AOI21_X1 U15413 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(n13687) );
  INV_X1 U15414 ( .A(n13687), .ZN(n13688) );
  OAI22_X1 U15415 ( .A1(n13692), .A2(keyinput_17), .B1(keyinput_16), .B2(
        SI_16_), .ZN(n13691) );
  AOI221_X1 U15416 ( .B1(n13692), .B2(keyinput_17), .C1(SI_16_), .C2(
        keyinput_16), .A(n13691), .ZN(n13693) );
  OAI21_X1 U15417 ( .B1(keyinput_18), .B2(SI_14_), .A(n13693), .ZN(n13694) );
  AOI22_X1 U15418 ( .A1(n13699), .A2(keyinput_20), .B1(keyinput_21), .B2(
        n13698), .ZN(n13697) );
  OAI221_X1 U15419 ( .B1(n13699), .B2(keyinput_20), .C1(n13698), .C2(
        keyinput_21), .A(n13697), .ZN(n13700) );
  XNOR2_X1 U15420 ( .A(n13702), .B(keyinput_22), .ZN(n13704) );
  XNOR2_X1 U15421 ( .A(SI_9_), .B(keyinput_23), .ZN(n13703) );
  INV_X1 U15422 ( .A(keyinput_25), .ZN(n13708) );
  XNOR2_X1 U15423 ( .A(SI_6_), .B(keyinput_26), .ZN(n13707) );
  XNOR2_X1 U15424 ( .A(n13705), .B(keyinput_24), .ZN(n13706) );
  AOI211_X1 U15425 ( .C1(SI_7_), .C2(n13708), .A(n13707), .B(n13706), .ZN(
        n13709) );
  NAND2_X1 U15426 ( .A1(keyinput_30), .A2(SI_2_), .ZN(n13712) );
  AOI22_X1 U15427 ( .A1(SI_1_), .A2(keyinput_31), .B1(n13715), .B2(keyinput_29), .ZN(n13714) );
  OAI221_X1 U15428 ( .B1(SI_1_), .B2(keyinput_31), .C1(n13715), .C2(
        keyinput_29), .A(n13714), .ZN(n13716) );
  OAI22_X1 U15429 ( .A1(P3_U3151), .A2(keyinput_34), .B1(n13718), .B2(
        keyinput_32), .ZN(n13717) );
  AOI221_X1 U15430 ( .B1(P3_U3151), .B2(keyinput_34), .C1(keyinput_32), .C2(
        n13718), .A(n13717), .ZN(n13721) );
  OAI22_X1 U15431 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_35), .B1(
        keyinput_33), .B2(P3_RD_REG_SCAN_IN), .ZN(n13719) );
  AOI221_X1 U15432 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(
        P3_RD_REG_SCAN_IN), .C2(keyinput_33), .A(n13719), .ZN(n13720) );
  INV_X1 U15433 ( .A(keyinput_36), .ZN(n13722) );
  OAI22_X1 U15434 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_38), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .ZN(n13728) );
  AOI221_X1 U15435 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        keyinput_37), .C2(P3_REG3_REG_14__SCAN_IN), .A(n13728), .ZN(n13730) );
  AOI21_X1 U15436 ( .B1(n13731), .B2(n13730), .A(n13729), .ZN(n13732) );
  INV_X1 U15437 ( .A(n13732), .ZN(n13733) );
  AOI22_X1 U15438 ( .A1(n13738), .A2(keyinput_46), .B1(keyinput_43), .B2(
        n13737), .ZN(n13736) );
  OAI221_X1 U15439 ( .B1(n13738), .B2(keyinput_46), .C1(n13737), .C2(
        keyinput_43), .A(n13736), .ZN(n13742) );
  AOI22_X1 U15440 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_44), .B1(n13740), 
        .B2(keyinput_45), .ZN(n13739) );
  OAI221_X1 U15441 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(n13740), .C2(keyinput_45), .A(n13739), .ZN(n13741) );
  AOI22_X1 U15442 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_48), .B1(n13745), .B2(keyinput_49), .ZN(n13744) );
  OAI221_X1 U15443 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .C1(
        n13745), .C2(keyinput_49), .A(n13744), .ZN(n13746) );
  OAI221_X1 U15444 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(n13749), .C1(n13748), 
        .C2(keyinput_50), .A(n13747), .ZN(n13754) );
  INV_X1 U15445 ( .A(keyinput_51), .ZN(n13750) );
  INV_X1 U15446 ( .A(n13752), .ZN(n13753) );
  INV_X1 U15447 ( .A(keyinput_52), .ZN(n13755) );
  AOI22_X1 U15448 ( .A1(n13761), .A2(keyinput_57), .B1(keyinput_56), .B2(
        n13555), .ZN(n13760) );
  OAI221_X1 U15449 ( .B1(n13761), .B2(keyinput_57), .C1(n13555), .C2(
        keyinput_56), .A(n13760), .ZN(n13764) );
  AOI22_X1 U15450 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput_55), .B1(n15904), .B2(keyinput_54), .ZN(n13762) );
  OAI221_X1 U15451 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        n15904), .C2(keyinput_54), .A(n13762), .ZN(n13763) );
  AOI211_X1 U15452 ( .C1(n13766), .C2(n13765), .A(n13764), .B(n13763), .ZN(
        n13769) );
  AOI22_X1 U15453 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .ZN(n13767) );
  OAI221_X1 U15454 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_58), .A(n13767), .ZN(n13768) );
  OAI22_X1 U15455 ( .A1(n13769), .A2(n13768), .B1(keyinput_60), .B2(
        P3_REG3_REG_18__SCAN_IN), .ZN(n13770) );
  AOI21_X1 U15456 ( .B1(keyinput_60), .B2(P3_REG3_REG_18__SCAN_IN), .A(n13770), 
        .ZN(n13785) );
  AOI22_X1 U15457 ( .A1(n13773), .A2(keyinput_65), .B1(n13772), .B2(
        keyinput_62), .ZN(n13771) );
  OAI221_X1 U15458 ( .B1(n13773), .B2(keyinput_65), .C1(n13772), .C2(
        keyinput_62), .A(n13771), .ZN(n13777) );
  AOI22_X1 U15459 ( .A1(P3_B_REG_SCAN_IN), .A2(keyinput_64), .B1(n13775), .B2(
        keyinput_63), .ZN(n13774) );
  OAI221_X1 U15460 ( .B1(P3_B_REG_SCAN_IN), .B2(keyinput_64), .C1(n13775), 
        .C2(keyinput_63), .A(n13774), .ZN(n13776) );
  AOI211_X1 U15461 ( .C1(keyinput_61), .C2(P3_REG3_REG_6__SCAN_IN), .A(n13777), 
        .B(n13776), .ZN(n13778) );
  OAI21_X1 U15462 ( .B1(keyinput_61), .B2(P3_REG3_REG_6__SCAN_IN), .A(n13778), 
        .ZN(n13784) );
  OAI22_X1 U15463 ( .A1(n13780), .A2(keyinput_68), .B1(
        P3_DATAO_REG_29__SCAN_IN), .B2(keyinput_67), .ZN(n13779) );
  AOI221_X1 U15464 ( .B1(n13780), .B2(keyinput_68), .C1(keyinput_67), .C2(
        P3_DATAO_REG_29__SCAN_IN), .A(n13779), .ZN(n13783) );
  OAI22_X1 U15465 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(keyinput_69), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(keyinput_66), .ZN(n13781) );
  AOI221_X1 U15466 ( .B1(P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_69), .C1(
        keyinput_66), .C2(P3_DATAO_REG_30__SCAN_IN), .A(n13781), .ZN(n13782)
         );
  OAI211_X1 U15467 ( .C1(n13785), .C2(n13784), .A(n13783), .B(n13782), .ZN(
        n13786) );
  AOI22_X1 U15468 ( .A1(keyinput_71), .A2(P3_DATAO_REG_25__SCAN_IN), .B1(
        n13787), .B2(n13786), .ZN(n13794) );
  INV_X1 U15469 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n13789) );
  INV_X1 U15470 ( .A(keyinput_71), .ZN(n13788) );
  NAND2_X1 U15471 ( .A1(n13789), .A2(n13788), .ZN(n13793) );
  INV_X1 U15472 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n13791) );
  AOI22_X1 U15473 ( .A1(P3_DATAO_REG_24__SCAN_IN), .A2(keyinput_72), .B1(
        n13791), .B2(keyinput_73), .ZN(n13790) );
  OAI221_X1 U15474 ( .B1(P3_DATAO_REG_24__SCAN_IN), .B2(keyinput_72), .C1(
        n13791), .C2(keyinput_73), .A(n13790), .ZN(n13792) );
  INV_X1 U15475 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n13796) );
  AOI22_X1 U15476 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_75), .B1(
        n13796), .B2(keyinput_74), .ZN(n13795) );
  OAI221_X1 U15477 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_75), .C1(
        n13796), .C2(keyinput_74), .A(n13795), .ZN(n13802) );
  INV_X1 U15478 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n13798) );
  NAND2_X1 U15479 ( .A1(P3_DATAO_REG_20__SCAN_IN), .A2(keyinput_76), .ZN(
        n13799) );
  XOR2_X1 U15480 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n13807)
         );
  AOI22_X1 U15481 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput_79), .B1(
        n13805), .B2(keyinput_80), .ZN(n13804) );
  OAI221_X1 U15482 ( .B1(P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_79), .C1(
        n13805), .C2(keyinput_80), .A(n13804), .ZN(n13806) );
  AOI211_X1 U15483 ( .C1(n13809), .C2(n13808), .A(n13807), .B(n13806), .ZN(
        n13810) );
  INV_X1 U15484 ( .A(n13810), .ZN(n13816) );
  AOI22_X1 U15485 ( .A1(keyinput_82), .A2(P3_DATAO_REG_14__SCAN_IN), .B1(
        n13812), .B2(keyinput_83), .ZN(n13811) );
  OAI221_X1 U15486 ( .B1(keyinput_82), .B2(P3_DATAO_REG_14__SCAN_IN), .C1(
        n13812), .C2(keyinput_83), .A(n13811), .ZN(n13814) );
  NAND2_X1 U15487 ( .A1(n13816), .A2(n13815), .ZN(n13820) );
  INV_X1 U15488 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n13818) );
  AOI22_X1 U15489 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput_87), .B1(n13818), .B2(keyinput_86), .ZN(n13817) );
  OAI221_X1 U15490 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_87), .C1(
        n13818), .C2(keyinput_86), .A(n13817), .ZN(n13819) );
  AOI22_X1 U15491 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput_92), .B1(
        P3_DATAO_REG_5__SCAN_IN), .B2(keyinput_91), .ZN(n13828) );
  OAI221_X1 U15492 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput_92), .C1(
        P3_DATAO_REG_5__SCAN_IN), .C2(keyinput_91), .A(n13828), .ZN(n13834) );
  OAI22_X1 U15493 ( .A1(n13831), .A2(keyinput_94), .B1(n13830), .B2(
        keyinput_95), .ZN(n13829) );
  AOI221_X1 U15494 ( .B1(n13831), .B2(keyinput_94), .C1(keyinput_95), .C2(
        n13830), .A(n13829), .ZN(n13833) );
  XNOR2_X1 U15495 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n13832)
         );
  OAI211_X1 U15496 ( .C1(n13835), .C2(n13834), .A(n13833), .B(n13832), .ZN(
        n13836) );
  OAI221_X1 U15497 ( .B1(keyinput_96), .B2(n13838), .C1(n13837), .C2(
        P3_DATAO_REG_0__SCAN_IN), .A(n13836), .ZN(n13844) );
  AOI22_X1 U15498 ( .A1(n15982), .A2(keyinput_103), .B1(n15806), .B2(
        keyinput_106), .ZN(n13839) );
  OAI221_X1 U15499 ( .B1(n15982), .B2(keyinput_103), .C1(n15806), .C2(
        keyinput_106), .A(n13839), .ZN(n13843) );
  INV_X1 U15500 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U15501 ( .A1(n15772), .A2(keyinput_102), .B1(n13841), .B2(
        keyinput_104), .ZN(n13840) );
  OAI221_X1 U15502 ( .B1(n15772), .B2(keyinput_102), .C1(n13841), .C2(
        keyinput_104), .A(n13840), .ZN(n13842) );
  AOI211_X1 U15503 ( .C1(n13845), .C2(n13844), .A(n13843), .B(n13842), .ZN(
        n13851) );
  INV_X1 U15504 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15796) );
  XNOR2_X1 U15505 ( .A(keyinput_105), .B(n15796), .ZN(n13850) );
  XOR2_X1 U15506 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_108), .Z(n13849) );
  XOR2_X1 U15507 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_109), .Z(n13847) );
  XNOR2_X1 U15508 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_107), .ZN(n13846) );
  NAND2_X1 U15509 ( .A1(n13847), .A2(n13846), .ZN(n13848) );
  XOR2_X1 U15510 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_110), .Z(n13853) );
  XOR2_X1 U15511 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_111), .Z(n13852) );
  OAI21_X1 U15512 ( .B1(n13854), .B2(n13853), .A(n13852), .ZN(n13860) );
  INV_X1 U15513 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n13856) );
  OAI22_X1 U15514 ( .A1(n13856), .A2(keyinput_113), .B1(P1_IR_REG_5__SCAN_IN), 
        .B2(keyinput_112), .ZN(n13855) );
  AOI221_X1 U15515 ( .B1(n13856), .B2(keyinput_113), .C1(keyinput_112), .C2(
        P1_IR_REG_5__SCAN_IN), .A(n13855), .ZN(n13859) );
  XOR2_X1 U15516 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_114), .Z(n13858) );
  XNOR2_X1 U15517 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_115), .ZN(n13857) );
  AOI211_X1 U15518 ( .C1(n13860), .C2(n13859), .A(n13858), .B(n13857), .ZN(
        n13866) );
  AOI22_X1 U15519 ( .A1(n13862), .A2(keyinput_118), .B1(n9289), .B2(
        keyinput_119), .ZN(n13861) );
  OAI221_X1 U15520 ( .B1(n13862), .B2(keyinput_118), .C1(n9289), .C2(
        keyinput_119), .A(n13861), .ZN(n13865) );
  XOR2_X1 U15521 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_116), .Z(n13864) );
  XOR2_X1 U15522 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_117), .Z(n13863) );
  OR4_X1 U15523 ( .A1(n13866), .A2(n13865), .A3(n13864), .A4(n13863), .ZN(
        n13874) );
  AOI22_X1 U15524 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_121), .B1(n13868), 
        .B2(keyinput_120), .ZN(n13867) );
  OAI221_X1 U15525 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_121), .C1(n13868), .C2(keyinput_120), .A(n13867), .ZN(n13869) );
  INV_X1 U15526 ( .A(n13869), .ZN(n13873) );
  NAND2_X1 U15527 ( .A1(n13871), .A2(keyinput_122), .ZN(n13870) );
  OAI21_X1 U15528 ( .B1(n13871), .B2(keyinput_122), .A(n13870), .ZN(n13872) );
  AOI21_X1 U15529 ( .B1(n13874), .B2(n13873), .A(n13872), .ZN(n13884) );
  XOR2_X1 U15530 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_123), .Z(n13883) );
  INV_X1 U15531 ( .A(keyinput_127), .ZN(n13881) );
  OAI22_X1 U15532 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_126), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_125), .ZN(n13880) );
  AOI22_X1 U15533 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_125), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_126), .ZN(n13877) );
  AOI22_X1 U15534 ( .A1(n13875), .A2(keyinput_127), .B1(keyinput_124), .B2(
        n13878), .ZN(n13876) );
  OAI211_X1 U15535 ( .C1(n13878), .C2(keyinput_124), .A(n13877), .B(n13876), 
        .ZN(n13879) );
  AOI211_X1 U15536 ( .C1(P1_IR_REG_20__SCAN_IN), .C2(n13881), .A(n13880), .B(
        n13879), .ZN(n13882) );
  XNOR2_X1 U15537 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_254), .ZN(n13888)
         );
  XNOR2_X1 U15538 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_253), .ZN(n13887)
         );
  XNOR2_X1 U15539 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_252), .ZN(n13886)
         );
  XNOR2_X1 U15540 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n13885)
         );
  NOR4_X1 U15541 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n13889) );
  OAI211_X1 U15542 ( .C1(n13892), .C2(n13891), .A(n13890), .B(n13889), .ZN(
        n13895) );
  MUX2_X1 U15543 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n13893), .S(P3_U3897), .Z(
        n13894) );
  XNOR2_X1 U15544 ( .A(n13895), .B(n13894), .ZN(P3_U3491) );
  INV_X1 U15545 ( .A(n13896), .ZN(n13897) );
  AOI21_X1 U15546 ( .B1(n13899), .B2(n13898), .A(n13897), .ZN(n13916) );
  XNOR2_X1 U15547 ( .A(n13901), .B(n13900), .ZN(n13914) );
  NAND2_X1 U15548 ( .A1(n13902), .A2(n16052), .ZN(n13912) );
  AOI21_X1 U15549 ( .B1(n13905), .B2(n13904), .A(n13903), .ZN(n13911) );
  INV_X1 U15550 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n13906) );
  NOR2_X1 U15551 ( .A1(n15981), .A2(n13906), .ZN(n13907) );
  AOI211_X1 U15552 ( .C1(n16043), .C2(n13909), .A(n13908), .B(n13907), .ZN(
        n13910) );
  OAI21_X1 U15553 ( .B1(n13912), .B2(n13911), .A(n13910), .ZN(n13913) );
  AOI21_X1 U15554 ( .B1(n13914), .B2(n16079), .A(n13913), .ZN(n13915) );
  OAI21_X1 U15555 ( .B1(n13916), .B2(n16082), .A(n13915), .ZN(P3_U3196) );
  AOI21_X1 U15556 ( .B1(n13919), .B2(n13918), .A(n13917), .ZN(n13933) );
  OAI21_X1 U15557 ( .B1(n13922), .B2(n13921), .A(n13920), .ZN(n13931) );
  OAI21_X1 U15558 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n13924), .A(n13923), 
        .ZN(n13925) );
  NAND2_X1 U15559 ( .A1(n13925), .A2(n16079), .ZN(n13928) );
  AOI21_X1 U15560 ( .B1(n16073), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13926), 
        .ZN(n13927) );
  OAI211_X1 U15561 ( .C1(n16076), .C2(n13929), .A(n13928), .B(n13927), .ZN(
        n13930) );
  AOI21_X1 U15562 ( .B1(n16052), .B2(n13931), .A(n13930), .ZN(n13932) );
  OAI21_X1 U15563 ( .B1(n13933), .B2(n16082), .A(n13932), .ZN(P3_U3197) );
  AND3_X1 U15564 ( .A1(n16061), .A2(n13935), .A3(n13934), .ZN(n13936) );
  OAI21_X1 U15565 ( .B1(n13937), .B2(n13936), .A(n16054), .ZN(n13953) );
  OAI21_X1 U15566 ( .B1(n13940), .B2(n13939), .A(n13938), .ZN(n13951) );
  NAND2_X1 U15567 ( .A1(n16073), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13941) );
  OAI211_X1 U15568 ( .C1(n16076), .C2(n13943), .A(n13942), .B(n13941), .ZN(
        n13950) );
  INV_X1 U15569 ( .A(n13944), .ZN(n13945) );
  NAND3_X1 U15570 ( .A1(n13946), .A2(n16065), .A3(n13945), .ZN(n13947) );
  AOI21_X1 U15571 ( .B1(n13948), .B2(n13947), .A(n15969), .ZN(n13949) );
  AOI211_X1 U15572 ( .C1(n16052), .C2(n13951), .A(n13950), .B(n13949), .ZN(
        n13952) );
  NAND2_X1 U15573 ( .A1(n13953), .A2(n13952), .ZN(P3_U3200) );
  NAND2_X1 U15574 ( .A1(n13961), .A2(n14163), .ZN(n13956) );
  NAND2_X1 U15575 ( .A1(n13955), .A2(n13954), .ZN(n16561) );
  NAND3_X1 U15576 ( .A1(n14169), .A2(n13956), .A3(n16561), .ZN(n13958) );
  OAI21_X1 U15577 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n14169), .A(n13958), 
        .ZN(n13957) );
  OAI21_X1 U15578 ( .B1(n14173), .B2(n14166), .A(n13957), .ZN(P3_U3202) );
  OAI21_X1 U15579 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n14169), .A(n13958), 
        .ZN(n13959) );
  OAI21_X1 U15580 ( .B1(n14176), .B2(n14166), .A(n13959), .ZN(P3_U3203) );
  INV_X1 U15581 ( .A(n13960), .ZN(n13967) );
  AOI22_X1 U15582 ( .A1(n13961), .A2(n14163), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n14164), .ZN(n13962) );
  OAI21_X1 U15583 ( .B1(n13963), .B2(n14166), .A(n13962), .ZN(n13964) );
  AOI21_X1 U15584 ( .B1(n13965), .B2(n14100), .A(n13964), .ZN(n13966) );
  OAI21_X1 U15585 ( .B1(n13967), .B2(n14164), .A(n13966), .ZN(P3_U3204) );
  NAND2_X1 U15586 ( .A1(n13969), .A2(n13968), .ZN(n13970) );
  NAND2_X1 U15587 ( .A1(n13970), .A2(n13977), .ZN(n13971) );
  NAND2_X1 U15588 ( .A1(n13971), .A2(n16183), .ZN(n13972) );
  OAI22_X1 U15589 ( .A1(n13999), .A2(n14161), .B1(n13974), .B2(n14159), .ZN(
        n13975) );
  INV_X1 U15590 ( .A(n13975), .ZN(n13976) );
  INV_X1 U15591 ( .A(n14179), .ZN(n13985) );
  OR2_X1 U15592 ( .A1(n13978), .A2(n13977), .ZN(n13979) );
  NAND2_X1 U15593 ( .A1(n13980), .A2(n13979), .ZN(n14177) );
  AOI22_X1 U15594 ( .A1(n13981), .A2(n14163), .B1(n14164), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13982) );
  OAI21_X1 U15595 ( .B1(n14247), .B2(n14166), .A(n13982), .ZN(n13983) );
  AOI21_X1 U15596 ( .B1(n14177), .B2(n14100), .A(n13983), .ZN(n13984) );
  OAI21_X1 U15597 ( .B1(n13985), .B2(n14164), .A(n13984), .ZN(P3_U3205) );
  MUX2_X1 U15598 ( .A(n14248), .B(P3_REG2_REG_27__SCAN_IN), .S(n14164), .Z(
        n13990) );
  AOI22_X1 U15599 ( .A1(n13987), .A2(n14097), .B1(n14163), .B2(n13986), .ZN(
        n13988) );
  OAI21_X1 U15600 ( .B1(n14250), .B2(n14082), .A(n13988), .ZN(n13989) );
  NAND2_X1 U15601 ( .A1(n14017), .A2(n13992), .ZN(n13994) );
  NAND2_X1 U15602 ( .A1(n13994), .A2(n13993), .ZN(n13995) );
  NAND2_X1 U15603 ( .A1(n14006), .A2(n13996), .ZN(n13998) );
  XNOR2_X1 U15604 ( .A(n13998), .B(n13997), .ZN(n14001) );
  OAI22_X1 U15605 ( .A1(n13999), .A2(n14159), .B1(n14027), .B2(n14161), .ZN(
        n14000) );
  MUX2_X1 U15606 ( .A(n14002), .B(n14253), .S(n14169), .Z(n14005) );
  AOI22_X1 U15607 ( .A1(n14255), .A2(n14097), .B1(n14163), .B2(n14003), .ZN(
        n14004) );
  OAI211_X1 U15608 ( .C1(n14257), .C2(n14082), .A(n14005), .B(n14004), .ZN(
        P3_U3207) );
  OAI211_X1 U15609 ( .C1(n14008), .C2(n14007), .A(n14006), .B(n16183), .ZN(
        n14013) );
  OAI22_X1 U15610 ( .A1(n14010), .A2(n14159), .B1(n14009), .B2(n14161), .ZN(
        n14011) );
  INV_X1 U15611 ( .A(n14011), .ZN(n14012) );
  OR2_X1 U15612 ( .A1(n14015), .A2(n14014), .ZN(n14016) );
  NAND2_X1 U15613 ( .A1(n14017), .A2(n14016), .ZN(n14185) );
  INV_X1 U15614 ( .A(n14260), .ZN(n14020) );
  AOI22_X1 U15615 ( .A1(n14018), .A2(n14163), .B1(n14164), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n14019) );
  OAI21_X1 U15616 ( .B1(n14020), .B2(n14166), .A(n14019), .ZN(n14021) );
  AOI21_X1 U15617 ( .B1(n14185), .B2(n14100), .A(n14021), .ZN(n14022) );
  OAI21_X1 U15618 ( .B1(n14187), .B2(n14164), .A(n14022), .ZN(P3_U3208) );
  INV_X1 U15619 ( .A(n14023), .ZN(n14024) );
  AOI21_X1 U15620 ( .B1(n14030), .B2(n14025), .A(n14024), .ZN(n14026) );
  OAI222_X1 U15621 ( .A1(n14161), .A2(n14028), .B1(n14159), .B2(n14027), .C1(
        n14156), .C2(n14026), .ZN(n14191) );
  INV_X1 U15622 ( .A(n14191), .ZN(n14035) );
  OAI21_X1 U15623 ( .B1(n8339), .B2(n14030), .A(n14029), .ZN(n14192) );
  AOI22_X1 U15624 ( .A1(n14031), .A2(n14163), .B1(n14164), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n14032) );
  OAI21_X1 U15625 ( .B1(n14265), .B2(n14166), .A(n14032), .ZN(n14033) );
  AOI21_X1 U15626 ( .B1(n14192), .B2(n14100), .A(n14033), .ZN(n14034) );
  OAI21_X1 U15627 ( .B1(n14035), .B2(n14164), .A(n14034), .ZN(P3_U3209) );
  XOR2_X1 U15628 ( .A(n14038), .B(n14036), .Z(n14196) );
  INV_X1 U15629 ( .A(n14196), .ZN(n14049) );
  INV_X1 U15630 ( .A(n14037), .ZN(n14040) );
  OAI211_X1 U15631 ( .C1(n14040), .C2(n8013), .A(n14039), .B(n16183), .ZN(
        n14044) );
  AOI22_X1 U15632 ( .A1(n14042), .A2(n16178), .B1(n16180), .B2(n14041), .ZN(
        n14043) );
  NAND2_X1 U15633 ( .A1(n14044), .A2(n14043), .ZN(n14195) );
  AOI22_X1 U15634 ( .A1(n14164), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n14163), 
        .B2(n14045), .ZN(n14046) );
  OAI21_X1 U15635 ( .B1(n14269), .B2(n14166), .A(n14046), .ZN(n14047) );
  AOI21_X1 U15636 ( .B1(n14195), .B2(n14169), .A(n14047), .ZN(n14048) );
  OAI21_X1 U15637 ( .B1(n14171), .B2(n14049), .A(n14048), .ZN(P3_U3210) );
  NAND2_X1 U15638 ( .A1(n14068), .A2(n14050), .ZN(n14052) );
  NAND2_X1 U15639 ( .A1(n14052), .A2(n14051), .ZN(n14054) );
  NAND2_X1 U15640 ( .A1(n14054), .A2(n14053), .ZN(n14272) );
  AOI22_X1 U15641 ( .A1(n16178), .A2(n14056), .B1(n14055), .B2(n16180), .ZN(
        n14061) );
  XNOR2_X1 U15642 ( .A(n14058), .B(n14057), .ZN(n14059) );
  NAND2_X1 U15643 ( .A1(n14059), .A2(n16183), .ZN(n14060) );
  OAI211_X1 U15644 ( .C1(n14272), .C2(n16188), .A(n14061), .B(n14060), .ZN(
        n14270) );
  MUX2_X1 U15645 ( .A(n14270), .B(P3_REG2_REG_22__SCAN_IN), .S(n14164), .Z(
        n14062) );
  INV_X1 U15646 ( .A(n14062), .ZN(n14065) );
  AOI22_X1 U15647 ( .A1(n14199), .A2(n14097), .B1(n14163), .B2(n14063), .ZN(
        n14064) );
  OAI211_X1 U15648 ( .C1(n14272), .C2(n14082), .A(n14065), .B(n14064), .ZN(
        P3_U3211) );
  NAND2_X1 U15649 ( .A1(n14066), .A2(n14069), .ZN(n14067) );
  NAND2_X1 U15650 ( .A1(n14068), .A2(n14067), .ZN(n14072) );
  INV_X1 U15651 ( .A(n14072), .ZN(n14277) );
  XNOR2_X1 U15652 ( .A(n14070), .B(n7899), .ZN(n14071) );
  NAND2_X1 U15653 ( .A1(n14071), .A2(n16183), .ZN(n14077) );
  NAND2_X1 U15654 ( .A1(n14072), .A2(n16475), .ZN(n14076) );
  OAI22_X1 U15655 ( .A1(n14073), .A2(n14159), .B1(n14109), .B2(n14161), .ZN(
        n14074) );
  INV_X1 U15656 ( .A(n14074), .ZN(n14075) );
  NAND3_X1 U15657 ( .A1(n14077), .A2(n14076), .A3(n14075), .ZN(n14275) );
  MUX2_X1 U15658 ( .A(n14275), .B(P3_REG2_REG_21__SCAN_IN), .S(n14164), .Z(
        n14078) );
  INV_X1 U15659 ( .A(n14078), .ZN(n14081) );
  AOI22_X1 U15660 ( .A1(n14202), .A2(n14097), .B1(n14163), .B2(n14079), .ZN(
        n14080) );
  OAI211_X1 U15661 ( .C1(n14277), .C2(n14082), .A(n14081), .B(n14080), .ZN(
        P3_U3212) );
  NAND2_X1 U15662 ( .A1(n14119), .A2(n14083), .ZN(n14085) );
  AND2_X1 U15663 ( .A1(n14085), .A2(n14084), .ZN(n14086) );
  AOI21_X1 U15664 ( .B1(n14086), .B2(n14098), .A(n14156), .ZN(n14092) );
  AND2_X1 U15665 ( .A1(n14088), .A2(n14087), .ZN(n14091) );
  OAI22_X1 U15666 ( .A1(n14089), .A2(n14159), .B1(n14122), .B2(n14161), .ZN(
        n14090) );
  AOI21_X1 U15667 ( .B1(n14092), .B2(n14091), .A(n14090), .ZN(n14208) );
  INV_X1 U15668 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n14095) );
  INV_X1 U15669 ( .A(n14093), .ZN(n14094) );
  OAI22_X1 U15670 ( .A1(n14169), .A2(n14095), .B1(n14094), .B2(n16194), .ZN(
        n14096) );
  AOI21_X1 U15671 ( .B1(n14205), .B2(n14097), .A(n14096), .ZN(n14102) );
  XNOR2_X1 U15672 ( .A(n14099), .B(n9929), .ZN(n14206) );
  NAND2_X1 U15673 ( .A1(n14206), .A2(n14100), .ZN(n14101) );
  OAI211_X1 U15674 ( .C1(n14208), .C2(n14164), .A(n14102), .B(n14101), .ZN(
        P3_U3213) );
  XOR2_X1 U15675 ( .A(n14106), .B(n14103), .Z(n14212) );
  INV_X1 U15676 ( .A(n14212), .ZN(n14114) );
  NAND2_X1 U15677 ( .A1(n14119), .A2(n14104), .ZN(n14105) );
  XOR2_X1 U15678 ( .A(n14106), .B(n14105), .Z(n14107) );
  OAI222_X1 U15679 ( .A1(n14159), .A2(n14109), .B1(n14161), .B2(n14108), .C1(
        n14156), .C2(n14107), .ZN(n14211) );
  AOI22_X1 U15680 ( .A1(n14164), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14163), 
        .B2(n14110), .ZN(n14111) );
  OAI21_X1 U15681 ( .B1(n14287), .B2(n14166), .A(n14111), .ZN(n14112) );
  AOI21_X1 U15682 ( .B1(n14211), .B2(n14169), .A(n14112), .ZN(n14113) );
  OAI21_X1 U15683 ( .B1(n14171), .B2(n14114), .A(n14113), .ZN(P3_U3214) );
  XNOR2_X1 U15684 ( .A(n14115), .B(n14116), .ZN(n14216) );
  INV_X1 U15685 ( .A(n14216), .ZN(n14127) );
  INV_X1 U15686 ( .A(n14129), .ZN(n14118) );
  OAI21_X1 U15687 ( .B1(n14118), .B2(n14117), .A(n14116), .ZN(n14120) );
  AND2_X1 U15688 ( .A1(n14120), .A2(n14119), .ZN(n14121) );
  OAI222_X1 U15689 ( .A1(n14159), .A2(n14122), .B1(n14161), .B2(n14147), .C1(
        n14156), .C2(n14121), .ZN(n14215) );
  AOI22_X1 U15690 ( .A1(n14164), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n14163), 
        .B2(n14123), .ZN(n14124) );
  OAI21_X1 U15691 ( .B1(n14291), .B2(n14166), .A(n14124), .ZN(n14125) );
  AOI21_X1 U15692 ( .B1(n14215), .B2(n14169), .A(n14125), .ZN(n14126) );
  OAI21_X1 U15693 ( .B1(n14171), .B2(n14127), .A(n14126), .ZN(P3_U3215) );
  XNOR2_X1 U15694 ( .A(n14128), .B(n14130), .ZN(n14222) );
  OAI211_X1 U15695 ( .C1(n7500), .C2(n14130), .A(n14129), .B(n16183), .ZN(
        n14134) );
  AOI22_X1 U15696 ( .A1(n14132), .A2(n16178), .B1(n16180), .B2(n14131), .ZN(
        n14133) );
  NAND2_X1 U15697 ( .A1(n14134), .A2(n14133), .ZN(n14219) );
  INV_X1 U15698 ( .A(n14220), .ZN(n14137) );
  AOI22_X1 U15699 ( .A1(n14164), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n14163), 
        .B2(n14135), .ZN(n14136) );
  OAI21_X1 U15700 ( .B1(n14137), .B2(n14166), .A(n14136), .ZN(n14138) );
  AOI21_X1 U15701 ( .B1(n14219), .B2(n14169), .A(n14138), .ZN(n14139) );
  OAI21_X1 U15702 ( .B1(n14171), .B2(n14222), .A(n14139), .ZN(P3_U3216) );
  XNOR2_X1 U15703 ( .A(n14140), .B(n14144), .ZN(n14224) );
  INV_X1 U15704 ( .A(n14224), .ZN(n14152) );
  INV_X1 U15705 ( .A(n14141), .ZN(n14142) );
  AOI21_X1 U15706 ( .B1(n14144), .B2(n14143), .A(n14142), .ZN(n14145) );
  OAI222_X1 U15707 ( .A1(n14159), .A2(n14147), .B1(n14161), .B2(n14146), .C1(
        n14156), .C2(n14145), .ZN(n14223) );
  AOI22_X1 U15708 ( .A1(n14164), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14163), 
        .B2(n14148), .ZN(n14149) );
  OAI21_X1 U15709 ( .B1(n14297), .B2(n14166), .A(n14149), .ZN(n14150) );
  AOI21_X1 U15710 ( .B1(n14223), .B2(n14169), .A(n14150), .ZN(n14151) );
  OAI21_X1 U15711 ( .B1(n14152), .B2(n14171), .A(n14151), .ZN(P3_U3217) );
  XNOR2_X1 U15712 ( .A(n14153), .B(n14154), .ZN(n14231) );
  XNOR2_X1 U15713 ( .A(n14155), .B(n14154), .ZN(n14157) );
  OAI222_X1 U15714 ( .A1(n14161), .A2(n14160), .B1(n14159), .B2(n14158), .C1(
        n14157), .C2(n14156), .ZN(n14228) );
  AOI22_X1 U15715 ( .A1(n14164), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n14163), 
        .B2(n14162), .ZN(n14165) );
  OAI21_X1 U15716 ( .B1(n14167), .B2(n14166), .A(n14165), .ZN(n14168) );
  AOI21_X1 U15717 ( .B1(n14228), .B2(n14169), .A(n14168), .ZN(n14170) );
  OAI21_X1 U15718 ( .B1(n14171), .B2(n14231), .A(n14170), .ZN(P3_U3218) );
  NOR2_X1 U15719 ( .A1(n16470), .A2(n16561), .ZN(n14174) );
  AOI21_X1 U15720 ( .B1(n16470), .B2(P3_REG1_REG_31__SCAN_IN), .A(n14174), 
        .ZN(n14172) );
  OAI21_X1 U15721 ( .B1(n14173), .B2(n14227), .A(n14172), .ZN(P3_U3490) );
  AOI21_X1 U15722 ( .B1(n16470), .B2(P3_REG1_REG_30__SCAN_IN), .A(n14174), 
        .ZN(n14175) );
  OAI21_X1 U15723 ( .B1(n14176), .B2(n14227), .A(n14175), .ZN(P3_U3489) );
  INV_X1 U15724 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n14180) );
  AND2_X1 U15725 ( .A1(n14177), .A2(n16469), .ZN(n14178) );
  NOR2_X1 U15726 ( .A1(n14179), .A2(n14178), .ZN(n14244) );
  MUX2_X1 U15727 ( .A(n14180), .B(n14244), .S(n16473), .Z(n14181) );
  INV_X1 U15728 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n14182) );
  MUX2_X1 U15729 ( .A(n14182), .B(n14253), .S(n16473), .Z(n14184) );
  NAND2_X1 U15730 ( .A1(n14255), .A2(n14189), .ZN(n14183) );
  OAI211_X1 U15731 ( .C1(n14257), .C2(n14243), .A(n14184), .B(n14183), .ZN(
        P3_U3485) );
  NAND2_X1 U15732 ( .A1(n14185), .A2(n16469), .ZN(n14186) );
  NAND2_X1 U15733 ( .A1(n14187), .A2(n14186), .ZN(n14258) );
  MUX2_X1 U15734 ( .A(n14258), .B(P3_REG1_REG_25__SCAN_IN), .S(n16470), .Z(
        n14188) );
  AOI21_X1 U15735 ( .B1(n14189), .B2(n14260), .A(n14188), .ZN(n14190) );
  INV_X1 U15736 ( .A(n14190), .ZN(P3_U3484) );
  INV_X1 U15737 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n14193) );
  AOI21_X1 U15738 ( .B1(n16469), .B2(n14192), .A(n14191), .ZN(n14262) );
  MUX2_X1 U15739 ( .A(n14193), .B(n14262), .S(n16473), .Z(n14194) );
  OAI21_X1 U15740 ( .B1(n14265), .B2(n14227), .A(n14194), .ZN(P3_U3483) );
  INV_X1 U15741 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n14197) );
  AOI21_X1 U15742 ( .B1(n14196), .B2(n16469), .A(n14195), .ZN(n14266) );
  MUX2_X1 U15743 ( .A(n14197), .B(n14266), .S(n16473), .Z(n14198) );
  OAI21_X1 U15744 ( .B1(n14269), .B2(n14227), .A(n14198), .ZN(P3_U3482) );
  MUX2_X1 U15745 ( .A(n14270), .B(P3_REG1_REG_22__SCAN_IN), .S(n16470), .Z(
        n14201) );
  INV_X1 U15746 ( .A(n14199), .ZN(n14271) );
  OAI22_X1 U15747 ( .A1(n14272), .A2(n14243), .B1(n14271), .B2(n14227), .ZN(
        n14200) );
  OR2_X1 U15748 ( .A1(n14201), .A2(n14200), .ZN(P3_U3481) );
  MUX2_X1 U15749 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n14275), .S(n16473), .Z(
        n14204) );
  INV_X1 U15750 ( .A(n14202), .ZN(n14276) );
  OAI22_X1 U15751 ( .A1(n14277), .A2(n14243), .B1(n14276), .B2(n14227), .ZN(
        n14203) );
  OR2_X1 U15752 ( .A1(n14204), .A2(n14203), .ZN(P3_U3480) );
  INV_X1 U15753 ( .A(n14205), .ZN(n14283) );
  INV_X1 U15754 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n14209) );
  NAND2_X1 U15755 ( .A1(n14206), .A2(n16469), .ZN(n14207) );
  AND2_X1 U15756 ( .A1(n14208), .A2(n14207), .ZN(n14280) );
  MUX2_X1 U15757 ( .A(n14209), .B(n14280), .S(n16473), .Z(n14210) );
  OAI21_X1 U15758 ( .B1(n14283), .B2(n14227), .A(n14210), .ZN(P3_U3479) );
  AOI21_X1 U15759 ( .B1(n14212), .B2(n16469), .A(n14211), .ZN(n14284) );
  MUX2_X1 U15760 ( .A(n14213), .B(n14284), .S(n16473), .Z(n14214) );
  OAI21_X1 U15761 ( .B1(n14227), .B2(n14287), .A(n14214), .ZN(P3_U3478) );
  AOI21_X1 U15762 ( .B1(n14216), .B2(n16469), .A(n14215), .ZN(n14288) );
  MUX2_X1 U15763 ( .A(n14217), .B(n14288), .S(n16473), .Z(n14218) );
  OAI21_X1 U15764 ( .B1(n14291), .B2(n14227), .A(n14218), .ZN(P3_U3477) );
  INV_X1 U15765 ( .A(n16469), .ZN(n14232) );
  AOI21_X1 U15766 ( .B1(n16410), .B2(n14220), .A(n14219), .ZN(n14221) );
  OAI21_X1 U15767 ( .B1(n14232), .B2(n14222), .A(n14221), .ZN(n14292) );
  MUX2_X1 U15768 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n14292), .S(n16473), .Z(
        P3_U3476) );
  AOI21_X1 U15769 ( .B1(n16469), .B2(n14224), .A(n14223), .ZN(n14293) );
  MUX2_X1 U15770 ( .A(n14225), .B(n14293), .S(n16473), .Z(n14226) );
  OAI21_X1 U15771 ( .B1(n14297), .B2(n14227), .A(n14226), .ZN(P3_U3475) );
  AOI21_X1 U15772 ( .B1(n16410), .B2(n14229), .A(n14228), .ZN(n14230) );
  OAI21_X1 U15773 ( .B1(n14232), .B2(n14231), .A(n14230), .ZN(n14298) );
  MUX2_X1 U15774 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n14298), .S(n16473), .Z(
        P3_U3474) );
  NAND2_X1 U15775 ( .A1(n14233), .A2(n16469), .ZN(n14234) );
  OAI211_X1 U15776 ( .C1(n16467), .C2(n14236), .A(n14235), .B(n14234), .ZN(
        n14299) );
  MUX2_X1 U15777 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n14299), .S(n16473), .Z(
        P3_U3473) );
  INV_X1 U15778 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14241) );
  OAI21_X1 U15779 ( .B1(n14238), .B2(n16467), .A(n14237), .ZN(n14239) );
  AOI21_X1 U15780 ( .B1(n14240), .B2(n16475), .A(n14239), .ZN(n14300) );
  MUX2_X1 U15781 ( .A(n14241), .B(n14300), .S(n16473), .Z(n14242) );
  OAI21_X1 U15782 ( .B1(n14304), .B2(n14243), .A(n14242), .ZN(P3_U3472) );
  INV_X1 U15783 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n14245) );
  MUX2_X1 U15784 ( .A(n14245), .B(n14244), .S(n16447), .Z(n14246) );
  MUX2_X1 U15785 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n14248), .S(n16447), .Z(
        n14252) );
  OAI22_X1 U15786 ( .A1(n14250), .A2(n14303), .B1(n14249), .B2(n14296), .ZN(
        n14251) );
  INV_X1 U15787 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14254) );
  INV_X1 U15788 ( .A(n14296), .ZN(n16558) );
  NAND2_X1 U15789 ( .A1(n14255), .A2(n16558), .ZN(n14256) );
  MUX2_X1 U15790 ( .A(n14258), .B(P3_REG0_REG_25__SCAN_IN), .S(n16562), .Z(
        n14259) );
  AOI21_X1 U15791 ( .B1(n16558), .B2(n14260), .A(n14259), .ZN(n14261) );
  INV_X1 U15792 ( .A(n14261), .ZN(P3_U3452) );
  INV_X1 U15793 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14263) );
  MUX2_X1 U15794 ( .A(n14263), .B(n14262), .S(n16447), .Z(n14264) );
  OAI21_X1 U15795 ( .B1(n14265), .B2(n14296), .A(n14264), .ZN(P3_U3451) );
  MUX2_X1 U15796 ( .A(n14267), .B(n14266), .S(n16447), .Z(n14268) );
  OAI21_X1 U15797 ( .B1(n14269), .B2(n14296), .A(n14268), .ZN(P3_U3450) );
  MUX2_X1 U15798 ( .A(n14270), .B(P3_REG0_REG_22__SCAN_IN), .S(n16562), .Z(
        n14274) );
  OAI22_X1 U15799 ( .A1(n14272), .A2(n14303), .B1(n14271), .B2(n14296), .ZN(
        n14273) );
  OR2_X1 U15800 ( .A1(n14274), .A2(n14273), .ZN(P3_U3449) );
  MUX2_X1 U15801 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n14275), .S(n16447), .Z(
        n14279) );
  OAI22_X1 U15802 ( .A1(n14277), .A2(n14303), .B1(n14276), .B2(n14296), .ZN(
        n14278) );
  OR2_X1 U15803 ( .A1(n14279), .A2(n14278), .ZN(P3_U3448) );
  INV_X1 U15804 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n14281) );
  MUX2_X1 U15805 ( .A(n14281), .B(n14280), .S(n16447), .Z(n14282) );
  OAI21_X1 U15806 ( .B1(n14283), .B2(n14296), .A(n14282), .ZN(P3_U3447) );
  INV_X1 U15807 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14285) );
  MUX2_X1 U15808 ( .A(n14285), .B(n14284), .S(n16447), .Z(n14286) );
  OAI21_X1 U15809 ( .B1(n14296), .B2(n14287), .A(n14286), .ZN(P3_U3446) );
  INV_X1 U15810 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n14289) );
  MUX2_X1 U15811 ( .A(n14289), .B(n14288), .S(n16447), .Z(n14290) );
  OAI21_X1 U15812 ( .B1(n14291), .B2(n14296), .A(n14290), .ZN(P3_U3444) );
  MUX2_X1 U15813 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n14292), .S(n16447), .Z(
        P3_U3441) );
  INV_X1 U15814 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n14294) );
  MUX2_X1 U15815 ( .A(n14294), .B(n14293), .S(n16447), .Z(n14295) );
  OAI21_X1 U15816 ( .B1(n14297), .B2(n14296), .A(n14295), .ZN(P3_U3438) );
  MUX2_X1 U15817 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n14298), .S(n16447), .Z(
        P3_U3435) );
  MUX2_X1 U15818 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n14299), .S(n16447), .Z(
        P3_U3432) );
  INV_X1 U15819 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14301) );
  MUX2_X1 U15820 ( .A(n14301), .B(n14300), .S(n16447), .Z(n14302) );
  OAI21_X1 U15821 ( .B1(n14304), .B2(n14303), .A(n14302), .ZN(P3_U3429) );
  MUX2_X1 U15822 ( .A(n14305), .B(P3_D_REG_1__SCAN_IN), .S(n14306), .Z(
        P3_U3377) );
  MUX2_X1 U15823 ( .A(n14307), .B(P3_D_REG_0__SCAN_IN), .S(n14306), .Z(
        P3_U3376) );
  INV_X1 U15824 ( .A(n14308), .ZN(n14313) );
  NOR4_X1 U15825 ( .A1(n9618), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n8405), .ZN(n14309) );
  AOI21_X1 U15826 ( .B1(n14310), .B2(SI_31_), .A(n14309), .ZN(n14311) );
  OAI21_X1 U15827 ( .B1(n14313), .B2(n14312), .A(n14311), .ZN(P3_U3264) );
  INV_X1 U15828 ( .A(n14314), .ZN(n14318) );
  OAI222_X1 U15829 ( .A1(n14312), .A2(n14318), .B1(n14317), .B2(P3_U3151), 
        .C1(n14316), .C2(n14315), .ZN(P3_U3266) );
  XNOR2_X1 U15830 ( .A(n10455), .B(n10853), .ZN(n14331) );
  INV_X1 U15831 ( .A(n14331), .ZN(n14333) );
  NAND2_X1 U15832 ( .A1(n14454), .A2(n14491), .ZN(n14332) );
  INV_X1 U15833 ( .A(n14319), .ZN(n14322) );
  INV_X1 U15834 ( .A(n14320), .ZN(n14321) );
  NAND2_X1 U15835 ( .A1(n14322), .A2(n14321), .ZN(n14323) );
  XNOR2_X1 U15836 ( .A(n14585), .B(n10853), .ZN(n14326) );
  NOR2_X1 U15837 ( .A1(n14597), .A2(n16261), .ZN(n14410) );
  XNOR2_X1 U15838 ( .A(n14721), .B(n10853), .ZN(n14327) );
  XNOR2_X1 U15839 ( .A(n14329), .B(n14327), .ZN(n14348) );
  NAND2_X1 U15840 ( .A1(n14558), .A2(n14491), .ZN(n14347) );
  INV_X1 U15841 ( .A(n14327), .ZN(n14328) );
  AND2_X1 U15842 ( .A1(n14329), .A2(n14328), .ZN(n14330) );
  XNOR2_X1 U15843 ( .A(n14331), .B(n14332), .ZN(n14391) );
  NAND2_X1 U15844 ( .A1(n14392), .A2(n14391), .ZN(n14390) );
  XNOR2_X1 U15845 ( .A(n14768), .B(n10853), .ZN(n14335) );
  NAND2_X1 U15846 ( .A1(n14559), .A2(n14491), .ZN(n14334) );
  NAND2_X1 U15847 ( .A1(n14335), .A2(n14334), .ZN(n14379) );
  NOR2_X1 U15848 ( .A1(n14335), .A2(n14334), .ZN(n14381) );
  AND2_X1 U15849 ( .A1(n14453), .A2(n14491), .ZN(n14337) );
  XNOR2_X1 U15850 ( .A(n14705), .B(n10853), .ZN(n14336) );
  NOR2_X1 U15851 ( .A1(n14336), .A2(n14337), .ZN(n14338) );
  AOI21_X1 U15852 ( .B1(n14337), .B2(n14336), .A(n14338), .ZN(n14436) );
  INV_X1 U15853 ( .A(n14338), .ZN(n14339) );
  XNOR2_X1 U15854 ( .A(n14511), .B(n10853), .ZN(n14367) );
  NAND2_X1 U15855 ( .A1(n14452), .A2(n14491), .ZN(n14366) );
  XNOR2_X1 U15856 ( .A(n14367), .B(n14366), .ZN(n14368) );
  OAI22_X1 U15857 ( .A1(n14369), .A2(n16108), .B1(n14340), .B2(n14652), .ZN(
        n14505) );
  INV_X1 U15858 ( .A(n14509), .ZN(n14342) );
  OAI22_X1 U15859 ( .A1(n14342), .A2(n14442), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14341), .ZN(n14343) );
  AOI21_X1 U15860 ( .B1(n14505), .B2(n14445), .A(n14343), .ZN(n14345) );
  NAND2_X1 U15861 ( .A1(n14700), .A2(n14432), .ZN(n14344) );
  OAI211_X1 U15862 ( .C1(n14346), .C2(n14427), .A(n14345), .B(n14344), .ZN(
        P2_U3186) );
  NAND2_X1 U15863 ( .A1(n14411), .A2(n14558), .ZN(n14350) );
  NAND2_X1 U15864 ( .A1(n14347), .A2(n14437), .ZN(n14349) );
  MUX2_X1 U15865 ( .A(n14350), .B(n14349), .S(n14348), .Z(n14354) );
  AOI22_X1 U15866 ( .A1(n14420), .A2(n14574), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14353) );
  AOI22_X1 U15867 ( .A1(n14424), .A2(n14455), .B1(n14423), .B2(n14454), .ZN(
        n14352) );
  NAND2_X1 U15868 ( .A1(n14721), .A2(n14432), .ZN(n14351) );
  NAND4_X1 U15869 ( .A1(n14354), .A2(n14353), .A3(n14352), .A4(n14351), .ZN(
        P2_U3188) );
  INV_X1 U15870 ( .A(n14401), .ZN(n14355) );
  AOI21_X1 U15871 ( .B1(n7489), .B2(n14359), .A(n14355), .ZN(n14365) );
  NAND2_X1 U15872 ( .A1(n14420), .A2(n14634), .ZN(n14356) );
  OAI211_X1 U15873 ( .C1(n14417), .C2(n14596), .A(n14357), .B(n14356), .ZN(
        n14363) );
  NAND3_X1 U15874 ( .A1(n14359), .A2(n14411), .A3(n14358), .ZN(n14361) );
  AOI21_X1 U15875 ( .B1(n14361), .B2(n14416), .A(n14360), .ZN(n14362) );
  AOI211_X1 U15876 ( .C1(n14742), .C2(n14432), .A(n14363), .B(n14362), .ZN(
        n14364) );
  OAI21_X1 U15877 ( .B1(n14365), .B2(n14408), .A(n14364), .ZN(P2_U3191) );
  NOR2_X1 U15878 ( .A1(n14369), .A2(n16261), .ZN(n14370) );
  XNOR2_X1 U15879 ( .A(n14370), .B(n10853), .ZN(n14371) );
  XNOR2_X1 U15880 ( .A(n14493), .B(n14371), .ZN(n14372) );
  OAI22_X1 U15881 ( .A1(n14440), .A2(n14652), .B1(n14373), .B2(n16108), .ZN(
        n14487) );
  OAI22_X1 U15882 ( .A1(n14495), .A2(n14442), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14374), .ZN(n14375) );
  AOI21_X1 U15883 ( .B1(n14487), .B2(n14445), .A(n14375), .ZN(n14377) );
  NAND2_X1 U15884 ( .A1(n14695), .A2(n14432), .ZN(n14376) );
  INV_X1 U15885 ( .A(n14379), .ZN(n14380) );
  NOR2_X1 U15886 ( .A1(n14381), .A2(n14380), .ZN(n14382) );
  XNOR2_X1 U15887 ( .A(n14383), .B(n14382), .ZN(n14389) );
  AOI22_X1 U15888 ( .A1(n14453), .A2(n14628), .B1(n14627), .B2(n14454), .ZN(
        n14536) );
  INV_X1 U15889 ( .A(n14384), .ZN(n14541) );
  AOI22_X1 U15890 ( .A1(n14541), .A2(n14420), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14385) );
  OAI21_X1 U15891 ( .B1(n14536), .B2(n14386), .A(n14385), .ZN(n14387) );
  AOI21_X1 U15892 ( .B1(n7754), .B2(n14432), .A(n14387), .ZN(n14388) );
  OAI21_X1 U15893 ( .B1(n14389), .B2(n14408), .A(n14388), .ZN(P2_U3197) );
  OAI211_X1 U15894 ( .C1(n14392), .C2(n14391), .A(n14390), .B(n14437), .ZN(
        n14396) );
  NOR2_X1 U15895 ( .A1(n14551), .A2(n14442), .ZN(n14394) );
  OAI22_X1 U15896 ( .A1(n14439), .A2(n14417), .B1(n14582), .B2(n14416), .ZN(
        n14393) );
  AOI211_X1 U15897 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3088), .A(n14394), 
        .B(n14393), .ZN(n14395) );
  OAI211_X1 U15898 ( .C1(n14772), .C2(n14448), .A(n14396), .B(n14395), .ZN(
        P2_U3201) );
  INV_X1 U15899 ( .A(n14397), .ZN(n14402) );
  OAI22_X1 U15900 ( .A1(n14399), .A2(n14408), .B1(n14654), .B2(n14398), .ZN(
        n14400) );
  NAND3_X1 U15901 ( .A1(n14402), .A2(n14401), .A3(n14400), .ZN(n14407) );
  AOI22_X1 U15902 ( .A1(n14456), .A2(n14628), .B1(n14627), .B2(n14457), .ZN(
        n14610) );
  INV_X1 U15903 ( .A(n14610), .ZN(n14403) );
  AOI22_X1 U15904 ( .A1(n14403), .A2(n14445), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14404) );
  OAI21_X1 U15905 ( .B1(n14613), .B2(n14442), .A(n14404), .ZN(n14405) );
  AOI21_X1 U15906 ( .B1(n14739), .B2(n14432), .A(n14405), .ZN(n14406) );
  OAI211_X1 U15907 ( .C1(n14409), .C2(n14408), .A(n14407), .B(n14406), .ZN(
        P2_U3205) );
  OR2_X1 U15908 ( .A1(n14410), .A2(n14427), .ZN(n14414) );
  NAND2_X1 U15909 ( .A1(n14411), .A2(n14455), .ZN(n14413) );
  MUX2_X1 U15910 ( .A(n14414), .B(n14413), .S(n14412), .Z(n14422) );
  NOR2_X1 U15911 ( .A1(n14415), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14419) );
  OAI22_X1 U15912 ( .A1(n14582), .A2(n14417), .B1(n14416), .B2(n14581), .ZN(
        n14418) );
  AOI211_X1 U15913 ( .C1(n14420), .C2(n14586), .A(n14419), .B(n14418), .ZN(
        n14421) );
  OAI211_X1 U15914 ( .C1(n14777), .C2(n14448), .A(n14422), .B(n14421), .ZN(
        P2_U3207) );
  INV_X1 U15915 ( .A(n14646), .ZN(n14426) );
  AOI22_X1 U15916 ( .A1(n14424), .A2(n14458), .B1(n14423), .B2(n14457), .ZN(
        n14425) );
  NAND2_X1 U15917 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n15679)
         );
  OAI211_X1 U15918 ( .C1(n14426), .C2(n14442), .A(n14425), .B(n15679), .ZN(
        n14431) );
  AOI211_X1 U15919 ( .C1(n14429), .C2(n14428), .A(n14427), .B(n7489), .ZN(
        n14430) );
  AOI211_X1 U15920 ( .C1(n14645), .C2(n14432), .A(n14431), .B(n14430), .ZN(
        n14433) );
  INV_X1 U15921 ( .A(n14433), .ZN(P2_U3210) );
  OAI21_X1 U15922 ( .B1(n14436), .B2(n14435), .A(n14434), .ZN(n14438) );
  NAND2_X1 U15923 ( .A1(n14438), .A2(n14437), .ZN(n14447) );
  OAI22_X1 U15924 ( .A1(n14440), .A2(n16108), .B1(n14439), .B2(n14652), .ZN(
        n14519) );
  INV_X1 U15925 ( .A(n14524), .ZN(n14443) );
  OAI22_X1 U15926 ( .A1(n14443), .A2(n14442), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14441), .ZN(n14444) );
  AOI21_X1 U15927 ( .B1(n14519), .B2(n14445), .A(n14444), .ZN(n14446) );
  OAI211_X1 U15928 ( .C1(n14521), .C2(n14448), .A(n14447), .B(n14446), .ZN(
        P2_U3212) );
  MUX2_X1 U15929 ( .A(n14449), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14474), .Z(
        P2_U3561) );
  INV_X2 U15930 ( .A(P2_U3947), .ZN(n14474) );
  MUX2_X1 U15931 ( .A(n14450), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14474), .Z(
        P2_U3560) );
  MUX2_X1 U15932 ( .A(n14451), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14474), .Z(
        P2_U3559) );
  MUX2_X1 U15933 ( .A(n14452), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14474), .Z(
        P2_U3558) );
  MUX2_X1 U15934 ( .A(n14453), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14474), .Z(
        P2_U3557) );
  MUX2_X1 U15935 ( .A(n14559), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14474), .Z(
        P2_U3556) );
  MUX2_X1 U15936 ( .A(n14454), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14474), .Z(
        P2_U3555) );
  MUX2_X1 U15937 ( .A(n14558), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14474), .Z(
        P2_U3554) );
  MUX2_X1 U15938 ( .A(n14455), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14474), .Z(
        P2_U3553) );
  MUX2_X1 U15939 ( .A(n14456), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14474), .Z(
        P2_U3552) );
  MUX2_X1 U15940 ( .A(n14629), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14474), .Z(
        P2_U3551) );
  MUX2_X1 U15941 ( .A(n14457), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14474), .Z(
        P2_U3550) );
  MUX2_X1 U15942 ( .A(n14626), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14474), .Z(
        P2_U3549) );
  MUX2_X1 U15943 ( .A(n14458), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14474), .Z(
        P2_U3548) );
  MUX2_X1 U15944 ( .A(n14459), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14474), .Z(
        P2_U3547) );
  MUX2_X1 U15945 ( .A(n14460), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14474), .Z(
        P2_U3546) );
  MUX2_X1 U15946 ( .A(n14461), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14474), .Z(
        P2_U3545) );
  MUX2_X1 U15947 ( .A(n14462), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14474), .Z(
        P2_U3543) );
  MUX2_X1 U15948 ( .A(n14463), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14474), .Z(
        P2_U3542) );
  MUX2_X1 U15949 ( .A(n14464), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14474), .Z(
        P2_U3541) );
  MUX2_X1 U15950 ( .A(n14465), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14474), .Z(
        P2_U3540) );
  MUX2_X1 U15951 ( .A(n14466), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14474), .Z(
        P2_U3539) );
  MUX2_X1 U15952 ( .A(n14467), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14474), .Z(
        P2_U3538) );
  MUX2_X1 U15953 ( .A(n14468), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14474), .Z(
        P2_U3537) );
  MUX2_X1 U15954 ( .A(n14469), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14474), .Z(
        P2_U3536) );
  MUX2_X1 U15955 ( .A(n14470), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14474), .Z(
        P2_U3535) );
  MUX2_X1 U15956 ( .A(n14471), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14474), .Z(
        P2_U3534) );
  MUX2_X1 U15957 ( .A(n14472), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14474), .Z(
        P2_U3533) );
  MUX2_X1 U15958 ( .A(n14473), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14474), .Z(
        P2_U3532) );
  MUX2_X1 U15959 ( .A(n14475), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14474), .Z(
        P2_U3531) );
  NOR2_X1 U15960 ( .A1(n14675), .A2(n14476), .ZN(n14477) );
  NOR2_X1 U15961 ( .A1(n16408), .A2(n14688), .ZN(n14484) );
  AOI211_X1 U15962 ( .C1(n14687), .C2(n16399), .A(n14477), .B(n14484), .ZN(
        n14478) );
  OAI21_X1 U15963 ( .B1(n14479), .B2(n16228), .A(n14478), .ZN(P2_U3234) );
  AOI21_X1 U15964 ( .B1(n14480), .B2(n14691), .A(n14491), .ZN(n14482) );
  NAND2_X1 U15965 ( .A1(n14482), .A2(n14481), .ZN(n14689) );
  NOR2_X1 U15966 ( .A1(n8926), .A2(n14648), .ZN(n14483) );
  AOI211_X1 U15967 ( .C1(n16408), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14484), 
        .B(n14483), .ZN(n14485) );
  OAI21_X1 U15968 ( .B1(n14689), .B2(n16228), .A(n14485), .ZN(P2_U3235) );
  AOI21_X1 U15969 ( .B1(n14486), .B2(n14499), .A(n16256), .ZN(n14489) );
  AOI21_X1 U15970 ( .B1(n14489), .B2(n14488), .A(n14487), .ZN(n14696) );
  INV_X1 U15971 ( .A(n14507), .ZN(n14492) );
  AOI211_X1 U15972 ( .C1(n14695), .C2(n14492), .A(n14491), .B(n8912), .ZN(
        n14694) );
  NOR2_X1 U15973 ( .A1(n14493), .A2(n14648), .ZN(n14497) );
  OAI22_X1 U15974 ( .A1(n14495), .A2(n16117), .B1(n14494), .B2(n14675), .ZN(
        n14496) );
  AOI211_X1 U15975 ( .C1(n14694), .C2(n16403), .A(n14497), .B(n14496), .ZN(
        n14502) );
  NAND2_X1 U15976 ( .A1(n14693), .A2(n14678), .ZN(n14501) );
  OAI211_X1 U15977 ( .C1(n16408), .C2(n14696), .A(n14502), .B(n14501), .ZN(
        P2_U3237) );
  XNOR2_X1 U15978 ( .A(n14504), .B(n14503), .ZN(n14506) );
  AOI21_X1 U15979 ( .B1(n14506), .B2(n16107), .A(n14505), .ZN(n14701) );
  INV_X1 U15980 ( .A(n14523), .ZN(n14508) );
  AOI211_X1 U15981 ( .C1(n14700), .C2(n14508), .A(n14491), .B(n14507), .ZN(
        n14699) );
  AOI22_X1 U15982 ( .A1(n14509), .A2(n16397), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n16408), .ZN(n14510) );
  OAI21_X1 U15983 ( .B1(n14511), .B2(n14648), .A(n14510), .ZN(n14516) );
  OAI21_X1 U15984 ( .B1(n14514), .B2(n14513), .A(n14512), .ZN(n14703) );
  NOR2_X1 U15985 ( .A1(n14703), .A2(n14620), .ZN(n14515) );
  AOI211_X1 U15986 ( .C1(n14699), .C2(n16403), .A(n14516), .B(n14515), .ZN(
        n14517) );
  OAI21_X1 U15987 ( .B1(n16408), .B2(n14701), .A(n14517), .ZN(P2_U3238) );
  XNOR2_X1 U15988 ( .A(n14518), .B(n14529), .ZN(n14520) );
  AOI21_X1 U15989 ( .B1(n14520), .B2(n16107), .A(n14519), .ZN(n14708) );
  NOR2_X1 U15990 ( .A1(n7410), .A2(n14521), .ZN(n14522) );
  NAND2_X1 U15991 ( .A1(n14524), .A2(n16397), .ZN(n14525) );
  OAI21_X1 U15992 ( .B1(n14675), .B2(n14526), .A(n14525), .ZN(n14527) );
  AOI21_X1 U15993 ( .B1(n14705), .B2(n16399), .A(n14527), .ZN(n14532) );
  NAND2_X1 U15994 ( .A1(n14530), .A2(n14529), .ZN(n14704) );
  NAND3_X1 U15995 ( .A1(n14528), .A2(n14678), .A3(n14704), .ZN(n14531) );
  OAI211_X1 U15996 ( .C1(n14707), .C2(n16228), .A(n14532), .B(n14531), .ZN(
        n14533) );
  INV_X1 U15997 ( .A(n14533), .ZN(n14534) );
  OAI21_X1 U15998 ( .B1(n14708), .B2(n16408), .A(n14534), .ZN(P2_U3239) );
  XNOR2_X1 U15999 ( .A(n14538), .B(n14535), .ZN(n14537) );
  OAI21_X1 U16000 ( .B1(n14537), .B2(n16256), .A(n14536), .ZN(n14710) );
  INV_X1 U16001 ( .A(n14710), .ZN(n14546) );
  XOR2_X1 U16002 ( .A(n14539), .B(n14538), .Z(n14712) );
  INV_X1 U16003 ( .A(n14549), .ZN(n14540) );
  AOI211_X1 U16004 ( .C1(n7754), .C2(n14540), .A(n14491), .B(n7410), .ZN(
        n14711) );
  NAND2_X1 U16005 ( .A1(n14711), .A2(n16403), .ZN(n14543) );
  AOI22_X1 U16006 ( .A1(n14541), .A2(n16397), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n16408), .ZN(n14542) );
  OAI211_X1 U16007 ( .C1(n14768), .C2(n14648), .A(n14543), .B(n14542), .ZN(
        n14544) );
  AOI21_X1 U16008 ( .B1(n14678), .B2(n14712), .A(n14544), .ZN(n14545) );
  OAI21_X1 U16009 ( .B1(n16408), .B2(n14546), .A(n14545), .ZN(P2_U3240) );
  INV_X1 U16010 ( .A(n14547), .ZN(n14548) );
  XNOR2_X1 U16011 ( .A(n14557), .B(n14548), .ZN(n14717) );
  INV_X1 U16012 ( .A(n14717), .ZN(n14565) );
  INV_X1 U16013 ( .A(n16401), .ZN(n14660) );
  AOI211_X1 U16014 ( .C1(n10455), .C2(n14573), .A(n14491), .B(n14549), .ZN(
        n14716) );
  NOR2_X1 U16015 ( .A1(n14772), .A2(n14648), .ZN(n14553) );
  OAI22_X1 U16016 ( .A1(n14551), .A2(n16117), .B1(n14550), .B2(n14675), .ZN(
        n14552) );
  AOI211_X1 U16017 ( .C1(n14716), .C2(n16403), .A(n14553), .B(n14552), .ZN(
        n14564) );
  INV_X1 U16018 ( .A(n14554), .ZN(n14555) );
  AOI21_X1 U16019 ( .B1(n14557), .B2(n14556), .A(n14555), .ZN(n14562) );
  AOI22_X1 U16020 ( .A1(n14559), .A2(n14628), .B1(n14627), .B2(n14558), .ZN(
        n14561) );
  NAND2_X1 U16021 ( .A1(n14717), .A2(n16259), .ZN(n14560) );
  OAI211_X1 U16022 ( .C1(n14562), .C2(n16256), .A(n14561), .B(n14560), .ZN(
        n14715) );
  NAND2_X1 U16023 ( .A1(n14715), .A2(n14675), .ZN(n14563) );
  OAI211_X1 U16024 ( .C1(n14565), .C2(n14660), .A(n14564), .B(n14563), .ZN(
        P2_U3241) );
  XOR2_X1 U16025 ( .A(n14566), .B(n14569), .Z(n14572) );
  OAI22_X1 U16026 ( .A1(n14567), .A2(n16108), .B1(n14597), .B2(n14652), .ZN(
        n14571) );
  XNOR2_X1 U16027 ( .A(n14568), .B(n14569), .ZN(n14724) );
  NOR2_X1 U16028 ( .A1(n14724), .A2(n16431), .ZN(n14570) );
  AOI211_X1 U16029 ( .C1(n14572), .C2(n16107), .A(n14571), .B(n14570), .ZN(
        n14723) );
  AOI211_X1 U16030 ( .C1(n14721), .C2(n14584), .A(n14491), .B(n7752), .ZN(
        n14720) );
  AOI22_X1 U16031 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(n16408), .B1(n14574), 
        .B2(n16397), .ZN(n14575) );
  OAI21_X1 U16032 ( .B1(n8873), .B2(n14648), .A(n14575), .ZN(n14577) );
  NOR2_X1 U16033 ( .A1(n14724), .A2(n14660), .ZN(n14576) );
  AOI211_X1 U16034 ( .C1(n14720), .C2(n16403), .A(n14577), .B(n14576), .ZN(
        n14578) );
  OAI21_X1 U16035 ( .B1(n14723), .B2(n16408), .A(n14578), .ZN(P2_U3242) );
  XNOR2_X1 U16036 ( .A(n14583), .B(n14579), .ZN(n14580) );
  OAI222_X1 U16037 ( .A1(n16108), .A2(n14582), .B1(n14652), .B2(n14581), .C1(
        n16256), .C2(n14580), .ZN(n14725) );
  INV_X1 U16038 ( .A(n14725), .ZN(n14591) );
  XOR2_X1 U16039 ( .A(n7408), .B(n14583), .Z(n14727) );
  AOI211_X1 U16040 ( .C1(n14585), .C2(n14598), .A(n14491), .B(n8872), .ZN(
        n14726) );
  NAND2_X1 U16041 ( .A1(n14726), .A2(n16403), .ZN(n14588) );
  AOI22_X1 U16042 ( .A1(n16408), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14586), 
        .B2(n16397), .ZN(n14587) );
  OAI211_X1 U16043 ( .C1(n14777), .C2(n14648), .A(n14588), .B(n14587), .ZN(
        n14589) );
  AOI21_X1 U16044 ( .B1(n14678), .B2(n14727), .A(n14589), .ZN(n14590) );
  OAI21_X1 U16045 ( .B1(n16408), .B2(n14591), .A(n14590), .ZN(P2_U3243) );
  XNOR2_X1 U16046 ( .A(n14593), .B(n14592), .ZN(n14734) );
  XOR2_X1 U16047 ( .A(n14594), .B(n14593), .Z(n14595) );
  OAI222_X1 U16048 ( .A1(n16108), .A2(n14597), .B1(n14652), .B2(n14596), .C1(
        n16256), .C2(n14595), .ZN(n14730) );
  NAND2_X1 U16049 ( .A1(n14730), .A2(n14675), .ZN(n14604) );
  AOI211_X1 U16050 ( .C1(n14732), .C2(n14612), .A(n14491), .B(n8871), .ZN(
        n14731) );
  NOR2_X1 U16051 ( .A1(n7743), .A2(n14648), .ZN(n14602) );
  OAI22_X1 U16052 ( .A1(n14675), .A2(n14600), .B1(n14599), .B2(n16117), .ZN(
        n14601) );
  AOI211_X1 U16053 ( .C1(n14731), .C2(n16403), .A(n14602), .B(n14601), .ZN(
        n14603) );
  OAI211_X1 U16054 ( .C1(n14734), .C2(n14620), .A(n14604), .B(n14603), .ZN(
        P2_U3244) );
  XNOR2_X1 U16055 ( .A(n14605), .B(n14606), .ZN(n14737) );
  OAI211_X1 U16056 ( .C1(n14609), .C2(n14608), .A(n14607), .B(n16107), .ZN(
        n14611) );
  AND2_X1 U16057 ( .A1(n14611), .A2(n14610), .ZN(n14736) );
  INV_X1 U16058 ( .A(n14736), .ZN(n14618) );
  OAI211_X1 U16059 ( .C1(n14782), .C2(n14633), .A(n16261), .B(n14612), .ZN(
        n14735) );
  OAI22_X1 U16060 ( .A1(n14675), .A2(n14614), .B1(n14613), .B2(n16117), .ZN(
        n14615) );
  AOI21_X1 U16061 ( .B1(n14739), .B2(n16399), .A(n14615), .ZN(n14616) );
  OAI21_X1 U16062 ( .B1(n14735), .B2(n16228), .A(n14616), .ZN(n14617) );
  AOI21_X1 U16063 ( .B1(n14618), .B2(n14675), .A(n14617), .ZN(n14619) );
  OAI21_X1 U16064 ( .B1(n14620), .B2(n14737), .A(n14619), .ZN(P2_U3245) );
  XNOR2_X1 U16065 ( .A(n14621), .B(n14623), .ZN(n14632) );
  NAND2_X1 U16066 ( .A1(n14623), .A2(n14622), .ZN(n14624) );
  NAND2_X1 U16067 ( .A1(n14625), .A2(n14624), .ZN(n14745) );
  AOI22_X1 U16068 ( .A1(n14629), .A2(n14628), .B1(n14627), .B2(n14626), .ZN(
        n14630) );
  OAI21_X1 U16069 ( .B1(n14745), .B2(n16431), .A(n14630), .ZN(n14631) );
  AOI21_X1 U16070 ( .B1(n14632), .B2(n16107), .A(n14631), .ZN(n14743) );
  AOI211_X1 U16071 ( .C1(n14742), .C2(n14642), .A(n14491), .B(n14633), .ZN(
        n14741) );
  INV_X1 U16072 ( .A(n14742), .ZN(n14636) );
  AOI22_X1 U16073 ( .A1(n16408), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14634), 
        .B2(n16397), .ZN(n14635) );
  OAI21_X1 U16074 ( .B1(n14636), .B2(n14648), .A(n14635), .ZN(n14638) );
  NOR2_X1 U16075 ( .A1(n14745), .A2(n14660), .ZN(n14637) );
  AOI211_X1 U16076 ( .C1(n14741), .C2(n16403), .A(n14638), .B(n14637), .ZN(
        n14639) );
  OAI21_X1 U16077 ( .B1(n16408), .B2(n14743), .A(n14639), .ZN(P2_U3246) );
  OAI21_X1 U16078 ( .B1(n14650), .B2(n14641), .A(n14640), .ZN(n14748) );
  INV_X1 U16079 ( .A(n14748), .ZN(n14661) );
  INV_X1 U16080 ( .A(n14642), .ZN(n14643) );
  AOI211_X1 U16081 ( .C1(n7745), .C2(n14644), .A(n14491), .B(n14643), .ZN(
        n14746) );
  AOI22_X1 U16082 ( .A1(n16408), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14646), 
        .B2(n16397), .ZN(n14647) );
  OAI21_X1 U16083 ( .B1(n14788), .B2(n14648), .A(n14647), .ZN(n14649) );
  AOI21_X1 U16084 ( .B1(n14746), .B2(n16403), .A(n14649), .ZN(n14659) );
  XOR2_X1 U16085 ( .A(n14651), .B(n14650), .Z(n14657) );
  OAI22_X1 U16086 ( .A1(n14654), .A2(n16108), .B1(n14653), .B2(n14652), .ZN(
        n14655) );
  AOI21_X1 U16087 ( .B1(n14748), .B2(n16259), .A(n14655), .ZN(n14656) );
  OAI21_X1 U16088 ( .B1(n14657), .B2(n16256), .A(n14656), .ZN(n14747) );
  NAND2_X1 U16089 ( .A1(n14747), .A2(n14675), .ZN(n14658) );
  OAI211_X1 U16090 ( .C1(n14661), .C2(n14660), .A(n14659), .B(n14658), .ZN(
        P2_U3247) );
  NAND2_X1 U16091 ( .A1(n14662), .A2(n14675), .ZN(n14672) );
  OAI22_X1 U16092 ( .A1(n14675), .A2(n14664), .B1(n14663), .B2(n16117), .ZN(
        n14665) );
  AOI21_X1 U16093 ( .B1(n14666), .B2(n16399), .A(n14665), .ZN(n14671) );
  NAND2_X1 U16094 ( .A1(n14667), .A2(n14678), .ZN(n14670) );
  NAND2_X1 U16095 ( .A1(n14668), .A2(n16403), .ZN(n14669) );
  NAND4_X1 U16096 ( .A1(n14672), .A2(n14671), .A3(n14670), .A4(n14669), .ZN(
        P2_U3251) );
  NAND2_X1 U16097 ( .A1(n14673), .A2(n14675), .ZN(n14684) );
  OAI22_X1 U16098 ( .A1(n14675), .A2(n11542), .B1(n14674), .B2(n16117), .ZN(
        n14676) );
  AOI21_X1 U16099 ( .B1(n14677), .B2(n16399), .A(n14676), .ZN(n14683) );
  NAND2_X1 U16100 ( .A1(n14679), .A2(n14678), .ZN(n14682) );
  NAND2_X1 U16101 ( .A1(n14680), .A2(n16403), .ZN(n14681) );
  NAND4_X1 U16102 ( .A1(n14684), .A2(n14683), .A3(n14682), .A4(n14681), .ZN(
        P2_U3253) );
  NAND2_X1 U16103 ( .A1(n14689), .A2(n14688), .ZN(n14759) );
  MUX2_X1 U16104 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14759), .S(n16512), .Z(
        n14690) );
  AOI21_X1 U16105 ( .B1(n14757), .B2(n14691), .A(n14690), .ZN(n14692) );
  INV_X1 U16106 ( .A(n14692), .ZN(P2_U3529) );
  INV_X1 U16107 ( .A(n14693), .ZN(n14698) );
  AOI21_X1 U16108 ( .B1(n16265), .B2(n14695), .A(n14694), .ZN(n14697) );
  OAI211_X1 U16109 ( .C1(n16456), .C2(n14698), .A(n14697), .B(n14696), .ZN(
        n14762) );
  MUX2_X1 U16110 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14762), .S(n16512), .Z(
        P2_U3527) );
  AOI21_X1 U16111 ( .B1(n16265), .B2(n14700), .A(n14699), .ZN(n14702) );
  OAI211_X1 U16112 ( .C1(n16456), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14763) );
  MUX2_X1 U16113 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14763), .S(n16512), .Z(
        P2_U3526) );
  NAND3_X1 U16114 ( .A1(n14528), .A2(n14751), .A3(n14704), .ZN(n14709) );
  NAND2_X1 U16115 ( .A1(n14705), .A2(n16265), .ZN(n14706) );
  NAND4_X1 U16116 ( .A1(n14709), .A2(n14708), .A3(n14707), .A4(n14706), .ZN(
        n14764) );
  MUX2_X1 U16117 ( .A(n14764), .B(P2_REG1_REG_26__SCAN_IN), .S(n16510), .Z(
        P2_U3525) );
  INV_X1 U16118 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14713) );
  AOI211_X1 U16119 ( .C1(n14751), .C2(n14712), .A(n14711), .B(n14710), .ZN(
        n14765) );
  MUX2_X1 U16120 ( .A(n14713), .B(n14765), .S(n16512), .Z(n14714) );
  OAI21_X1 U16121 ( .B1(n14768), .B2(n14750), .A(n14714), .ZN(P2_U3524) );
  INV_X1 U16122 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14718) );
  AOI211_X1 U16123 ( .C1(n14717), .C2(n16509), .A(n14716), .B(n14715), .ZN(
        n14769) );
  MUX2_X1 U16124 ( .A(n14718), .B(n14769), .S(n16512), .Z(n14719) );
  OAI21_X1 U16125 ( .B1(n14772), .B2(n14750), .A(n14719), .ZN(P2_U3523) );
  AOI21_X1 U16126 ( .B1(n16265), .B2(n14721), .A(n14720), .ZN(n14722) );
  OAI211_X1 U16127 ( .C1(n14724), .C2(n16430), .A(n14723), .B(n14722), .ZN(
        n14773) );
  MUX2_X1 U16128 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14773), .S(n16512), .Z(
        P2_U3522) );
  INV_X1 U16129 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14728) );
  AOI211_X1 U16130 ( .C1(n14751), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14774) );
  MUX2_X1 U16131 ( .A(n14728), .B(n14774), .S(n16512), .Z(n14729) );
  OAI21_X1 U16132 ( .B1(n14777), .B2(n14750), .A(n14729), .ZN(P2_U3521) );
  AOI211_X1 U16133 ( .C1(n16265), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        n14733) );
  OAI21_X1 U16134 ( .B1(n16456), .B2(n14734), .A(n14733), .ZN(n14778) );
  MUX2_X1 U16135 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14778), .S(n16512), .Z(
        P2_U3520) );
  OAI211_X1 U16136 ( .C1(n16456), .C2(n14737), .A(n14736), .B(n14735), .ZN(
        n14779) );
  MUX2_X1 U16137 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14779), .S(n16512), .Z(
        n14738) );
  AOI21_X1 U16138 ( .B1(n14757), .B2(n14739), .A(n14738), .ZN(n14740) );
  INV_X1 U16139 ( .A(n14740), .ZN(P2_U3519) );
  AOI21_X1 U16140 ( .B1(n16265), .B2(n14742), .A(n14741), .ZN(n14744) );
  OAI211_X1 U16141 ( .C1(n16430), .C2(n14745), .A(n14744), .B(n14743), .ZN(
        n14783) );
  MUX2_X1 U16142 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14783), .S(n16512), .Z(
        P2_U3518) );
  AOI211_X1 U16143 ( .C1(n16509), .C2(n14748), .A(n14747), .B(n14746), .ZN(
        n14784) );
  MUX2_X1 U16144 ( .A(n15675), .B(n14784), .S(n16512), .Z(n14749) );
  OAI21_X1 U16145 ( .B1(n14788), .B2(n14750), .A(n14749), .ZN(P2_U3517) );
  NAND2_X1 U16146 ( .A1(n14752), .A2(n14751), .ZN(n14755) );
  NAND3_X1 U16147 ( .A1(n14755), .A2(n14754), .A3(n14753), .ZN(n14789) );
  MUX2_X1 U16148 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14789), .S(n16512), .Z(
        n14756) );
  AOI21_X1 U16149 ( .B1(n14757), .B2(n14791), .A(n14756), .ZN(n14758) );
  INV_X1 U16150 ( .A(n14758), .ZN(P2_U3516) );
  MUX2_X1 U16151 ( .A(n14759), .B(P2_REG0_REG_30__SCAN_IN), .S(n16513), .Z(
        n14760) );
  INV_X1 U16152 ( .A(n14760), .ZN(n14761) );
  OAI21_X1 U16153 ( .B1(n8926), .B2(n14787), .A(n14761), .ZN(P2_U3497) );
  MUX2_X1 U16154 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14762), .S(n16516), .Z(
        P2_U3495) );
  MUX2_X1 U16155 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14763), .S(n16516), .Z(
        P2_U3494) );
  MUX2_X1 U16156 ( .A(n14764), .B(P2_REG0_REG_26__SCAN_IN), .S(n16513), .Z(
        P2_U3493) );
  INV_X1 U16157 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14766) );
  MUX2_X1 U16158 ( .A(n14766), .B(n14765), .S(n16516), .Z(n14767) );
  OAI21_X1 U16159 ( .B1(n14768), .B2(n14787), .A(n14767), .ZN(P2_U3492) );
  INV_X1 U16160 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14770) );
  MUX2_X1 U16161 ( .A(n14770), .B(n14769), .S(n16516), .Z(n14771) );
  OAI21_X1 U16162 ( .B1(n14772), .B2(n14787), .A(n14771), .ZN(P2_U3491) );
  MUX2_X1 U16163 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14773), .S(n16516), .Z(
        P2_U3490) );
  INV_X1 U16164 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14775) );
  MUX2_X1 U16165 ( .A(n14775), .B(n14774), .S(n16516), .Z(n14776) );
  OAI21_X1 U16166 ( .B1(n14777), .B2(n14787), .A(n14776), .ZN(P2_U3489) );
  MUX2_X1 U16167 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14778), .S(n16516), .Z(
        P2_U3488) );
  MUX2_X1 U16168 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14779), .S(n16516), .Z(
        n14780) );
  INV_X1 U16169 ( .A(n14780), .ZN(n14781) );
  OAI21_X1 U16170 ( .B1(n14782), .B2(n14787), .A(n14781), .ZN(P2_U3487) );
  MUX2_X1 U16171 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14783), .S(n16516), .Z(
        P2_U3486) );
  INV_X1 U16172 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14785) );
  MUX2_X1 U16173 ( .A(n14785), .B(n14784), .S(n16516), .Z(n14786) );
  OAI21_X1 U16174 ( .B1(n14788), .B2(n14787), .A(n14786), .ZN(P2_U3484) );
  MUX2_X1 U16175 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14789), .S(n16516), .Z(
        n14790) );
  AOI21_X1 U16176 ( .B1(n14792), .B2(n14791), .A(n14790), .ZN(n14793) );
  INV_X1 U16177 ( .A(n14793), .ZN(P2_U3481) );
  INV_X1 U16178 ( .A(n14794), .ZN(n15547) );
  NOR4_X1 U16179 ( .A1(n14796), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14795), .A4(
        P2_U3088), .ZN(n14797) );
  AOI21_X1 U16180 ( .B1(n14798), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14797), 
        .ZN(n14799) );
  OAI21_X1 U16181 ( .B1(n15547), .B2(n14819), .A(n14799), .ZN(P2_U3296) );
  OAI222_X1 U16182 ( .A1(n14802), .A2(P2_U3088), .B1(n14819), .B2(n14801), 
        .C1(n14800), .C2(n14821), .ZN(P2_U3298) );
  NAND2_X1 U16183 ( .A1(n14804), .A2(n14803), .ZN(n14806) );
  OAI211_X1 U16184 ( .C1(n14821), .C2(n14807), .A(n14806), .B(n14805), .ZN(
        P2_U3299) );
  OAI222_X1 U16185 ( .A1(n14821), .A2(n14810), .B1(n14819), .B2(n14809), .C1(
        P2_U3088), .C2(n14808), .ZN(P2_U3300) );
  INV_X1 U16186 ( .A(n14811), .ZN(n15549) );
  OAI222_X1 U16187 ( .A1(n14813), .A2(P2_U3088), .B1(n14819), .B2(n15549), 
        .C1(n14812), .C2(n14821), .ZN(P2_U3301) );
  INV_X1 U16188 ( .A(n14814), .ZN(n15552) );
  OAI222_X1 U16189 ( .A1(n14821), .A2(n14816), .B1(n14819), .B2(n15552), .C1(
        n14815), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U16190 ( .A(n14817), .ZN(n15555) );
  OAI222_X1 U16191 ( .A1(n14821), .A2(n14820), .B1(n14819), .B2(n15555), .C1(
        n14818), .C2(P2_U3088), .ZN(P2_U3303) );
  MUX2_X1 U16192 ( .A(n14822), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U16193 ( .A1(n15436), .A2(n14950), .ZN(n14824) );
  NAND2_X1 U16194 ( .A1(n8086), .A2(n14954), .ZN(n14823) );
  NAND2_X1 U16195 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  XNOR2_X1 U16196 ( .A(n14825), .B(n15001), .ZN(n14829) );
  NAND2_X1 U16197 ( .A1(n15436), .A2(n14954), .ZN(n14827) );
  NAND2_X1 U16198 ( .A1(n8086), .A2(n14955), .ZN(n14826) );
  NAND2_X1 U16199 ( .A1(n14827), .A2(n14826), .ZN(n14828) );
  NOR2_X1 U16200 ( .A1(n14829), .A2(n14828), .ZN(n14998) );
  AOI21_X1 U16201 ( .B1(n14829), .B2(n14828), .A(n14998), .ZN(n14963) );
  NAND2_X1 U16202 ( .A1(n15457), .A2(n14950), .ZN(n14831) );
  NAND2_X1 U16203 ( .A1(n15122), .A2(n14954), .ZN(n14830) );
  NAND2_X1 U16204 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  XNOR2_X1 U16205 ( .A(n14832), .B(n14925), .ZN(n14935) );
  NOR2_X1 U16206 ( .A1(n14833), .A2(n15003), .ZN(n14834) );
  AOI21_X1 U16207 ( .B1(n15457), .B2(n14900), .A(n14834), .ZN(n14936) );
  NAND2_X1 U16208 ( .A1(n14935), .A2(n14936), .ZN(n14940) );
  INV_X1 U16209 ( .A(n14940), .ZN(n15026) );
  AND2_X1 U16210 ( .A1(n14837), .A2(n14838), .ZN(n14835) );
  INV_X1 U16211 ( .A(n14837), .ZN(n14840) );
  INV_X1 U16212 ( .A(n14838), .ZN(n14839) );
  NAND2_X1 U16213 ( .A1(n14840), .A2(n14839), .ZN(n14841) );
  NAND2_X1 U16214 ( .A1(n16523), .A2(n14950), .ZN(n14843) );
  NAND2_X1 U16215 ( .A1(n15132), .A2(n14954), .ZN(n14842) );
  NAND2_X1 U16216 ( .A1(n14843), .A2(n14842), .ZN(n14844) );
  XNOR2_X1 U16217 ( .A(n14844), .B(n14925), .ZN(n14846) );
  AND2_X1 U16218 ( .A1(n14955), .A2(n15132), .ZN(n14845) );
  AOI21_X1 U16219 ( .B1(n16523), .B2(n14900), .A(n14845), .ZN(n14847) );
  NAND2_X1 U16220 ( .A1(n14846), .A2(n14847), .ZN(n14852) );
  INV_X1 U16221 ( .A(n14846), .ZN(n14849) );
  INV_X1 U16222 ( .A(n14847), .ZN(n14848) );
  NAND2_X1 U16223 ( .A1(n14849), .A2(n14848), .ZN(n14850) );
  NAND2_X1 U16224 ( .A1(n14852), .A2(n14850), .ZN(n16517) );
  INV_X1 U16225 ( .A(n16517), .ZN(n14851) );
  NAND2_X1 U16226 ( .A1(n16529), .A2(n14950), .ZN(n14854) );
  NAND2_X1 U16227 ( .A1(n15131), .A2(n14954), .ZN(n14853) );
  NAND2_X1 U16228 ( .A1(n14854), .A2(n14853), .ZN(n14855) );
  XNOR2_X1 U16229 ( .A(n14855), .B(n15001), .ZN(n14858) );
  XNOR2_X1 U16230 ( .A(n14860), .B(n14858), .ZN(n15110) );
  NAND2_X1 U16231 ( .A1(n16529), .A2(n14954), .ZN(n14857) );
  NAND2_X1 U16232 ( .A1(n15131), .A2(n14955), .ZN(n14856) );
  NAND2_X1 U16233 ( .A1(n14857), .A2(n14856), .ZN(n15109) );
  INV_X1 U16234 ( .A(n14858), .ZN(n14859) );
  NOR2_X1 U16235 ( .A1(n14860), .A2(n14859), .ZN(n14861) );
  AOI21_X1 U16236 ( .B1(n15110), .B2(n15109), .A(n14861), .ZN(n16544) );
  NAND2_X1 U16237 ( .A1(n16550), .A2(n14950), .ZN(n14863) );
  NAND2_X1 U16238 ( .A1(n15130), .A2(n14954), .ZN(n14862) );
  NAND2_X1 U16239 ( .A1(n14863), .A2(n14862), .ZN(n14864) );
  XNOR2_X1 U16240 ( .A(n14864), .B(n14925), .ZN(n14866) );
  AND2_X1 U16241 ( .A1(n15130), .A2(n14955), .ZN(n14865) );
  AOI21_X1 U16242 ( .B1(n16550), .B2(n14954), .A(n14865), .ZN(n14867) );
  NAND2_X1 U16243 ( .A1(n14866), .A2(n14867), .ZN(n15038) );
  INV_X1 U16244 ( .A(n14866), .ZN(n14869) );
  INV_X1 U16245 ( .A(n14867), .ZN(n14868) );
  NAND2_X1 U16246 ( .A1(n14869), .A2(n14868), .ZN(n14870) );
  AND2_X1 U16247 ( .A1(n15038), .A2(n14870), .ZN(n16545) );
  NAND2_X1 U16248 ( .A1(n16544), .A2(n16545), .ZN(n15037) );
  NAND2_X1 U16249 ( .A1(n15037), .A2(n15038), .ZN(n14880) );
  NAND2_X1 U16250 ( .A1(n15508), .A2(n14950), .ZN(n14872) );
  NAND2_X1 U16251 ( .A1(n15129), .A2(n14954), .ZN(n14871) );
  NAND2_X1 U16252 ( .A1(n14872), .A2(n14871), .ZN(n14873) );
  XNOR2_X1 U16253 ( .A(n14873), .B(n14925), .ZN(n14875) );
  AND2_X1 U16254 ( .A1(n15129), .A2(n14955), .ZN(n14874) );
  AOI21_X1 U16255 ( .B1(n15508), .B2(n14900), .A(n14874), .ZN(n14876) );
  NAND2_X1 U16256 ( .A1(n14875), .A2(n14876), .ZN(n15081) );
  INV_X1 U16257 ( .A(n14875), .ZN(n14878) );
  INV_X1 U16258 ( .A(n14876), .ZN(n14877) );
  NAND2_X1 U16259 ( .A1(n14878), .A2(n14877), .ZN(n14879) );
  AND2_X1 U16260 ( .A1(n15081), .A2(n14879), .ZN(n15039) );
  NAND2_X1 U16261 ( .A1(n14880), .A2(n15039), .ZN(n15042) );
  NAND2_X1 U16262 ( .A1(n15042), .A2(n15081), .ZN(n14890) );
  NAND2_X1 U16263 ( .A1(n15500), .A2(n14950), .ZN(n14882) );
  NAND2_X1 U16264 ( .A1(n15128), .A2(n14954), .ZN(n14881) );
  NAND2_X1 U16265 ( .A1(n14882), .A2(n14881), .ZN(n14883) );
  XNOR2_X1 U16266 ( .A(n14883), .B(n14925), .ZN(n14885) );
  AND2_X1 U16267 ( .A1(n15128), .A2(n14955), .ZN(n14884) );
  AOI21_X1 U16268 ( .B1(n15500), .B2(n14900), .A(n14884), .ZN(n14886) );
  NAND2_X1 U16269 ( .A1(n14885), .A2(n14886), .ZN(n14891) );
  INV_X1 U16270 ( .A(n14885), .ZN(n14888) );
  INV_X1 U16271 ( .A(n14886), .ZN(n14887) );
  NAND2_X1 U16272 ( .A1(n14888), .A2(n14887), .ZN(n14889) );
  AND2_X1 U16273 ( .A1(n14891), .A2(n14889), .ZN(n15082) );
  NAND2_X1 U16274 ( .A1(n14890), .A2(n15082), .ZN(n15085) );
  NAND2_X1 U16275 ( .A1(n15370), .A2(n14950), .ZN(n14893) );
  OR2_X1 U16276 ( .A1(n15088), .A2(n15005), .ZN(n14892) );
  NAND2_X1 U16277 ( .A1(n14893), .A2(n14892), .ZN(n14894) );
  XNOR2_X1 U16278 ( .A(n14894), .B(n15001), .ZN(n14901) );
  NOR2_X1 U16279 ( .A1(n15088), .A2(n15003), .ZN(n14895) );
  AOI21_X1 U16280 ( .B1(n15370), .B2(n14954), .A(n14895), .ZN(n14902) );
  XNOR2_X1 U16281 ( .A(n14901), .B(n14902), .ZN(n14992) );
  NAND2_X1 U16282 ( .A1(n15484), .A2(n14950), .ZN(n14897) );
  NAND2_X1 U16283 ( .A1(n15126), .A2(n14954), .ZN(n14896) );
  NAND2_X1 U16284 ( .A1(n14897), .A2(n14896), .ZN(n14898) );
  XNOR2_X1 U16285 ( .A(n14898), .B(n15001), .ZN(n14916) );
  AND2_X1 U16286 ( .A1(n15126), .A2(n14955), .ZN(n14899) );
  AOI21_X1 U16287 ( .B1(n15484), .B2(n14900), .A(n14899), .ZN(n14914) );
  XNOR2_X1 U16288 ( .A(n14916), .B(n14914), .ZN(n15063) );
  INV_X1 U16289 ( .A(n14901), .ZN(n14903) );
  NAND2_X1 U16290 ( .A1(n14903), .A2(n14902), .ZN(n15064) );
  AND2_X1 U16291 ( .A1(n15063), .A2(n15064), .ZN(n14904) );
  NAND2_X1 U16292 ( .A1(n15334), .A2(n14950), .ZN(n14906) );
  NAND2_X1 U16293 ( .A1(n15125), .A2(n14954), .ZN(n14905) );
  NAND2_X1 U16294 ( .A1(n14906), .A2(n14905), .ZN(n14907) );
  XNOR2_X1 U16295 ( .A(n14907), .B(n14925), .ZN(n14909) );
  AND2_X1 U16296 ( .A1(n15125), .A2(n14955), .ZN(n14908) );
  AOI21_X1 U16297 ( .B1(n15334), .B2(n14954), .A(n14908), .ZN(n14910) );
  NAND2_X1 U16298 ( .A1(n14909), .A2(n14910), .ZN(n15073) );
  INV_X1 U16299 ( .A(n14909), .ZN(n14912) );
  INV_X1 U16300 ( .A(n14910), .ZN(n14911) );
  NAND2_X1 U16301 ( .A1(n14912), .A2(n14911), .ZN(n14913) );
  NAND2_X1 U16302 ( .A1(n15073), .A2(n14913), .ZN(n15018) );
  INV_X1 U16303 ( .A(n14914), .ZN(n14915) );
  AND2_X1 U16304 ( .A1(n14916), .A2(n14915), .ZN(n15017) );
  NOR2_X1 U16305 ( .A1(n15018), .A2(n15017), .ZN(n14917) );
  OAI22_X1 U16306 ( .A1(n15326), .A2(n15000), .B1(n14919), .B2(n15005), .ZN(
        n14918) );
  XNOR2_X1 U16307 ( .A(n14918), .B(n15001), .ZN(n14921) );
  OAI22_X1 U16308 ( .A1(n15326), .A2(n15005), .B1(n14919), .B2(n15003), .ZN(
        n14920) );
  NAND2_X1 U16309 ( .A1(n14921), .A2(n14920), .ZN(n14922) );
  NAND2_X1 U16310 ( .A1(n14970), .A2(n14971), .ZN(n14934) );
  NAND2_X1 U16311 ( .A1(n14928), .A2(n14950), .ZN(n14924) );
  NAND2_X1 U16312 ( .A1(n15123), .A2(n14954), .ZN(n14923) );
  NAND2_X1 U16313 ( .A1(n14924), .A2(n14923), .ZN(n14926) );
  XNOR2_X1 U16314 ( .A(n14926), .B(n14925), .ZN(n14929) );
  NOR2_X1 U16315 ( .A1(n15057), .A2(n15003), .ZN(n14927) );
  AOI21_X1 U16316 ( .B1(n14928), .B2(n14954), .A(n14927), .ZN(n14930) );
  NAND2_X1 U16317 ( .A1(n14929), .A2(n14930), .ZN(n15051) );
  INV_X1 U16318 ( .A(n14929), .ZN(n14932) );
  INV_X1 U16319 ( .A(n14930), .ZN(n14931) );
  NAND2_X1 U16320 ( .A1(n14932), .A2(n14931), .ZN(n14933) );
  AND2_X1 U16321 ( .A1(n15051), .A2(n14933), .ZN(n14972) );
  INV_X1 U16322 ( .A(n14935), .ZN(n14938) );
  INV_X1 U16323 ( .A(n14936), .ZN(n14937) );
  NAND2_X1 U16324 ( .A1(n14938), .A2(n14937), .ZN(n14939) );
  AND2_X1 U16325 ( .A1(n14940), .A2(n14939), .ZN(n15052) );
  NAND2_X1 U16326 ( .A1(n9544), .A2(n11038), .ZN(n14942) );
  NAND2_X1 U16327 ( .A1(n15121), .A2(n14954), .ZN(n14941) );
  NAND2_X1 U16328 ( .A1(n14942), .A2(n14941), .ZN(n14943) );
  XNOR2_X1 U16329 ( .A(n14943), .B(n15001), .ZN(n14947) );
  NAND2_X1 U16330 ( .A1(n9544), .A2(n14954), .ZN(n14945) );
  NAND2_X1 U16331 ( .A1(n15121), .A2(n14955), .ZN(n14944) );
  NAND2_X1 U16332 ( .A1(n14945), .A2(n14944), .ZN(n14946) );
  NOR2_X1 U16333 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  AOI21_X1 U16334 ( .B1(n14947), .B2(n14946), .A(n14948), .ZN(n15027) );
  INV_X1 U16335 ( .A(n14948), .ZN(n14949) );
  NAND2_X1 U16336 ( .A1(n15274), .A2(n14950), .ZN(n14952) );
  NAND2_X1 U16337 ( .A1(n15120), .A2(n14954), .ZN(n14951) );
  NAND2_X1 U16338 ( .A1(n14952), .A2(n14951), .ZN(n14953) );
  XNOR2_X1 U16339 ( .A(n14953), .B(n15001), .ZN(n14959) );
  NAND2_X1 U16340 ( .A1(n15274), .A2(n14954), .ZN(n14957) );
  NAND2_X1 U16341 ( .A1(n14955), .A2(n15120), .ZN(n14956) );
  NAND2_X1 U16342 ( .A1(n14957), .A2(n14956), .ZN(n14958) );
  NOR2_X1 U16343 ( .A1(n14959), .A2(n14958), .ZN(n14960) );
  AOI21_X1 U16344 ( .B1(n14959), .B2(n14958), .A(n14960), .ZN(n15097) );
  NAND2_X1 U16345 ( .A1(n15096), .A2(n15097), .ZN(n15095) );
  INV_X1 U16346 ( .A(n14960), .ZN(n14961) );
  OAI21_X1 U16347 ( .B1(n14963), .B2(n14962), .A(n14999), .ZN(n14964) );
  INV_X1 U16348 ( .A(n14964), .ZN(n14969) );
  OAI22_X1 U16349 ( .A1(n14965), .A2(n15399), .B1(n15004), .B2(n15401), .ZN(
        n15249) );
  AOI22_X1 U16350 ( .A1(n16548), .A2(n15249), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14966) );
  OAI21_X1 U16351 ( .B1(n16555), .B2(n15254), .A(n14966), .ZN(n14967) );
  AOI21_X1 U16352 ( .B1(n15436), .B2(n16551), .A(n14967), .ZN(n14968) );
  OAI21_X1 U16353 ( .B1(n14969), .B2(n15115), .A(n14968), .ZN(P1_U3214) );
  INV_X1 U16354 ( .A(n14970), .ZN(n15075) );
  INV_X1 U16355 ( .A(n14971), .ZN(n14973) );
  NOR3_X1 U16356 ( .A1(n15075), .A2(n14973), .A3(n14972), .ZN(n14975) );
  INV_X1 U16357 ( .A(n15054), .ZN(n14974) );
  OAI21_X1 U16358 ( .B1(n14975), .B2(n14974), .A(n16546), .ZN(n14980) );
  INV_X1 U16359 ( .A(n14976), .ZN(n15309) );
  AOI22_X1 U16360 ( .A1(n15122), .A2(n15099), .B1(n15100), .B2(n15124), .ZN(
        n15462) );
  INV_X1 U16361 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14977) );
  OAI22_X1 U16362 ( .A1(n15462), .A2(n15102), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14977), .ZN(n14978) );
  AOI21_X1 U16363 ( .B1(n15104), .B2(n15309), .A(n14978), .ZN(n14979) );
  OAI211_X1 U16364 ( .C1(n15464), .C2(n15108), .A(n14980), .B(n14979), .ZN(
        P1_U3216) );
  AOI21_X1 U16365 ( .B1(n14982), .B2(n14981), .A(n15115), .ZN(n14984) );
  NAND2_X1 U16366 ( .A1(n14984), .A2(n14983), .ZN(n14990) );
  AOI22_X1 U16367 ( .A1(n16548), .A2(n14986), .B1(n16551), .B2(n14985), .ZN(
        n14989) );
  MUX2_X1 U16368 ( .A(P1_STATE_REG_SCAN_IN), .B(n16555), .S(n14987), .Z(n14988) );
  NAND3_X1 U16369 ( .A1(n14990), .A2(n14989), .A3(n14988), .ZN(P1_U3218) );
  OAI21_X1 U16370 ( .B1(n14992), .B2(n14991), .A(n15065), .ZN(n14993) );
  NAND2_X1 U16371 ( .A1(n14993), .A2(n16546), .ZN(n14997) );
  AOI22_X1 U16372 ( .A1(n15126), .A2(n15099), .B1(n15100), .B2(n15128), .ZN(
        n15492) );
  NAND2_X1 U16373 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15234)
         );
  OAI21_X1 U16374 ( .B1(n15492), .B2(n15102), .A(n15234), .ZN(n14994) );
  AOI21_X1 U16375 ( .B1(n14995), .B2(n15104), .A(n14994), .ZN(n14996) );
  OAI211_X1 U16376 ( .C1(n15494), .C2(n15108), .A(n14997), .B(n14996), .ZN(
        P1_U3219) );
  OAI22_X1 U16377 ( .A1(n15006), .A2(n15000), .B1(n15004), .B2(n15005), .ZN(
        n15002) );
  XNOR2_X1 U16378 ( .A(n15002), .B(n15001), .ZN(n15008) );
  OAI22_X1 U16379 ( .A1(n15006), .A2(n15005), .B1(n15004), .B2(n15003), .ZN(
        n15007) );
  XNOR2_X1 U16380 ( .A(n15008), .B(n15007), .ZN(n15009) );
  OAI22_X1 U16381 ( .A1(n15102), .A2(n15011), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15010), .ZN(n15012) );
  AOI21_X1 U16382 ( .B1(n15104), .B2(n15013), .A(n15012), .ZN(n15015) );
  NAND2_X1 U16383 ( .A1(n15428), .A2(n16551), .ZN(n15014) );
  OAI211_X1 U16384 ( .C1(n15016), .C2(n15115), .A(n15015), .B(n15014), .ZN(
        P1_U3220) );
  INV_X1 U16385 ( .A(n15334), .ZN(n15476) );
  INV_X1 U16386 ( .A(n15017), .ZN(n15020) );
  INV_X1 U16387 ( .A(n15018), .ZN(n15019) );
  AOI21_X1 U16388 ( .B1(n15062), .B2(n15020), .A(n15019), .ZN(n15021) );
  OAI21_X1 U16389 ( .B1(n7395), .B2(n15021), .A(n16546), .ZN(n15025) );
  AOI22_X1 U16390 ( .A1(n15126), .A2(n15100), .B1(n15099), .B2(n15124), .ZN(
        n15475) );
  INV_X1 U16391 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15022) );
  OAI22_X1 U16392 ( .A1(n15475), .A2(n15102), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15022), .ZN(n15023) );
  AOI21_X1 U16393 ( .B1(n15338), .B2(n15104), .A(n15023), .ZN(n15024) );
  OAI211_X1 U16394 ( .C1(n15476), .C2(n15108), .A(n15025), .B(n15024), .ZN(
        P1_U3223) );
  INV_X1 U16395 ( .A(n9544), .ZN(n15450) );
  NOR3_X1 U16396 ( .A1(n15027), .A2(n15026), .A3(n15053), .ZN(n15030) );
  INV_X1 U16397 ( .A(n15028), .ZN(n15029) );
  OAI21_X1 U16398 ( .B1(n15030), .B2(n15029), .A(n16546), .ZN(n15036) );
  INV_X1 U16399 ( .A(n15031), .ZN(n15285) );
  AND2_X1 U16400 ( .A1(n15120), .A2(n15099), .ZN(n15032) );
  AOI21_X1 U16401 ( .B1(n15122), .B2(n15100), .A(n15032), .ZN(n15448) );
  INV_X1 U16402 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15033) );
  OAI22_X1 U16403 ( .A1(n15448), .A2(n15102), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15033), .ZN(n15034) );
  AOI21_X1 U16404 ( .B1(n15104), .B2(n15285), .A(n15034), .ZN(n15035) );
  OAI211_X1 U16405 ( .C1(n15450), .C2(n15108), .A(n15036), .B(n15035), .ZN(
        P1_U3225) );
  INV_X1 U16406 ( .A(n15037), .ZN(n15041) );
  INV_X1 U16407 ( .A(n15038), .ZN(n15040) );
  NOR3_X1 U16408 ( .A1(n15041), .A2(n15040), .A3(n15039), .ZN(n15043) );
  INV_X1 U16409 ( .A(n15042), .ZN(n15084) );
  OAI21_X1 U16410 ( .B1(n15043), .B2(n15084), .A(n16546), .ZN(n15049) );
  INV_X1 U16411 ( .A(n15044), .ZN(n15047) );
  OAI21_X1 U16412 ( .B1(n15509), .B2(n15102), .A(n15045), .ZN(n15046) );
  AOI21_X1 U16413 ( .B1(n15047), .B2(n15104), .A(n15046), .ZN(n15048) );
  OAI211_X1 U16414 ( .C1(n15050), .C2(n15108), .A(n15049), .B(n15048), .ZN(
        P1_U3228) );
  NOR2_X1 U16415 ( .A1(n15052), .A2(n7687), .ZN(n15055) );
  AOI21_X1 U16416 ( .B1(n15055), .B2(n15054), .A(n15053), .ZN(n15061) );
  OAI22_X1 U16417 ( .A1(n15057), .A2(n15399), .B1(n15056), .B2(n15401), .ZN(
        n15456) );
  AOI22_X1 U16418 ( .A1(n16548), .A2(n15456), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15058) );
  OAI21_X1 U16419 ( .B1(n16555), .B2(n15295), .A(n15058), .ZN(n15059) );
  AOI21_X1 U16420 ( .B1(n15457), .B2(n16551), .A(n15059), .ZN(n15060) );
  OAI21_X1 U16421 ( .B1(n15061), .B2(n15115), .A(n15060), .ZN(P1_U3229) );
  NAND2_X1 U16422 ( .A1(n15062), .A2(n16546), .ZN(n15072) );
  AOI21_X1 U16423 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n15071) );
  NAND2_X1 U16424 ( .A1(n15125), .A2(n15099), .ZN(n15067) );
  OR2_X1 U16425 ( .A1(n15088), .A2(n15399), .ZN(n15066) );
  NAND2_X1 U16426 ( .A1(n15067), .A2(n15066), .ZN(n15483) );
  AOI22_X1 U16427 ( .A1(n15483), .A2(n16548), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15068) );
  OAI21_X1 U16428 ( .B1(n16555), .B2(n15350), .A(n15068), .ZN(n15069) );
  AOI21_X1 U16429 ( .B1(n15484), .B2(n16551), .A(n15069), .ZN(n15070) );
  OAI21_X1 U16430 ( .B1(n15072), .B2(n15071), .A(n15070), .ZN(P1_U3233) );
  NOR3_X1 U16431 ( .A1(n7395), .A2(n8150), .A3(n15074), .ZN(n15076) );
  OAI21_X1 U16432 ( .B1(n15076), .B2(n15075), .A(n16546), .ZN(n15080) );
  AOI22_X1 U16433 ( .A1(n15125), .A2(n15100), .B1(n15099), .B2(n15123), .ZN(
        n15319) );
  OAI22_X1 U16434 ( .A1(n15319), .A2(n15102), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15077), .ZN(n15078) );
  AOI21_X1 U16435 ( .B1(n15323), .B2(n15104), .A(n15078), .ZN(n15079) );
  OAI211_X1 U16436 ( .C1(n15108), .C2(n15326), .A(n15080), .B(n15079), .ZN(
        P1_U3235) );
  INV_X1 U16437 ( .A(n15081), .ZN(n15083) );
  NOR3_X1 U16438 ( .A1(n15084), .A2(n15083), .A3(n15082), .ZN(n15087) );
  INV_X1 U16439 ( .A(n15085), .ZN(n15086) );
  OAI21_X1 U16440 ( .B1(n15087), .B2(n15086), .A(n16546), .ZN(n15094) );
  OR2_X1 U16441 ( .A1(n15088), .A2(n15401), .ZN(n15090) );
  NAND2_X1 U16442 ( .A1(n15129), .A2(n15100), .ZN(n15089) );
  AND2_X1 U16443 ( .A1(n15090), .A2(n15089), .ZN(n15379) );
  OAI21_X1 U16444 ( .B1(n15379), .B2(n15102), .A(n15091), .ZN(n15092) );
  AOI21_X1 U16445 ( .B1(n15388), .B2(n15104), .A(n15092), .ZN(n15093) );
  OAI211_X1 U16446 ( .C1(n15391), .C2(n15108), .A(n15094), .B(n15093), .ZN(
        P1_U3238) );
  INV_X1 U16447 ( .A(n15274), .ZN(n15441) );
  OAI21_X1 U16448 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n15098) );
  NAND2_X1 U16449 ( .A1(n15098), .A2(n16546), .ZN(n15107) );
  INV_X1 U16450 ( .A(n15270), .ZN(n15105) );
  AOI22_X1 U16451 ( .A1(n15100), .A2(n15121), .B1(n8086), .B2(n15099), .ZN(
        n15440) );
  INV_X1 U16452 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n15101) );
  OAI22_X1 U16453 ( .A1(n15440), .A2(n15102), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15101), .ZN(n15103) );
  AOI21_X1 U16454 ( .B1(n15105), .B2(n15104), .A(n15103), .ZN(n15106) );
  OAI211_X1 U16455 ( .C1(n15441), .C2(n15108), .A(n15107), .B(n15106), .ZN(
        P1_U3240) );
  XNOR2_X1 U16456 ( .A(n15110), .B(n15109), .ZN(n15116) );
  NAND2_X1 U16457 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15710)
         );
  NAND2_X1 U16458 ( .A1(n16527), .A2(n16548), .ZN(n15111) );
  OAI211_X1 U16459 ( .C1(n16555), .C2(n15112), .A(n15710), .B(n15111), .ZN(
        n15113) );
  AOI21_X1 U16460 ( .B1(n16529), .B2(n16551), .A(n15113), .ZN(n15114) );
  OAI21_X1 U16461 ( .B1(n15116), .B2(n15115), .A(n15114), .ZN(P1_U3241) );
  MUX2_X1 U16462 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15238), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16463 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15117), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16464 ( .A(n15118), .B(P1_DATAO_REG_29__SCAN_IN), .S(n15142), .Z(
        P1_U3589) );
  MUX2_X1 U16465 ( .A(n15119), .B(P1_DATAO_REG_28__SCAN_IN), .S(n15142), .Z(
        P1_U3588) );
  MUX2_X1 U16466 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8086), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16467 ( .A(n15120), .B(P1_DATAO_REG_26__SCAN_IN), .S(n15142), .Z(
        P1_U3586) );
  MUX2_X1 U16468 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15121), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16469 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15122), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16470 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15123), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16471 ( .A(n15124), .B(P1_DATAO_REG_22__SCAN_IN), .S(n15142), .Z(
        P1_U3582) );
  MUX2_X1 U16472 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15125), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16473 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15126), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16474 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15127), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16475 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15128), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16476 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15129), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16477 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15130), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16478 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15131), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16479 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15132), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16480 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15133), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16481 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15134), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16482 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15135), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16483 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15136), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16484 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15137), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16485 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15138), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16486 ( .A(n15139), .B(P1_DATAO_REG_6__SCAN_IN), .S(n15142), .Z(
        P1_U3566) );
  MUX2_X1 U16487 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15140), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16488 ( .A(n15141), .B(P1_DATAO_REG_3__SCAN_IN), .S(n15142), .Z(
        P1_U3563) );
  MUX2_X1 U16489 ( .A(n11171), .B(P1_DATAO_REG_2__SCAN_IN), .S(n15142), .Z(
        P1_U3562) );
  MUX2_X1 U16490 ( .A(n15143), .B(P1_DATAO_REG_1__SCAN_IN), .S(n15142), .Z(
        P1_U3561) );
  OAI211_X1 U16491 ( .C1(n15146), .C2(n15145), .A(n7362), .B(n15144), .ZN(
        n15154) );
  AOI22_X1 U16492 ( .A1(n15696), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n15153) );
  OAI211_X1 U16493 ( .C1(n15149), .C2(n15148), .A(n15720), .B(n15147), .ZN(
        n15152) );
  NAND2_X1 U16494 ( .A1(n15722), .A2(n15150), .ZN(n15151) );
  NAND4_X1 U16495 ( .A1(n15154), .A2(n15153), .A3(n15152), .A4(n15151), .ZN(
        P1_U3244) );
  MUX2_X1 U16496 ( .A(n12051), .B(P1_REG2_REG_3__SCAN_IN), .S(n15163), .Z(
        n15155) );
  NAND3_X1 U16497 ( .A1(n15157), .A2(n15156), .A3(n15155), .ZN(n15158) );
  NAND3_X1 U16498 ( .A1(n7362), .A2(n15175), .A3(n15158), .ZN(n15167) );
  NOR2_X1 U16499 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14987), .ZN(n15159) );
  AOI21_X1 U16500 ( .B1(n15696), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n15159), .ZN(
        n15166) );
  OAI211_X1 U16501 ( .C1(n15162), .C2(n15161), .A(n15720), .B(n15160), .ZN(
        n15165) );
  NAND2_X1 U16502 ( .A1(n15722), .A2(n15163), .ZN(n15164) );
  NAND4_X1 U16503 ( .A1(n15167), .A2(n15166), .A3(n15165), .A4(n15164), .ZN(
        P1_U3246) );
  NAND2_X1 U16504 ( .A1(n15696), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n15168) );
  OAI211_X1 U16505 ( .C1(n15704), .C2(n15170), .A(n15169), .B(n15168), .ZN(
        n15171) );
  INV_X1 U16506 ( .A(n15171), .ZN(n15183) );
  MUX2_X1 U16507 ( .A(n11273), .B(P1_REG2_REG_4__SCAN_IN), .S(n15172), .Z(
        n15173) );
  NAND3_X1 U16508 ( .A1(n15175), .A2(n15174), .A3(n15173), .ZN(n15176) );
  NAND3_X1 U16509 ( .A1(n7362), .A2(n15177), .A3(n15176), .ZN(n15182) );
  OAI211_X1 U16510 ( .C1(n15180), .C2(n15179), .A(n15720), .B(n15178), .ZN(
        n15181) );
  NAND4_X1 U16511 ( .A1(n15184), .A2(n15183), .A3(n15182), .A4(n15181), .ZN(
        P1_U3247) );
  OAI21_X1 U16512 ( .B1(n15187), .B2(n15186), .A(n15185), .ZN(n15188) );
  NAND2_X1 U16513 ( .A1(n15188), .A2(n15720), .ZN(n15200) );
  AND2_X1 U16514 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n15189) );
  AOI21_X1 U16515 ( .B1(n15696), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n15189), .ZN(
        n15199) );
  INV_X1 U16516 ( .A(n15190), .ZN(n15192) );
  MUX2_X1 U16517 ( .A(n11316), .B(P1_REG2_REG_8__SCAN_IN), .S(n15196), .Z(
        n15191) );
  NAND2_X1 U16518 ( .A1(n15192), .A2(n15191), .ZN(n15194) );
  OAI211_X1 U16519 ( .C1(n15195), .C2(n15194), .A(n15193), .B(n7362), .ZN(
        n15198) );
  NAND2_X1 U16520 ( .A1(n15722), .A2(n15196), .ZN(n15197) );
  NAND4_X1 U16521 ( .A1(n15200), .A2(n15199), .A3(n15198), .A4(n15197), .ZN(
        P1_U3251) );
  INV_X1 U16522 ( .A(n15201), .ZN(n15203) );
  MUX2_X1 U16523 ( .A(n12266), .B(P1_REG2_REG_10__SCAN_IN), .S(n15212), .Z(
        n15202) );
  NAND2_X1 U16524 ( .A1(n15203), .A2(n15202), .ZN(n15205) );
  OAI211_X1 U16525 ( .C1(n15206), .C2(n15205), .A(n15204), .B(n7362), .ZN(
        n15216) );
  AOI21_X1 U16526 ( .B1(n15208), .B2(n15207), .A(n15227), .ZN(n15210) );
  NAND2_X1 U16527 ( .A1(n15210), .A2(n15209), .ZN(n15215) );
  AND2_X1 U16528 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n15211) );
  AOI21_X1 U16529 ( .B1(n15696), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n15211), 
        .ZN(n15214) );
  NAND2_X1 U16530 ( .A1(n15722), .A2(n15212), .ZN(n15213) );
  NAND4_X1 U16531 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        P1_U3253) );
  NOR2_X1 U16532 ( .A1(n15217), .A2(n7542), .ZN(n15218) );
  NOR2_X1 U16533 ( .A1(n15219), .A2(n15218), .ZN(n15220) );
  XNOR2_X1 U16534 ( .A(n15220), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n15228) );
  NAND2_X1 U16535 ( .A1(n15222), .A2(n15221), .ZN(n15224) );
  NAND2_X1 U16536 ( .A1(n15224), .A2(n15223), .ZN(n15225) );
  XOR2_X1 U16537 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n15225), .Z(n15226) );
  AOI22_X1 U16538 ( .A1(n15228), .A2(n15720), .B1(n7362), .B2(n15226), .ZN(
        n15233) );
  INV_X1 U16539 ( .A(n15226), .ZN(n15230) );
  NOR2_X1 U16540 ( .A1(n15228), .A2(n15227), .ZN(n15229) );
  AOI211_X1 U16541 ( .C1(n15231), .C2(n15230), .A(n15722), .B(n15229), .ZN(
        n15232) );
  MUX2_X1 U16542 ( .A(n15233), .B(n15232), .S(n7363), .Z(n15235) );
  OAI211_X1 U16543 ( .C1(n8581), .C2(n15728), .A(n15235), .B(n15234), .ZN(
        P1_U3262) );
  NAND2_X1 U16544 ( .A1(n15242), .A2(n15418), .ZN(n15236) );
  XNOR2_X1 U16545 ( .A(n15236), .B(n15415), .ZN(n15413) );
  NAND2_X1 U16546 ( .A1(n15413), .A2(n15387), .ZN(n15240) );
  NAND2_X1 U16547 ( .A1(n15238), .A2(n15237), .ZN(n15416) );
  NOR2_X1 U16548 ( .A1(n16153), .A2(n15416), .ZN(n15245) );
  AOI21_X1 U16549 ( .B1(n16153), .B2(P1_REG2_REG_31__SCAN_IN), .A(n15245), 
        .ZN(n15239) );
  OAI211_X1 U16550 ( .C1(n15415), .C2(n16156), .A(n15240), .B(n15239), .ZN(
        P1_U3263) );
  XNOR2_X1 U16551 ( .A(n15242), .B(n15241), .ZN(n15243) );
  NAND2_X1 U16552 ( .A1(n15243), .A2(n15501), .ZN(n15417) );
  NOR2_X1 U16553 ( .A1(n15418), .A2(n16156), .ZN(n15244) );
  AOI211_X1 U16554 ( .C1(n16153), .C2(P1_REG2_REG_30__SCAN_IN), .A(n15245), 
        .B(n15244), .ZN(n15246) );
  OAI21_X1 U16555 ( .B1(n15417), .B2(n15372), .A(n15246), .ZN(P1_U3264) );
  XNOR2_X1 U16556 ( .A(n15248), .B(n15247), .ZN(n15250) );
  AOI21_X1 U16557 ( .B1(n15250), .B2(n16248), .A(n15249), .ZN(n15438) );
  INV_X1 U16558 ( .A(n15268), .ZN(n15253) );
  INV_X1 U16559 ( .A(n15251), .ZN(n15252) );
  AOI211_X1 U16560 ( .C1(n15436), .C2(n15253), .A(n16495), .B(n15252), .ZN(
        n15435) );
  INV_X1 U16561 ( .A(n15254), .ZN(n15255) );
  AOI22_X1 U16562 ( .A1(n16153), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n15255), 
        .B2(n16312), .ZN(n15256) );
  OAI21_X1 U16563 ( .B1(n15257), .B2(n16156), .A(n15256), .ZN(n15264) );
  INV_X1 U16564 ( .A(n15260), .ZN(n15261) );
  AOI21_X1 U16565 ( .B1(n15262), .B2(n15259), .A(n15261), .ZN(n15439) );
  NOR2_X1 U16566 ( .A1(n15439), .A2(n15412), .ZN(n15263) );
  AOI211_X1 U16567 ( .C1(n15435), .C2(n16317), .A(n15264), .B(n15263), .ZN(
        n15265) );
  OAI21_X1 U16568 ( .B1(n16153), .B2(n15438), .A(n15265), .ZN(P1_U3266) );
  XNOR2_X1 U16569 ( .A(n15266), .B(n7726), .ZN(n15442) );
  XNOR2_X1 U16570 ( .A(n15267), .B(n7726), .ZN(n15447) );
  AOI21_X1 U16571 ( .B1(n15274), .B2(n15284), .A(n15268), .ZN(n15445) );
  INV_X1 U16572 ( .A(n15269), .ZN(n15407) );
  OAI21_X1 U16573 ( .B1(n15270), .B2(n16104), .A(n15440), .ZN(n15271) );
  AOI21_X1 U16574 ( .B1(n15445), .B2(n15407), .A(n15271), .ZN(n15272) );
  OAI21_X1 U16575 ( .B1(n15447), .B2(n15345), .A(n15272), .ZN(n15273) );
  NAND2_X1 U16576 ( .A1(n15273), .A2(n15352), .ZN(n15276) );
  AOI22_X1 U16577 ( .A1(n15274), .A2(n16313), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n16153), .ZN(n15275) );
  OAI211_X1 U16578 ( .C1(n15442), .C2(n15412), .A(n15276), .B(n15275), .ZN(
        P1_U3267) );
  OAI21_X1 U16579 ( .B1(n15278), .B2(n7380), .A(n15277), .ZN(n15279) );
  INV_X1 U16580 ( .A(n15279), .ZN(n15454) );
  INV_X1 U16581 ( .A(n15281), .ZN(n15282) );
  AOI21_X1 U16582 ( .B1(n7380), .B2(n15280), .A(n15282), .ZN(n15452) );
  NAND2_X1 U16583 ( .A1(n9544), .A2(n15293), .ZN(n15283) );
  NAND3_X1 U16584 ( .A1(n15284), .A2(n15501), .A3(n15283), .ZN(n15449) );
  NAND2_X1 U16585 ( .A1(n16312), .A2(n15285), .ZN(n15287) );
  NAND2_X1 U16586 ( .A1(n16153), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n15286) );
  OAI211_X1 U16587 ( .C1(n15448), .C2(n16153), .A(n15287), .B(n15286), .ZN(
        n15288) );
  AOI21_X1 U16588 ( .B1(n9544), .B2(n16313), .A(n15288), .ZN(n15289) );
  OAI21_X1 U16589 ( .B1(n15449), .B2(n15372), .A(n15289), .ZN(n15290) );
  AOI21_X1 U16590 ( .B1(n15452), .B2(n15393), .A(n15290), .ZN(n15291) );
  OAI21_X1 U16591 ( .B1(n15454), .B2(n15345), .A(n15291), .ZN(P1_U3268) );
  AOI21_X1 U16592 ( .B1(n15292), .B2(n7644), .A(n7426), .ZN(n15461) );
  INV_X1 U16593 ( .A(n15293), .ZN(n15294) );
  AOI211_X1 U16594 ( .C1(n15457), .C2(n15308), .A(n16495), .B(n15294), .ZN(
        n15455) );
  INV_X1 U16595 ( .A(n15456), .ZN(n15296) );
  OAI22_X1 U16596 ( .A1(n15296), .A2(n16153), .B1(n15295), .B2(n16104), .ZN(
        n15297) );
  AOI21_X1 U16597 ( .B1(P1_REG2_REG_24__SCAN_IN), .B2(n16153), .A(n15297), 
        .ZN(n15298) );
  OAI21_X1 U16598 ( .B1(n15299), .B2(n16156), .A(n15298), .ZN(n15300) );
  AOI21_X1 U16599 ( .B1(n15455), .B2(n16317), .A(n15300), .ZN(n15304) );
  NAND2_X1 U16600 ( .A1(n15302), .A2(n13055), .ZN(n15458) );
  NAND3_X1 U16601 ( .A1(n8266), .A2(n15374), .A3(n15458), .ZN(n15303) );
  OAI211_X1 U16602 ( .C1(n15412), .C2(n15461), .A(n15304), .B(n15303), .ZN(
        P1_U3269) );
  XOR2_X1 U16603 ( .A(n7387), .B(n15305), .Z(n15468) );
  XNOR2_X1 U16604 ( .A(n15306), .B(n15305), .ZN(n15466) );
  NAND2_X1 U16605 ( .A1(n15466), .A2(n15374), .ZN(n15316) );
  INV_X1 U16606 ( .A(n15307), .ZN(n15321) );
  OAI211_X1 U16607 ( .C1(n15464), .C2(n15321), .A(n15308), .B(n15501), .ZN(
        n15463) );
  NAND2_X1 U16608 ( .A1(n16312), .A2(n15309), .ZN(n15310) );
  OAI211_X1 U16609 ( .C1(n15463), .C2(n7363), .A(n15462), .B(n15310), .ZN(
        n15314) );
  INV_X1 U16610 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n15312) );
  OAI22_X1 U16611 ( .A1(n15464), .A2(n16156), .B1(n15352), .B2(n15312), .ZN(
        n15313) );
  AOI21_X1 U16612 ( .B1(n15314), .B2(n15352), .A(n15313), .ZN(n15315) );
  OAI211_X1 U16613 ( .C1(n15468), .C2(n15412), .A(n15316), .B(n15315), .ZN(
        P1_U3270) );
  XNOR2_X1 U16614 ( .A(n15318), .B(n7460), .ZN(n15474) );
  AOI21_X1 U16615 ( .B1(n15318), .B2(n15317), .A(n7441), .ZN(n15320) );
  OAI21_X1 U16616 ( .B1(n15320), .B2(n16532), .A(n15319), .ZN(n15469) );
  INV_X1 U16617 ( .A(n15337), .ZN(n15322) );
  AOI21_X1 U16618 ( .B1(n15470), .B2(n15322), .A(n15321), .ZN(n15471) );
  NAND2_X1 U16619 ( .A1(n15471), .A2(n15387), .ZN(n15325) );
  AOI22_X1 U16620 ( .A1(n16153), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n15323), 
        .B2(n16312), .ZN(n15324) );
  OAI211_X1 U16621 ( .C1(n16156), .C2(n15326), .A(n15325), .B(n15324), .ZN(
        n15327) );
  AOI21_X1 U16622 ( .B1(n15469), .B2(n15352), .A(n15327), .ZN(n15328) );
  OAI21_X1 U16623 ( .B1(n15474), .B2(n15412), .A(n15328), .ZN(P1_U3271) );
  OAI21_X1 U16624 ( .B1(n15331), .B2(n15330), .A(n15329), .ZN(n15481) );
  NAND2_X1 U16625 ( .A1(n15334), .A2(n15349), .ZN(n15335) );
  NAND2_X1 U16626 ( .A1(n15335), .A2(n15501), .ZN(n15336) );
  NOR2_X1 U16627 ( .A1(n15337), .A2(n15336), .ZN(n15477) );
  NAND2_X1 U16628 ( .A1(n15477), .A2(n16317), .ZN(n15342) );
  INV_X1 U16629 ( .A(n15338), .ZN(n15339) );
  OAI22_X1 U16630 ( .A1(n15475), .A2(n16153), .B1(n15339), .B2(n16104), .ZN(
        n15340) );
  AOI21_X1 U16631 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(n16153), .A(n15340), 
        .ZN(n15341) );
  OAI211_X1 U16632 ( .C1(n15476), .C2(n16156), .A(n15342), .B(n15341), .ZN(
        n15343) );
  AOI21_X1 U16633 ( .B1(n15393), .B2(n15479), .A(n15343), .ZN(n15344) );
  OAI21_X1 U16634 ( .B1(n15345), .B2(n15481), .A(n15344), .ZN(P1_U3272) );
  OR2_X1 U16635 ( .A1(n15346), .A2(n15359), .ZN(n15482) );
  NAND3_X1 U16636 ( .A1(n15482), .A2(n15374), .A3(n15347), .ZN(n15362) );
  NAND2_X1 U16637 ( .A1(n15484), .A2(n15365), .ZN(n15348) );
  NAND2_X1 U16638 ( .A1(n15484), .A2(n16313), .ZN(n15354) );
  INV_X1 U16639 ( .A(n15350), .ZN(n15351) );
  AOI22_X1 U16640 ( .A1(n15483), .A2(n15352), .B1(n15351), .B2(n16312), .ZN(
        n15353) );
  OAI211_X1 U16641 ( .C1(n15356), .C2(n15355), .A(n15354), .B(n15353), .ZN(
        n15357) );
  AOI21_X1 U16642 ( .B1(n15487), .B2(n15387), .A(n15357), .ZN(n15361) );
  NAND2_X1 U16643 ( .A1(n15359), .A2(n15358), .ZN(n15485) );
  NAND3_X1 U16644 ( .A1(n15486), .A2(n15485), .A3(n15393), .ZN(n15360) );
  NAND3_X1 U16645 ( .A1(n15362), .A2(n15361), .A3(n15360), .ZN(P1_U3273) );
  XNOR2_X1 U16646 ( .A(n15364), .B(n15363), .ZN(n15498) );
  OAI21_X1 U16647 ( .B1(n7389), .B2(n15364), .A(n7491), .ZN(n15496) );
  OAI211_X1 U16648 ( .C1(n15494), .C2(n15386), .A(n15501), .B(n15365), .ZN(
        n15493) );
  NOR2_X1 U16649 ( .A1(n15352), .A2(n15366), .ZN(n15369) );
  OAI22_X1 U16650 ( .A1(n15492), .A2(n16153), .B1(n15367), .B2(n16104), .ZN(
        n15368) );
  AOI211_X1 U16651 ( .C1(n15370), .C2(n16313), .A(n15369), .B(n15368), .ZN(
        n15371) );
  OAI21_X1 U16652 ( .B1(n15493), .B2(n15372), .A(n15371), .ZN(n15373) );
  AOI21_X1 U16653 ( .B1(n15496), .B2(n15374), .A(n15373), .ZN(n15375) );
  OAI21_X1 U16654 ( .B1(n15412), .B2(n15498), .A(n15375), .ZN(P1_U3274) );
  OAI211_X1 U16655 ( .C1(n15378), .C2(n15377), .A(n15376), .B(n16248), .ZN(
        n15380) );
  OAI21_X1 U16656 ( .B1(n15383), .B2(n15382), .A(n15381), .ZN(n15499) );
  AND2_X1 U16657 ( .A1(n15500), .A2(n15384), .ZN(n15385) );
  NOR2_X1 U16658 ( .A1(n15386), .A2(n15385), .ZN(n15502) );
  NAND2_X1 U16659 ( .A1(n15502), .A2(n15387), .ZN(n15390) );
  AOI22_X1 U16660 ( .A1(n16153), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15388), 
        .B2(n16312), .ZN(n15389) );
  OAI211_X1 U16661 ( .C1(n15391), .C2(n16156), .A(n15390), .B(n15389), .ZN(
        n15392) );
  AOI21_X1 U16662 ( .B1(n15393), .B2(n15499), .A(n15392), .ZN(n15394) );
  OAI21_X1 U16663 ( .B1(n16153), .B2(n15504), .A(n15394), .ZN(P1_U3275) );
  XOR2_X1 U16664 ( .A(n15395), .B(n15397), .Z(n15519) );
  OAI22_X1 U16665 ( .A1(n15352), .A2(n15396), .B1(n16554), .B2(n16104), .ZN(
        n15410) );
  OAI21_X1 U16666 ( .B1(n7498), .B2(n12956), .A(n15398), .ZN(n15403) );
  OAI22_X1 U16667 ( .A1(n15402), .A2(n15401), .B1(n15400), .B2(n15399), .ZN(
        n16549) );
  AOI21_X1 U16668 ( .B1(n15403), .B2(n16248), .A(n16549), .ZN(n15518) );
  INV_X1 U16669 ( .A(n15404), .ZN(n15405) );
  AOI21_X1 U16670 ( .B1(n16550), .B2(n15406), .A(n15405), .ZN(n15516) );
  NAND2_X1 U16671 ( .A1(n15516), .A2(n15407), .ZN(n15408) );
  AOI21_X1 U16672 ( .B1(n15518), .B2(n15408), .A(n16153), .ZN(n15409) );
  AOI211_X1 U16673 ( .C1(n16313), .C2(n16550), .A(n15410), .B(n15409), .ZN(
        n15411) );
  OAI21_X1 U16674 ( .B1(n15412), .B2(n15519), .A(n15411), .ZN(P1_U3277) );
  NAND2_X1 U16675 ( .A1(n15413), .A2(n15501), .ZN(n15414) );
  OAI211_X1 U16676 ( .C1(n16448), .C2(n15415), .A(n15414), .B(n15416), .ZN(
        n15525) );
  MUX2_X1 U16677 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15525), .S(n16539), .Z(
        P1_U3559) );
  OAI211_X1 U16678 ( .C1(n16448), .C2(n15418), .A(n15417), .B(n15416), .ZN(
        n15526) );
  INV_X2 U16679 ( .A(n16537), .ZN(n16539) );
  MUX2_X1 U16680 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15526), .S(n16539), .Z(
        P1_U3558) );
  NAND2_X1 U16681 ( .A1(n15419), .A2(n16248), .ZN(n15427) );
  OAI211_X1 U16682 ( .C1(n15422), .C2(n16448), .A(n15421), .B(n15420), .ZN(
        n15423) );
  AOI21_X1 U16683 ( .B1(n15424), .B2(n15501), .A(n15423), .ZN(n15425) );
  AOI22_X1 U16684 ( .A1(n15429), .A2(n15501), .B1(n15428), .B2(n16528), .ZN(
        n15430) );
  AOI21_X1 U16685 ( .B1(n15436), .B2(n16528), .A(n15435), .ZN(n15437) );
  OAI211_X1 U16686 ( .C1(n16243), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        n15528) );
  MUX2_X1 U16687 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15528), .S(n16539), .Z(
        P1_U3555) );
  OAI21_X1 U16688 ( .B1(n15441), .B2(n16448), .A(n15440), .ZN(n15444) );
  NOR2_X1 U16689 ( .A1(n15442), .A2(n16243), .ZN(n15443) );
  AOI211_X1 U16690 ( .C1(n15501), .C2(n15445), .A(n15444), .B(n15443), .ZN(
        n15446) );
  OAI21_X1 U16691 ( .B1(n16532), .B2(n15447), .A(n15446), .ZN(n15529) );
  MUX2_X1 U16692 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15529), .S(n16539), .Z(
        P1_U3554) );
  OAI211_X1 U16693 ( .C1(n15450), .C2(n16448), .A(n15449), .B(n15448), .ZN(
        n15451) );
  AOI21_X1 U16694 ( .B1(n15452), .B2(n16536), .A(n15451), .ZN(n15453) );
  OAI21_X1 U16695 ( .B1(n15454), .B2(n16532), .A(n15453), .ZN(n15530) );
  MUX2_X1 U16696 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15530), .S(n16539), .Z(
        P1_U3553) );
  AOI211_X1 U16697 ( .C1(n15457), .C2(n16528), .A(n15456), .B(n15455), .ZN(
        n15460) );
  NAND3_X1 U16698 ( .A1(n8266), .A2(n16248), .A3(n15458), .ZN(n15459) );
  OAI211_X1 U16699 ( .C1(n16243), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        n15531) );
  MUX2_X1 U16700 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15531), .S(n16539), .Z(
        P1_U3552) );
  OAI211_X1 U16701 ( .C1(n15464), .C2(n16448), .A(n15463), .B(n15462), .ZN(
        n15465) );
  AOI21_X1 U16702 ( .B1(n15466), .B2(n16248), .A(n15465), .ZN(n15467) );
  OAI21_X1 U16703 ( .B1(n16243), .B2(n15468), .A(n15467), .ZN(n15532) );
  MUX2_X1 U16704 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15532), .S(n16539), .Z(
        P1_U3551) );
  INV_X1 U16705 ( .A(n15469), .ZN(n15473) );
  AOI22_X1 U16706 ( .A1(n15471), .A2(n15501), .B1(n15470), .B2(n16528), .ZN(
        n15472) );
  OAI211_X1 U16707 ( .C1(n16243), .C2(n15474), .A(n15473), .B(n15472), .ZN(
        n15533) );
  MUX2_X1 U16708 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15533), .S(n16539), .Z(
        P1_U3550) );
  OAI21_X1 U16709 ( .B1(n15476), .B2(n16448), .A(n15475), .ZN(n15478) );
  AOI211_X1 U16710 ( .C1(n15479), .C2(n16536), .A(n15478), .B(n15477), .ZN(
        n15480) );
  OAI21_X1 U16711 ( .B1(n16532), .B2(n15481), .A(n15480), .ZN(n15534) );
  MUX2_X1 U16712 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15534), .S(n16539), .Z(
        P1_U3549) );
  NAND3_X1 U16713 ( .A1(n15482), .A2(n16248), .A3(n15347), .ZN(n15491) );
  AOI21_X1 U16714 ( .B1(n15484), .B2(n16528), .A(n15483), .ZN(n15490) );
  NAND3_X1 U16715 ( .A1(n15486), .A2(n16536), .A3(n15485), .ZN(n15489) );
  NAND2_X1 U16716 ( .A1(n15487), .A2(n15501), .ZN(n15488) );
  NAND4_X1 U16717 ( .A1(n15491), .A2(n15490), .A3(n15489), .A4(n15488), .ZN(
        n15535) );
  MUX2_X1 U16718 ( .A(n15535), .B(P1_REG1_REG_20__SCAN_IN), .S(n16537), .Z(
        P1_U3548) );
  OAI211_X1 U16719 ( .C1(n15494), .C2(n16448), .A(n15493), .B(n15492), .ZN(
        n15495) );
  AOI21_X1 U16720 ( .B1(n15496), .B2(n16248), .A(n15495), .ZN(n15497) );
  OAI21_X1 U16721 ( .B1(n16243), .B2(n15498), .A(n15497), .ZN(n15536) );
  MUX2_X1 U16722 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15536), .S(n16539), .Z(
        P1_U3547) );
  INV_X1 U16723 ( .A(n15499), .ZN(n15505) );
  AOI22_X1 U16724 ( .A1(n15502), .A2(n15501), .B1(n15500), .B2(n16528), .ZN(
        n15503) );
  OAI211_X1 U16725 ( .C1(n16243), .C2(n15505), .A(n15504), .B(n15503), .ZN(
        n15537) );
  MUX2_X1 U16726 ( .A(n15537), .B(P1_REG1_REG_18__SCAN_IN), .S(n16537), .Z(
        P1_U3546) );
  NAND3_X1 U16727 ( .A1(n15507), .A2(n16248), .A3(n15506), .ZN(n15514) );
  NAND2_X1 U16728 ( .A1(n15508), .A2(n16528), .ZN(n15510) );
  NAND2_X1 U16729 ( .A1(n15510), .A2(n15509), .ZN(n15511) );
  AOI21_X1 U16730 ( .B1(n15512), .B2(n15501), .A(n15511), .ZN(n15513) );
  OAI211_X1 U16731 ( .C1(n16243), .C2(n15515), .A(n15514), .B(n15513), .ZN(
        n15538) );
  MUX2_X1 U16732 ( .A(n15538), .B(P1_REG1_REG_17__SCAN_IN), .S(n16537), .Z(
        P1_U3545) );
  AOI22_X1 U16733 ( .A1(n15516), .A2(n15501), .B1(n16550), .B2(n16528), .ZN(
        n15517) );
  OAI211_X1 U16734 ( .C1(n16243), .C2(n15519), .A(n15518), .B(n15517), .ZN(
        n15539) );
  MUX2_X1 U16735 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15539), .S(n16539), .Z(
        P1_U3544) );
  AOI211_X1 U16736 ( .C1(n16523), .C2(n16528), .A(n16522), .B(n15520), .ZN(
        n15523) );
  NAND3_X1 U16737 ( .A1(n12714), .A2(n15521), .A3(n16536), .ZN(n15522) );
  OAI211_X1 U16738 ( .C1(n15524), .C2(n16532), .A(n15523), .B(n15522), .ZN(
        n15540) );
  MUX2_X1 U16739 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15540), .S(n16539), .Z(
        P1_U3542) );
  MUX2_X1 U16740 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15525), .S(n16543), .Z(
        P1_U3527) );
  INV_X2 U16741 ( .A(n16540), .ZN(n16543) );
  MUX2_X1 U16742 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15526), .S(n16543), .Z(
        P1_U3526) );
  MUX2_X1 U16743 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15527), .S(n16543), .Z(
        P1_U3524) );
  MUX2_X1 U16744 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15528), .S(n16543), .Z(
        P1_U3523) );
  MUX2_X1 U16745 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15529), .S(n16543), .Z(
        P1_U3522) );
  MUX2_X1 U16746 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15530), .S(n16543), .Z(
        P1_U3521) );
  MUX2_X1 U16747 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15531), .S(n16543), .Z(
        P1_U3520) );
  MUX2_X1 U16748 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15532), .S(n16543), .Z(
        P1_U3519) );
  MUX2_X1 U16749 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15533), .S(n16543), .Z(
        P1_U3518) );
  MUX2_X1 U16750 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15534), .S(n16543), .Z(
        P1_U3517) );
  MUX2_X1 U16751 ( .A(n15535), .B(P1_REG0_REG_20__SCAN_IN), .S(n16540), .Z(
        P1_U3516) );
  MUX2_X1 U16752 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15536), .S(n16543), .Z(
        P1_U3515) );
  MUX2_X1 U16753 ( .A(n15537), .B(P1_REG0_REG_18__SCAN_IN), .S(n16540), .Z(
        P1_U3513) );
  MUX2_X1 U16754 ( .A(n15538), .B(P1_REG0_REG_17__SCAN_IN), .S(n16540), .Z(
        P1_U3510) );
  MUX2_X1 U16755 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15539), .S(n16543), .Z(
        P1_U3507) );
  MUX2_X1 U16756 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15540), .S(n16543), .Z(
        P1_U3501) );
  MUX2_X1 U16757 ( .A(n15541), .B(P1_D_REG_0__SCAN_IN), .S(n15563), .Z(
        P1_U3445) );
  NOR4_X1 U16758 ( .A1(n15543), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15542), .A4(
        P1_U3086), .ZN(n15544) );
  AOI21_X1 U16759 ( .B1(n15545), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15544), 
        .ZN(n15546) );
  OAI21_X1 U16760 ( .B1(n15547), .B2(n15556), .A(n15546), .ZN(P1_U3324) );
  OAI222_X1 U16761 ( .A1(P1_U3086), .A2(n15550), .B1(n15556), .B2(n15549), 
        .C1(n15548), .C2(n15558), .ZN(P1_U3329) );
  OAI222_X1 U16762 ( .A1(n15558), .A2(n15553), .B1(n15556), .B2(n15552), .C1(
        P1_U3086), .C2(n15551), .ZN(P1_U3330) );
  OAI222_X1 U16763 ( .A1(n15558), .A2(n15557), .B1(n15556), .B2(n15555), .C1(
        P1_U3086), .C2(n15554), .ZN(P1_U3331) );
  MUX2_X1 U16764 ( .A(n15560), .B(n15559), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16765 ( .A(n15561), .ZN(n15562) );
  MUX2_X1 U16766 ( .A(n15562), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16767 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15563), .ZN(P1_U3323) );
  AND2_X1 U16768 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15563), .ZN(P1_U3322) );
  AND2_X1 U16769 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15563), .ZN(P1_U3321) );
  AND2_X1 U16770 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15563), .ZN(P1_U3320) );
  AND2_X1 U16771 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15563), .ZN(P1_U3319) );
  AND2_X1 U16772 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15563), .ZN(P1_U3318) );
  AND2_X1 U16773 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15563), .ZN(P1_U3317) );
  AND2_X1 U16774 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15563), .ZN(P1_U3316) );
  AND2_X1 U16775 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15563), .ZN(P1_U3315) );
  AND2_X1 U16776 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15563), .ZN(P1_U3314) );
  AND2_X1 U16777 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15563), .ZN(P1_U3313) );
  AND2_X1 U16778 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15563), .ZN(P1_U3312) );
  AND2_X1 U16779 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15563), .ZN(P1_U3311) );
  AND2_X1 U16780 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15563), .ZN(P1_U3310) );
  AND2_X1 U16781 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15563), .ZN(P1_U3309) );
  AND2_X1 U16782 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15563), .ZN(P1_U3308) );
  AND2_X1 U16783 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15563), .ZN(P1_U3307) );
  AND2_X1 U16784 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15563), .ZN(P1_U3306) );
  AND2_X1 U16785 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15563), .ZN(P1_U3305) );
  AND2_X1 U16786 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15563), .ZN(P1_U3304) );
  AND2_X1 U16787 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15563), .ZN(P1_U3303) );
  AND2_X1 U16788 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15563), .ZN(P1_U3302) );
  AND2_X1 U16789 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15563), .ZN(P1_U3301) );
  AND2_X1 U16790 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15563), .ZN(P1_U3300) );
  AND2_X1 U16791 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15563), .ZN(P1_U3299) );
  AND2_X1 U16792 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15563), .ZN(P1_U3298) );
  AND2_X1 U16793 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15563), .ZN(P1_U3297) );
  AND2_X1 U16794 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15563), .ZN(P1_U3296) );
  AND2_X1 U16795 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15563), .ZN(P1_U3295) );
  AND2_X1 U16796 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15563), .ZN(P1_U3294) );
  INV_X1 U16797 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15565) );
  AOI21_X1 U16798 ( .B1(n15565), .B2(n15568), .A(n15564), .ZN(P2_U3417) );
  AND2_X1 U16799 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15567), .ZN(P2_U3295) );
  AND2_X1 U16800 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15567), .ZN(P2_U3294) );
  AND2_X1 U16801 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15567), .ZN(P2_U3293) );
  AND2_X1 U16802 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15567), .ZN(P2_U3292) );
  AND2_X1 U16803 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15567), .ZN(P2_U3291) );
  AND2_X1 U16804 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15567), .ZN(P2_U3290) );
  AND2_X1 U16805 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15567), .ZN(P2_U3289) );
  AND2_X1 U16806 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15567), .ZN(P2_U3288) );
  AND2_X1 U16807 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15567), .ZN(P2_U3287) );
  AND2_X1 U16808 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15567), .ZN(P2_U3286) );
  AND2_X1 U16809 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15567), .ZN(P2_U3285) );
  AND2_X1 U16810 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15567), .ZN(P2_U3284) );
  AND2_X1 U16811 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15567), .ZN(P2_U3283) );
  AND2_X1 U16812 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15567), .ZN(P2_U3282) );
  AND2_X1 U16813 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15567), .ZN(P2_U3281) );
  AND2_X1 U16814 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15567), .ZN(P2_U3280) );
  AND2_X1 U16815 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15567), .ZN(P2_U3279) );
  AND2_X1 U16816 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15567), .ZN(P2_U3278) );
  AND2_X1 U16817 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15567), .ZN(P2_U3277) );
  AND2_X1 U16818 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15567), .ZN(P2_U3276) );
  AND2_X1 U16819 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15567), .ZN(P2_U3275) );
  AND2_X1 U16820 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15567), .ZN(P2_U3274) );
  AND2_X1 U16821 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15567), .ZN(P2_U3273) );
  AND2_X1 U16822 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15567), .ZN(P2_U3272) );
  AND2_X1 U16823 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15567), .ZN(P2_U3271) );
  AND2_X1 U16824 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15567), .ZN(P2_U3270) );
  AND2_X1 U16825 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15567), .ZN(P2_U3269) );
  AND2_X1 U16826 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15567), .ZN(P2_U3268) );
  AND2_X1 U16827 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15567), .ZN(P2_U3267) );
  AND2_X1 U16828 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15567), .ZN(P2_U3266) );
  NOR2_X1 U16829 ( .A1(n15684), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16830 ( .A1(P3_U3897), .A2(n16073), .ZN(P3_U3150) );
  INV_X1 U16831 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15569) );
  AOI22_X1 U16832 ( .A1(n15571), .A2(n15570), .B1(n15569), .B2(n15568), .ZN(
        P2_U3416) );
  AOI22_X1 U16833 ( .A1(n15678), .A2(n15572), .B1(n15684), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n15582) );
  NAND2_X1 U16834 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n15581) );
  OAI211_X1 U16835 ( .C1(n15575), .C2(n15574), .A(n15661), .B(n15573), .ZN(
        n15580) );
  OAI211_X1 U16836 ( .C1(n15578), .C2(n15577), .A(n15668), .B(n15576), .ZN(
        n15579) );
  NAND4_X1 U16837 ( .A1(n15582), .A2(n15581), .A3(n15580), .A4(n15579), .ZN(
        P2_U3217) );
  AOI22_X1 U16838 ( .A1(n15678), .A2(n15583), .B1(n15684), .B2(
        P2_ADDR_REG_6__SCAN_IN), .ZN(n15593) );
  OAI211_X1 U16839 ( .C1(n15586), .C2(n15585), .A(n15661), .B(n15584), .ZN(
        n15591) );
  OAI211_X1 U16840 ( .C1(n15589), .C2(n15588), .A(n15587), .B(n15668), .ZN(
        n15590) );
  NAND4_X1 U16841 ( .A1(n15593), .A2(n15592), .A3(n15591), .A4(n15590), .ZN(
        P2_U3220) );
  AOI22_X1 U16842 ( .A1(n15678), .A2(n15594), .B1(n15684), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n15605) );
  NAND2_X1 U16843 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n15604) );
  AOI211_X1 U16844 ( .C1(n15597), .C2(n15596), .A(n15681), .B(n15595), .ZN(
        n15598) );
  INV_X1 U16845 ( .A(n15598), .ZN(n15603) );
  OAI211_X1 U16846 ( .C1(n15601), .C2(n15600), .A(n15599), .B(n15661), .ZN(
        n15602) );
  NAND4_X1 U16847 ( .A1(n15605), .A2(n15604), .A3(n15603), .A4(n15602), .ZN(
        P2_U3222) );
  AND2_X1 U16848 ( .A1(n15607), .A2(n15606), .ZN(n15608) );
  NOR2_X1 U16849 ( .A1(n15609), .A2(n15608), .ZN(n15620) );
  NOR2_X1 U16850 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15610), .ZN(n15613) );
  NOR2_X1 U16851 ( .A1(n15626), .A2(n15611), .ZN(n15612) );
  AOI211_X1 U16852 ( .C1(n15684), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n15613), 
        .B(n15612), .ZN(n15619) );
  AOI211_X1 U16853 ( .C1(n15616), .C2(n15615), .A(n15681), .B(n15614), .ZN(
        n15617) );
  INV_X1 U16854 ( .A(n15617), .ZN(n15618) );
  OAI211_X1 U16855 ( .C1(n15620), .C2(n15686), .A(n15619), .B(n15618), .ZN(
        P2_U3225) );
  AOI21_X1 U16856 ( .B1(n15623), .B2(n15622), .A(n15621), .ZN(n15634) );
  NOR2_X1 U16857 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15624), .ZN(n15628) );
  NOR2_X1 U16858 ( .A1(n15626), .A2(n15625), .ZN(n15627) );
  AOI211_X1 U16859 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n15684), .A(n15628), 
        .B(n15627), .ZN(n15633) );
  OAI211_X1 U16860 ( .C1(n15631), .C2(n15630), .A(n15629), .B(n15668), .ZN(
        n15632) );
  OAI211_X1 U16861 ( .C1(n15634), .C2(n15686), .A(n15633), .B(n15632), .ZN(
        P2_U3228) );
  AOI22_X1 U16862 ( .A1(n15684), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15643) );
  OAI211_X1 U16863 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15636), .A(n15661), 
        .B(n15635), .ZN(n15642) );
  NAND2_X1 U16864 ( .A1(n15678), .A2(n15637), .ZN(n15641) );
  OAI211_X1 U16865 ( .C1(n15639), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15668), 
        .B(n15638), .ZN(n15640) );
  NAND4_X1 U16866 ( .A1(n15643), .A2(n15642), .A3(n15641), .A4(n15640), .ZN(
        P2_U3229) );
  OAI21_X1 U16867 ( .B1(n15645), .B2(n15644), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15646) );
  OAI21_X1 U16868 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15646), .ZN(n15656) );
  OAI211_X1 U16869 ( .C1(n15649), .C2(n15648), .A(n15661), .B(n15647), .ZN(
        n15655) );
  NAND2_X1 U16870 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n15684), .ZN(n15654) );
  OAI211_X1 U16871 ( .C1(n15652), .C2(n15651), .A(n15650), .B(n15668), .ZN(
        n15653) );
  NAND4_X1 U16872 ( .A1(n15656), .A2(n15655), .A3(n15654), .A4(n15653), .ZN(
        P2_U3230) );
  AOI22_X1 U16873 ( .A1(n15684), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n15672) );
  MUX2_X1 U16874 ( .A(n15659), .B(P2_REG2_REG_17__SCAN_IN), .S(n15658), .Z(
        n15663) );
  NAND2_X1 U16875 ( .A1(n15662), .A2(n15663), .ZN(n15660) );
  OAI211_X1 U16876 ( .C1(n15663), .C2(n15662), .A(n15661), .B(n15660), .ZN(
        n15671) );
  NAND2_X1 U16877 ( .A1(n15678), .A2(n15664), .ZN(n15670) );
  XOR2_X1 U16878 ( .A(n15666), .B(n15665), .Z(n15667) );
  NAND2_X1 U16879 ( .A1(n15668), .A2(n15667), .ZN(n15669) );
  NAND4_X1 U16880 ( .A1(n15672), .A2(n15671), .A3(n15670), .A4(n15669), .ZN(
        P2_U3231) );
  AOI21_X1 U16881 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n15674), .A(n15673), 
        .ZN(n15687) );
  XNOR2_X1 U16882 ( .A(n15676), .B(n15675), .ZN(n15682) );
  NAND2_X1 U16883 ( .A1(n15678), .A2(n15677), .ZN(n15680) );
  OAI211_X1 U16884 ( .C1(n15682), .C2(n15681), .A(n15680), .B(n15679), .ZN(
        n15683) );
  AOI21_X1 U16885 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15684), .A(n15683), 
        .ZN(n15685) );
  OAI21_X1 U16886 ( .B1(n15687), .B2(n15686), .A(n15685), .ZN(P2_U3232) );
  INV_X1 U16887 ( .A(n15688), .ZN(n15690) );
  NAND2_X1 U16888 ( .A1(n15689), .A2(n11039), .ZN(n15692) );
  NAND2_X1 U16889 ( .A1(n15690), .A2(n15692), .ZN(n15693) );
  MUX2_X1 U16890 ( .A(n15693), .B(n15692), .S(n15691), .Z(n15695) );
  NAND2_X1 U16891 ( .A1(n15695), .A2(n15694), .ZN(n15698) );
  AOI22_X1 U16892 ( .A1(n15696), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15697) );
  OAI21_X1 U16893 ( .B1(n15699), .B2(n15698), .A(n15697), .ZN(P1_U3243) );
  INV_X1 U16894 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15855) );
  OAI21_X1 U16895 ( .B1(n15701), .B2(n16538), .A(n15700), .ZN(n15709) );
  AOI21_X1 U16896 ( .B1(n15703), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15702), 
        .ZN(n15707) );
  OAI22_X1 U16897 ( .A1(n15707), .A2(n16567), .B1(n15705), .B2(n15704), .ZN(
        n15708) );
  AOI21_X1 U16898 ( .B1(n15709), .B2(n15720), .A(n15708), .ZN(n15711) );
  OAI211_X1 U16899 ( .C1(n15855), .C2(n15728), .A(n15711), .B(n15710), .ZN(
        P1_U3258) );
  INV_X1 U16900 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15729) );
  OAI21_X1 U16901 ( .B1(n15714), .B2(n15713), .A(n15712), .ZN(n15725) );
  MUX2_X1 U16902 ( .A(n11606), .B(P1_REG1_REG_12__SCAN_IN), .S(n15723), .Z(
        n15715) );
  NAND3_X1 U16903 ( .A1(n15717), .A2(n15716), .A3(n15715), .ZN(n15718) );
  NAND2_X1 U16904 ( .A1(n15719), .A2(n15718), .ZN(n15721) );
  AOI222_X1 U16905 ( .A1(n15725), .A2(n7362), .B1(n15723), .B2(n15722), .C1(
        n15721), .C2(n15720), .ZN(n15727) );
  OAI211_X1 U16906 ( .C1(n15729), .C2(n15728), .A(n15727), .B(n15726), .ZN(
        P1_U3255) );
  AOI21_X1 U16907 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15730), .A(n15735), .ZN(
        n15732) );
  INV_X1 U16908 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15731) );
  NOR2_X1 U16909 ( .A1(n15732), .A2(n15731), .ZN(n15896) );
  AOI21_X1 U16910 ( .B1(n15732), .B2(n15731), .A(n15896), .ZN(SUB_1596_U53) );
  XNOR2_X1 U16911 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15741), .ZN(n15743) );
  NAND2_X1 U16912 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15736), .ZN(n15738) );
  NAND2_X1 U16913 ( .A1(n15897), .A2(n15896), .ZN(n15737) );
  NAND2_X1 U16914 ( .A1(n15738), .A2(n15737), .ZN(n15744) );
  NOR2_X1 U16915 ( .A1(n15744), .A2(n15743), .ZN(n15745) );
  AOI21_X1 U16916 ( .B1(n15743), .B2(n15744), .A(n15745), .ZN(n15739) );
  INV_X1 U16917 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15747) );
  XNOR2_X1 U16918 ( .A(n15739), .B(n15747), .ZN(SUB_1596_U61) );
  NAND2_X1 U16919 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n15740), .ZN(n15742) );
  XNOR2_X1 U16920 ( .A(n15749), .B(n15750), .ZN(n15752) );
  NAND2_X1 U16921 ( .A1(n15744), .A2(n15743), .ZN(n15746) );
  AOI21_X1 U16922 ( .B1(n15747), .B2(n15746), .A(n15745), .ZN(n15753) );
  XNOR2_X1 U16923 ( .A(n15753), .B(n15752), .ZN(n15754) );
  XNOR2_X1 U16924 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15754), .ZN(SUB_1596_U60)
         );
  NAND2_X1 U16925 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15748), .ZN(n15751) );
  NOR2_X1 U16926 ( .A1(n15753), .A2(n15752), .ZN(n15756) );
  NOR2_X1 U16927 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15754), .ZN(n15755) );
  NOR2_X1 U16928 ( .A1(n15756), .A2(n15755), .ZN(n15764) );
  XOR2_X1 U16929 ( .A(n15765), .B(n15764), .Z(SUB_1596_U59) );
  NAND2_X1 U16930 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n15757), .ZN(n15761) );
  NAND2_X1 U16931 ( .A1(n15759), .A2(n15758), .ZN(n15760) );
  NAND2_X1 U16932 ( .A1(n15761), .A2(n15760), .ZN(n15773) );
  XOR2_X1 U16933 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), .Z(
        n15762) );
  XOR2_X1 U16934 ( .A(n15773), .B(n15762), .Z(n15768) );
  NAND2_X1 U16935 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15763), .ZN(n15766) );
  XOR2_X1 U16936 ( .A(n15769), .B(P2_ADDR_REG_5__SCAN_IN), .Z(SUB_1596_U58) );
  NAND2_X1 U16937 ( .A1(n15768), .A2(n15767), .ZN(n15771) );
  NAND2_X1 U16938 ( .A1(n15769), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n15770) );
  XNOR2_X1 U16939 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n15776) );
  INV_X1 U16940 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15775) );
  NOR2_X1 U16941 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15772), .ZN(n15774) );
  XOR2_X1 U16942 ( .A(n15776), .B(n15777), .Z(n15893) );
  XNOR2_X1 U16943 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15779), .ZN(n15780) );
  XNOR2_X1 U16944 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n15780), .ZN(n15784) );
  XNOR2_X1 U16945 ( .A(n15785), .B(n15784), .ZN(SUB_1596_U56) );
  NAND2_X1 U16946 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15779), .ZN(n15782) );
  XOR2_X1 U16947 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n15794) );
  XOR2_X1 U16948 ( .A(n15793), .B(n15794), .Z(n15789) );
  NOR2_X1 U16949 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n15783), .ZN(n15787) );
  NOR2_X1 U16950 ( .A1(n15785), .A2(n15784), .ZN(n15786) );
  NOR2_X1 U16951 ( .A1(n15789), .A2(n15788), .ZN(n15792) );
  NOR2_X1 U16952 ( .A1(n15792), .A2(n15791), .ZN(n15790) );
  XOR2_X1 U16953 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n15790), .Z(SUB_1596_U55) );
  XNOR2_X1 U16954 ( .A(n15806), .B(P1_ADDR_REG_9__SCAN_IN), .ZN(n15803) );
  XOR2_X1 U16955 ( .A(n15804), .B(n15803), .Z(n15798) );
  NAND2_X1 U16956 ( .A1(n15799), .A2(n15798), .ZN(n15800) );
  OAI21_X1 U16957 ( .B1(n15799), .B2(n15798), .A(n15800), .ZN(n15797) );
  XNOR2_X1 U16958 ( .A(n15797), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  NOR2_X1 U16959 ( .A1(n15799), .A2(n15798), .ZN(n15802) );
  INV_X1 U16960 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15801) );
  XNOR2_X1 U16961 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n15811) );
  XNOR2_X1 U16962 ( .A(n15812), .B(n15811), .ZN(n15808) );
  XOR2_X1 U16963 ( .A(n15809), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  NAND2_X1 U16964 ( .A1(n15808), .A2(n15807), .ZN(n15810) );
  XNOR2_X1 U16965 ( .A(n15822), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n15820) );
  INV_X1 U16966 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15814) );
  NAND2_X1 U16967 ( .A1(n15812), .A2(n15811), .ZN(n15813) );
  XOR2_X1 U16968 ( .A(n15820), .B(n15819), .Z(n15817) );
  NAND2_X1 U16969 ( .A1(n15817), .A2(n15816), .ZN(n15818) );
  OAI21_X1 U16970 ( .B1(n15816), .B2(n15817), .A(n15818), .ZN(n15815) );
  XNOR2_X1 U16971 ( .A(n15815), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  XNOR2_X1 U16972 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n15826) );
  XNOR2_X1 U16973 ( .A(n15827), .B(n15826), .ZN(n15823) );
  XNOR2_X1 U16974 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n15825), .ZN(SUB_1596_U68)
         );
  XNOR2_X1 U16975 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n15830) );
  INV_X1 U16976 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15829) );
  NAND2_X1 U16977 ( .A1(n15827), .A2(n15826), .ZN(n15828) );
  XNOR2_X1 U16978 ( .A(n15830), .B(n15838), .ZN(n15833) );
  NOR2_X1 U16979 ( .A1(n15833), .A2(n15832), .ZN(n15834) );
  AOI21_X1 U16980 ( .B1(n15832), .B2(n15833), .A(n15834), .ZN(n15831) );
  XNOR2_X1 U16981 ( .A(n15831), .B(n11933), .ZN(SUB_1596_U67) );
  NAND2_X1 U16982 ( .A1(n15833), .A2(n15832), .ZN(n15835) );
  INV_X1 U16983 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15839) );
  NAND2_X1 U16984 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15836), .ZN(n15837) );
  XOR2_X1 U16985 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n15845) );
  XNOR2_X1 U16986 ( .A(n15846), .B(n15845), .ZN(n15841) );
  AOI21_X1 U16987 ( .B1(n15842), .B2(n15841), .A(n15843), .ZN(n15840) );
  INV_X1 U16988 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15844) );
  XNOR2_X1 U16989 ( .A(n15840), .B(n15844), .ZN(SUB_1596_U66) );
  INV_X1 U16990 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15848) );
  NOR2_X1 U16991 ( .A1(n15846), .A2(n15845), .ZN(n15847) );
  AOI21_X1 U16992 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15848), .A(n15847), 
        .ZN(n15857) );
  XOR2_X1 U16993 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .Z(n15849) );
  XNOR2_X1 U16994 ( .A(n15857), .B(n15849), .ZN(n15852) );
  AOI21_X1 U16995 ( .B1(n15851), .B2(n15852), .A(n7394), .ZN(n15850) );
  INV_X1 U16996 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15854) );
  XNOR2_X1 U16997 ( .A(n15850), .B(n15854), .ZN(SUB_1596_U65) );
  NAND2_X1 U16998 ( .A1(n15852), .A2(n15851), .ZN(n15853) );
  INV_X1 U16999 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15858) );
  NOR2_X1 U17000 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15855), .ZN(n15856) );
  OAI22_X1 U17001 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15858), .B1(n15857), 
        .B2(n15856), .ZN(n15861) );
  INV_X1 U17002 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15860) );
  XNOR2_X1 U17003 ( .A(n15861), .B(n15860), .ZN(n15862) );
  XOR2_X1 U17004 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15862), .Z(n15865) );
  NAND2_X1 U17005 ( .A1(n15866), .A2(n15865), .ZN(n15867) );
  OAI21_X1 U17006 ( .B1(n15866), .B2(n15865), .A(n15867), .ZN(n15859) );
  XNOR2_X1 U17007 ( .A(n15859), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U17008 ( .A1(n15861), .A2(n15860), .ZN(n15864) );
  NOR2_X1 U17009 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15862), .ZN(n15863) );
  XOR2_X1 U17010 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n15870), .Z(n15871) );
  XNOR2_X1 U17011 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15871), .ZN(n15874) );
  XOR2_X1 U17012 ( .A(n15874), .B(P2_ADDR_REG_17__SCAN_IN), .Z(n15876) );
  NOR2_X1 U17013 ( .A1(n15866), .A2(n15865), .ZN(n15869) );
  INV_X1 U17014 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15868) );
  XOR2_X1 U17015 ( .A(n15875), .B(n15876), .Z(SUB_1596_U63) );
  NOR2_X1 U17016 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15870), .ZN(n15873) );
  AND2_X1 U17017 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15871), .ZN(n15872) );
  NOR2_X1 U17018 ( .A1(n15873), .A2(n15872), .ZN(n15884) );
  XOR2_X1 U17019 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n15883) );
  XNOR2_X1 U17020 ( .A(n15884), .B(n15883), .ZN(n15879) );
  NAND2_X1 U17021 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n15874), .ZN(n15877) );
  XOR2_X1 U17022 ( .A(n15878), .B(P2_ADDR_REG_18__SCAN_IN), .Z(SUB_1596_U62)
         );
  NAND2_X1 U17023 ( .A1(n15878), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15882) );
  NAND2_X1 U17024 ( .A1(n15880), .A2(n15879), .ZN(n15881) );
  NAND2_X1 U17025 ( .A1(n15882), .A2(n15881), .ZN(n15891) );
  NOR2_X1 U17026 ( .A1(n15884), .A2(n15883), .ZN(n15885) );
  AOI21_X1 U17027 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n12968), .A(n15885), 
        .ZN(n15889) );
  XNOR2_X1 U17028 ( .A(n15886), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n15887) );
  XNOR2_X1 U17029 ( .A(n15887), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15888) );
  XNOR2_X1 U17030 ( .A(n15889), .B(n15888), .ZN(n15890) );
  XNOR2_X1 U17031 ( .A(n15891), .B(n15890), .ZN(SUB_1596_U4) );
  OAI21_X1 U17032 ( .B1(n15894), .B2(n15893), .A(n15892), .ZN(n15895) );
  XNOR2_X1 U17033 ( .A(n15895), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(SUB_1596_U57)
         );
  XOR2_X1 U17034 ( .A(n15897), .B(n15896), .Z(SUB_1596_U5) );
  NAND3_X1 U17035 ( .A1(n16082), .A2(n15969), .A3(n16069), .ZN(n15901) );
  OAI21_X1 U17036 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n15899), .A(n15898), .ZN(
        n15900) );
  NAND2_X1 U17037 ( .A1(n15901), .A2(n15900), .ZN(n15903) );
  AOI22_X1 U17038 ( .A1(n16043), .A2(P3_IR_REG_0__SCAN_IN), .B1(n16073), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n15902) );
  OAI211_X1 U17039 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n15904), .A(n15903), .B(
        n15902), .ZN(P3_U3182) );
  NOR2_X1 U17040 ( .A1(n15905), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n15907) );
  NOR2_X1 U17041 ( .A1(n15907), .A2(n15906), .ZN(n15922) );
  INV_X1 U17042 ( .A(n15908), .ZN(n15909) );
  OAI21_X1 U17043 ( .B1(n15981), .B2(n8038), .A(n15909), .ZN(n15916) );
  INV_X1 U17044 ( .A(n15910), .ZN(n15911) );
  NAND3_X1 U17045 ( .A1(n15913), .A2(n15912), .A3(n15911), .ZN(n15914) );
  AOI21_X1 U17046 ( .B1(n15930), .B2(n15914), .A(n16069), .ZN(n15915) );
  AOI211_X1 U17047 ( .C1(n16043), .C2(n15917), .A(n15916), .B(n15915), .ZN(
        n15921) );
  XNOR2_X1 U17048 ( .A(n15918), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15919) );
  NAND2_X1 U17049 ( .A1(n16079), .A2(n15919), .ZN(n15920) );
  OAI211_X1 U17050 ( .C1(n15922), .C2(n16082), .A(n15921), .B(n15920), .ZN(
        P3_U3185) );
  AOI21_X1 U17051 ( .B1(n15925), .B2(n15924), .A(n15923), .ZN(n15942) );
  INV_X1 U17052 ( .A(n15926), .ZN(n15927) );
  NOR2_X1 U17053 ( .A1(n15928), .A2(n15927), .ZN(n15931) );
  INV_X1 U17054 ( .A(n15950), .ZN(n15929) );
  AOI21_X1 U17055 ( .B1(n15931), .B2(n15930), .A(n15929), .ZN(n15933) );
  OAI22_X1 U17056 ( .A1(n15933), .A2(n16069), .B1(n15932), .B2(n16076), .ZN(
        n15934) );
  AOI211_X1 U17057 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n16073), .A(n15935), .B(
        n15934), .ZN(n15941) );
  AOI21_X1 U17058 ( .B1(n15938), .B2(n15937), .A(n15936), .ZN(n15939) );
  OR2_X1 U17059 ( .A1(n15969), .A2(n15939), .ZN(n15940) );
  OAI211_X1 U17060 ( .C1(n15942), .C2(n16082), .A(n15941), .B(n15940), .ZN(
        P3_U3186) );
  AOI21_X1 U17061 ( .B1(n15945), .B2(n15944), .A(n15943), .ZN(n15961) );
  INV_X1 U17062 ( .A(n15946), .ZN(n15947) );
  NOR2_X1 U17063 ( .A1(n15948), .A2(n15947), .ZN(n15951) );
  INV_X1 U17064 ( .A(n15974), .ZN(n15949) );
  AOI21_X1 U17065 ( .B1(n15951), .B2(n15950), .A(n15949), .ZN(n15953) );
  OAI22_X1 U17066 ( .A1(n15953), .A2(n16069), .B1(n15952), .B2(n16076), .ZN(
        n15954) );
  AOI211_X1 U17067 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n16073), .A(n15955), .B(
        n15954), .ZN(n15960) );
  OAI21_X1 U17068 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15957), .A(n15956), .ZN(
        n15958) );
  NAND2_X1 U17069 ( .A1(n16079), .A2(n15958), .ZN(n15959) );
  OAI211_X1 U17070 ( .C1(n15961), .C2(n16082), .A(n15960), .B(n15959), .ZN(
        P3_U3187) );
  AOI21_X1 U17071 ( .B1(n15964), .B2(n15963), .A(n15962), .ZN(n15970) );
  AOI21_X1 U17072 ( .B1(n15967), .B2(n15966), .A(n15965), .ZN(n15968) );
  OAI22_X1 U17073 ( .A1(n15970), .A2(n15969), .B1(n16082), .B2(n15968), .ZN(
        n15977) );
  INV_X1 U17074 ( .A(n15971), .ZN(n15972) );
  NAND3_X1 U17075 ( .A1(n15974), .A2(n15973), .A3(n15972), .ZN(n15975) );
  AOI21_X1 U17076 ( .B1(n15990), .B2(n15975), .A(n16069), .ZN(n15976) );
  AOI211_X1 U17077 ( .C1(n16043), .C2(n15978), .A(n15977), .B(n15976), .ZN(
        n15980) );
  OAI211_X1 U17078 ( .C1(n15982), .C2(n15981), .A(n15980), .B(n15979), .ZN(
        P3_U3188) );
  AOI21_X1 U17079 ( .B1(n15985), .B2(n15984), .A(n15983), .ZN(n16001) );
  INV_X1 U17080 ( .A(n15986), .ZN(n15987) );
  NOR2_X1 U17081 ( .A1(n15988), .A2(n15987), .ZN(n15991) );
  INV_X1 U17082 ( .A(n16009), .ZN(n15989) );
  AOI21_X1 U17083 ( .B1(n15991), .B2(n15990), .A(n15989), .ZN(n15993) );
  OAI22_X1 U17084 ( .A1(n15993), .A2(n16069), .B1(n15992), .B2(n16076), .ZN(
        n15994) );
  AOI211_X1 U17085 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n16073), .A(n15995), .B(
        n15994), .ZN(n16000) );
  OAI21_X1 U17086 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n15997), .A(n15996), .ZN(
        n15998) );
  NAND2_X1 U17087 ( .A1(n15998), .A2(n16079), .ZN(n15999) );
  OAI211_X1 U17088 ( .C1(n16001), .C2(n16082), .A(n16000), .B(n15999), .ZN(
        P3_U3189) );
  AOI21_X1 U17089 ( .B1(n16004), .B2(n16003), .A(n16002), .ZN(n16021) );
  INV_X1 U17090 ( .A(n16005), .ZN(n16006) );
  NOR2_X1 U17091 ( .A1(n16007), .A2(n16006), .ZN(n16010) );
  INV_X1 U17092 ( .A(n16030), .ZN(n16008) );
  AOI21_X1 U17093 ( .B1(n16010), .B2(n16009), .A(n16008), .ZN(n16012) );
  OAI22_X1 U17094 ( .A1(n16012), .A2(n16069), .B1(n16011), .B2(n16076), .ZN(
        n16013) );
  AOI211_X1 U17095 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n16073), .A(n16014), .B(
        n16013), .ZN(n16020) );
  OAI21_X1 U17096 ( .B1(n16017), .B2(n16016), .A(n16015), .ZN(n16018) );
  NAND2_X1 U17097 ( .A1(n16018), .A2(n16079), .ZN(n16019) );
  OAI211_X1 U17098 ( .C1(n16021), .C2(n16082), .A(n16020), .B(n16019), .ZN(
        P3_U3190) );
  AOI21_X1 U17099 ( .B1(n16024), .B2(n16023), .A(n16022), .ZN(n16041) );
  INV_X1 U17100 ( .A(n16025), .ZN(n16026) );
  NOR2_X1 U17101 ( .A1(n16027), .A2(n16026), .ZN(n16031) );
  INV_X1 U17102 ( .A(n16028), .ZN(n16029) );
  AOI21_X1 U17103 ( .B1(n16031), .B2(n16030), .A(n16029), .ZN(n16033) );
  OAI22_X1 U17104 ( .A1(n16033), .A2(n16069), .B1(n16032), .B2(n16076), .ZN(
        n16034) );
  AOI211_X1 U17105 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n16073), .A(n16035), .B(
        n16034), .ZN(n16040) );
  OAI21_X1 U17106 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n16037), .A(n16036), .ZN(
        n16038) );
  NAND2_X1 U17107 ( .A1(n16038), .A2(n16079), .ZN(n16039) );
  OAI211_X1 U17108 ( .C1(n16041), .C2(n16082), .A(n16040), .B(n16039), .ZN(
        P3_U3191) );
  AOI22_X1 U17109 ( .A1(n16043), .A2(n16042), .B1(n16073), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n16060) );
  OAI21_X1 U17110 ( .B1(n16046), .B2(n16045), .A(n16044), .ZN(n16053) );
  NAND2_X1 U17111 ( .A1(n16048), .A2(n16047), .ZN(n16050) );
  XOR2_X1 U17112 ( .A(n16050), .B(n16049), .Z(n16051) );
  AOI22_X1 U17113 ( .A1(n16053), .A2(n16079), .B1(n16052), .B2(n16051), .ZN(
        n16059) );
  OAI221_X1 U17114 ( .B1(n16056), .B2(n7435), .C1(n16056), .C2(n16055), .A(
        n16054), .ZN(n16057) );
  NAND4_X1 U17115 ( .A1(n16060), .A2(n16059), .A3(n16058), .A4(n16057), .ZN(
        P3_U3198) );
  INV_X1 U17116 ( .A(n16061), .ZN(n16062) );
  AOI21_X1 U17117 ( .B1(n16064), .B2(n16063), .A(n16062), .ZN(n16083) );
  OAI21_X1 U17118 ( .B1(n16066), .B2(P3_REG1_REG_17__SCAN_IN), .A(n16065), 
        .ZN(n16080) );
  INV_X1 U17119 ( .A(n16067), .ZN(n16068) );
  AOI211_X1 U17120 ( .C1(n16071), .C2(n16070), .A(n16069), .B(n16068), .ZN(
        n16078) );
  AOI21_X1 U17121 ( .B1(n16073), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n16072), 
        .ZN(n16074) );
  OAI21_X1 U17122 ( .B1(n16076), .B2(n16075), .A(n16074), .ZN(n16077) );
  AOI211_X1 U17123 ( .C1(n16080), .C2(n16079), .A(n16078), .B(n16077), .ZN(
        n16081) );
  OAI21_X1 U17124 ( .B1(n16083), .B2(n16082), .A(n16081), .ZN(P3_U3199) );
  AOI21_X1 U17125 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n16084) );
  OAI21_X1 U17126 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n16084), 
        .ZN(U29) );
  NAND2_X1 U17127 ( .A1(n16085), .A2(n16532), .ZN(n16095) );
  AOI21_X1 U17128 ( .B1(n16086), .B2(n9047), .A(n16092), .ZN(n16087) );
  OAI21_X1 U17129 ( .B1(n16088), .B2(n16485), .A(n16087), .ZN(n16089) );
  AOI21_X1 U17130 ( .B1(n16094), .B2(n16095), .A(n16089), .ZN(n16091) );
  AOI22_X1 U17131 ( .A1(n16539), .A2(n16091), .B1(n11039), .B2(n16537), .ZN(
        P1_U3528) );
  INV_X1 U17132 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n16090) );
  AOI22_X1 U17133 ( .A1(n16543), .A2(n16091), .B1(n16090), .B2(n16540), .ZN(
        P1_U3459) );
  INV_X1 U17134 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n16103) );
  INV_X1 U17135 ( .A(n16092), .ZN(n16098) );
  INV_X1 U17136 ( .A(n16093), .ZN(n16096) );
  OAI21_X1 U17137 ( .B1(n16096), .B2(n16095), .A(n16094), .ZN(n16097) );
  AOI21_X1 U17138 ( .B1(n16098), .B2(n16097), .A(n16153), .ZN(n16101) );
  AOI21_X1 U17139 ( .B1(n16156), .B2(n16099), .A(n16142), .ZN(n16100) );
  AOI211_X1 U17140 ( .C1(n16153), .C2(P1_REG2_REG_0__SCAN_IN), .A(n16101), .B(
        n16100), .ZN(n16102) );
  OAI21_X1 U17141 ( .B1(n16104), .B2(n16103), .A(n16102), .ZN(P1_U3293) );
  INV_X1 U17142 ( .A(n16111), .ZN(n16121) );
  NAND2_X1 U17143 ( .A1(n16106), .A2(n16105), .ZN(n16116) );
  INV_X1 U17144 ( .A(n16116), .ZN(n16112) );
  NOR2_X1 U17145 ( .A1(n16259), .A2(n16107), .ZN(n16110) );
  OAI22_X1 U17146 ( .A1(n16111), .A2(n16110), .B1(n16109), .B2(n16108), .ZN(
        n16119) );
  AOI211_X1 U17147 ( .C1(n16509), .C2(n16121), .A(n16112), .B(n16119), .ZN(
        n16115) );
  AOI22_X1 U17148 ( .A1(n16512), .A2(n16115), .B1(n16113), .B2(n16510), .ZN(
        P2_U3499) );
  INV_X1 U17149 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n16114) );
  AOI22_X1 U17150 ( .A1(n16516), .A2(n16115), .B1(n16114), .B2(n16513), .ZN(
        P2_U3430) );
  INV_X1 U17151 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n16118) );
  OAI22_X1 U17152 ( .A1(n16118), .A2(n16117), .B1(n16116), .B2(n8334), .ZN(
        n16120) );
  AOI211_X1 U17153 ( .C1(n16122), .C2(n16121), .A(n16120), .B(n16119), .ZN(
        n16123) );
  AOI22_X1 U17154 ( .A1(n16408), .A2(n16124), .B1(n16123), .B2(n14675), .ZN(
        P2_U3265) );
  INV_X1 U17155 ( .A(n16135), .ZN(n16125) );
  NOR2_X1 U17156 ( .A1(n16125), .A2(n16413), .ZN(n16126) );
  OAI21_X1 U17157 ( .B1(n16127), .B2(n16126), .A(n16473), .ZN(n16128) );
  OAI21_X1 U17158 ( .B1(n16473), .B2(n8495), .A(n16128), .ZN(P3_U3460) );
  INV_X1 U17159 ( .A(n16129), .ZN(n16195) );
  OAI22_X1 U17160 ( .A1(n16194), .A2(n16131), .B1(n16130), .B2(n16195), .ZN(
        n16134) );
  INV_X1 U17161 ( .A(n16132), .ZN(n16133) );
  AOI211_X1 U17162 ( .C1(n16200), .C2(n16135), .A(n16134), .B(n16133), .ZN(
        n16136) );
  AOI22_X1 U17163 ( .A1(n14164), .A2(n16137), .B1(n16136), .B2(n14169), .ZN(
        P3_U3232) );
  INV_X1 U17164 ( .A(n16485), .ZN(n16391) );
  XNOR2_X1 U17165 ( .A(n16139), .B(n16138), .ZN(n16160) );
  INV_X1 U17166 ( .A(n16140), .ZN(n16141) );
  OAI211_X1 U17167 ( .C1(n16155), .C2(n16142), .A(n16141), .B(n15501), .ZN(
        n16158) );
  OAI21_X1 U17168 ( .B1(n16155), .B2(n16448), .A(n16158), .ZN(n16149) );
  XNOR2_X1 U17169 ( .A(n16144), .B(n16143), .ZN(n16145) );
  NOR2_X1 U17170 ( .A1(n16145), .A2(n16532), .ZN(n16146) );
  AOI211_X1 U17171 ( .C1(n16488), .C2(n16160), .A(n16147), .B(n16146), .ZN(
        n16163) );
  INV_X1 U17172 ( .A(n16163), .ZN(n16148) );
  AOI211_X1 U17173 ( .C1(n16391), .C2(n16160), .A(n16149), .B(n16148), .ZN(
        n16152) );
  AOI22_X1 U17174 ( .A1(n16539), .A2(n16152), .B1(n16150), .B2(n16537), .ZN(
        P1_U3529) );
  INV_X1 U17175 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n16151) );
  AOI22_X1 U17176 ( .A1(n16543), .A2(n16152), .B1(n16151), .B2(n16540), .ZN(
        P1_U3462) );
  AOI22_X1 U17177 ( .A1(n16153), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n16312), .ZN(n16154) );
  OAI21_X1 U17178 ( .B1(n16156), .B2(n16155), .A(n16154), .ZN(n16157) );
  INV_X1 U17179 ( .A(n16157), .ZN(n16162) );
  INV_X1 U17180 ( .A(n16158), .ZN(n16159) );
  AOI22_X1 U17181 ( .A1(n16315), .A2(n16160), .B1(n16317), .B2(n16159), .ZN(
        n16161) );
  OAI211_X1 U17182 ( .C1(n16153), .C2(n16163), .A(n16162), .B(n16161), .ZN(
        P1_U3292) );
  INV_X1 U17183 ( .A(n16164), .ZN(n16165) );
  AOI21_X1 U17184 ( .B1(n16431), .B2(n16430), .A(n16165), .ZN(n16170) );
  OAI211_X1 U17185 ( .C1(n16168), .C2(n16504), .A(n16167), .B(n16166), .ZN(
        n16169) );
  NOR2_X1 U17186 ( .A1(n16170), .A2(n16169), .ZN(n16173) );
  AOI22_X1 U17187 ( .A1(n16512), .A2(n16173), .B1(n16171), .B2(n16510), .ZN(
        P2_U3500) );
  INV_X1 U17188 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n16172) );
  AOI22_X1 U17189 ( .A1(n16516), .A2(n16173), .B1(n16172), .B2(n16513), .ZN(
        P2_U3433) );
  INV_X1 U17190 ( .A(n16174), .ZN(n16175) );
  AOI21_X1 U17191 ( .B1(n16177), .B2(n16176), .A(n16175), .ZN(n16192) );
  AOI22_X1 U17192 ( .A1(n16180), .A2(n11308), .B1(n16179), .B2(n16178), .ZN(
        n16187) );
  AND3_X1 U17193 ( .A1(n16182), .A2(n10066), .A3(n16181), .ZN(n16184) );
  OAI21_X1 U17194 ( .B1(n16185), .B2(n16184), .A(n16183), .ZN(n16186) );
  OAI211_X1 U17195 ( .C1(n16192), .C2(n16188), .A(n16187), .B(n16186), .ZN(
        n16197) );
  OAI22_X1 U17196 ( .A1(n16192), .A2(n16413), .B1(n16196), .B2(n16467), .ZN(
        n16189) );
  NOR2_X1 U17197 ( .A1(n16197), .A2(n16189), .ZN(n16191) );
  AOI22_X1 U17198 ( .A1(n16473), .A2(n16191), .B1(n8499), .B2(n16470), .ZN(
        P3_U3461) );
  INV_X1 U17199 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n16190) );
  AOI22_X1 U17200 ( .A1(n16447), .A2(n16191), .B1(n16190), .B2(n16562), .ZN(
        P3_U3396) );
  INV_X1 U17201 ( .A(n16192), .ZN(n16199) );
  OAI22_X1 U17202 ( .A1(n16196), .A2(n16195), .B1(n16194), .B2(n16193), .ZN(
        n16198) );
  AOI211_X1 U17203 ( .C1(n16200), .C2(n16199), .A(n16198), .B(n16197), .ZN(
        n16201) );
  AOI22_X1 U17204 ( .A1(n14164), .A2(n16202), .B1(n16201), .B2(n14169), .ZN(
        P3_U3231) );
  INV_X1 U17205 ( .A(n16203), .ZN(n16208) );
  OAI22_X1 U17206 ( .A1(n16205), .A2(n16495), .B1(n16204), .B2(n16448), .ZN(
        n16207) );
  AOI211_X1 U17207 ( .C1(n16391), .C2(n16208), .A(n16207), .B(n16206), .ZN(
        n16211) );
  AOI22_X1 U17208 ( .A1(n16539), .A2(n16211), .B1(n16209), .B2(n16537), .ZN(
        P1_U3530) );
  INV_X1 U17209 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n16210) );
  AOI22_X1 U17210 ( .A1(n16543), .A2(n16211), .B1(n16210), .B2(n16540), .ZN(
        P1_U3465) );
  XNOR2_X1 U17211 ( .A(n16212), .B(n16216), .ZN(n16224) );
  OAI211_X1 U17212 ( .C1(n16214), .C2(n16213), .A(n16261), .B(n16260), .ZN(
        n16229) );
  OAI21_X1 U17213 ( .B1(n16214), .B2(n16504), .A(n16229), .ZN(n16221) );
  XNOR2_X1 U17214 ( .A(n16216), .B(n16215), .ZN(n16218) );
  OAI21_X1 U17215 ( .B1(n16218), .B2(n16256), .A(n16217), .ZN(n16219) );
  AOI21_X1 U17216 ( .B1(n16259), .B2(n16224), .A(n16219), .ZN(n16233) );
  INV_X1 U17217 ( .A(n16233), .ZN(n16220) );
  AOI211_X1 U17218 ( .C1(n16509), .C2(n16224), .A(n16221), .B(n16220), .ZN(
        n16223) );
  AOI22_X1 U17219 ( .A1(n16512), .A2(n16223), .B1(n11094), .B2(n16510), .ZN(
        P2_U3501) );
  INV_X1 U17220 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n16222) );
  AOI22_X1 U17221 ( .A1(n16516), .A2(n16223), .B1(n16222), .B2(n16513), .ZN(
        P2_U3436) );
  AOI22_X1 U17222 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n16408), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n16397), .ZN(n16232) );
  NAND2_X1 U17223 ( .A1(n16401), .A2(n16224), .ZN(n16227) );
  NAND2_X1 U17224 ( .A1(n16399), .A2(n16225), .ZN(n16226) );
  OAI211_X1 U17225 ( .C1(n16229), .C2(n16228), .A(n16227), .B(n16226), .ZN(
        n16230) );
  INV_X1 U17226 ( .A(n16230), .ZN(n16231) );
  OAI211_X1 U17227 ( .C1(n16408), .C2(n16233), .A(n16232), .B(n16231), .ZN(
        P2_U3263) );
  NOR2_X1 U17228 ( .A1(n16234), .A2(n16467), .ZN(n16236) );
  AOI211_X1 U17229 ( .C1(n16382), .C2(n16237), .A(n16236), .B(n16235), .ZN(
        n16239) );
  AOI22_X1 U17230 ( .A1(n16473), .A2(n16239), .B1(n8505), .B2(n16470), .ZN(
        P3_U3462) );
  INV_X1 U17231 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n16238) );
  AOI22_X1 U17232 ( .A1(n16447), .A2(n16239), .B1(n16238), .B2(n16562), .ZN(
        P3_U3399) );
  OAI211_X1 U17233 ( .C1(n16242), .C2(n16448), .A(n16241), .B(n16240), .ZN(
        n16246) );
  NOR2_X1 U17234 ( .A1(n16244), .A2(n16243), .ZN(n16245) );
  AOI211_X1 U17235 ( .C1(n16248), .C2(n16247), .A(n16246), .B(n16245), .ZN(
        n16251) );
  AOI22_X1 U17236 ( .A1(n16539), .A2(n16251), .B1(n16249), .B2(n16537), .ZN(
        P1_U3531) );
  INV_X1 U17237 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n16250) );
  AOI22_X1 U17238 ( .A1(n16543), .A2(n16251), .B1(n16250), .B2(n16540), .ZN(
        P1_U3468) );
  XNOR2_X1 U17239 ( .A(n16252), .B(n16254), .ZN(n16274) );
  XOR2_X1 U17240 ( .A(n16254), .B(n16253), .Z(n16257) );
  OAI21_X1 U17241 ( .B1(n16257), .B2(n16256), .A(n16255), .ZN(n16258) );
  AOI21_X1 U17242 ( .B1(n16259), .B2(n16274), .A(n16258), .ZN(n16277) );
  NAND2_X1 U17243 ( .A1(n16270), .A2(n16260), .ZN(n16262) );
  NAND2_X1 U17244 ( .A1(n16262), .A2(n16261), .ZN(n16263) );
  OR2_X1 U17245 ( .A1(n16264), .A2(n16263), .ZN(n16272) );
  NAND2_X1 U17246 ( .A1(n16274), .A2(n16509), .ZN(n16267) );
  NAND2_X1 U17247 ( .A1(n16270), .A2(n16265), .ZN(n16266) );
  AOI22_X1 U17248 ( .A1(n16512), .A2(n16269), .B1(n11095), .B2(n16510), .ZN(
        P2_U3502) );
  INV_X1 U17249 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n16268) );
  AOI22_X1 U17250 ( .A1(n16516), .A2(n16269), .B1(n16268), .B2(n16513), .ZN(
        P2_U3439) );
  AOI222_X1 U17251 ( .A1(n16271), .A2(n16397), .B1(n16408), .B2(
        P2_REG2_REG_3__SCAN_IN), .C1(n16270), .C2(n16399), .ZN(n16276) );
  INV_X1 U17252 ( .A(n16272), .ZN(n16273) );
  AOI22_X1 U17253 ( .A1(n16274), .A2(n16401), .B1(n16403), .B2(n16273), .ZN(
        n16275) );
  OAI211_X1 U17254 ( .C1(n16408), .C2(n16277), .A(n16276), .B(n16275), .ZN(
        P2_U3262) );
  NOR2_X1 U17255 ( .A1(n16278), .A2(n16467), .ZN(n16280) );
  AOI211_X1 U17256 ( .C1(n16382), .C2(n16281), .A(n16280), .B(n16279), .ZN(
        n16284) );
  AOI22_X1 U17257 ( .A1(n16473), .A2(n16284), .B1(n16282), .B2(n16470), .ZN(
        P3_U3463) );
  INV_X1 U17258 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n16283) );
  AOI22_X1 U17259 ( .A1(n16447), .A2(n16284), .B1(n16283), .B2(n16562), .ZN(
        P3_U3402) );
  INV_X1 U17260 ( .A(n16285), .ZN(n16291) );
  OAI211_X1 U17261 ( .C1(n16288), .C2(n16448), .A(n16287), .B(n16286), .ZN(
        n16290) );
  AOI211_X1 U17262 ( .C1(n16291), .C2(n16536), .A(n16290), .B(n16289), .ZN(
        n16294) );
  AOI22_X1 U17263 ( .A1(n16539), .A2(n16294), .B1(n16292), .B2(n16537), .ZN(
        P1_U3532) );
  INV_X1 U17264 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16293) );
  AOI22_X1 U17265 ( .A1(n16543), .A2(n16294), .B1(n16293), .B2(n16540), .ZN(
        P1_U3471) );
  INV_X1 U17266 ( .A(n16295), .ZN(n16297) );
  OAI211_X1 U17267 ( .C1(n16298), .C2(n16504), .A(n16297), .B(n16296), .ZN(
        n16301) );
  AOI21_X1 U17268 ( .B1(n16431), .B2(n16430), .A(n16299), .ZN(n16300) );
  NOR2_X1 U17269 ( .A1(n16301), .A2(n16300), .ZN(n16304) );
  AOI22_X1 U17270 ( .A1(n16512), .A2(n16304), .B1(n16302), .B2(n16510), .ZN(
        P2_U3503) );
  INV_X1 U17271 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n16303) );
  AOI22_X1 U17272 ( .A1(n16516), .A2(n16304), .B1(n16303), .B2(n16513), .ZN(
        P2_U3442) );
  OAI22_X1 U17273 ( .A1(n16306), .A2(n16413), .B1(n16305), .B2(n16467), .ZN(
        n16308) );
  NOR2_X1 U17274 ( .A1(n16308), .A2(n16307), .ZN(n16310) );
  AOI22_X1 U17275 ( .A1(n16473), .A2(n16310), .B1(n8517), .B2(n16470), .ZN(
        P3_U3464) );
  INV_X1 U17276 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n16309) );
  AOI22_X1 U17277 ( .A1(n16447), .A2(n16310), .B1(n16309), .B2(n16562), .ZN(
        P3_U3405) );
  AOI222_X1 U17278 ( .A1(n16314), .A2(n16313), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n16153), .C1(n16312), .C2(n16311), .ZN(n16320) );
  AOI22_X1 U17279 ( .A1(n16318), .A2(n16317), .B1(n16316), .B2(n16315), .ZN(
        n16319) );
  OAI211_X1 U17280 ( .C1(n16153), .C2(n16321), .A(n16320), .B(n16319), .ZN(
        P1_U3288) );
  OAI21_X1 U17281 ( .B1(n16323), .B2(n16504), .A(n16322), .ZN(n16325) );
  AOI211_X1 U17282 ( .C1(n16509), .C2(n16326), .A(n16325), .B(n16324), .ZN(
        n16329) );
  AOI22_X1 U17283 ( .A1(n16512), .A2(n16329), .B1(n16327), .B2(n16510), .ZN(
        P2_U3504) );
  INV_X1 U17284 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n16328) );
  AOI22_X1 U17285 ( .A1(n16516), .A2(n16329), .B1(n16328), .B2(n16513), .ZN(
        P2_U3445) );
  NOR2_X1 U17286 ( .A1(n16330), .A2(n16413), .ZN(n16331) );
  AOI211_X1 U17287 ( .C1(n16410), .C2(n16333), .A(n16332), .B(n16331), .ZN(
        n16336) );
  AOI22_X1 U17288 ( .A1(n16473), .A2(n16336), .B1(n16334), .B2(n16470), .ZN(
        P3_U3465) );
  INV_X1 U17289 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n16335) );
  AOI22_X1 U17290 ( .A1(n16447), .A2(n16336), .B1(n16335), .B2(n16562), .ZN(
        P3_U3408) );
  OAI21_X1 U17291 ( .B1(n16338), .B2(n16448), .A(n16337), .ZN(n16340) );
  AOI211_X1 U17292 ( .C1(n16391), .C2(n16341), .A(n16340), .B(n16339), .ZN(
        n16344) );
  INV_X1 U17293 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n16342) );
  AOI22_X1 U17294 ( .A1(n16539), .A2(n16344), .B1(n16342), .B2(n16537), .ZN(
        P1_U3534) );
  INV_X1 U17295 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n16343) );
  AOI22_X1 U17296 ( .A1(n16543), .A2(n16344), .B1(n16343), .B2(n16540), .ZN(
        P1_U3477) );
  OAI22_X1 U17297 ( .A1(n16346), .A2(n16413), .B1(n16345), .B2(n16467), .ZN(
        n16348) );
  NOR2_X1 U17298 ( .A1(n16348), .A2(n16347), .ZN(n16350) );
  AOI22_X1 U17299 ( .A1(n16473), .A2(n16350), .B1(n8527), .B2(n16470), .ZN(
        P3_U3466) );
  INV_X1 U17300 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n16349) );
  AOI22_X1 U17301 ( .A1(n16447), .A2(n16350), .B1(n16349), .B2(n16562), .ZN(
        P3_U3411) );
  OAI22_X1 U17302 ( .A1(n16352), .A2(n16495), .B1(n16351), .B2(n16448), .ZN(
        n16354) );
  AOI211_X1 U17303 ( .C1(n16391), .C2(n16355), .A(n16354), .B(n16353), .ZN(
        n16358) );
  AOI22_X1 U17304 ( .A1(n16539), .A2(n16358), .B1(n16356), .B2(n16537), .ZN(
        P1_U3535) );
  INV_X1 U17305 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n16357) );
  AOI22_X1 U17306 ( .A1(n16543), .A2(n16358), .B1(n16357), .B2(n16540), .ZN(
        P1_U3480) );
  OAI21_X1 U17307 ( .B1(n16360), .B2(n16504), .A(n16359), .ZN(n16362) );
  AOI211_X1 U17308 ( .C1(n16509), .C2(n16363), .A(n16362), .B(n16361), .ZN(
        n16366) );
  AOI22_X1 U17309 ( .A1(n16512), .A2(n16366), .B1(n16364), .B2(n16510), .ZN(
        P2_U3506) );
  INV_X1 U17310 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n16365) );
  AOI22_X1 U17311 ( .A1(n16516), .A2(n16366), .B1(n16365), .B2(n16513), .ZN(
        P2_U3451) );
  OAI21_X1 U17312 ( .B1(n16368), .B2(n16467), .A(n16367), .ZN(n16369) );
  AOI21_X1 U17313 ( .B1(n16469), .B2(n16370), .A(n16369), .ZN(n16373) );
  AOI22_X1 U17314 ( .A1(n16473), .A2(n16373), .B1(n16371), .B2(n16470), .ZN(
        P3_U3467) );
  INV_X1 U17315 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n16372) );
  AOI22_X1 U17316 ( .A1(n16447), .A2(n16373), .B1(n16372), .B2(n16562), .ZN(
        P3_U3414) );
  OAI22_X1 U17317 ( .A1(n16375), .A2(n16495), .B1(n16374), .B2(n16448), .ZN(
        n16377) );
  AOI211_X1 U17318 ( .C1(n16391), .C2(n16378), .A(n16377), .B(n16376), .ZN(
        n16380) );
  AOI22_X1 U17319 ( .A1(n16539), .A2(n16380), .B1(n11325), .B2(n16537), .ZN(
        P1_U3536) );
  INV_X1 U17320 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n16379) );
  AOI22_X1 U17321 ( .A1(n16543), .A2(n16380), .B1(n16379), .B2(n16540), .ZN(
        P1_U3483) );
  AOI22_X1 U17322 ( .A1(n16383), .A2(n16382), .B1(n16381), .B2(n16410), .ZN(
        n16384) );
  AOI22_X1 U17323 ( .A1(n16473), .A2(n16387), .B1(n8536), .B2(n16470), .ZN(
        P3_U3468) );
  INV_X1 U17324 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16386) );
  AOI22_X1 U17325 ( .A1(n16447), .A2(n16387), .B1(n16386), .B2(n16562), .ZN(
        P3_U3417) );
  OAI22_X1 U17326 ( .A1(n16389), .A2(n16495), .B1(n7765), .B2(n16448), .ZN(
        n16390) );
  AOI21_X1 U17327 ( .B1(n16392), .B2(n16391), .A(n16390), .ZN(n16393) );
  AOI22_X1 U17328 ( .A1(n16539), .A2(n16396), .B1(n11321), .B2(n16537), .ZN(
        P1_U3537) );
  INV_X1 U17329 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16395) );
  AOI22_X1 U17330 ( .A1(n16543), .A2(n16396), .B1(n16395), .B2(n16540), .ZN(
        P1_U3486) );
  AOI222_X1 U17331 ( .A1(n16400), .A2(n16399), .B1(P2_REG2_REG_9__SCAN_IN), 
        .B2(n16408), .C1(n16398), .C2(n16397), .ZN(n16406) );
  AOI22_X1 U17332 ( .A1(n16404), .A2(n16403), .B1(n16402), .B2(n16401), .ZN(
        n16405) );
  OAI211_X1 U17333 ( .C1(n16408), .C2(n16407), .A(n16406), .B(n16405), .ZN(
        P2_U3256) );
  INV_X1 U17334 ( .A(n16414), .ZN(n16416) );
  AOI21_X1 U17335 ( .B1(n16411), .B2(n16410), .A(n16409), .ZN(n16412) );
  OAI21_X1 U17336 ( .B1(n16414), .B2(n16413), .A(n16412), .ZN(n16415) );
  AOI21_X1 U17337 ( .B1(n16475), .B2(n16416), .A(n16415), .ZN(n16418) );
  AOI22_X1 U17338 ( .A1(n16473), .A2(n16418), .B1(n8542), .B2(n16470), .ZN(
        P3_U3469) );
  INV_X1 U17339 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n16417) );
  AOI22_X1 U17340 ( .A1(n16447), .A2(n16418), .B1(n16417), .B2(n16562), .ZN(
        P3_U3420) );
  INV_X1 U17341 ( .A(n16419), .ZN(n16426) );
  AOI21_X1 U17342 ( .B1(n16421), .B2(n16528), .A(n16420), .ZN(n16423) );
  NAND3_X1 U17343 ( .A1(n16424), .A2(n16423), .A3(n16422), .ZN(n16425) );
  AOI21_X1 U17344 ( .B1(n16426), .B2(n16536), .A(n16425), .ZN(n16428) );
  AOI22_X1 U17345 ( .A1(n16539), .A2(n16428), .B1(n11359), .B2(n16537), .ZN(
        P1_U3538) );
  INV_X1 U17346 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n16427) );
  AOI22_X1 U17347 ( .A1(n16543), .A2(n16428), .B1(n16427), .B2(n16540), .ZN(
        P1_U3489) );
  AOI21_X1 U17348 ( .B1(n16431), .B2(n16430), .A(n16429), .ZN(n16436) );
  OAI211_X1 U17349 ( .C1(n16434), .C2(n16504), .A(n16433), .B(n16432), .ZN(
        n16435) );
  NOR2_X1 U17350 ( .A1(n16436), .A2(n16435), .ZN(n16439) );
  AOI22_X1 U17351 ( .A1(n16512), .A2(n16439), .B1(n16437), .B2(n16510), .ZN(
        P2_U3509) );
  INV_X1 U17352 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n16438) );
  AOI22_X1 U17353 ( .A1(n16516), .A2(n16439), .B1(n16438), .B2(n16513), .ZN(
        P2_U3460) );
  OAI21_X1 U17354 ( .B1(n16441), .B2(n16467), .A(n16440), .ZN(n16442) );
  AOI21_X1 U17355 ( .B1(n16443), .B2(n16469), .A(n16442), .ZN(n16446) );
  INV_X1 U17356 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U17357 ( .A1(n16473), .A2(n16446), .B1(n16444), .B2(n16470), .ZN(
        P3_U3470) );
  INV_X1 U17358 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16445) );
  AOI22_X1 U17359 ( .A1(n16447), .A2(n16446), .B1(n16445), .B2(n16562), .ZN(
        P3_U3423) );
  OAI22_X1 U17360 ( .A1(n16450), .A2(n16495), .B1(n16449), .B2(n16448), .ZN(
        n16452) );
  AOI211_X1 U17361 ( .C1(n16453), .C2(n16536), .A(n16452), .B(n16451), .ZN(
        n16455) );
  AOI22_X1 U17362 ( .A1(n16539), .A2(n16455), .B1(n11361), .B2(n16537), .ZN(
        P1_U3539) );
  INV_X1 U17363 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n16454) );
  AOI22_X1 U17364 ( .A1(n16543), .A2(n16455), .B1(n16454), .B2(n16540), .ZN(
        P1_U3492) );
  NOR2_X1 U17365 ( .A1(n16457), .A2(n16456), .ZN(n16462) );
  OAI21_X1 U17366 ( .B1(n16459), .B2(n16504), .A(n16458), .ZN(n16461) );
  AOI211_X1 U17367 ( .C1(n16462), .C2(n12257), .A(n16461), .B(n16460), .ZN(
        n16465) );
  AOI22_X1 U17368 ( .A1(n16512), .A2(n16465), .B1(n16463), .B2(n16510), .ZN(
        P2_U3510) );
  INV_X1 U17369 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n16464) );
  AOI22_X1 U17370 ( .A1(n16516), .A2(n16465), .B1(n16464), .B2(n16513), .ZN(
        P2_U3463) );
  OAI21_X1 U17371 ( .B1(n16468), .B2(n16467), .A(n16466), .ZN(n16474) );
  AOI21_X1 U17372 ( .B1(n16469), .B2(n16477), .A(n16474), .ZN(n16472) );
  INV_X1 U17373 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n16471) );
  AOI22_X1 U17374 ( .A1(n16473), .A2(n16472), .B1(n16471), .B2(n16470), .ZN(
        P3_U3471) );
  AOI21_X1 U17375 ( .B1(n16475), .B2(n16477), .A(n16474), .ZN(n16479) );
  AOI22_X1 U17376 ( .A1(n16477), .A2(n16476), .B1(P3_REG0_REG_12__SCAN_IN), 
        .B2(n16562), .ZN(n16478) );
  OAI21_X1 U17377 ( .B1(n16479), .B2(n16562), .A(n16478), .ZN(P3_U3426) );
  INV_X1 U17378 ( .A(n16484), .ZN(n16487) );
  AOI211_X1 U17379 ( .C1(n16482), .C2(n16528), .A(n16481), .B(n16480), .ZN(
        n16483) );
  OAI21_X1 U17380 ( .B1(n16485), .B2(n16484), .A(n16483), .ZN(n16486) );
  AOI21_X1 U17381 ( .B1(n16488), .B2(n16487), .A(n16486), .ZN(n16490) );
  AOI22_X1 U17382 ( .A1(n16539), .A2(n16490), .B1(n11606), .B2(n16537), .ZN(
        P1_U3540) );
  INV_X1 U17383 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U17384 ( .A1(n16543), .A2(n16490), .B1(n16489), .B2(n16540), .ZN(
        P1_U3495) );
  INV_X1 U17385 ( .A(n16491), .ZN(n16492) );
  AOI21_X1 U17386 ( .B1(n16493), .B2(n16528), .A(n16492), .ZN(n16494) );
  OAI21_X1 U17387 ( .B1(n16496), .B2(n16495), .A(n16494), .ZN(n16499) );
  NOR2_X1 U17388 ( .A1(n16497), .A2(n16532), .ZN(n16498) );
  AOI211_X1 U17389 ( .C1(n16500), .C2(n16536), .A(n16499), .B(n16498), .ZN(
        n16502) );
  AOI22_X1 U17390 ( .A1(n16539), .A2(n16502), .B1(n11610), .B2(n16537), .ZN(
        P1_U3541) );
  INV_X1 U17391 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n16501) );
  AOI22_X1 U17392 ( .A1(n16543), .A2(n16502), .B1(n16501), .B2(n16540), .ZN(
        P1_U3498) );
  OAI21_X1 U17393 ( .B1(n16505), .B2(n16504), .A(n16503), .ZN(n16507) );
  AOI211_X1 U17394 ( .C1(n16509), .C2(n16508), .A(n16507), .B(n16506), .ZN(
        n16515) );
  AOI22_X1 U17395 ( .A1(n16512), .A2(n16515), .B1(n16511), .B2(n16510), .ZN(
        P2_U3512) );
  INV_X1 U17396 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n16514) );
  AOI22_X1 U17397 ( .A1(n16516), .A2(n16515), .B1(n16514), .B2(n16513), .ZN(
        P2_U3469) );
  NAND2_X1 U17398 ( .A1(n16518), .A2(n16517), .ZN(n16519) );
  NAND2_X1 U17399 ( .A1(n16520), .A2(n16519), .ZN(n16521) );
  AOI222_X1 U17400 ( .A1(n16551), .A2(n16523), .B1(n16522), .B2(n16548), .C1(
        n16521), .C2(n16546), .ZN(n16525) );
  OAI211_X1 U17401 ( .C1(n16555), .C2(n16526), .A(n16525), .B(n16524), .ZN(
        P1_U3215) );
  AOI21_X1 U17402 ( .B1(n16529), .B2(n16528), .A(n16527), .ZN(n16531) );
  OAI211_X1 U17403 ( .C1(n16533), .C2(n16532), .A(n16531), .B(n16530), .ZN(
        n16534) );
  AOI21_X1 U17404 ( .B1(n16536), .B2(n16535), .A(n16534), .ZN(n16542) );
  AOI22_X1 U17405 ( .A1(n16539), .A2(n16542), .B1(n16538), .B2(n16537), .ZN(
        P1_U3543) );
  INV_X1 U17406 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n16541) );
  AOI22_X1 U17407 ( .A1(n16543), .A2(n16542), .B1(n16541), .B2(n16540), .ZN(
        P1_U3504) );
  OAI21_X1 U17408 ( .B1(n16545), .B2(n16544), .A(n15037), .ZN(n16547) );
  AOI222_X1 U17409 ( .A1(n16551), .A2(n16550), .B1(n16549), .B2(n16548), .C1(
        n16547), .C2(n16546), .ZN(n16553) );
  OAI211_X1 U17410 ( .C1(n16555), .C2(n16554), .A(n16553), .B(n16552), .ZN(
        P1_U3226) );
  AOI22_X1 U17411 ( .A1(n16558), .A2(n16556), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n16562), .ZN(n16557) );
  OAI21_X1 U17412 ( .B1(n16562), .B2(n16561), .A(n16557), .ZN(P3_U3457) );
  AOI22_X1 U17413 ( .A1(n16559), .A2(n16558), .B1(P3_REG0_REG_31__SCAN_IN), 
        .B2(n16562), .ZN(n16560) );
  OAI21_X1 U17414 ( .B1(n16562), .B2(n16561), .A(n16560), .ZN(P3_U3458) );
  AOI21_X1 U17415 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16563) );
  OAI21_X1 U17416 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16563), 
        .ZN(U28) );
  NAND2_X1 U7505 ( .A1(n8299), .A2(n8298), .ZN(n11565) );
  CLKBUF_X3 U7470 ( .A(n8827), .Z(n10830) );
  BUF_X1 U7472 ( .A(n9358), .Z(n7365) );
  CLKBUF_X1 U7474 ( .A(n10296), .Z(n10505) );
  CLKBUF_X1 U7483 ( .A(n8862), .Z(n8933) );
  OAI211_X1 U7484 ( .C1(n9009), .C2(n7781), .A(n7778), .B(n7776), .ZN(n9015)
         );
  CLKBUF_X1 U7501 ( .A(n15311), .Z(n7363) );
  OR2_X1 U7511 ( .A1(n11281), .A2(n9598), .ZN(n16567) );
endmodule

