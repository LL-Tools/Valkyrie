

module b15_C_AntiSAT_k_256_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3200, n3201, n3202,
         n3203, n3204, n3206, n3207, n3208, n3209, n3210, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032;

  CLKBUF_X2 U3639 ( .A(n5969), .Z(n3197) );
  OAI221_X1 U3640 ( .B1(n6766), .B2(keyinput155), .C1(n6765), .C2(keyinput171), 
        .A(n6764), .ZN(n6774) );
  INV_X2 U3641 ( .A(n3725), .ZN(n5754) );
  BUF_X2 U3642 ( .A(n3483), .Z(n3444) );
  CLKBUF_X2 U3643 ( .A(n3463), .Z(n4431) );
  CLKBUF_X2 U3644 ( .A(n3383), .Z(n3561) );
  CLKBUF_X2 U3645 ( .A(n3371), .Z(n4299) );
  CLKBUF_X2 U3646 ( .A(n3452), .Z(n4408) );
  BUF_X1 U3648 ( .A(n3337), .Z(n4441) );
  AND4_X1 U3650 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3332)
         );
  AND2_X2 U3651 ( .A1(n3317), .A2(n5337), .ZN(n3629) );
  AOI22_X1 U3652 ( .A1(n6872), .A2(keyinput135), .B1(n6780), .B2(keyinput192), 
        .ZN(n6779) );
  AOI22_X1 U3653 ( .A1(n6766), .A2(keyinput155), .B1(n6765), .B2(keyinput171), 
        .ZN(n6764) );
  CLKBUF_X2 U3654 ( .A(n3360), .Z(n3446) );
  CLKBUF_X2 U3655 ( .A(n3629), .Z(n3206) );
  AOI22_X1 U3656 ( .A1(n6913), .A2(keyinput89), .B1(keyinput69), .B2(n6912), 
        .ZN(n6911) );
  OAI221_X1 U3657 ( .B1(n6872), .B2(keyinput135), .C1(n6780), .C2(keyinput192), 
        .A(n6779), .ZN(n6785) );
  OAI221_X1 U3659 ( .B1(n6913), .B2(keyinput89), .C1(n6912), .C2(keyinput69), 
        .A(n6911), .ZN(n6925) );
  AND2_X2 U3660 ( .A1(n3767), .A2(n3801), .ZN(n3755) );
  NAND2_X1 U3661 ( .A1(n4717), .A2(n3834), .ZN(n3916) );
  NAND2_X1 U3663 ( .A1(n3441), .A2(n3938), .ZN(n3514) );
  INV_X1 U3664 ( .A(n3478), .ZN(n3192) );
  INV_X1 U3665 ( .A(n3834), .ZN(n3472) );
  AND2_X1 U3666 ( .A1(n4699), .A2(n4698), .ZN(n4700) );
  INV_X1 U3667 ( .A(n4530), .ZN(n6075) );
  NAND2_X2 U3668 ( .A1(n3530), .A2(n3529), .ZN(n6308) );
  AND2_X1 U3669 ( .A1(n4533), .A2(n4565), .ZN(n6081) );
  NAND2_X1 U3670 ( .A1(n5479), .A2(n5480), .ZN(n4467) );
  NAND2_X2 U3671 ( .A1(n3652), .A2(n3651), .ZN(n4788) );
  NAND2_X2 U3672 ( .A1(n3332), .A2(n3331), .ZN(n3412) );
  AND4_X2 U3673 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3331)
         );
  AND4_X2 U3674 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3213)
         );
  NAND3_X2 U3675 ( .A1(n3322), .A2(n3321), .A3(n3320), .ZN(n3411) );
  AND4_X2 U3676 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3322)
         );
  NAND2_X2 U3677 ( .A1(n3257), .A2(n3540), .ZN(n6187) );
  NAND2_X2 U3678 ( .A1(n4906), .A2(n4599), .ZN(n3376) );
  AND3_X2 U3679 ( .A1(n3316), .A2(n3315), .A3(n3314), .ZN(n3321) );
  INV_X4 U3680 ( .A(n3348), .ZN(n3678) );
  OR2_X4 U3681 ( .A1(n3382), .A2(n3381), .ZN(n3834) );
  INV_X1 U3682 ( .A(n5754), .ZN(n5756) );
  INV_X2 U3683 ( .A(n6002), .ZN(n6017) );
  AND2_X1 U3684 ( .A1(n3598), .A2(n3597), .ZN(n3798) );
  BUF_X2 U3685 ( .A(n3408), .Z(n4528) );
  AND2_X1 U3686 ( .A1(n3531), .A2(n3827), .ZN(n5544) );
  INV_X2 U3687 ( .A(n3412), .ZN(n4993) );
  NAND2_X1 U3688 ( .A1(n3393), .A2(n3392), .ZN(n3531) );
  NOR2_X4 U3690 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4901) );
  AOI21_X1 U3691 ( .B1(n6189), .B2(n5738), .A(n5737), .ZN(n5740) );
  OAI22_X1 U3692 ( .A1(n5503), .A2(n4480), .B1(n5423), .B2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4482) );
  XNOR2_X1 U3693 ( .A(n5503), .B(n3272), .ZN(n5732) );
  NOR2_X1 U3694 ( .A1(n5515), .A2(n5514), .ZN(n5513) );
  AOI21_X1 U3695 ( .B1(n3273), .B2(n3214), .A(n3233), .ZN(n5430) );
  AOI21_X1 U3696 ( .B1(n4398), .B2(n6189), .A(n4397), .ZN(n4399) );
  AOI221_X1 U3697 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5624), .C1(n5623), .C2(
        n5624), .A(n5622), .ZN(n5625) );
  OR2_X1 U3698 ( .A1(n5686), .A2(n6203), .ZN(n4559) );
  XNOR2_X1 U3699 ( .A(n4461), .B(n4460), .ZN(n4569) );
  AND2_X1 U3700 ( .A1(n4558), .A2(n4557), .ZN(n4461) );
  INV_X1 U3701 ( .A(n5418), .ZN(n5691) );
  AND2_X1 U3702 ( .A1(n5369), .A2(n5368), .ZN(n5727) );
  NAND2_X1 U3703 ( .A1(n3726), .A2(n6158), .ZN(n5444) );
  AOI21_X1 U3704 ( .B1(n3265), .B2(n3267), .A(n3226), .ZN(n3264) );
  NAND2_X1 U3705 ( .A1(n3675), .A2(n3674), .ZN(n4746) );
  NOR2_X1 U3706 ( .A1(n4752), .A2(n3231), .ZN(n3278) );
  AND2_X1 U3707 ( .A1(n4032), .A2(n4031), .ZN(n4752) );
  NAND2_X1 U3708 ( .A1(n3621), .A2(n3620), .ZN(n4697) );
  OAI21_X1 U3709 ( .B1(n4017), .B2(n3648), .A(n3647), .ZN(n3650) );
  XNOR2_X1 U3710 ( .A(n3707), .B(n3706), .ZN(n4033) );
  XNOR2_X1 U3711 ( .A(n3619), .B(n4880), .ZN(n4708) );
  NAND2_X1 U3712 ( .A1(n3693), .A2(n3692), .ZN(n3707) );
  CLKBUF_X1 U3713 ( .A(n3997), .Z(n6271) );
  AND2_X1 U3714 ( .A1(n3677), .A2(n3676), .ZN(n3693) );
  NOR2_X1 U3715 ( .A1(n3639), .A2(n3638), .ZN(n3677) );
  CLKBUF_X1 U3716 ( .A(n5329), .Z(n6088) );
  NAND2_X1 U3717 ( .A1(n3613), .A2(n3612), .ZN(n4732) );
  AND2_X1 U3718 ( .A1(n5965), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5299) );
  CLKBUF_X1 U3719 ( .A(n4719), .Z(n5058) );
  NAND2_X2 U3720 ( .A1(n6616), .A2(n4496), .ZN(n5965) );
  NAND2_X1 U3721 ( .A1(n4638), .A2(n3989), .ZN(n5143) );
  BUF_X1 U3722 ( .A(n3593), .Z(n4895) );
  OR2_X1 U3723 ( .A1(n4635), .A2(n4636), .ZN(n4638) );
  AND2_X1 U3724 ( .A1(n3987), .A2(n3986), .ZN(n4635) );
  NAND2_X1 U3725 ( .A1(n3596), .A2(n3595), .ZN(n4894) );
  CLKBUF_X1 U3726 ( .A(n3820), .Z(n4619) );
  AND2_X1 U3727 ( .A1(n3437), .A2(n3440), .ZN(n3938) );
  AND3_X1 U3728 ( .A1(n4909), .A2(n3431), .A3(n3430), .ZN(n3436) );
  NAND2_X1 U3729 ( .A1(n3825), .A2(n5544), .ZN(n3940) );
  NAND2_X1 U3730 ( .A1(n3438), .A2(n3531), .ZN(n3932) );
  OR2_X1 U3731 ( .A1(n3471), .A2(n3470), .ZN(n3532) );
  OR2_X1 U3732 ( .A1(n3458), .A2(n3457), .ZN(n3716) );
  CLKBUF_X1 U3734 ( .A(n3759), .Z(n5038) );
  BUF_X2 U3735 ( .A(n3412), .Z(n5327) );
  NOR2_X1 U3736 ( .A1(n5952), .A2(n4039), .ZN(n4066) );
  INV_X2 U3737 ( .A(n3419), .ZN(n4999) );
  NAND3_X2 U3738 ( .A1(n3369), .A2(n3368), .A3(n3301), .ZN(n3827) );
  NAND3_X1 U3739 ( .A1(n3305), .A2(n3344), .A3(n3343), .ZN(n3419) );
  AND4_X1 U3740 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3392)
         );
  AND4_X1 U3741 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3393)
         );
  AND4_X1 U3742 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3368)
         );
  NOR2_X1 U3743 ( .A1(n6203), .A2(n4931), .ZN(n6394) );
  NOR2_X2 U3744 ( .A1(n6203), .A2(n5000), .ZN(n5001) );
  AND3_X1 U3745 ( .A1(n3342), .A2(n3341), .A3(n3340), .ZN(n3343) );
  CLKBUF_X2 U3746 ( .A(n3605), .Z(n3484) );
  NOR2_X2 U3747 ( .A1(n6203), .A2(n5042), .ZN(n5043) );
  INV_X1 U3748 ( .A(n3337), .ZN(n4069) );
  OR2_X2 U3749 ( .A1(n6536), .A2(n6617), .ZN(n6203) );
  INV_X1 U3750 ( .A(n3445), .ZN(n3485) );
  INV_X2 U3751 ( .A(n6631), .ZN(n6629) );
  INV_X2 U3752 ( .A(n3445), .ZN(n3202) );
  INV_X2 U3753 ( .A(n6619), .ZN(n3193) );
  NAND2_X2 U3754 ( .A1(n4900), .A2(n4599), .ZN(n3445) );
  AND2_X2 U3755 ( .A1(n3306), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5333)
         );
  AND2_X2 U3756 ( .A1(n3308), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5337)
         );
  NOR2_X2 U3757 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4458) );
  AND2_X2 U3758 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4900) );
  CLKBUF_X1 U3759 ( .A(n6170), .Z(n3194) );
  CLKBUF_X1 U3760 ( .A(n5095), .Z(n3195) );
  NAND2_X1 U3761 ( .A1(n3703), .A2(n3702), .ZN(n6170) );
  NAND2_X1 U3762 ( .A1(n3713), .A2(n3712), .ZN(n5095) );
  CLKBUF_X1 U3763 ( .A(n3427), .Z(n4988) );
  INV_X2 U3764 ( .A(n4438), .ZN(n4414) );
  NAND2_X2 U3766 ( .A1(n5337), .A2(n4901), .ZN(n3337) );
  AND2_X1 U3767 ( .A1(n3429), .A2(n4857), .ZN(n3415) );
  AND2_X4 U3768 ( .A1(n3759), .A2(n3834), .ZN(n4588) );
  AND2_X1 U3769 ( .A1(n3834), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3767) );
  AND2_X2 U3770 ( .A1(n5333), .A2(n4901), .ZN(n4340) );
  INV_X1 U3771 ( .A(n3376), .ZN(n3443) );
  AND2_X2 U3772 ( .A1(n5337), .A2(n4900), .ZN(n3483) );
  AND2_X2 U3773 ( .A1(n4906), .A2(n5337), .ZN(n3442) );
  AND2_X1 U3774 ( .A1(n4900), .A2(n5333), .ZN(n3196) );
  AND2_X2 U3775 ( .A1(n4900), .A2(n5333), .ZN(n3605) );
  NAND2_X4 U3776 ( .A1(n3317), .A2(n4921), .ZN(n3348) );
  OAI21_X1 U3777 ( .B1(n3409), .B2(n4999), .A(n3410), .ZN(n3416) );
  INV_X1 U3778 ( .A(n3206), .ZN(n3198) );
  NAND2_X2 U3779 ( .A1(n5403), .A2(n3282), .ZN(n5394) );
  NAND2_X2 U3780 ( .A1(n4131), .A2(n4130), .ZN(n5403) );
  NOR2_X4 U3782 ( .A1(n5394), .A2(n5762), .ZN(n5387) );
  XNOR2_X2 U3783 ( .A(n3576), .B(n3575), .ZN(n3578) );
  NAND2_X1 U3784 ( .A1(n3639), .A2(n3615), .ZN(n5577) );
  AND2_X2 U3785 ( .A1(n3243), .A2(n3242), .ZN(n3227) );
  OR2_X4 U3786 ( .A1(n3715), .A2(n3476), .ZN(n3725) );
  NAND2_X2 U3787 ( .A1(n4390), .A2(n4389), .ZN(n5618) );
  AOI21_X1 U3788 ( .B1(n3262), .B2(n3723), .A(n3260), .ZN(n3259) );
  NOR2_X1 U3789 ( .A1(n5765), .A2(n3735), .ZN(n5757) );
  OAI21_X1 U3790 ( .B1(n5577), .B2(n4160), .A(n4009), .ZN(n4711) );
  NAND2_X2 U3791 ( .A1(n3722), .A2(n3721), .ZN(n6164) );
  AND2_X1 U3792 ( .A1(n3834), .A2(n3827), .ZN(n4530) );
  INV_X1 U3793 ( .A(n3376), .ZN(n3200) );
  INV_X1 U3794 ( .A(n3445), .ZN(n3201) );
  INV_X1 U3795 ( .A(n3202), .ZN(n3203) );
  NOR2_X2 U3796 ( .A1(n5388), .A2(n3286), .ZN(n5374) );
  NAND2_X2 U3797 ( .A1(n5387), .A2(n5390), .ZN(n5388) );
  AND2_X2 U3799 ( .A1(n4599), .A2(n3317), .ZN(n3478) );
  INV_X1 U3800 ( .A(n3348), .ZN(n3207) );
  INV_X2 U3801 ( .A(n3348), .ZN(n3208) );
  INV_X1 U3802 ( .A(n3192), .ZN(n3209) );
  INV_X1 U3803 ( .A(n3192), .ZN(n3210) );
  NAND2_X1 U3806 ( .A1(n3358), .A2(n4857), .ZN(n3803) );
  OR2_X1 U3807 ( .A1(n3418), .A2(n3801), .ZN(n3420) );
  AND2_X1 U3808 ( .A1(n4528), .A2(n4857), .ZN(n3421) );
  NAND2_X1 U3809 ( .A1(n6092), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3598) );
  NAND2_X1 U3810 ( .A1(n4999), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3597) );
  OR2_X1 U3811 ( .A1(n4857), .A2(n6403), .ZN(n3298) );
  NAND2_X1 U3812 ( .A1(n3835), .A2(n6075), .ZN(n3908) );
  OR2_X1 U3813 ( .A1(n4858), .A2(n3802), .ZN(n4173) );
  NAND2_X1 U3814 ( .A1(n3755), .A2(n3786), .ZN(n3800) );
  INV_X1 U3815 ( .A(n3754), .ZN(n3813) );
  AOI221_X1 U3816 ( .B1(n3756), .B2(n5840), .C1(n3756), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n3753), .ZN(n3754) );
  OR2_X1 U3817 ( .A1(n4578), .A2(n4580), .ZN(n4584) );
  INV_X1 U3818 ( .A(n6529), .ZN(n4565) );
  AND2_X1 U3819 ( .A1(n4606), .A2(n4565), .ZN(n5597) );
  NAND2_X1 U3820 ( .A1(n4479), .A2(n3294), .ZN(n5503) );
  AND2_X1 U3821 ( .A1(n5790), .A2(n5547), .ZN(n5525) );
  INV_X1 U3822 ( .A(n3669), .ZN(n3694) );
  INV_X1 U3823 ( .A(n3645), .ZN(n3643) );
  INV_X1 U3824 ( .A(n3520), .ZN(n3517) );
  OR2_X1 U3825 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  OR2_X1 U3826 ( .A1(n3611), .A2(n3610), .ZN(n3641) );
  AND2_X1 U3827 ( .A1(n5374), .A2(n5375), .ZN(n4486) );
  NOR2_X1 U3828 ( .A1(n3288), .A2(n5384), .ZN(n3287) );
  NOR2_X2 U3829 ( .A1(n4173), .A2(n6523), .ZN(n4455) );
  INV_X1 U3830 ( .A(n4751), .ZN(n3279) );
  NAND2_X1 U3831 ( .A1(n5725), .A2(n5726), .ZN(n3971) );
  INV_X1 U3832 ( .A(n5516), .ZN(n3251) );
  INV_X1 U3833 ( .A(n5269), .ZN(n3260) );
  NAND2_X1 U3834 ( .A1(n3837), .A2(n3220), .ZN(n3841) );
  NAND2_X1 U3835 ( .A1(n3204), .A2(n4530), .ZN(n3917) );
  INV_X1 U3836 ( .A(n3573), .ZN(n3586) );
  XNOR2_X1 U3837 ( .A(n4895), .B(n4894), .ZN(n4719) );
  OR2_X1 U3838 ( .A1(n3807), .A2(n3808), .ZN(n4580) );
  AND2_X1 U3839 ( .A1(n3947), .A2(n3943), .ZN(n4623) );
  INV_X1 U3840 ( .A(n6543), .ZN(n5596) );
  OR2_X1 U3841 ( .A1(n4470), .A2(n5600), .ZN(n4472) );
  NAND2_X1 U3842 ( .A1(n4403), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4470)
         );
  NOR2_X2 U3843 ( .A1(n6913), .A2(n4333), .ZN(n4354) );
  NAND2_X1 U3844 ( .A1(n4264), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4313)
         );
  NAND2_X1 U3845 ( .A1(n5433), .A2(n3289), .ZN(n3288) );
  INV_X1 U3846 ( .A(n5682), .ZN(n3289) );
  CLKBUF_X1 U3847 ( .A(n5249), .Z(n5250) );
  INV_X1 U3848 ( .A(n5409), .ZN(n3742) );
  OR2_X1 U3849 ( .A1(n4543), .A2(n4544), .ZN(n5638) );
  NAND2_X1 U3850 ( .A1(n5525), .A2(n3215), .ZN(n5519) );
  NOR2_X1 U3851 ( .A1(n5816), .A2(n3885), .ZN(n5790) );
  NAND2_X1 U3852 ( .A1(n5215), .A2(n3244), .ZN(n5963) );
  NOR2_X1 U3853 ( .A1(n3246), .A2(n3245), .ZN(n3244) );
  OR2_X1 U3854 ( .A1(n5960), .A2(n5961), .ZN(n3246) );
  INV_X1 U3855 ( .A(n4796), .ZN(n3245) );
  NOR2_X1 U3856 ( .A1(n5214), .A2(n5213), .ZN(n5215) );
  NAND2_X1 U3857 ( .A1(n5837), .A2(n6523), .ZN(n6618) );
  INV_X1 U3858 ( .A(n3954), .ZN(n3949) );
  NOR2_X1 U3859 ( .A1(n4580), .A2(n5038), .ZN(n5594) );
  OR2_X1 U3860 ( .A1(n6271), .A2(n4732), .ZN(n6310) );
  INV_X2 U3861 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6403) );
  NOR2_X1 U3862 ( .A1(n3796), .A2(n3795), .ZN(n3797) );
  NAND2_X1 U3863 ( .A1(n3296), .A2(n3351), .ZN(n3357) );
  AND2_X1 U3864 ( .A1(n4669), .A2(n4567), .ZN(n6089) );
  INV_X1 U3865 ( .A(n6089), .ZN(n5405) );
  INV_X1 U3866 ( .A(n5618), .ZN(n4398) );
  NAND2_X1 U3867 ( .A1(n6198), .A2(n5731), .ZN(n3269) );
  OR2_X1 U3868 ( .A1(n5734), .A2(n6203), .ZN(n3270) );
  INV_X1 U3869 ( .A(n5741), .ZN(n6194) );
  AND2_X1 U3870 ( .A1(n5741), .A2(n4639), .ZN(n6198) );
  AND2_X1 U3871 ( .A1(n5597), .A2(n4577), .ZN(n6199) );
  XNOR2_X1 U3872 ( .A(n4520), .B(n4519), .ZN(n6025) );
  INV_X1 U3873 ( .A(n5504), .ZN(n3272) );
  INV_X1 U3874 ( .A(n4716), .ZN(n6309) );
  NAND2_X1 U3875 ( .A1(n3408), .A2(n4999), .ZN(n3413) );
  NAND2_X1 U3876 ( .A1(n3409), .A2(n3933), .ZN(n3410) );
  XNOR2_X1 U3877 ( .A(n3750), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3757)
         );
  AND2_X1 U3878 ( .A1(n3498), .A2(n3497), .ZN(n3511) );
  AOI22_X1 U3879 ( .A1(n3629), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U3880 ( .A1(n3605), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U3881 ( .A1(n4340), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U3882 ( .A1(n3409), .A2(n4993), .ZN(n3408) );
  INV_X1 U3883 ( .A(n5115), .ZN(n3281) );
  OR2_X1 U3884 ( .A1(n3798), .A2(n3694), .ZN(n3667) );
  AND2_X1 U3885 ( .A1(n3637), .A2(n3636), .ZN(n3638) );
  OR2_X1 U3886 ( .A1(n3688), .A2(n3687), .ZN(n3696) );
  OR2_X1 U3887 ( .A1(n3665), .A2(n3664), .ZN(n3669) );
  OR2_X1 U3888 ( .A1(n3635), .A2(n3634), .ZN(n3645) );
  INV_X1 U3889 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U3890 ( .A1(n4340), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U3891 ( .A1(n4340), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3485), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3342) );
  INV_X1 U3892 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U3893 ( .A1(n3629), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3328) );
  NOR2_X1 U3894 ( .A1(n3505), .A2(n3763), .ZN(n3783) );
  AOI21_X1 U3895 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n4948), .A(n3752), 
        .ZN(n3756) );
  NOR2_X1 U3896 ( .A1(n3751), .A2(n3757), .ZN(n3752) );
  INV_X1 U3897 ( .A(n3758), .ZN(n3751) );
  NAND2_X1 U3898 ( .A1(n3500), .A2(n3499), .ZN(n3820) );
  INV_X1 U3899 ( .A(n3803), .ZN(n3500) );
  INV_X1 U3900 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4249) );
  AND2_X1 U3901 ( .A1(n3283), .A2(n5395), .ZN(n3282) );
  INV_X1 U3902 ( .A(n4129), .ZN(n4114) );
  NAND2_X1 U3903 ( .A1(n5525), .A2(n3237), .ZN(n4543) );
  INV_X1 U3904 ( .A(n3239), .ZN(n3250) );
  NAND2_X1 U3905 ( .A1(n4477), .A2(n3276), .ZN(n3275) );
  INV_X1 U3906 ( .A(n3737), .ZN(n3276) );
  NOR2_X1 U3907 ( .A1(n3735), .A2(n3222), .ZN(n3277) );
  INV_X1 U3908 ( .A(n3266), .ZN(n3265) );
  OAI21_X1 U3909 ( .B1(n3730), .B2(n3267), .A(n3733), .ZN(n3266) );
  INV_X1 U3910 ( .A(n3732), .ZN(n3267) );
  NOR2_X1 U3911 ( .A1(n4621), .A2(n3941), .ZN(n3947) );
  INV_X1 U3912 ( .A(n5440), .ZN(n3730) );
  NOR2_X1 U3913 ( .A1(n3204), .A2(n6075), .ZN(n4512) );
  XNOR2_X1 U3914 ( .A(n3841), .B(n3241), .ZN(n3840) );
  INV_X1 U3915 ( .A(n4647), .ZN(n3241) );
  AND2_X1 U3916 ( .A1(n5327), .A2(n3827), .ZN(n3786) );
  AND2_X1 U3917 ( .A1(n3805), .A2(n3806), .ZN(n3826) );
  OAI211_X1 U3918 ( .C1(n3517), .C2(n3598), .A(n3494), .B(n3493), .ZN(n3580)
         );
  NAND2_X1 U3919 ( .A1(n3555), .A2(n3554), .ZN(n3558) );
  AND2_X2 U3920 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4599) );
  AND2_X1 U3921 ( .A1(n5577), .A2(n6271), .ZN(n4941) );
  NAND2_X1 U3922 ( .A1(n4719), .A2(n6523), .ZN(n3613) );
  INV_X1 U3923 ( .A(n3827), .ZN(n3759) );
  AOI21_X1 U3924 ( .B1(n6535), .B2(n5592), .A(n5343), .ZN(n4723) );
  INV_X1 U3925 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6506) );
  AND4_X1 U3926 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n4609), .ZN(n4613)
         );
  INV_X1 U3927 ( .A(n4588), .ZN(n6623) );
  NOR2_X1 U3928 ( .A1(n4619), .A2(n6092), .ZN(n4583) );
  NOR2_X1 U3929 ( .A1(n6579), .A2(n5669), .ZN(n5658) );
  NOR2_X1 U3930 ( .A1(n6574), .A2(n5872), .ZN(n5865) );
  OR2_X1 U3931 ( .A1(n4573), .A2(READY_N), .ZN(n4592) );
  NOR2_X1 U3932 ( .A1(n4402), .A2(n4401), .ZN(n4403) );
  AND2_X1 U3933 ( .A1(n4428), .A2(n4427), .ZN(n4538) );
  OR2_X1 U3934 ( .A1(n5608), .A2(n4493), .ZN(n4428) );
  AOI22_X1 U3935 ( .A1(n4458), .A2(n5719), .B1(n4353), .B2(n4352), .ZN(n5364)
         );
  NOR2_X1 U3936 ( .A1(n4313), .A2(n4484), .ZN(n4314) );
  NAND2_X1 U3937 ( .A1(n4314), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4333)
         );
  NOR2_X1 U3938 ( .A1(n4250), .A2(n4249), .ZN(n4264) );
  AND2_X1 U3939 ( .A1(n4290), .A2(n4289), .ZN(n5375) );
  OR2_X1 U3940 ( .A1(n5650), .A2(n4493), .ZN(n4290) );
  NAND2_X1 U3941 ( .A1(n5381), .A2(n3287), .ZN(n3286) );
  CLKBUF_X1 U3942 ( .A(n4486), .Z(n4487) );
  INV_X1 U3943 ( .A(n3287), .ZN(n3285) );
  NOR2_X1 U3944 ( .A1(n6780), .A2(n4222), .ZN(n4235) );
  NOR2_X1 U3945 ( .A1(n4207), .A2(n5867), .ZN(n4208) );
  CLKBUF_X1 U3946 ( .A(n5388), .Z(n5389) );
  NAND2_X1 U3947 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n4178), .ZN(n4207)
         );
  INV_X1 U3948 ( .A(n4163), .ZN(n4164) );
  INV_X1 U3949 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6766) );
  NOR2_X1 U3950 ( .A1(n6766), .A2(n4164), .ZN(n4178) );
  NOR2_X1 U3951 ( .A1(n5400), .A2(n3284), .ZN(n3283) );
  INV_X1 U3952 ( .A(n5404), .ZN(n3284) );
  NAND2_X1 U3953 ( .A1(n4146), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4147)
         );
  NOR2_X1 U3954 ( .A1(n6933), .A2(n4147), .ZN(n4163) );
  AND2_X1 U3955 ( .A1(n4132), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4146)
         );
  INV_X1 U3956 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5916) );
  NOR2_X1 U3957 ( .A1(n5916), .A2(n4096), .ZN(n4132) );
  NAND2_X1 U3958 ( .A1(n4066), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4067)
         );
  NOR2_X1 U3959 ( .A1(n6771), .A2(n4067), .ZN(n4095) );
  AND2_X1 U3960 ( .A1(n5252), .A2(n5251), .ZN(n5935) );
  CLKBUF_X1 U3961 ( .A(n5113), .Z(n5114) );
  INV_X1 U3962 ( .A(n5133), .ZN(n3280) );
  NAND2_X1 U3963 ( .A1(n4034), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4039)
         );
  INV_X1 U3964 ( .A(n4019), .ZN(n4020) );
  NAND2_X1 U3965 ( .A1(n4020), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4027)
         );
  CLKBUF_X1 U3966 ( .A(n4700), .Z(n4701) );
  NOR2_X1 U3967 ( .A1(n4003), .A2(n6011), .ZN(n4013) );
  NAND2_X1 U3968 ( .A1(n4716), .A2(n4141), .ZN(n3994) );
  NAND2_X1 U3969 ( .A1(n5484), .A2(n3254), .ZN(n4536) );
  NOR2_X1 U3970 ( .A1(n3256), .A2(n3255), .ZN(n3254) );
  INV_X1 U3971 ( .A(n3974), .ZN(n3255) );
  AND2_X1 U3972 ( .A1(n3252), .A2(n3253), .ZN(n5484) );
  INV_X1 U3973 ( .A(n5485), .ZN(n3252) );
  AND2_X1 U3974 ( .A1(n5484), .A2(n5471), .ZN(n5469) );
  OAI21_X1 U3975 ( .B1(n5540), .B2(n3740), .A(n3739), .ZN(n5725) );
  AOI22_X1 U3976 ( .A1(n5430), .A2(n5431), .B1(n3725), .B2(n4478), .ZN(n5515)
         );
  INV_X1 U3977 ( .A(n3204), .ZN(n5526) );
  OR3_X1 U3978 ( .A1(n5925), .A2(n3229), .A3(n3248), .ZN(n3247) );
  INV_X1 U3979 ( .A(n5568), .ZN(n3248) );
  NAND2_X1 U3980 ( .A1(n3731), .A2(n3730), .ZN(n5437) );
  AND3_X1 U3981 ( .A1(n3869), .A2(n3908), .A3(n3868), .ZN(n5914) );
  NOR3_X1 U3982 ( .A1(n5924), .A2(n5925), .A3(n3229), .ZN(n5822) );
  NOR2_X1 U3983 ( .A1(n5924), .A2(n5925), .ZN(n5923) );
  AND2_X1 U3984 ( .A1(n3238), .A2(n3724), .ZN(n3262) );
  OR2_X1 U3985 ( .A1(n5945), .A2(n5274), .ZN(n5924) );
  NAND2_X1 U3986 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  AND3_X1 U3987 ( .A1(n3859), .A2(n3908), .A3(n3858), .ZN(n5100) );
  NOR2_X1 U3988 ( .A1(n5963), .A2(n5100), .ZN(n5944) );
  AND3_X1 U3989 ( .A1(n3854), .A2(n3908), .A3(n3853), .ZN(n5961) );
  NAND2_X1 U3990 ( .A1(n5215), .A2(n4796), .ZN(n5962) );
  NOR2_X1 U3991 ( .A1(n6243), .A2(n4848), .ZN(n4794) );
  INV_X1 U3992 ( .A(n6255), .ZN(n5804) );
  OR2_X1 U3993 ( .A1(n5301), .A2(n3848), .ZN(n5214) );
  INV_X1 U3994 ( .A(n3840), .ZN(n6076) );
  AND2_X1 U3995 ( .A1(n3539), .A2(n3540), .ZN(n6195) );
  NAND2_X1 U3996 ( .A1(n6196), .A2(n6195), .ZN(n3257) );
  AND2_X1 U3997 ( .A1(n3826), .A2(n3505), .ZN(n4622) );
  NAND2_X1 U3998 ( .A1(n5526), .A2(n3916), .ZN(n4645) );
  AND2_X1 U3999 ( .A1(n3824), .A2(n3823), .ZN(n3954) );
  NAND3_X1 U4000 ( .A1(n3577), .A2(n3578), .A3(n4732), .ZN(n3639) );
  CLKBUF_X1 U4001 ( .A(n4599), .Z(n4600) );
  NOR2_X1 U4002 ( .A1(n6310), .A2(n6390), .ZN(n4738) );
  NOR2_X1 U4003 ( .A1(n6396), .A2(n6308), .ZN(n6391) );
  INV_X1 U4004 ( .A(n3531), .ZN(n4717) );
  INV_X1 U4005 ( .A(n6308), .ZN(n4942) );
  OR2_X1 U4006 ( .A1(n6604), .A2(n4723), .ZN(n5039) );
  INV_X1 U4007 ( .A(n6400), .ZN(n6315) );
  AND2_X1 U4008 ( .A1(n5334), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3818) );
  INV_X1 U4009 ( .A(n4458), .ZN(n4493) );
  OR2_X1 U4010 ( .A1(n4619), .A2(n6623), .ZN(n6519) );
  NAND2_X1 U4011 ( .A1(n5597), .A2(n4583), .ZN(n4573) );
  INV_X1 U4012 ( .A(n4584), .ZN(n4492) );
  OR2_X1 U4013 ( .A1(n4502), .A2(n4501), .ZN(n4503) );
  OR2_X1 U4014 ( .A1(n5292), .A2(n5290), .ZN(n5969) );
  INV_X1 U4015 ( .A(n3197), .ZN(n5978) );
  INV_X1 U4016 ( .A(n5997), .ZN(n5993) );
  INV_X1 U4017 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6011) );
  CLKBUF_X1 U4018 ( .A(n4720), .Z(n4721) );
  NAND2_X1 U4019 ( .A1(n5965), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6012) );
  INV_X1 U4020 ( .A(n6012), .ZN(n6000) );
  AND2_X1 U4021 ( .A1(n5292), .A2(n5291), .ZN(n6002) );
  INV_X1 U4022 ( .A(n6081), .ZN(n6068) );
  INV_X1 U4023 ( .A(n5727), .ZN(n5697) );
  INV_X1 U4024 ( .A(n5407), .ZN(n6086) );
  NAND2_X1 U4025 ( .A1(n5405), .A2(n4860), .ZN(n5406) );
  INV_X1 U4026 ( .A(n6086), .ZN(n5398) );
  OR2_X1 U4027 ( .A1(n5592), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6619) );
  AND3_X1 U4028 ( .A1(n5597), .A2(n5596), .A3(n5595), .ZN(n6136) );
  INV_X1 U4029 ( .A(n4669), .ZN(n6153) );
  CLKBUF_X1 U4030 ( .A(n5765), .Z(n5766) );
  INV_X1 U4031 ( .A(n6198), .ZN(n6193) );
  OR2_X1 U4032 ( .A1(n6199), .A2(n4391), .ZN(n5741) );
  INV_X1 U4033 ( .A(n6199), .ZN(n6179) );
  XNOR2_X1 U4034 ( .A(n3745), .B(n6898), .ZN(n4556) );
  NAND2_X1 U4035 ( .A1(n3744), .A2(n3743), .ZN(n3745) );
  NAND2_X1 U4036 ( .A1(n5525), .A2(n3898), .ZN(n5517) );
  OR2_X1 U4037 ( .A1(n6164), .A2(n3723), .ZN(n3258) );
  OR2_X1 U4038 ( .A1(n5103), .A2(n5102), .ZN(n6234) );
  OR2_X1 U4039 ( .A1(n5561), .A2(n5828), .ZN(n6255) );
  INV_X1 U4040 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6902) );
  INV_X1 U4041 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6500) );
  CLKBUF_X1 U4042 ( .A(n4616), .Z(n4617) );
  INV_X1 U4043 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6265) );
  OAI21_X1 U4044 ( .B1(n4923), .B2(n6603), .A(n6353), .ZN(n6264) );
  INV_X1 U4045 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5334) );
  INV_X1 U4046 ( .A(n6524), .ZN(n5343) );
  NOR2_X1 U4047 ( .A1(n5836), .A2(n4615), .ZN(n5586) );
  INV_X1 U4048 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5840) );
  NOR2_X1 U4049 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5837) );
  INV_X1 U4050 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5184) );
  INV_X1 U4051 ( .A(n4947), .ZN(n5239) );
  OAI21_X1 U4052 ( .B1(n5228), .B2(n6605), .A(n5066), .ZN(n5226) );
  INV_X1 U4053 ( .A(n7024), .ZN(n5195) );
  OR2_X1 U4054 ( .A1(n6355), .A2(n6354), .ZN(n6372) );
  INV_X1 U4055 ( .A(n5282), .ZN(n6384) );
  NOR2_X1 U4056 ( .A1(n4724), .A2(n4942), .ZN(n6491) );
  NAND2_X1 U4057 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4606), .ZN(n6524) );
  NAND2_X1 U4058 ( .A1(n3818), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6529) );
  NOR2_X1 U4059 ( .A1(n6089), .A2(n4857), .ZN(n4568) );
  OR2_X1 U4060 ( .A1(n3230), .A2(n4396), .ZN(n4397) );
  NAND2_X1 U4061 ( .A1(n3271), .A2(n3224), .ZN(U2964) );
  NAND2_X1 U4062 ( .A1(n5732), .A2(n6199), .ZN(n3271) );
  AND2_X1 U4063 ( .A1(n5733), .A2(n3269), .ZN(n3268) );
  OAI21_X1 U4064 ( .B1(n6025), .B2(n6258), .A(n3227), .ZN(U2987) );
  AND2_X1 U4065 ( .A1(n5456), .A2(n5457), .ZN(n3242) );
  NOR2_X1 U4066 ( .A1(n4550), .A2(n4549), .ZN(n4551) );
  NOR2_X1 U4067 ( .A1(n5388), .A2(n3285), .ZN(n5379) );
  NAND2_X1 U4068 ( .A1(n5403), .A2(n5404), .ZN(n5399) );
  AND2_X1 U4069 ( .A1(n4750), .A2(n3234), .ZN(n5112) );
  NAND2_X1 U4070 ( .A1(n4750), .A2(n5148), .ZN(n5132) );
  AND2_X1 U4071 ( .A1(n3277), .A2(n4477), .ZN(n3214) );
  AND2_X1 U4072 ( .A1(n3898), .A2(n3251), .ZN(n3215) );
  AND2_X1 U4073 ( .A1(n3215), .A2(n3240), .ZN(n3216) );
  INV_X1 U4074 ( .A(n3442), .ZN(n3464) );
  AND2_X2 U4075 ( .A1(n4921), .A2(n4901), .ZN(n3452) );
  NOR2_X1 U4077 ( .A1(n5388), .A2(n5682), .ZN(n5432) );
  OR2_X1 U4078 ( .A1(n5924), .A2(n3247), .ZN(n3217) );
  AND4_X1 U4079 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3218)
         );
  NAND2_X1 U4080 ( .A1(n5437), .A2(n3732), .ZN(n5554) );
  XNOR2_X1 U4081 ( .A(n4558), .B(n4557), .ZN(n5686) );
  AND2_X1 U4082 ( .A1(n5358), .A2(n4388), .ZN(n4537) );
  AND2_X2 U4083 ( .A1(n3317), .A2(n5333), .ZN(n3463) );
  OR2_X1 U4084 ( .A1(n5388), .A2(n3288), .ZN(n3219) );
  XNOR2_X1 U4085 ( .A(n3668), .B(n3676), .ZN(n4018) );
  AND2_X1 U4086 ( .A1(n3908), .A2(n3836), .ZN(n3220) );
  AND3_X1 U4087 ( .A1(n3474), .A2(STATE2_REG_0__SCAN_IN), .A3(n3473), .ZN(
        n3221) );
  AND2_X1 U4088 ( .A1(n3725), .A2(n3736), .ZN(n3222) );
  OR2_X1 U4089 ( .A1(n4558), .A2(n4539), .ZN(n3223) );
  AND2_X1 U4090 ( .A1(n3270), .A2(n3268), .ZN(n3224) );
  NOR2_X1 U4091 ( .A1(n3425), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3225)
         );
  AND2_X1 U4092 ( .A1(n3725), .A2(n5567), .ZN(n3226) );
  NAND2_X1 U4093 ( .A1(n3741), .A2(n3303), .ZN(n5409) );
  NAND2_X1 U4094 ( .A1(n4038), .A2(n4037), .ZN(n5148) );
  NAND2_X1 U4095 ( .A1(n5525), .A2(n3216), .ZN(n3228) );
  OR2_X1 U4096 ( .A1(n5914), .A2(n5821), .ZN(n3229) );
  NOR2_X1 U4097 ( .A1(n4751), .A2(n4752), .ZN(n4750) );
  NAND2_X1 U4098 ( .A1(n3261), .A2(n3259), .ZN(n6156) );
  NAND2_X1 U4099 ( .A1(n3258), .A2(n3724), .ZN(n5268) );
  AND2_X1 U4100 ( .A1(n5614), .A2(n6198), .ZN(n3230) );
  AND2_X1 U4101 ( .A1(n5403), .A2(n3283), .ZN(n5393) );
  OR2_X1 U4102 ( .A1(n5133), .A2(n3281), .ZN(n3231) );
  NAND2_X1 U4103 ( .A1(n5754), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3232) );
  NOR2_X1 U4104 ( .A1(n5638), .A2(n5637), .ZN(n3253) );
  NAND2_X1 U4105 ( .A1(n3275), .A2(n3232), .ZN(n3233) );
  AND2_X1 U4106 ( .A1(n5148), .A2(n3280), .ZN(n3234) );
  AND2_X1 U4107 ( .A1(n4538), .A2(n4388), .ZN(n3235) );
  NOR2_X1 U4108 ( .A1(n5791), .A2(n5790), .ZN(n3236) );
  NAND2_X1 U4109 ( .A1(n4988), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4160) );
  NAND2_X1 U4110 ( .A1(n5146), .A2(n3998), .ZN(n5150) );
  NOR2_X1 U4111 ( .A1(n3217), .A2(n5814), .ZN(n3249) );
  OAI21_X1 U4112 ( .B1(n4017), .B2(n4160), .A(n4016), .ZN(n4698) );
  AND2_X1 U4113 ( .A1(n3216), .A2(n3250), .ZN(n3237) );
  NAND2_X1 U4114 ( .A1(n3725), .A2(n3863), .ZN(n3238) );
  OR2_X1 U4115 ( .A1(n3906), .A2(n3905), .ZN(n3239) );
  AND2_X2 U4116 ( .A1(n3307), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4906)
         );
  NAND3_X1 U4117 ( .A1(n3904), .A2(n3908), .A3(n3903), .ZN(n3240) );
  OR2_X1 U4118 ( .A1(n6618), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6256) );
  INV_X1 U4119 ( .A(n3277), .ZN(n3274) );
  AND2_X2 U4120 ( .A1(n4921), .A2(n4900), .ZN(n3371) );
  NOR2_X4 U4121 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4921) );
  OR2_X2 U4122 ( .A1(n5458), .A2(n6208), .ZN(n3243) );
  INV_X1 U4123 ( .A(n3249), .ZN(n5816) );
  INV_X1 U4124 ( .A(n3253), .ZN(n5636) );
  INV_X1 U4125 ( .A(n5471), .ZN(n3256) );
  OAI21_X1 U4126 ( .B1(n6196), .B2(n6195), .A(n3257), .ZN(n6197) );
  XNOR2_X2 U4127 ( .A(n3519), .B(n3542), .ZN(n4716) );
  NAND2_X1 U4128 ( .A1(n6164), .A2(n3262), .ZN(n3261) );
  NAND2_X1 U4129 ( .A1(n6156), .A2(n6157), .ZN(n3726) );
  NAND2_X1 U4130 ( .A1(n3731), .A2(n3265), .ZN(n3263) );
  NAND2_X1 U4131 ( .A1(n3263), .A2(n3264), .ZN(n5588) );
  INV_X1 U4132 ( .A(n5765), .ZN(n3273) );
  OR2_X2 U4133 ( .A1(n5765), .A2(n3274), .ZN(n5425) );
  NAND2_X2 U4134 ( .A1(n5425), .A2(n3737), .ZN(n5540) );
  NAND3_X1 U4135 ( .A1(n5148), .A2(n3279), .A3(n3278), .ZN(n5113) );
  AND2_X1 U4136 ( .A1(n5358), .A2(n3235), .ZN(n4558) );
  INV_X1 U4137 ( .A(n4732), .ZN(n4715) );
  NAND2_X1 U4138 ( .A1(n3577), .A2(n3578), .ZN(n3614) );
  INV_X1 U4139 ( .A(n3971), .ZN(n4464) );
  XNOR2_X1 U4140 ( .A(n3673), .B(n4849), .ZN(n4789) );
  NAND2_X1 U4141 ( .A1(n3981), .A2(n6199), .ZN(n4400) );
  NAND2_X1 U4142 ( .A1(n4556), .A2(n3833), .ZN(n3970) );
  AND2_X2 U4143 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n3309), .ZN(n3317)
         );
  AOI22_X1 U4144 ( .A1(n3678), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3387) );
  INV_X1 U4145 ( .A(n3413), .ZN(n3358) );
  INV_X1 U4146 ( .A(n3411), .ZN(n3427) );
  BUF_X1 U4147 ( .A(n3502), .Z(n3807) );
  OR2_X1 U4148 ( .A1(n3597), .A2(n3517), .ZN(n3290) );
  AND2_X1 U4149 ( .A1(n3477), .A2(n3476), .ZN(n3291) );
  NAND2_X1 U4150 ( .A1(n3542), .A2(n3543), .ZN(n3579) );
  NOR2_X1 U4151 ( .A1(n6434), .A2(n4718), .ZN(n3292) );
  INV_X1 U4152 ( .A(n4857), .ZN(n5328) );
  NAND2_X1 U4153 ( .A1(n3725), .A2(n5778), .ZN(n3293) );
  OR2_X1 U4154 ( .A1(n5754), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3294)
         );
  OR2_X1 U4155 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3295)
         );
  AND3_X1 U4156 ( .A1(n3347), .A2(n3346), .A3(n3345), .ZN(n3296) );
  OR2_X1 U4157 ( .A1(n5617), .A2(REIP_REG_28__SCAN_IN), .ZN(n3297) );
  OR2_X1 U4158 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3299)
         );
  OR2_X1 U4159 ( .A1(n3512), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3300)
         );
  INV_X1 U4160 ( .A(n6083), .ZN(n6072) );
  INV_X1 U4161 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6780) );
  INV_X1 U4162 ( .A(n3982), .ZN(n6312) );
  INV_X1 U4163 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5952) );
  AND3_X1 U4164 ( .A1(n3367), .A2(n3366), .A3(n3365), .ZN(n3301) );
  INV_X1 U4165 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4656) );
  AND3_X1 U4166 ( .A1(n4465), .A2(n5461), .A3(n6898), .ZN(n3302) );
  AND2_X1 U4167 ( .A1(n5481), .A2(n4465), .ZN(n3303) );
  OR2_X1 U4168 ( .A1(n4618), .A2(n4570), .ZN(n3304) );
  INV_X1 U4169 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6771) );
  AND4_X1 U4170 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3305)
         );
  INV_X1 U4171 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6921) );
  INV_X1 U4172 ( .A(n6617), .ZN(n6442) );
  NAND2_X1 U4173 ( .A1(n6403), .A2(n6605), .ZN(n6617) );
  INV_X1 U4174 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3750) );
  AND2_X2 U4175 ( .A1(n4906), .A2(n5333), .ZN(n3383) );
  NAND2_X1 U4176 ( .A1(n4002), .A2(n4001), .ZN(n4710) );
  NOR2_X1 U4177 ( .A1(n3827), .A2(n3810), .ZN(n3506) );
  INV_X1 U4178 ( .A(n3543), .ZN(n3544) );
  OR2_X1 U4179 ( .A1(n3798), .A2(n3782), .ZN(n3784) );
  OR2_X1 U4180 ( .A1(n3798), .A2(n3643), .ZN(n3637) );
  NAND2_X1 U4181 ( .A1(n3532), .A2(n3472), .ZN(n3473) );
  OR2_X1 U4182 ( .A1(n3491), .A2(n3490), .ZN(n3520) );
  AND2_X1 U4183 ( .A1(n3402), .A2(n3401), .ZN(n3403) );
  AND2_X1 U4184 ( .A1(n6902), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3764)
         );
  NAND2_X1 U4185 ( .A1(n3749), .A2(n3748), .ZN(n3758) );
  OR2_X1 U4186 ( .A1(n3798), .A2(n3689), .ZN(n3691) );
  AND2_X2 U4187 ( .A1(n4906), .A2(n4921), .ZN(n3370) );
  AOI22_X1 U4188 ( .A1(n3463), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3315) );
  INV_X1 U4189 ( .A(n3755), .ZN(n3793) );
  NAND2_X1 U4190 ( .A1(n3691), .A2(n3690), .ZN(n3692) );
  INV_X1 U4191 ( .A(n3558), .ZN(n3556) );
  AND4_X1 U4192 ( .A1(n3472), .A2(n4988), .A3(n4857), .A4(n3801), .ZN(n3428)
         );
  AOI22_X1 U4193 ( .A1(n3605), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3200), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4194 ( .A1(n3629), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3380) );
  OR2_X1 U4195 ( .A1(n4305), .A2(n4304), .ZN(n4315) );
  NAND2_X1 U4196 ( .A1(n3412), .A2(n3427), .ZN(n3418) );
  OR4_X1 U4197 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(n4355) );
  NAND2_X1 U4198 ( .A1(n4527), .A2(n3428), .ZN(n4909) );
  NAND2_X1 U4199 ( .A1(n3475), .A2(n3221), .ZN(n3526) );
  NAND2_X1 U4200 ( .A1(n4235), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4250)
         );
  INV_X1 U4201 ( .A(n4160), .ZN(n4141) );
  AND2_X1 U4202 ( .A1(n3866), .A2(n3865), .ZN(n5274) );
  INV_X1 U4203 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4948) );
  OAI21_X1 U4204 ( .B1(n3798), .B2(n3813), .A(n3797), .ZN(n3799) );
  NAND2_X1 U4205 ( .A1(n4095), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4096)
         );
  NAND2_X1 U4206 ( .A1(n4013), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4019)
         );
  OR2_X1 U4207 ( .A1(n5644), .A2(n4493), .ZN(n4312) );
  OR2_X1 U4208 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  INV_X1 U4209 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5867) );
  INV_X1 U4210 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6933) );
  NOR2_X1 U4212 ( .A1(n6921), .A2(n4027), .ZN(n4034) );
  AND2_X1 U4213 ( .A1(n5779), .A2(n3965), .ZN(n5454) );
  INV_X1 U4214 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4481) );
  NOR2_X1 U4215 ( .A1(n5565), .A2(n6205), .ZN(n5801) );
  OAI21_X1 U4216 ( .B1(n6187), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6185), 
        .ZN(n3592) );
  INV_X1 U4217 ( .A(n6245), .ZN(n6258) );
  NOR2_X1 U4218 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4723), .ZN(n4867) );
  OR2_X1 U4219 ( .A1(n4833), .A2(n6390), .ZN(n4839) );
  NAND2_X1 U4220 ( .A1(n4941), .A2(n6390), .ZN(n5060) );
  NAND2_X1 U4221 ( .A1(n6391), .A2(n6309), .ZN(n5282) );
  OR2_X1 U4222 ( .A1(n5577), .A2(n4800), .ZN(n6396) );
  OR2_X1 U4223 ( .A1(n4757), .A2(n6390), .ZN(n4724) );
  OR2_X1 U4224 ( .A1(n4757), .A2(n6309), .ZN(n4776) );
  OAI21_X1 U4225 ( .B1(n3813), .B2(n3800), .A(n3799), .ZN(n4606) );
  NAND2_X1 U4226 ( .A1(n4354), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4402)
         );
  NOR2_X1 U4227 ( .A1(n6874), .A2(n5660), .ZN(n5654) );
  AND2_X1 U4228 ( .A1(n5299), .A2(n4521), .ZN(n5983) );
  XNOR2_X1 U4229 ( .A(n4472), .B(n4471), .ZN(n5292) );
  INV_X1 U4230 ( .A(n5984), .ZN(n5999) );
  NOR2_X2 U4231 ( .A1(n4857), .A2(n6068), .ZN(n6071) );
  NOR2_X2 U4232 ( .A1(n6089), .A2(n4570), .ZN(n6085) );
  NOR2_X1 U4233 ( .A1(n6092), .A2(n6146), .ZN(n6110) );
  OR2_X1 U4234 ( .A1(n4592), .A2(n5038), .ZN(n4669) );
  NAND2_X1 U4235 ( .A1(n4208), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4222)
         );
  NAND2_X1 U4236 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4003) );
  INV_X1 U4237 ( .A(n6208), .ZN(n3833) );
  NOR2_X1 U4238 ( .A1(n3944), .A2(n5098), .ZN(n5565) );
  NOR2_X1 U4239 ( .A1(n5825), .A2(n4793), .ZN(n6205) );
  NAND2_X1 U4240 ( .A1(n3949), .A2(n4623), .ZN(n6243) );
  INV_X1 U4241 ( .A(n4867), .ZN(n6353) );
  NOR2_X2 U4242 ( .A1(n4839), .A2(n4942), .ZN(n5243) );
  NOR2_X1 U4243 ( .A1(n4739), .A2(n4942), .ZN(n5197) );
  INV_X1 U4244 ( .A(n6343), .ZN(n7021) );
  AND2_X1 U4245 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6316), .ZN(n6338)
         );
  INV_X1 U4246 ( .A(n6349), .ZN(n6383) );
  INV_X1 U4247 ( .A(n6432), .ZN(n6421) );
  INV_X1 U4248 ( .A(n6495), .ZN(n6441) );
  INV_X1 U4249 ( .A(n6309), .ZN(n6390) );
  INV_X1 U4250 ( .A(n6203), .ZN(n6189) );
  INV_X1 U4251 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6523) );
  INV_X1 U4252 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6554) );
  AND2_X1 U4253 ( .A1(n4575), .A2(n4573), .ZN(n6616) );
  NAND2_X1 U4254 ( .A1(n4522), .A2(n5983), .ZN(n4523) );
  INV_X1 U4255 ( .A(n5983), .ZN(n6015) );
  INV_X1 U4256 ( .A(n6021), .ZN(n5951) );
  INV_X1 U4257 ( .A(n5935), .ZN(n6051) );
  NAND2_X1 U4258 ( .A1(n5405), .A2(n4859), .ZN(n5407) );
  INV_X1 U4259 ( .A(n6126), .ZN(n6144) );
  INV_X1 U4260 ( .A(n6110), .ZN(n6117) );
  OR2_X1 U4261 ( .A1(n3193), .A2(n6136), .ZN(n6126) );
  INV_X1 U4262 ( .A(n6136), .ZN(n6146) );
  OR2_X1 U4263 ( .A1(n5458), .A2(n6179), .ZN(n4475) );
  NAND2_X1 U4264 ( .A1(n4569), .A2(n6189), .ZN(n4476) );
  OR2_X1 U4265 ( .A1(n5699), .A2(n6203), .ZN(n4490) );
  INV_X1 U4266 ( .A(n5904), .ZN(n6044) );
  AND2_X1 U4267 ( .A1(n5493), .A2(n3963), .ZN(n5779) );
  NAND2_X1 U4268 ( .A1(n3949), .A2(n3832), .ZN(n6208) );
  INV_X1 U4269 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6818) );
  AND2_X1 U4270 ( .A1(n4870), .A2(n4869), .ZN(n5247) );
  INV_X1 U4271 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5238) );
  INV_X1 U4272 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5176) );
  INV_X1 U4273 ( .A(n5197), .ZN(n5232) );
  INV_X1 U4274 ( .A(n4734), .ZN(n5200) );
  INV_X1 U4275 ( .A(n4824), .ZN(n7030) );
  OR3_X1 U4276 ( .A1(n6310), .A2(n4942), .A3(n6309), .ZN(n6343) );
  OR3_X1 U4277 ( .A1(n6310), .A2(n6309), .A3(n6308), .ZN(n6375) );
  INV_X1 U4278 ( .A(n4808), .ZN(n5287) );
  NAND2_X1 U4279 ( .A1(n4802), .A2(n4801), .ZN(n6432) );
  NAND2_X1 U4280 ( .A1(n6391), .A2(n6390), .ZN(n6495) );
  INV_X1 U4281 ( .A(n6491), .ZN(n5212) );
  INV_X1 U4282 ( .A(n4761), .ZN(n5124) );
  AOI21_X1 U4283 ( .B1(n4775), .B2(n4777), .A(n4774), .ZN(n5131) );
  INV_X1 U4284 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6605) );
  INV_X1 U4285 ( .A(n6602), .ZN(n6600) );
  INV_X1 U4286 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6544) );
  INV_X1 U4287 ( .A(n6591), .ZN(n6587) );
  OAI222_X1 U4288 ( .A1(n4541), .A2(n4540), .B1(n4513), .B2(n6081), .C1(n3223), 
        .C2(n6083), .ZN(U2830) );
  INV_X1 U4289 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3306) );
  INV_X1 U4290 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3307) );
  INV_X1 U4291 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4292 ( .A1(n3483), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3312) );
  INV_X1 U4293 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4294 ( .A1(n3478), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3311) );
  AND2_X2 U4295 ( .A1(n4901), .A2(n4599), .ZN(n3360) );
  AOI22_X1 U4296 ( .A1(n3442), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3314) );
  INV_X1 U4297 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3318) );
  OAI22_X1 U4298 ( .A1(n3348), .A2(n3318), .B1(n3337), .B2(n5176), .ZN(n3319)
         );
  INV_X1 U4299 ( .A(n3319), .ZN(n3320) );
  BUF_X2 U4300 ( .A(n3411), .Z(n3409) );
  AOI22_X1 U4301 ( .A1(n3207), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4302 ( .A1(n4069), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4303 ( .A1(n3371), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4304 ( .A1(n3478), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3200), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4305 ( .A1(n3370), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4306 ( .A1(n4340), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4307 ( .A1(n3463), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4308 ( .A1(n3605), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3200), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4309 ( .A1(n3483), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4310 ( .A1(n3478), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4311 ( .A1(n3629), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3333) );
  OAI22_X1 U4312 ( .A1(n3348), .A2(n3338), .B1(n3337), .B2(n5184), .ZN(n3339)
         );
  INV_X1 U4313 ( .A(n3339), .ZN(n3344) );
  AOI22_X1 U4314 ( .A1(n3442), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4315 ( .A1(n3463), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4316 ( .A1(n4340), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3485), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4317 ( .A1(n3442), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4318 ( .A1(n3463), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3345) );
  INV_X1 U4319 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3349) );
  INV_X1 U4320 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4955) );
  OAI22_X1 U4321 ( .A1(n3349), .A2(n3348), .B1(n3337), .B2(n4955), .ZN(n3350)
         );
  INV_X1 U4322 ( .A(n3350), .ZN(n3351) );
  AOI22_X1 U4323 ( .A1(n3629), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4324 ( .A1(n3483), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4325 ( .A1(n3478), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4326 ( .A1(n3605), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3352) );
  NAND4_X1 U4327 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3356)
         );
  OR2_X2 U4328 ( .A1(n3357), .A2(n3356), .ZN(n4857) );
  OAI22_X1 U4329 ( .A1(n3348), .A2(n6831), .B1(n3337), .B2(n5238), .ZN(n3359)
         );
  INV_X1 U4330 ( .A(n3359), .ZN(n3369) );
  AOI22_X1 U4331 ( .A1(n3605), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4332 ( .A1(n3483), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4333 ( .A1(n3478), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4334 ( .A1(n3629), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4335 ( .A1(n4340), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3201), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4336 ( .A1(n3442), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4337 ( .A1(n3463), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4338 ( .A1(n3463), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4340), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4339 ( .A1(n3208), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4340 ( .A1(n4069), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4341 ( .A1(n3478), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3372) );
  NAND4_X1 U4342 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3382)
         );
  AOI22_X1 U4343 ( .A1(n3442), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4344 ( .A1(n3383), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3485), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3377) );
  NAND4_X1 U4345 ( .A1(n3380), .A2(n3379), .A3(n3378), .A4(n3377), .ZN(n3381)
         );
  NAND2_X1 U4346 ( .A1(n3803), .A2(n4588), .ZN(n3394) );
  AND2_X2 U4347 ( .A1(n4999), .A2(n5327), .ZN(n3825) );
  AOI22_X1 U4348 ( .A1(n4340), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3485), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4349 ( .A1(n3442), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4350 ( .A1(n3463), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4351 ( .A1(n3478), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4352 ( .A1(n3629), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4353 ( .A1(n3483), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4354 ( .A1(n3605), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3200), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3388) );
  AND2_X2 U4355 ( .A1(n3394), .A2(n3940), .ZN(n3434) );
  NOR2_X1 U4356 ( .A1(n6544), .A2(n6554), .ZN(n6547) );
  INV_X1 U4357 ( .A(n6547), .ZN(n3395) );
  OAI21_X1 U4358 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n3395), .ZN(n3396) );
  INV_X1 U4359 ( .A(n3396), .ZN(n3810) );
  AOI22_X1 U4360 ( .A1(n3463), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4361 ( .A1(n3442), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3370), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4362 ( .A1(n4069), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4363 ( .A1(n3605), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4364 ( .A1(n3629), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4365 ( .A1(n3478), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4366 ( .A1(n3678), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U4367 ( .A1(n3485), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3401)
         );
  NAND2_X2 U4368 ( .A1(n3218), .A2(n3213), .ZN(n3933) );
  INV_X2 U4369 ( .A(n3933), .ZN(n3438) );
  INV_X1 U4370 ( .A(n3932), .ZN(n3521) );
  NAND2_X1 U4371 ( .A1(n3472), .A2(n3827), .ZN(n4587) );
  OAI211_X1 U4372 ( .C1(n3506), .C2(n5327), .A(n3521), .B(n4587), .ZN(n3407)
         );
  INV_X1 U4373 ( .A(n3407), .ZN(n3422) );
  INV_X1 U4374 ( .A(n4528), .ZN(n3417) );
  NAND2_X1 U4375 ( .A1(n3418), .A2(n3531), .ZN(n3429) );
  NAND2_X1 U4376 ( .A1(n3413), .A2(n3933), .ZN(n3414) );
  OAI211_X2 U4377 ( .C1(n3417), .C2(n3416), .A(n3415), .B(n3414), .ZN(n3502)
         );
  NAND2_X1 U4378 ( .A1(n3502), .A2(n3505), .ZN(n3437) );
  AND2_X2 U4379 ( .A1(n3421), .A2(n3420), .ZN(n3805) );
  NAND4_X1 U4380 ( .A1(n3434), .A2(n3422), .A3(n3437), .A4(n3805), .ZN(n3423)
         );
  NAND2_X1 U4381 ( .A1(n3423), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U4382 ( .A1(n3755), .A2(n4858), .ZN(n3495) );
  MUX2_X1 U4383 ( .A(n3818), .B(n6618), .S(n6902), .Z(n3424) );
  AND2_X1 U4384 ( .A1(n3495), .A2(n3424), .ZN(n3426) );
  INV_X1 U4385 ( .A(n3424), .ZN(n3425) );
  AOI21_X2 U4386 ( .B1(n3496), .B2(n3426), .A(n3225), .ZN(n3515) );
  NOR2_X1 U4387 ( .A1(n3531), .A2(n3933), .ZN(n4527) );
  NAND2_X1 U4388 ( .A1(n3429), .A2(n4588), .ZN(n3431) );
  NAND2_X1 U4389 ( .A1(n5837), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6530) );
  INV_X1 U4390 ( .A(n6530), .ZN(n3430) );
  AOI21_X1 U4391 ( .B1(n4858), .B2(n3801), .A(n4717), .ZN(n3432) );
  NAND2_X1 U4392 ( .A1(n3805), .A2(n3432), .ZN(n3433) );
  NAND2_X1 U4393 ( .A1(n3433), .A2(n3827), .ZN(n3435) );
  AND3_X2 U4394 ( .A1(n3436), .A2(n3435), .A3(n3434), .ZN(n3441) );
  OAI22_X1 U4395 ( .A1(n3825), .A2(n4587), .B1(n6092), .B2(n3438), .ZN(n3439)
         );
  INV_X1 U4396 ( .A(n3439), .ZN(n3440) );
  XNOR2_X2 U4397 ( .A(n3515), .B(n3514), .ZN(n3982) );
  OR2_X2 U4398 ( .A1(n3982), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3530) );
  INV_X2 U4399 ( .A(n3464), .ZN(n4407) );
  AOI22_X1 U4400 ( .A1(n4431), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4401 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n3444), .B1(n4414), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3449) );
  INV_X2 U4402 ( .A(n4343), .ZN(n4415) );
  AOI22_X1 U4403 ( .A1(n4415), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4404 ( .A1(n3629), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3447) );
  NAND4_X1 U4405 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3458)
         );
  INV_X1 U4406 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4437) );
  INV_X1 U4407 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4436) );
  OAI22_X1 U4408 ( .A1(n4437), .A2(n4442), .B1(n4441), .B2(n4436), .ZN(n3451)
         );
  INV_X1 U4409 ( .A(n3451), .ZN(n3456) );
  INV_X1 U4410 ( .A(n3370), .ZN(n3465) );
  INV_X2 U4411 ( .A(n3465), .ZN(n4439) );
  AOI22_X1 U4412 ( .A1(n3561), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4413 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n3605), .B1(n4408), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4414 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n3209), .B1(n4299), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3453) );
  NAND4_X1 U4415 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3457)
         );
  NAND2_X1 U4416 ( .A1(n4999), .A2(n3716), .ZN(n3475) );
  NOR2_X1 U4417 ( .A1(n3475), .A2(n6523), .ZN(n3714) );
  NOR2_X1 U4418 ( .A1(n3597), .A2(n3716), .ZN(n3492) );
  AOI22_X1 U4419 ( .A1(n3605), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4420 ( .A1(n3208), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4421 ( .A1(n3629), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4422 ( .A1(n4415), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3459) );
  NAND4_X1 U4423 ( .A1(n3462), .A2(n3461), .A3(n3460), .A4(n3459), .ZN(n3471)
         );
  AOI22_X1 U4424 ( .A1(n4431), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4425 ( .A1(n4413), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4426 ( .A1(n4407), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3467) );
  INV_X1 U4427 ( .A(n3443), .ZN(n4438) );
  AOI22_X1 U4428 ( .A1(n4414), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4429 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3470)
         );
  MUX2_X1 U4430 ( .A(n3714), .B(n3492), .S(n3532), .Z(n3528) );
  NAND2_X1 U4431 ( .A1(n3755), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3474) );
  NAND2_X1 U4432 ( .A1(n3528), .A2(n3526), .ZN(n3477) );
  INV_X1 U4433 ( .A(n3714), .ZN(n3476) );
  NAND2_X2 U4434 ( .A1(n3530), .A2(n3291), .ZN(n3543) );
  AOI22_X1 U4435 ( .A1(n4415), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4436 ( .A1(n4413), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4437 ( .A1(n3206), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4438 ( .A1(n3678), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3479) );
  NAND4_X1 U4439 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3491)
         );
  AOI22_X1 U4440 ( .A1(n4407), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4441 ( .A1(n3605), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4442 ( .A1(n4439), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4443 ( .A1(n4299), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3486) );
  NAND4_X1 U4444 ( .A1(n3489), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(n3490)
         );
  NAND2_X1 U4445 ( .A1(n3755), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3494) );
  INV_X1 U4446 ( .A(n3492), .ZN(n3493) );
  XNOR2_X2 U4447 ( .A(n3543), .B(n3580), .ZN(n3519) );
  NAND2_X1 U4448 ( .A1(n3496), .A2(n3495), .ZN(n3551) );
  NAND2_X1 U4449 ( .A1(n3551), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3509) );
  INV_X1 U4450 ( .A(n6618), .ZN(n3553) );
  XNOR2_X1 U4451 ( .A(n6902), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6347)
         );
  NAND2_X1 U4452 ( .A1(n3553), .A2(n6347), .ZN(n3498) );
  INV_X1 U4453 ( .A(n3818), .ZN(n3552) );
  NAND2_X1 U4454 ( .A1(n3552), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3497) );
  NOR2_X1 U4455 ( .A1(n3932), .A2(n5327), .ZN(n3499) );
  INV_X1 U4456 ( .A(n3820), .ZN(n3501) );
  NAND2_X1 U4457 ( .A1(n3501), .A2(n3834), .ZN(n3507) );
  INV_X1 U4458 ( .A(n3807), .ZN(n3504) );
  AND2_X1 U4459 ( .A1(n3825), .A2(n3505), .ZN(n3503) );
  NAND2_X2 U4460 ( .A1(n3504), .A2(n3503), .ZN(n3829) );
  NAND3_X1 U4461 ( .A1(n3505), .A2(n4993), .A3(n4527), .ZN(n4618) );
  NAND2_X1 U4462 ( .A1(n4857), .A2(n3411), .ZN(n4570) );
  OAI211_X1 U4463 ( .C1(n3507), .C2(n3506), .A(n3829), .B(n3304), .ZN(n3508)
         );
  NAND2_X1 U4464 ( .A1(n3508), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3510) );
  NAND3_X1 U4465 ( .A1(n3509), .A2(n3511), .A3(n3510), .ZN(n3547) );
  INV_X1 U4466 ( .A(n3510), .ZN(n3513) );
  INV_X1 U4467 ( .A(n3511), .ZN(n3512) );
  NAND2_X1 U4468 ( .A1(n3513), .A2(n3300), .ZN(n3549) );
  NAND2_X1 U4469 ( .A1(n3547), .A2(n3549), .ZN(n3516) );
  AND2_X2 U4470 ( .A1(n3515), .A2(n3514), .ZN(n3548) );
  XNOR2_X1 U4471 ( .A(n3516), .B(n3548), .ZN(n4720) );
  NAND2_X1 U4472 ( .A1(n4720), .A2(n6523), .ZN(n3518) );
  NAND2_X2 U4473 ( .A1(n3518), .A2(n3290), .ZN(n3542) );
  NAND2_X1 U4474 ( .A1(n4716), .A2(n3786), .ZN(n3525) );
  NAND2_X1 U4475 ( .A1(n3520), .A2(n3532), .ZN(n3585) );
  OAI21_X1 U4476 ( .B1(n3520), .B2(n3532), .A(n3585), .ZN(n3522) );
  OAI211_X1 U4477 ( .C1(n3522), .C2(n6623), .A(n3521), .B(n5327), .ZN(n3523)
         );
  INV_X1 U4478 ( .A(n3523), .ZN(n3524) );
  NAND2_X1 U4479 ( .A1(n3525), .A2(n3524), .ZN(n6196) );
  INV_X1 U4480 ( .A(n3526), .ZN(n3527) );
  XNOR2_X1 U4481 ( .A(n3528), .B(n3527), .ZN(n3529) );
  INV_X1 U4482 ( .A(n3786), .ZN(n3648) );
  OR2_X2 U4483 ( .A1(n6308), .A2(n3648), .ZN(n3535) );
  NAND2_X1 U4484 ( .A1(n6092), .A2(n3531), .ZN(n3587) );
  OAI21_X1 U4485 ( .B1(n6623), .B2(n3532), .A(n3587), .ZN(n3533) );
  INV_X1 U4486 ( .A(n3533), .ZN(n3534) );
  NAND2_X1 U4487 ( .A1(n3535), .A2(n3534), .ZN(n4634) );
  NAND2_X1 U4488 ( .A1(n4634), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3537)
         );
  INV_X1 U4489 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3536) );
  NAND2_X1 U4490 ( .A1(n3537), .A2(n3536), .ZN(n3539) );
  NAND2_X1 U4491 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6240) );
  INV_X1 U4492 ( .A(n6240), .ZN(n3538) );
  NAND2_X1 U4493 ( .A1(n4634), .A2(n3538), .ZN(n3540) );
  INV_X1 U4494 ( .A(n3580), .ZN(n3541) );
  NAND2_X1 U4495 ( .A1(n3579), .A2(n3541), .ZN(n3546) );
  INV_X1 U4496 ( .A(n3542), .ZN(n3545) );
  NAND2_X1 U4497 ( .A1(n3545), .A2(n3544), .ZN(n3581) );
  AND2_X2 U4498 ( .A1(n3546), .A2(n3581), .ZN(n3577) );
  NAND2_X1 U4499 ( .A1(n3548), .A2(n3547), .ZN(n3550) );
  NAND2_X1 U4500 ( .A1(n3550), .A2(n3549), .ZN(n3559) );
  INV_X1 U4501 ( .A(n3559), .ZN(n3557) );
  NAND2_X1 U4502 ( .A1(n3551), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3555) );
  NAND2_X1 U4503 ( .A1(n6500), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6434) );
  NOR2_X1 U4504 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6500), .ZN(n4940)
         );
  NAND2_X1 U4505 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4940), .ZN(n6392) );
  OAI211_X1 U4506 ( .C1(n6506), .C2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n6434), .B(n6392), .ZN(n4762) );
  AOI22_X1 U4507 ( .A1(n3553), .A2(n4762), .B1(n3552), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3554) );
  NAND2_X1 U4508 ( .A1(n3557), .A2(n3556), .ZN(n3560) );
  NAND2_X1 U4509 ( .A1(n3559), .A2(n3558), .ZN(n3593) );
  NAND2_X1 U4510 ( .A1(n3560), .A2(n3593), .ZN(n4616) );
  AOI22_X1 U4511 ( .A1(n4431), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3566) );
  INV_X1 U4512 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4318) );
  INV_X1 U4513 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4317) );
  OAI22_X1 U4514 ( .A1(n4442), .A2(n4318), .B1(n4441), .B2(n4317), .ZN(n3562)
         );
  INV_X1 U4515 ( .A(n3562), .ZN(n3565) );
  AOI22_X1 U4516 ( .A1(n4407), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4517 ( .A1(n4415), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4518 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3572)
         );
  AOI22_X1 U4519 ( .A1(n3484), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4520 ( .A1(n3444), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4521 ( .A1(n3210), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4522 ( .A1(n3206), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4523 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3571)
         );
  OAI22_X2 U4524 ( .A1(n4616), .A2(STATE2_REG_0__SCAN_IN), .B1(n3586), .B2(
        n3597), .ZN(n3576) );
  INV_X1 U4525 ( .A(n3598), .ZN(n3574) );
  AOI22_X1 U4526 ( .A1(n3755), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3574), 
        .B2(n3573), .ZN(n3575) );
  INV_X1 U4527 ( .A(n3578), .ZN(n3583) );
  NAND2_X1 U4528 ( .A1(n3581), .A2(n3580), .ZN(n3582) );
  NAND3_X1 U4529 ( .A1(n3583), .A2(n3579), .A3(n3582), .ZN(n3584) );
  NAND2_X1 U4530 ( .A1(n3614), .A2(n3584), .ZN(n3997) );
  NAND2_X1 U4531 ( .A1(n3585), .A2(n3586), .ZN(n3642) );
  OAI21_X1 U4532 ( .B1(n3586), .B2(n3585), .A(n3642), .ZN(n3589) );
  INV_X1 U4533 ( .A(n3587), .ZN(n3588) );
  AOI21_X1 U4534 ( .B1(n3589), .B2(n4588), .A(n3588), .ZN(n3590) );
  OAI21_X1 U4535 ( .B1(n3997), .B2(n3648), .A(n3590), .ZN(n6185) );
  NAND2_X1 U4536 ( .A1(n6187), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3591)
         );
  NAND2_X1 U4537 ( .A1(n3592), .A2(n3591), .ZN(n4709) );
  NAND2_X1 U4538 ( .A1(n3551), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3596) );
  NAND3_X1 U4539 ( .A1(n4948), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6318) );
  INV_X1 U4540 ( .A(n6318), .ZN(n6316) );
  NAND3_X1 U4541 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4756) );
  INV_X1 U4542 ( .A(n4756), .ZN(n4779) );
  NAND2_X1 U4543 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4779), .ZN(n4771) );
  OAI21_X1 U4544 ( .B1(n6338), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n4771), 
        .ZN(n6346) );
  OAI22_X1 U4545 ( .A1(n6346), .A2(n6618), .B1(n3818), .B2(n4948), .ZN(n3594)
         );
  INV_X1 U4546 ( .A(n3594), .ZN(n3595) );
  INV_X1 U4547 ( .A(n3798), .ZN(n3772) );
  AOI22_X1 U4548 ( .A1(n4431), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3604) );
  INV_X1 U4549 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4344) );
  INV_X1 U4550 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3599) );
  OAI22_X1 U4551 ( .A1(n4344), .A2(n4442), .B1(n4441), .B2(n3599), .ZN(n3600)
         );
  INV_X1 U4552 ( .A(n3600), .ZN(n3603) );
  AOI22_X1 U4553 ( .A1(n4407), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4554 ( .A1(n4415), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3601) );
  NAND4_X1 U4555 ( .A1(n3604), .A2(n3603), .A3(n3602), .A4(n3601), .ZN(n3611)
         );
  AOI22_X1 U4556 ( .A1(n3484), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4557 ( .A1(n3444), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4558 ( .A1(n3209), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4559 ( .A1(n3206), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3606) );
  NAND4_X1 U4560 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(n3610)
         );
  AOI22_X1 U4561 ( .A1(n3772), .A2(n3641), .B1(n3755), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3612) );
  NAND2_X1 U4562 ( .A1(n3614), .A2(n4715), .ZN(n3615) );
  INV_X1 U4563 ( .A(n3641), .ZN(n3616) );
  XNOR2_X1 U4564 ( .A(n3642), .B(n3616), .ZN(n3617) );
  NAND2_X1 U4565 ( .A1(n3617), .A2(n4588), .ZN(n3618) );
  OAI21_X2 U4566 ( .B1(n5577), .B2(n3648), .A(n3618), .ZN(n3619) );
  INV_X1 U4567 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U4568 ( .A1(n4709), .A2(n4708), .ZN(n3621) );
  NAND2_X1 U4569 ( .A1(n3619), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3620)
         );
  AOI22_X1 U4570 ( .A1(n4431), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3628) );
  INV_X1 U4571 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3623) );
  INV_X1 U4572 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3622) );
  OAI22_X1 U4573 ( .A1(n4442), .A2(n3623), .B1(n4441), .B2(n3622), .ZN(n3624)
         );
  INV_X1 U4574 ( .A(n3624), .ZN(n3627) );
  AOI22_X1 U4575 ( .A1(n4407), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4576 ( .A1(n4415), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3625) );
  NAND4_X1 U4577 ( .A1(n3628), .A2(n3627), .A3(n3626), .A4(n3625), .ZN(n3635)
         );
  AOI22_X1 U4578 ( .A1(n3484), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4579 ( .A1(n3444), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4580 ( .A1(n3210), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4581 ( .A1(n3206), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3630) );
  NAND4_X1 U4582 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3634)
         );
  NAND2_X1 U4583 ( .A1(n3755), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3636) );
  INV_X1 U4584 ( .A(n3677), .ZN(n3668) );
  NAND2_X1 U4585 ( .A1(n3639), .A2(n3638), .ZN(n3640) );
  NAND2_X1 U4586 ( .A1(n3668), .A2(n3640), .ZN(n4017) );
  NAND2_X1 U4587 ( .A1(n3642), .A2(n3641), .ZN(n3644) );
  INV_X1 U4588 ( .A(n3644), .ZN(n3646) );
  OR2_X1 U4589 ( .A1(n3644), .A2(n3643), .ZN(n3695) );
  OAI211_X1 U4590 ( .C1(n3646), .C2(n3645), .A(n4588), .B(n3695), .ZN(n3647)
         );
  INV_X1 U4591 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3649) );
  XNOR2_X1 U4592 ( .A(n3650), .B(n3649), .ZN(n4696) );
  NAND2_X1 U4593 ( .A1(n4697), .A2(n4696), .ZN(n3652) );
  NAND2_X1 U4594 ( .A1(n3650), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3651)
         );
  AOI22_X1 U4595 ( .A1(n4431), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3659) );
  INV_X1 U4596 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3654) );
  INV_X1 U4597 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3653) );
  OAI22_X1 U4598 ( .A1(n4442), .A2(n3654), .B1(n4441), .B2(n3653), .ZN(n3655)
         );
  INV_X1 U4599 ( .A(n3655), .ZN(n3658) );
  AOI22_X1 U4600 ( .A1(n4407), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4601 ( .A1(n4415), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3656) );
  NAND4_X1 U4602 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3665)
         );
  AOI22_X1 U4603 ( .A1(n3484), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4604 ( .A1(n3444), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4605 ( .A1(n3209), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4606 ( .A1(n3206), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3660) );
  NAND4_X1 U4607 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3664)
         );
  NAND2_X1 U4608 ( .A1(n3755), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4609 ( .A1(n3667), .A2(n3666), .ZN(n3676) );
  NAND2_X1 U4610 ( .A1(n4018), .A2(n3786), .ZN(n3672) );
  XNOR2_X1 U4611 ( .A(n3695), .B(n3669), .ZN(n3670) );
  NAND2_X1 U4612 ( .A1(n3670), .A2(n4588), .ZN(n3671) );
  NAND2_X1 U4613 ( .A1(n3672), .A2(n3671), .ZN(n3673) );
  INV_X1 U4614 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4849) );
  NAND2_X1 U4615 ( .A1(n4788), .A2(n4789), .ZN(n3675) );
  NAND2_X1 U4616 ( .A1(n3673), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3674)
         );
  AOI22_X1 U4617 ( .A1(n4431), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4618 ( .A1(n3208), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4619 ( .A1(n4415), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4620 ( .A1(n3209), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3679) );
  NAND4_X1 U4621 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n3688)
         );
  AOI22_X1 U4622 ( .A1(n4413), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4623 ( .A1(n3484), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4624 ( .A1(n3444), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4625 ( .A1(n3206), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3683) );
  NAND4_X1 U4626 ( .A1(n3686), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(n3687)
         );
  INV_X1 U4627 ( .A(n3696), .ZN(n3689) );
  NAND2_X1 U4628 ( .A1(n3755), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3690) );
  NAND2_X1 U4629 ( .A1(n3707), .A2(n3786), .ZN(n3715) );
  NOR2_X1 U4630 ( .A1(n3693), .A2(n3692), .ZN(n4025) );
  OR2_X1 U4631 ( .A1(n3715), .A2(n4025), .ZN(n3699) );
  NOR2_X1 U4632 ( .A1(n3695), .A2(n3694), .ZN(n3697) );
  NAND2_X1 U4633 ( .A1(n3697), .A2(n3696), .ZN(n3718) );
  OAI211_X1 U4634 ( .C1(n3697), .C2(n3696), .A(n3718), .B(n4588), .ZN(n3698)
         );
  NAND2_X1 U4635 ( .A1(n3699), .A2(n3698), .ZN(n3701) );
  INV_X1 U4636 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3700) );
  XNOR2_X1 U4637 ( .A(n3701), .B(n3700), .ZN(n4747) );
  NAND2_X1 U4638 ( .A1(n4746), .A2(n4747), .ZN(n3703) );
  NAND2_X1 U4639 ( .A1(n3701), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3702)
         );
  INV_X1 U4640 ( .A(n3716), .ZN(n3705) );
  NAND2_X1 U4641 ( .A1(n3755), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3704) );
  OAI21_X1 U4642 ( .B1(n3798), .B2(n3705), .A(n3704), .ZN(n3706) );
  NAND2_X1 U4643 ( .A1(n4033), .A2(n3786), .ZN(n3710) );
  XNOR2_X1 U4644 ( .A(n3718), .B(n3716), .ZN(n3708) );
  NAND2_X1 U4645 ( .A1(n3708), .A2(n4588), .ZN(n3709) );
  NAND2_X1 U4646 ( .A1(n3710), .A2(n3709), .ZN(n3711) );
  INV_X1 U4647 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6237) );
  XNOR2_X1 U4648 ( .A(n3711), .B(n6237), .ZN(n6171) );
  NAND2_X1 U4649 ( .A1(n6170), .A2(n6171), .ZN(n3713) );
  NAND2_X1 U4650 ( .A1(n3711), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3712)
         );
  NAND2_X1 U4651 ( .A1(n4588), .A2(n3716), .ZN(n3717) );
  OR2_X1 U4652 ( .A1(n3718), .A2(n3717), .ZN(n3719) );
  NAND2_X1 U4653 ( .A1(n3725), .A2(n3719), .ZN(n3720) );
  INV_X1 U4654 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6757) );
  XNOR2_X1 U4655 ( .A(n3720), .B(n6757), .ZN(n5096) );
  NAND2_X1 U4656 ( .A1(n5095), .A2(n5096), .ZN(n3722) );
  NAND2_X1 U4657 ( .A1(n3720), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3721)
         );
  INV_X1 U4658 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6227) );
  NOR2_X1 U4659 ( .A1(n5756), .A2(n6227), .ZN(n3723) );
  NAND2_X1 U4660 ( .A1(n3725), .A2(n6227), .ZN(n3724) );
  INV_X1 U4661 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4662 ( .A1(n5754), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5269) );
  INV_X1 U4663 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U4664 ( .A1(n5756), .A2(n6765), .ZN(n6157) );
  NAND2_X1 U4665 ( .A1(n5754), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6158) );
  INV_X1 U4666 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U4667 ( .A1(n3725), .A2(n6966), .ZN(n3727) );
  NAND2_X1 U4668 ( .A1(n5444), .A2(n3727), .ZN(n3729) );
  NAND2_X1 U4669 ( .A1(n5754), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4670 ( .A1(n3729), .A2(n3728), .ZN(n5439) );
  INV_X1 U4671 ( .A(n5439), .ZN(n3731) );
  INV_X1 U4672 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6752) );
  XNOR2_X1 U4673 ( .A(n5756), .B(n6752), .ZN(n5440) );
  NAND2_X1 U4674 ( .A1(n5756), .A2(n6752), .ZN(n3732) );
  NAND2_X1 U4675 ( .A1(n5754), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3733) );
  INV_X1 U4676 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U4677 ( .A(n5756), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5589)
         );
  NAND2_X2 U4678 ( .A1(n5588), .A2(n5589), .ZN(n5750) );
  INV_X1 U4679 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3950) );
  NAND2_X1 U4680 ( .A1(n3725), .A2(n3950), .ZN(n3734) );
  NAND2_X2 U4681 ( .A1(n5750), .A2(n3734), .ZN(n5765) );
  INV_X1 U4682 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5805) );
  AND2_X1 U4683 ( .A1(n3725), .A2(n5805), .ZN(n3735) );
  NAND2_X1 U4684 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3736) );
  INV_X1 U4685 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U4686 ( .A1(n5805), .A2(n5795), .ZN(n5749) );
  OAI21_X1 U4687 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5749), .A(n5754), 
        .ZN(n3737) );
  NOR2_X1 U4688 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5530) );
  NOR2_X1 U4689 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4548) );
  NOR2_X1 U4690 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5508) );
  AND3_X1 U4691 ( .A1(n5530), .A2(n4548), .A3(n5508), .ZN(n3738) );
  NOR2_X1 U4692 ( .A1(n3725), .A2(n3738), .ZN(n3740) );
  AND2_X1 U4693 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5531) );
  AND2_X1 U4694 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5507) );
  AND2_X1 U4695 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3960) );
  NAND3_X1 U4696 ( .A1(n5531), .A2(n5507), .A3(n3960), .ZN(n3951) );
  NAND2_X1 U4697 ( .A1(n3725), .A2(n3951), .ZN(n3739) );
  XNOR2_X1 U4698 ( .A(n3725), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5726)
         );
  INV_X1 U4699 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5778) );
  AND2_X2 U4700 ( .A1(n3971), .A2(n3293), .ZN(n5479) );
  AND2_X1 U4701 ( .A1(n3725), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5480)
         );
  AND2_X1 U4702 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4463) );
  INV_X1 U4703 ( .A(n4463), .ZN(n5462) );
  NOR2_X2 U4704 ( .A1(n4467), .A2(n5462), .ZN(n5408) );
  NAND2_X1 U4705 ( .A1(n5408), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3744) );
  INV_X1 U4706 ( .A(n5479), .ZN(n3741) );
  NOR2_X1 U4707 ( .A1(n3725), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5481)
         );
  NOR2_X1 U4708 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4465) );
  NAND2_X1 U4709 ( .A1(n3742), .A2(n5461), .ZN(n3743) );
  INV_X1 U4710 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6898) );
  XNOR2_X1 U4711 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U4712 ( .A1(n3764), .A2(n3761), .ZN(n3747) );
  NAND2_X1 U4713 ( .A1(n6500), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4714 ( .A1(n3747), .A2(n3746), .ZN(n3781) );
  XNOR2_X1 U4715 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U4716 ( .A1(n3781), .A2(n3779), .ZN(n3749) );
  NAND2_X1 U4717 ( .A1(n6506), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3748) );
  NOR2_X1 U4718 ( .A1(n6265), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3753)
         );
  NAND3_X1 U4719 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3756), .A3(n5840), .ZN(n3794) );
  XNOR2_X1 U4720 ( .A(n3758), .B(n3757), .ZN(n3785) );
  NAND2_X1 U4721 ( .A1(n3794), .A2(n3785), .ZN(n3815) );
  OR2_X1 U4722 ( .A1(n3798), .A2(n5038), .ZN(n3760) );
  AND2_X1 U4723 ( .A1(n3760), .A2(n5327), .ZN(n3778) );
  INV_X1 U4724 ( .A(n3761), .ZN(n3762) );
  XNOR2_X1 U4725 ( .A(n3762), .B(n3764), .ZN(n3811) );
  NAND2_X1 U4726 ( .A1(n3811), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3777) );
  INV_X1 U4727 ( .A(n3811), .ZN(n3770) );
  AND2_X1 U4728 ( .A1(n5038), .A2(n5327), .ZN(n3763) );
  INV_X1 U4729 ( .A(n3764), .ZN(n3766) );
  NAND2_X1 U4730 ( .A1(n4656), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3765) );
  NAND2_X1 U4731 ( .A1(n3766), .A2(n3765), .ZN(n3771) );
  OAI21_X1 U4732 ( .B1(n3825), .B2(n3771), .A(n3767), .ZN(n3768) );
  AOI22_X1 U4733 ( .A1(n3778), .A2(n3777), .B1(n3783), .B2(n3768), .ZN(n3773)
         );
  INV_X1 U4734 ( .A(n3800), .ZN(n3769) );
  OAI21_X1 U4735 ( .B1(n3770), .B2(n3773), .A(n3769), .ZN(n3776) );
  INV_X1 U4736 ( .A(n3771), .ZN(n3774) );
  NAND3_X1 U4737 ( .A1(n3774), .A2(n3773), .A3(n3772), .ZN(n3775) );
  OAI211_X1 U4738 ( .C1(n3778), .C2(n3777), .A(n3776), .B(n3775), .ZN(n3791)
         );
  INV_X1 U4739 ( .A(n3779), .ZN(n3780) );
  XNOR2_X1 U4740 ( .A(n3781), .B(n3780), .ZN(n3812) );
  INV_X1 U4741 ( .A(n3812), .ZN(n3782) );
  OAI211_X1 U4742 ( .C1(n3812), .C2(n3793), .A(n3783), .B(n3784), .ZN(n3790)
         );
  INV_X1 U4743 ( .A(n3783), .ZN(n3789) );
  INV_X1 U4744 ( .A(n3784), .ZN(n3788) );
  INV_X1 U4745 ( .A(n3785), .ZN(n3787) );
  AOI222_X1 U4746 ( .A1(n3791), .A2(n3790), .B1(n3789), .B2(n3788), .C1(n3787), 
        .C2(n3786), .ZN(n3792) );
  AOI21_X1 U4747 ( .B1(n3793), .B2(n3815), .A(n3792), .ZN(n3796) );
  OAI22_X1 U4748 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5840), .B1(n3794), .B2(
        n3800), .ZN(n3795) );
  NAND2_X1 U4749 ( .A1(n4857), .A2(n3801), .ZN(n3802) );
  INV_X1 U4750 ( .A(n4173), .ZN(n5336) );
  NAND2_X1 U4751 ( .A1(n5336), .A2(n3827), .ZN(n3942) );
  NAND2_X1 U4752 ( .A1(n3803), .A2(n3834), .ZN(n3804) );
  MUX2_X1 U4753 ( .A(n6623), .B(n3804), .S(n4858), .Z(n3939) );
  AOI21_X1 U4754 ( .B1(n4173), .B2(n6092), .A(n3932), .ZN(n3806) );
  NAND2_X1 U4755 ( .A1(n3939), .A2(n3826), .ZN(n3809) );
  NAND2_X1 U4756 ( .A1(n3825), .A2(n6092), .ZN(n3808) );
  NAND2_X1 U4757 ( .A1(n3809), .A2(n4580), .ZN(n4610) );
  INV_X1 U4758 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U4759 ( .A1(n3810), .A2(n6545), .ZN(n6543) );
  NAND2_X1 U4760 ( .A1(n3827), .A2(n6543), .ZN(n3816) );
  NAND2_X1 U4761 ( .A1(n3812), .A2(n3811), .ZN(n3814) );
  OAI21_X1 U4762 ( .B1(n3815), .B2(n3814), .A(n3813), .ZN(n4578) );
  NOR2_X1 U4763 ( .A1(READY_N), .A2(n4578), .ZN(n4561) );
  NAND3_X1 U4764 ( .A1(n3816), .A2(n4561), .A3(n3933), .ZN(n3817) );
  OAI211_X1 U4765 ( .C1(n4606), .C2(n3942), .A(n4610), .B(n3817), .ZN(n3819)
         );
  NAND2_X1 U4766 ( .A1(n3819), .A2(n4565), .ZN(n3824) );
  INV_X1 U4767 ( .A(READY_N), .ZN(n3821) );
  OAI21_X1 U4768 ( .B1(n3827), .B2(n5596), .A(n3821), .ZN(n4605) );
  OAI211_X1 U4769 ( .C1(n4619), .C2(n4605), .A(n3834), .B(n4570), .ZN(n3822)
         );
  NAND3_X1 U4770 ( .A1(n5597), .A2(n3438), .A3(n3822), .ZN(n3823) );
  AND2_X1 U4771 ( .A1(n3826), .A2(n3825), .ZN(n4577) );
  INV_X1 U4772 ( .A(n4577), .ZN(n6511) );
  INV_X1 U4773 ( .A(n4622), .ZN(n3831) );
  OAI22_X1 U4774 ( .A1(n4619), .A2(n6075), .B1(n4999), .B2(n3304), .ZN(n3828)
         );
  INV_X1 U4775 ( .A(n3828), .ZN(n3830) );
  NAND4_X1 U4776 ( .A1(n6511), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3832)
         );
  MUX2_X1 U4777 ( .A(n3917), .B(n3916), .S(EBX_REG_1__SCAN_IN), .Z(n3837) );
  INV_X1 U4778 ( .A(n3916), .ZN(n3835) );
  NAND2_X1 U4779 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3836)
         );
  INV_X1 U4780 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U4781 ( .A1(n5526), .A2(n6082), .ZN(n3839) );
  NAND2_X1 U4782 ( .A1(n3916), .A2(EBX_REG_0__SCAN_IN), .ZN(n3838) );
  AND2_X1 U4783 ( .A1(n3839), .A2(n3838), .ZN(n4647) );
  NAND2_X1 U4784 ( .A1(n3840), .A2(n4530), .ZN(n6078) );
  NAND2_X1 U4785 ( .A1(n6078), .A2(n3841), .ZN(n5301) );
  MUX2_X1 U4786 ( .A(n4512), .B(n3204), .S(EBX_REG_3__SCAN_IN), .Z(n3843) );
  NOR2_X1 U4787 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3842)
         );
  NOR2_X1 U4788 ( .A1(n3843), .A2(n3842), .ZN(n4881) );
  INV_X1 U4789 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3844) );
  NAND2_X1 U4790 ( .A1(n3916), .A2(n3844), .ZN(n3846) );
  INV_X1 U4791 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U4792 ( .A1(n4530), .A2(n6074), .ZN(n3845) );
  NAND3_X1 U4793 ( .A1(n3846), .A2(n5526), .A3(n3845), .ZN(n3847) );
  OAI21_X1 U4794 ( .B1(n3917), .B2(EBX_REG_2__SCAN_IN), .A(n3847), .ZN(n5300)
         );
  NAND2_X1 U4795 ( .A1(n4881), .A2(n5300), .ZN(n3848) );
  MUX2_X1 U4796 ( .A(n3917), .B(n3916), .S(EBX_REG_4__SCAN_IN), .Z(n3850) );
  NAND2_X1 U4797 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3849)
         );
  AND3_X1 U4798 ( .A1(n3850), .A2(n3908), .A3(n3849), .ZN(n5213) );
  MUX2_X1 U4799 ( .A(n4512), .B(n3204), .S(EBX_REG_5__SCAN_IN), .Z(n3852) );
  NOR2_X1 U4800 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3851)
         );
  NOR2_X1 U4801 ( .A1(n3852), .A2(n3851), .ZN(n4796) );
  MUX2_X1 U4802 ( .A(n3917), .B(n3916), .S(EBX_REG_6__SCAN_IN), .Z(n3854) );
  NAND2_X1 U4803 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6075), .ZN(n3853)
         );
  INV_X1 U4804 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U4805 ( .A1(n4512), .A2(n6058), .ZN(n3857) );
  NAND2_X1 U4806 ( .A1(n4530), .A2(n6058), .ZN(n3855) );
  OAI211_X1 U4807 ( .C1(n3204), .C2(n6237), .A(n3855), .B(n3916), .ZN(n3856)
         );
  NAND2_X1 U4808 ( .A1(n3857), .A2(n3856), .ZN(n5960) );
  MUX2_X1 U4809 ( .A(n3917), .B(n3916), .S(EBX_REG_8__SCAN_IN), .Z(n3859) );
  NAND2_X1 U4810 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3858)
         );
  INV_X1 U4811 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U4812 ( .A1(n4512), .A2(n6053), .ZN(n3862) );
  NAND2_X1 U4813 ( .A1(n4530), .A2(n6053), .ZN(n3860) );
  OAI211_X1 U4814 ( .C1(n3204), .C2(n6227), .A(n3860), .B(n3916), .ZN(n3861)
         );
  AND2_X1 U4815 ( .A1(n3862), .A2(n3861), .ZN(n5943) );
  INV_X1 U4816 ( .A(n3917), .ZN(n3886) );
  INV_X1 U4817 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U4818 ( .A1(n3886), .A2(n6050), .ZN(n3866) );
  NAND2_X1 U4819 ( .A1(n3916), .A2(n3863), .ZN(n3864) );
  OAI211_X1 U4820 ( .C1(n6075), .C2(EBX_REG_10__SCAN_IN), .A(n3864), .B(n5526), 
        .ZN(n3865) );
  INV_X1 U4821 ( .A(n4512), .ZN(n3910) );
  MUX2_X1 U4822 ( .A(n3910), .B(n5526), .S(EBX_REG_11__SCAN_IN), .Z(n3867) );
  NAND2_X1 U4823 ( .A1(n3299), .A2(n3867), .ZN(n5925) );
  MUX2_X1 U4824 ( .A(n3917), .B(n3916), .S(EBX_REG_12__SCAN_IN), .Z(n3869) );
  NAND2_X1 U4825 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6075), .ZN(n3868) );
  INV_X1 U4826 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U4827 ( .A1(n4512), .A2(n6043), .ZN(n3872) );
  NAND2_X1 U4828 ( .A1(n4530), .A2(n6043), .ZN(n3870) );
  OAI211_X1 U4829 ( .C1(n3204), .C2(n6752), .A(n3870), .B(n3916), .ZN(n3871)
         );
  NAND2_X1 U4830 ( .A1(n3872), .A2(n3871), .ZN(n5821) );
  MUX2_X1 U4831 ( .A(n3917), .B(n3916), .S(EBX_REG_14__SCAN_IN), .Z(n3875) );
  NAND2_X1 U4832 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3873) );
  AND2_X1 U4833 ( .A1(n3908), .A2(n3873), .ZN(n3874) );
  NAND2_X1 U4834 ( .A1(n3875), .A2(n3874), .ZN(n5568) );
  INV_X1 U4835 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U4836 ( .A1(n4512), .A2(n6037), .ZN(n3878) );
  NAND2_X1 U4837 ( .A1(n4530), .A2(n6037), .ZN(n3876) );
  OAI211_X1 U4838 ( .C1(n3204), .C2(n3950), .A(n3876), .B(n3916), .ZN(n3877)
         );
  NAND2_X1 U4839 ( .A1(n3878), .A2(n3877), .ZN(n5814) );
  MUX2_X1 U4840 ( .A(n3917), .B(n3916), .S(EBX_REG_16__SCAN_IN), .Z(n3881) );
  NAND2_X1 U4841 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6075), .ZN(n3879) );
  AND2_X1 U4842 ( .A1(n3908), .A2(n3879), .ZN(n3880) );
  NAND2_X1 U4843 ( .A1(n3881), .A2(n3880), .ZN(n5799) );
  INV_X1 U4844 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U4845 ( .A1(n4512), .A2(n6031), .ZN(n3884) );
  NAND2_X1 U4846 ( .A1(n4530), .A2(n6031), .ZN(n3882) );
  OAI211_X1 U4847 ( .C1(n3204), .C2(n5795), .A(n3882), .B(n3916), .ZN(n3883)
         );
  AND2_X1 U4848 ( .A1(n3884), .A2(n3883), .ZN(n5789) );
  NAND2_X1 U4849 ( .A1(n5799), .A2(n5789), .ZN(n3885) );
  INV_X1 U4850 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U4851 ( .A1(n3886), .A2(n5712), .ZN(n3889) );
  INV_X1 U4852 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U4853 ( .A1(n3916), .A2(n5541), .ZN(n3887) );
  OAI211_X1 U4854 ( .C1(n6075), .C2(EBX_REG_19__SCAN_IN), .A(n3887), .B(n5526), 
        .ZN(n3888) );
  NAND2_X1 U4855 ( .A1(n3889), .A2(n3888), .ZN(n5547) );
  OR2_X1 U4856 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3892)
         );
  INV_X1 U4857 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4858 ( .A1(n4530), .A2(n3890), .ZN(n3891) );
  AND2_X1 U4859 ( .A1(n3892), .A2(n3891), .ZN(n5527) );
  OR2_X1 U4860 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3894)
         );
  INV_X1 U4861 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3893) );
  NAND2_X1 U4862 ( .A1(n4530), .A2(n3893), .ZN(n5545) );
  NAND2_X1 U4863 ( .A1(n3894), .A2(n5545), .ZN(n5546) );
  NAND2_X1 U4864 ( .A1(n3204), .A2(EBX_REG_20__SCAN_IN), .ZN(n3896) );
  NAND2_X1 U4865 ( .A1(n5546), .A2(n5526), .ZN(n3895) );
  OAI211_X1 U4866 ( .C1(n5527), .C2(n5546), .A(n3896), .B(n3895), .ZN(n3897)
         );
  INV_X1 U4867 ( .A(n3897), .ZN(n3898) );
  INV_X1 U4868 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U4869 ( .A1(n4512), .A2(n5707), .ZN(n3902) );
  INV_X1 U4870 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3900) );
  NAND2_X1 U4871 ( .A1(n4530), .A2(n5707), .ZN(n3899) );
  OAI211_X1 U4872 ( .C1(n3204), .C2(n3900), .A(n3899), .B(n3916), .ZN(n3901)
         );
  NAND2_X1 U4873 ( .A1(n3902), .A2(n3901), .ZN(n5516) );
  MUX2_X1 U4874 ( .A(n3917), .B(n3916), .S(EBX_REG_22__SCAN_IN), .Z(n3904) );
  NAND2_X1 U4875 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3903) );
  MUX2_X1 U4876 ( .A(n4512), .B(n3204), .S(EBX_REG_23__SCAN_IN), .Z(n3906) );
  NOR2_X1 U4877 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3905)
         );
  MUX2_X1 U4878 ( .A(n3917), .B(n3916), .S(EBX_REG_24__SCAN_IN), .Z(n3909) );
  NAND2_X1 U4879 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3907) );
  AND3_X1 U4880 ( .A1(n3909), .A2(n3908), .A3(n3907), .ZN(n4544) );
  MUX2_X1 U4881 ( .A(n3910), .B(n5526), .S(EBX_REG_25__SCAN_IN), .Z(n3911) );
  NAND2_X1 U4882 ( .A1(n3295), .A2(n3911), .ZN(n5637) );
  NAND2_X1 U4883 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3913) );
  MUX2_X1 U4884 ( .A(n3917), .B(n3916), .S(EBX_REG_26__SCAN_IN), .Z(n3912) );
  AND2_X1 U4885 ( .A1(n3913), .A2(n3912), .ZN(n5485) );
  MUX2_X1 U4886 ( .A(n4512), .B(n3204), .S(EBX_REG_27__SCAN_IN), .Z(n3915) );
  NOR2_X1 U4887 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3914)
         );
  NOR2_X1 U4888 ( .A1(n3915), .A2(n3914), .ZN(n5471) );
  MUX2_X1 U4889 ( .A(n3917), .B(n3916), .S(EBX_REG_28__SCAN_IN), .Z(n3919) );
  NAND2_X1 U4890 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3918) );
  NAND2_X1 U4891 ( .A1(n3919), .A2(n3918), .ZN(n3974) );
  OR2_X1 U4892 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4511)
         );
  OAI21_X1 U4893 ( .B1(EBX_REG_29__SCAN_IN), .B2(n6075), .A(n4511), .ZN(n3920)
         );
  NOR2_X1 U4894 ( .A1(n4536), .A2(n3920), .ZN(n3925) );
  INV_X1 U4895 ( .A(n3925), .ZN(n3924) );
  INV_X1 U4896 ( .A(n4536), .ZN(n3923) );
  NAND2_X1 U4897 ( .A1(n4645), .A2(EBX_REG_30__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4898 ( .A1(n6075), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3921) );
  NAND2_X1 U4899 ( .A1(n3922), .A2(n3921), .ZN(n3926) );
  INV_X1 U4900 ( .A(n3926), .ZN(n4516) );
  AOI21_X1 U4901 ( .B1(n3924), .B2(n3923), .A(n4516), .ZN(n3928) );
  NAND2_X1 U4902 ( .A1(n3924), .A2(n5526), .ZN(n4517) );
  AOI211_X1 U4903 ( .C1(n3204), .C2(n4536), .A(n3926), .B(n3925), .ZN(n3927)
         );
  AOI21_X1 U4904 ( .B1(n3928), .B2(n4517), .A(n3927), .ZN(n5687) );
  INV_X1 U4905 ( .A(n3304), .ZN(n3929) );
  NAND2_X1 U4906 ( .A1(n3929), .A2(n4999), .ZN(n3930) );
  AND2_X1 U4907 ( .A1(n6519), .A2(n3930), .ZN(n3931) );
  NOR2_X2 U4908 ( .A1(n3954), .A2(n3931), .ZN(n6245) );
  INV_X2 U4909 ( .A(n6256), .ZN(n6221) );
  NAND2_X1 U4910 ( .A1(n6221), .A2(REIP_REG_30__SCAN_IN), .ZN(n4553) );
  INV_X1 U4911 ( .A(n4553), .ZN(n3953) );
  NAND2_X1 U4912 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U4913 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5273) );
  NOR2_X1 U4914 ( .A1(n5272), .A2(n5273), .ZN(n3946) );
  INV_X1 U4915 ( .A(n3946), .ZN(n3944) );
  NOR2_X1 U4916 ( .A1(n4587), .A2(n3933), .ZN(n4602) );
  OAI21_X1 U4917 ( .B1(n4602), .B2(n4645), .A(n3932), .ZN(n3935) );
  NAND2_X1 U4918 ( .A1(n4570), .A2(n3933), .ZN(n3934) );
  OAI211_X1 U4919 ( .C1(n3805), .C2(n5526), .A(n3935), .B(n3934), .ZN(n3936)
         );
  INV_X1 U4920 ( .A(n3936), .ZN(n3937) );
  NAND3_X1 U4921 ( .A1(n3939), .A2(n3938), .A3(n3937), .ZN(n4621) );
  OAI21_X1 U4922 ( .B1(n3940), .B2(n3834), .A(n4909), .ZN(n3941) );
  INV_X1 U4923 ( .A(n3942), .ZN(n3943) );
  NAND2_X1 U4924 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5220) );
  INV_X1 U4925 ( .A(n5220), .ZN(n3945) );
  NAND2_X1 U4926 ( .A1(n3844), .A2(n6240), .ZN(n6239) );
  NAND2_X1 U4927 ( .A1(n3945), .A2(n6239), .ZN(n4848) );
  NAND3_X1 U4928 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4794), .ZN(n5098) );
  NAND3_X1 U4929 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n3945), .ZN(n5103) );
  NOR3_X1 U4930 ( .A1(n3844), .A2(n3536), .A3(n5103), .ZN(n5097) );
  NAND2_X1 U4931 ( .A1(n5097), .A2(n3946), .ZN(n5825) );
  NAND2_X1 U4932 ( .A1(n3949), .A2(n5594), .ZN(n5559) );
  INV_X1 U4933 ( .A(n3947), .ZN(n3948) );
  NAND2_X1 U4934 ( .A1(n3949), .A2(n3948), .ZN(n5563) );
  NAND2_X1 U4935 ( .A1(n5559), .A2(n5563), .ZN(n5558) );
  INV_X1 U4936 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U4937 ( .A1(n5559), .A2(n5562), .ZN(n6254) );
  NAND2_X1 U4938 ( .A1(n5558), .A2(n6254), .ZN(n4793) );
  NAND2_X1 U4939 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6204) );
  NOR2_X1 U4940 ( .A1(n6752), .A2(n6204), .ZN(n5566) );
  NAND2_X1 U4941 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5566), .ZN(n5802) );
  NOR2_X1 U4942 ( .A1(n3950), .A2(n5802), .ZN(n5806) );
  NAND2_X1 U4943 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5806), .ZN(n3955) );
  NOR2_X1 U4944 ( .A1(n5801), .A2(n3955), .ZN(n5796) );
  NAND3_X1 U4945 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5796), .ZN(n5543) );
  NOR2_X1 U4946 ( .A1(n5543), .A2(n3951), .ZN(n5773) );
  AND2_X1 U4947 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U4948 ( .A1(n5773), .A2(n5483), .ZN(n5463) );
  INV_X1 U4949 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5461) );
  NOR4_X1 U4950 ( .A1(n5463), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5462), 
        .A4(n5461), .ZN(n3952) );
  AOI211_X1 U4951 ( .C1(n5687), .C2(n6245), .A(n3953), .B(n3952), .ZN(n3968)
         );
  NAND2_X1 U4952 ( .A1(n6243), .A2(n5563), .ZN(n5561) );
  INV_X1 U4953 ( .A(n5559), .ZN(n5828) );
  OAI21_X1 U4954 ( .B1(n5825), .B2(n3955), .A(n5558), .ZN(n5535) );
  AND2_X1 U4955 ( .A1(n6256), .A2(n3954), .ZN(n4651) );
  AND2_X1 U4956 ( .A1(n5562), .A2(n5561), .ZN(n4648) );
  NOR2_X1 U4957 ( .A1(n4651), .A2(n4648), .ZN(n6262) );
  NAND2_X1 U4958 ( .A1(n6262), .A2(n6243), .ZN(n5557) );
  NAND3_X1 U4959 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5531), .ZN(n3956) );
  INV_X1 U4960 ( .A(n5565), .ZN(n5556) );
  OR2_X1 U4961 ( .A1(n3955), .A2(n5556), .ZN(n5534) );
  AOI222_X1 U4962 ( .A1(n5557), .A2(n3956), .B1(n5557), .B2(n5534), .C1(n3956), 
        .C2(n5558), .ZN(n3957) );
  NAND2_X1 U4963 ( .A1(n5535), .A2(n3957), .ZN(n5523) );
  INV_X1 U4964 ( .A(n5507), .ZN(n3958) );
  AND2_X1 U4965 ( .A1(n6255), .A2(n3958), .ZN(n3959) );
  NOR2_X1 U4966 ( .A1(n5523), .A2(n3959), .ZN(n5493) );
  NAND2_X1 U4967 ( .A1(n4793), .A2(n6243), .ZN(n3962) );
  INV_X1 U4968 ( .A(n3960), .ZN(n3961) );
  NAND2_X1 U4969 ( .A1(n3962), .A2(n3961), .ZN(n3963) );
  INV_X1 U4970 ( .A(n5779), .ZN(n3966) );
  INV_X1 U4971 ( .A(n5483), .ZN(n3964) );
  NAND2_X1 U4972 ( .A1(n6255), .A2(n3964), .ZN(n3965) );
  OAI211_X1 U4973 ( .C1(n4463), .C2(n5804), .A(n5454), .B(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5465) );
  OAI211_X1 U4974 ( .C1(n6255), .C2(n3966), .A(n5465), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3967) );
  AND2_X1 U4975 ( .A1(n3968), .A2(n3967), .ZN(n3969) );
  NAND2_X1 U4976 ( .A1(n3970), .A2(n3969), .ZN(U2988) );
  INV_X1 U4977 ( .A(n4467), .ZN(n5416) );
  INV_X1 U4978 ( .A(n4464), .ZN(n5724) );
  NOR3_X1 U4979 ( .A1(n5724), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n3725), 
        .ZN(n3972) );
  INV_X1 U4980 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5492) );
  OAI22_X1 U4981 ( .A1(n5416), .A2(n3972), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5492), .ZN(n3973) );
  XNOR2_X1 U4982 ( .A(n3973), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3981)
         );
  NAND2_X1 U4983 ( .A1(n3981), .A2(n3833), .ZN(n3980) );
  INV_X1 U4984 ( .A(n5454), .ZN(n5475) );
  OR2_X1 U4985 ( .A1(n5469), .A2(n3974), .ZN(n3975) );
  NAND2_X1 U4986 ( .A1(n4536), .A2(n3975), .ZN(n5690) );
  NOR3_X1 U4987 ( .A1(n4463), .A2(n4465), .A3(n5463), .ZN(n3976) );
  AOI21_X1 U4988 ( .B1(n6221), .B2(REIP_REG_28__SCAN_IN), .A(n3976), .ZN(n3977) );
  OAI21_X1 U4989 ( .B1(n5690), .B2(n6258), .A(n3977), .ZN(n3978) );
  AOI21_X1 U4990 ( .B1(n5475), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n3978), 
        .ZN(n3979) );
  NAND2_X1 U4991 ( .A1(n3980), .A2(n3979), .ZN(U2990) );
  OR2_X1 U4992 ( .A1(n3982), .A2(n4160), .ZN(n3987) );
  INV_X1 U4993 ( .A(n4570), .ZN(n3983) );
  NAND2_X1 U4994 ( .A1(n3983), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4007) );
  INV_X1 U4995 ( .A(n4007), .ZN(n4010) );
  INV_X1 U4996 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4640) );
  INV_X2 U4997 ( .A(n3298), .ZN(n4306) );
  NAND2_X1 U4998 ( .A1(n4306), .A2(EAX_REG_0__SCAN_IN), .ZN(n3984) );
  OAI21_X1 U4999 ( .B1(n4640), .B2(STATE2_REG_2__SCAN_IN), .A(n3984), .ZN(
        n3985) );
  AOI21_X1 U5000 ( .B1(n4010), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n3985), 
        .ZN(n3986) );
  NAND2_X1 U5001 ( .A1(n6308), .A2(n4988), .ZN(n3988) );
  NAND2_X1 U5002 ( .A1(n3988), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4636) );
  NAND2_X1 U5003 ( .A1(n4635), .A2(n4458), .ZN(n3989) );
  NAND2_X1 U5004 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6403), .ZN(n3991)
         );
  NAND2_X1 U5005 ( .A1(n4306), .A2(EAX_REG_1__SCAN_IN), .ZN(n3990) );
  OAI211_X1 U5006 ( .C1(n4007), .C2(n6818), .A(n3991), .B(n3990), .ZN(n3992)
         );
  INV_X1 U5007 ( .A(n3992), .ZN(n3993) );
  NAND2_X1 U5008 ( .A1(n3994), .A2(n3993), .ZN(n5144) );
  NAND2_X1 U5009 ( .A1(n5143), .A2(n5144), .ZN(n5146) );
  NOR2_X2 U5010 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4392), .ZN(n4459) );
  AOI22_X1 U5011 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_2__SCAN_IN), .ZN(n3996) );
  OAI21_X1 U5012 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4003), .ZN(n6192) );
  AOI22_X1 U5013 ( .A1(n4010), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(n4458), .B2(n6192), .ZN(n3995) );
  AND2_X1 U5014 ( .A1(n3996), .A2(n3995), .ZN(n3998) );
  INV_X1 U5015 ( .A(n4459), .ZN(n4112) );
  OAI21_X2 U5016 ( .B1(n3997), .B2(n4160), .A(n4112), .ZN(n5151) );
  NAND2_X1 U5017 ( .A1(n5150), .A2(n5151), .ZN(n4002) );
  INV_X1 U5018 ( .A(n5146), .ZN(n4000) );
  INV_X1 U5019 ( .A(n3998), .ZN(n3999) );
  NAND2_X1 U5020 ( .A1(n4000), .A2(n3999), .ZN(n4001) );
  AOI21_X1 U5021 ( .B1(n4003), .B2(n6011), .A(n4013), .ZN(n4004) );
  INV_X1 U5022 ( .A(n4004), .ZN(n6016) );
  AOI22_X1 U5023 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4459), .B1(n4458), 
        .B2(n6016), .ZN(n4006) );
  NAND2_X1 U5024 ( .A1(n4306), .A2(EAX_REG_3__SCAN_IN), .ZN(n4005) );
  OAI211_X1 U5025 ( .C1(n4007), .C2(n3750), .A(n4006), .B(n4005), .ZN(n4008)
         );
  INV_X1 U5026 ( .A(n4008), .ZN(n4009) );
  AND2_X2 U5027 ( .A1(n4710), .A2(n4711), .ZN(n4699) );
  AOI22_X1 U5028 ( .A1(n4306), .A2(EAX_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6403), .ZN(n4012) );
  NAND2_X1 U5029 ( .A1(n4010), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4011) );
  NAND2_X1 U5030 ( .A1(n4012), .A2(n4011), .ZN(n4015) );
  OAI21_X1 U5031 ( .B1(n4013), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4019), 
        .ZN(n6001) );
  AND2_X1 U5032 ( .A1(n6001), .A2(n4458), .ZN(n4014) );
  AOI21_X1 U5033 ( .B1(n4015), .B2(n4493), .A(n4014), .ZN(n4016) );
  NAND2_X1 U5034 ( .A1(n4018), .A2(n4141), .ZN(n4024) );
  AOI22_X1 U5035 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_5__SCAN_IN), .ZN(n4022) );
  OAI21_X1 U5036 ( .B1(n4020), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4027), 
        .ZN(n6178) );
  NAND2_X1 U5037 ( .A1(n4458), .A2(n6178), .ZN(n4021) );
  AND2_X1 U5038 ( .A1(n4022), .A2(n4021), .ZN(n4023) );
  NAND2_X1 U5039 ( .A1(n4024), .A2(n4023), .ZN(n5140) );
  NAND2_X1 U5040 ( .A1(n4700), .A2(n5140), .ZN(n4751) );
  INV_X1 U5041 ( .A(n4025), .ZN(n4026) );
  NAND2_X1 U5042 ( .A1(n4026), .A2(n4141), .ZN(n4032) );
  AOI21_X1 U5043 ( .B1(n6921), .B2(n4027), .A(n4034), .ZN(n5979) );
  INV_X1 U5044 ( .A(n5979), .ZN(n4028) );
  NAND2_X1 U5045 ( .A1(n4458), .A2(n4028), .ZN(n4030) );
  AOI22_X1 U5046 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_6__SCAN_IN), .ZN(n4029) );
  AND2_X1 U5047 ( .A1(n4030), .A2(n4029), .ZN(n4031) );
  NAND2_X1 U5048 ( .A1(n4033), .A2(n4141), .ZN(n4038) );
  NAND2_X1 U5049 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n4459), .ZN(n4036)
         );
  OAI21_X1 U5050 ( .B1(n4034), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4039), 
        .ZN(n6173) );
  AOI22_X1 U5051 ( .A1(n4458), .A2(n6173), .B1(n4306), .B2(EAX_REG_7__SCAN_IN), 
        .ZN(n4035) );
  AND2_X1 U5052 ( .A1(n4036), .A2(n4035), .ZN(n4037) );
  AOI21_X1 U5053 ( .B1(n5952), .B2(n4039), .A(n4066), .ZN(n5957) );
  AOI22_X1 U5054 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_8__SCAN_IN), .ZN(n4040) );
  OAI21_X1 U5055 ( .B1(n5957), .B2(n4493), .A(n4040), .ZN(n4053) );
  AOI22_X1 U5056 ( .A1(n3561), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5057 ( .A1(n3678), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5058 ( .A1(n3484), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5059 ( .A1(n3206), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U5060 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4050)
         );
  AOI22_X1 U5061 ( .A1(n4431), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5062 ( .A1(n4413), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5063 ( .A1(n3210), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5064 ( .A1(n4415), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U5065 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4049)
         );
  NOR2_X1 U5066 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  NOR2_X1 U5067 ( .A1(n4160), .A2(n4051), .ZN(n4052) );
  NOR2_X1 U5068 ( .A1(n4053), .A2(n4052), .ZN(n5133) );
  XOR2_X1 U5069 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4066), .Z(n6166) );
  AOI22_X1 U5070 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_9__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5071 ( .A1(n4407), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5072 ( .A1(n3484), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5073 ( .A1(n4413), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5074 ( .A1(n4415), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4054) );
  NAND4_X1 U5075 ( .A1(n4057), .A2(n4056), .A3(n4055), .A4(n4054), .ZN(n4063)
         );
  AOI22_X1 U5076 ( .A1(n4431), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5077 ( .A1(n3208), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5078 ( .A1(n3209), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5079 ( .A1(n3206), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5080 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4062)
         );
  OAI21_X1 U5081 ( .B1(n4063), .B2(n4062), .A(n4141), .ZN(n4064) );
  OAI211_X1 U5082 ( .C1(n6166), .C2(n4493), .A(n4065), .B(n4064), .ZN(n5115)
         );
  AOI21_X1 U5083 ( .B1(n6771), .B2(n4067), .A(n4095), .ZN(n5936) );
  AOI22_X1 U5084 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_10__SCAN_IN), .ZN(n4068) );
  OAI21_X1 U5085 ( .B1(n5936), .B2(n4493), .A(n4068), .ZN(n4082) );
  AOI22_X1 U5086 ( .A1(n4415), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5087 ( .A1(n4413), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5088 ( .A1(n3678), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5089 ( .A1(n3484), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4070) );
  NAND4_X1 U5090 ( .A1(n4073), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4079)
         );
  AOI22_X1 U5091 ( .A1(n3444), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5092 ( .A1(n3209), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5093 ( .A1(n4431), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5094 ( .A1(n3206), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4074) );
  NAND4_X1 U5095 ( .A1(n4077), .A2(n4076), .A3(n4075), .A4(n4074), .ZN(n4078)
         );
  NOR2_X1 U5096 ( .A1(n4079), .A2(n4078), .ZN(n4080) );
  NOR2_X1 U5097 ( .A1(n4160), .A2(n4080), .ZN(n4081) );
  NOR2_X1 U5098 ( .A1(n4082), .A2(n4081), .ZN(n5248) );
  NOR2_X2 U5099 ( .A1(n5113), .A2(n5248), .ZN(n5249) );
  INV_X1 U5100 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5927) );
  XNOR2_X1 U5101 ( .A(n5927), .B(n4095), .ZN(n6160) );
  AOI22_X1 U5102 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_11__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5103 ( .A1(n4413), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5104 ( .A1(n4415), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5105 ( .A1(n4414), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5106 ( .A1(n3484), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4083) );
  NAND4_X1 U5107 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(n4092)
         );
  AOI22_X1 U5108 ( .A1(n3208), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5109 ( .A1(n3444), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5110 ( .A1(n3561), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5111 ( .A1(n3206), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4087) );
  NAND4_X1 U5112 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(n4091)
         );
  OAI21_X1 U5113 ( .B1(n4092), .B2(n4091), .A(n4141), .ZN(n4093) );
  OAI211_X1 U5114 ( .C1(n6160), .C2(n4493), .A(n4094), .B(n4093), .ZN(n5266)
         );
  NAND2_X1 U5115 ( .A1(n5249), .A2(n5266), .ZN(n5265) );
  AOI21_X1 U5116 ( .B1(n5916), .B2(n4096), .A(n4132), .ZN(n5918) );
  NAND2_X1 U5117 ( .A1(n4306), .A2(EAX_REG_12__SCAN_IN), .ZN(n4098) );
  OAI21_X1 U5118 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n4392), .A(n6403), 
        .ZN(n4097) );
  AOI22_X1 U5119 ( .A1(n4458), .A2(n5918), .B1(n4098), .B2(n4097), .ZN(n4111)
         );
  AOI22_X1 U5120 ( .A1(n4415), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5121 ( .A1(n3206), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5122 ( .A1(n4431), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5123 ( .A1(n4413), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U5124 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4108)
         );
  AOI22_X1 U5125 ( .A1(n3678), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5126 ( .A1(n3209), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5127 ( .A1(n4299), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5128 ( .A1(n4407), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4103) );
  NAND4_X1 U5129 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4107)
         );
  NOR2_X1 U5130 ( .A1(n4108), .A2(n4107), .ZN(n4109) );
  NOR2_X1 U5131 ( .A1(n4160), .A2(n4109), .ZN(n4110) );
  NOR2_X1 U5132 ( .A1(n4111), .A2(n4110), .ZN(n5312) );
  NOR2_X2 U5133 ( .A1(n5265), .A2(n5312), .ZN(n4128) );
  INV_X1 U5134 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6832) );
  INV_X1 U5135 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4113) );
  XNOR2_X1 U5136 ( .A(n4113), .B(n4132), .ZN(n5905) );
  OAI222_X1 U5137 ( .A1(n6832), .A2(n3298), .B1(n4493), .B2(n5905), .C1(n4113), 
        .C2(n4112), .ZN(n4129) );
  XNOR2_X1 U5138 ( .A(n4128), .B(n4114), .ZN(n5323) );
  AOI22_X1 U5139 ( .A1(n4431), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4120) );
  INV_X1 U5140 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4998) );
  INV_X1 U5141 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4115) );
  OAI22_X1 U5142 ( .A1(n4442), .A2(n4998), .B1(n4441), .B2(n4115), .ZN(n4116)
         );
  INV_X1 U5143 ( .A(n4116), .ZN(n4119) );
  AOI22_X1 U5144 ( .A1(n4407), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5145 ( .A1(n4415), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4117) );
  NAND4_X1 U5146 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4126)
         );
  AOI22_X1 U5147 ( .A1(n3484), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5148 ( .A1(n3444), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5149 ( .A1(n3210), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5150 ( .A1(n3206), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4121) );
  NAND4_X1 U5151 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4125)
         );
  NOR2_X1 U5152 ( .A1(n4126), .A2(n4125), .ZN(n4127) );
  NOR2_X1 U5153 ( .A1(n4160), .A2(n4127), .ZN(n5324) );
  NAND2_X1 U5154 ( .A1(n5323), .A2(n5324), .ZN(n4131) );
  NAND2_X1 U5155 ( .A1(n5311), .A2(n4129), .ZN(n4130) );
  XOR2_X1 U5156 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4146), .Z(n5901) );
  AOI22_X1 U5157 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_14__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5158 ( .A1(n3208), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5159 ( .A1(n4415), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5160 ( .A1(n3210), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5161 ( .A1(n3206), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U5162 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4143)
         );
  AOI22_X1 U5163 ( .A1(n4431), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5164 ( .A1(n3484), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U5165 ( .A1(n4413), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5166 ( .A1(n3561), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4137) );
  NAND4_X1 U5167 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4142)
         );
  OAI21_X1 U5168 ( .B1(n4143), .B2(n4142), .A(n4141), .ZN(n4144) );
  OAI211_X1 U5169 ( .C1(n5901), .C2(n4493), .A(n4145), .B(n4144), .ZN(n5404)
         );
  AOI21_X1 U5170 ( .B1(n6933), .B2(n4147), .A(n4163), .ZN(n5890) );
  AOI22_X1 U5171 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_15__SCAN_IN), .ZN(n4148) );
  OAI21_X1 U5172 ( .B1(n5890), .B2(n4493), .A(n4148), .ZN(n4162) );
  AOI22_X1 U5173 ( .A1(n4431), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5174 ( .A1(n3678), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5175 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n3209), .B1(n4408), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5176 ( .A1(n3206), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4149) );
  NAND4_X1 U5177 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4158)
         );
  AOI22_X1 U5178 ( .A1(n3561), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5179 ( .A1(n4413), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5180 ( .A1(n4415), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5181 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n3484), .B1(n4299), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4153) );
  NAND4_X1 U5182 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(n4157)
         );
  NOR2_X1 U5183 ( .A1(n4158), .A2(n4157), .ZN(n4159) );
  NOR2_X1 U5184 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  NOR2_X1 U5185 ( .A1(n4162), .A2(n4161), .ZN(n5400) );
  AOI21_X1 U5186 ( .B1(n6766), .B2(n4164), .A(n4178), .ZN(n5884) );
  AOI22_X1 U5187 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_16__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5188 ( .A1(n3484), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5189 ( .A1(n3444), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U5190 ( .A1(n4414), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U5191 ( .A1(n4431), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4165) );
  NAND4_X1 U5192 ( .A1(n4168), .A2(n4167), .A3(n4166), .A4(n4165), .ZN(n4175)
         );
  AOI22_X1 U5193 ( .A1(n4415), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5194 ( .A1(n4413), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5195 ( .A1(n3678), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5196 ( .A1(n3206), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4169) );
  NAND4_X1 U5197 ( .A1(n4172), .A2(n4171), .A3(n4170), .A4(n4169), .ZN(n4174)
         );
  OAI21_X1 U5198 ( .B1(n4175), .B2(n4174), .A(n4455), .ZN(n4176) );
  OAI211_X1 U5199 ( .C1(n5884), .C2(n4493), .A(n4177), .B(n4176), .ZN(n5395)
         );
  OAI21_X1 U5200 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4178), .A(n4207), 
        .ZN(n5878) );
  AOI22_X1 U5201 ( .A1(EAX_REG_17__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6403), .ZN(n4193) );
  AOI22_X1 U5202 ( .A1(n3561), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4185) );
  INV_X1 U5203 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4180) );
  INV_X1 U5204 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4179) );
  OAI22_X1 U5205 ( .A1(n4442), .A2(n4180), .B1(n4441), .B2(n4179), .ZN(n4181)
         );
  INV_X1 U5206 ( .A(n4181), .ZN(n4184) );
  AOI22_X1 U5207 ( .A1(n3444), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U5208 ( .A1(n4299), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4182) );
  NAND4_X1 U5209 ( .A1(n4185), .A2(n4184), .A3(n4183), .A4(n4182), .ZN(n4191)
         );
  AOI22_X1 U5210 ( .A1(n3206), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5211 ( .A1(n4431), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U5212 ( .A1(n3484), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5213 ( .A1(n4415), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4186) );
  NAND4_X1 U5214 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4190)
         );
  OAI21_X1 U5215 ( .B1(n4191), .B2(n4190), .A(n4455), .ZN(n4192) );
  NAND3_X1 U5216 ( .A1(n4493), .A2(n4193), .A3(n4192), .ZN(n4194) );
  OAI21_X1 U5217 ( .B1(n4493), .B2(n5878), .A(n4194), .ZN(n5762) );
  XNOR2_X1 U5218 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4207), .ZN(n5869)
         );
  AOI22_X1 U5219 ( .A1(EAX_REG_18__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6403), .ZN(n4206) );
  AOI22_X1 U5220 ( .A1(n4413), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5221 ( .A1(n3484), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U5222 ( .A1(n4431), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U5223 ( .A1(n3206), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4195) );
  NAND4_X1 U5224 ( .A1(n4198), .A2(n4197), .A3(n4196), .A4(n4195), .ZN(n4204)
         );
  AOI22_X1 U5225 ( .A1(n4415), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5226 ( .A1(n4407), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5227 ( .A1(n3208), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5228 ( .A1(n4414), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4199) );
  NAND4_X1 U5229 ( .A1(n4202), .A2(n4201), .A3(n4200), .A4(n4199), .ZN(n4203)
         );
  AOI221_X1 U5230 ( .B1(n4204), .B2(n4455), .C1(n4203), .C2(n4455), .A(n4458), 
        .ZN(n4205) );
  AOI22_X1 U5231 ( .A1(n4458), .A2(n5869), .B1(n4206), .B2(n4205), .ZN(n5390)
         );
  OAI21_X1 U5232 ( .B1(n4208), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n4222), 
        .ZN(n5747) );
  AOI22_X1 U5233 ( .A1(EAX_REG_19__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6403), .ZN(n4220) );
  AOI22_X1 U5234 ( .A1(n4431), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U5235 ( .A1(n3209), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U5236 ( .A1(n3208), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U5237 ( .A1(n4415), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4209) );
  NAND4_X1 U5238 ( .A1(n4212), .A2(n4211), .A3(n4210), .A4(n4209), .ZN(n4218)
         );
  AOI22_X1 U5239 ( .A1(n4413), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5240 ( .A1(n4407), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5241 ( .A1(n3484), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5242 ( .A1(n3206), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4213) );
  NAND4_X1 U5243 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4217)
         );
  OAI21_X1 U5244 ( .B1(n4218), .B2(n4217), .A(n4455), .ZN(n4219) );
  NAND3_X1 U5245 ( .A1(n4493), .A2(n4220), .A3(n4219), .ZN(n4221) );
  OAI21_X1 U5246 ( .B1(n4493), .B2(n5747), .A(n4221), .ZN(n5682) );
  AOI21_X1 U5247 ( .B1(n6780), .B2(n4222), .A(n4235), .ZN(n5672) );
  AOI22_X1 U5248 ( .A1(EAX_REG_20__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6403), .ZN(n4234) );
  AOI22_X1 U5249 ( .A1(n4413), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4226) );
  AOI22_X1 U5250 ( .A1(n3561), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4225) );
  AOI22_X1 U5251 ( .A1(n3209), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U5252 ( .A1(n4415), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4223) );
  NAND4_X1 U5253 ( .A1(n4226), .A2(n4225), .A3(n4224), .A4(n4223), .ZN(n4232)
         );
  AOI22_X1 U5254 ( .A1(n4431), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4230) );
  AOI22_X1 U5255 ( .A1(n3678), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U5256 ( .A1(n3484), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U5257 ( .A1(n3206), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4227) );
  NAND4_X1 U5258 ( .A1(n4230), .A2(n4229), .A3(n4228), .A4(n4227), .ZN(n4231)
         );
  AOI221_X1 U5259 ( .B1(n4232), .B2(n4455), .C1(n4231), .C2(n4455), .A(n4458), 
        .ZN(n4233) );
  AOI22_X1 U5260 ( .A1(n4458), .A2(n5672), .B1(n4234), .B2(n4233), .ZN(n5433)
         );
  OAI21_X1 U5261 ( .B1(n4235), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4250), 
        .ZN(n5735) );
  INV_X1 U5262 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6109) );
  AOI22_X1 U5263 ( .A1(n4431), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U5264 ( .A1(n3208), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U5265 ( .A1(n3210), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5266 ( .A1(n3206), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4236) );
  NAND4_X1 U5267 ( .A1(n4239), .A2(n4238), .A3(n4237), .A4(n4236), .ZN(n4245)
         );
  AOI22_X1 U5268 ( .A1(n3561), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U5269 ( .A1(n4413), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5270 ( .A1(n3484), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5271 ( .A1(n4415), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4240) );
  NAND4_X1 U5272 ( .A1(n4243), .A2(n4242), .A3(n4241), .A4(n4240), .ZN(n4244)
         );
  OAI21_X1 U5273 ( .B1(n4245), .B2(n4244), .A(n4455), .ZN(n4247) );
  OAI21_X1 U5274 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n4392), .A(n6403), 
        .ZN(n4246) );
  OAI211_X1 U5275 ( .C1(n3298), .C2(n6109), .A(n4247), .B(n4246), .ZN(n4248)
         );
  OAI21_X1 U5276 ( .B1(n5735), .B2(n4493), .A(n4248), .ZN(n5384) );
  AND2_X1 U5277 ( .A1(n4250), .A2(n4249), .ZN(n4251) );
  NOR2_X1 U5278 ( .A1(n4251), .A2(n4264), .ZN(n5731) );
  AOI22_X1 U5279 ( .A1(EAX_REG_22__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6403), .ZN(n4263) );
  AOI22_X1 U5280 ( .A1(n3678), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U5281 ( .A1(n4414), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5282 ( .A1(n3210), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5283 ( .A1(n4415), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4252) );
  NAND4_X1 U5284 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(n4261)
         );
  AOI22_X1 U5285 ( .A1(n4431), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4259) );
  AOI22_X1 U5286 ( .A1(n4413), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U5287 ( .A1(n4407), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U5288 ( .A1(n3206), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4256) );
  NAND4_X1 U5289 ( .A1(n4259), .A2(n4258), .A3(n4257), .A4(n4256), .ZN(n4260)
         );
  AOI221_X1 U5290 ( .B1(n4261), .B2(n4455), .C1(n4260), .C2(n4455), .A(n4458), 
        .ZN(n4262) );
  AOI22_X1 U5291 ( .A1(n4458), .A2(n5731), .B1(n4263), .B2(n4262), .ZN(n5381)
         );
  OR2_X1 U5292 ( .A1(n4264), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4265)
         );
  NAND2_X1 U5293 ( .A1(n4313), .A2(n4265), .ZN(n5650) );
  AOI22_X1 U5294 ( .A1(n3678), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4269) );
  AOI22_X1 U5295 ( .A1(n3444), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U5296 ( .A1(n3209), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U5297 ( .A1(n3206), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4266) );
  NAND4_X1 U5298 ( .A1(n4269), .A2(n4268), .A3(n4267), .A4(n4266), .ZN(n4275)
         );
  AOI22_X1 U5299 ( .A1(n4415), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U5300 ( .A1(n4413), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U5301 ( .A1(n4431), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U5302 ( .A1(n3484), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4270) );
  NAND4_X1 U5303 ( .A1(n4273), .A2(n4272), .A3(n4271), .A4(n4270), .ZN(n4274)
         );
  NOR2_X1 U5304 ( .A1(n4275), .A2(n4274), .ZN(n4291) );
  AOI22_X1 U5305 ( .A1(n4413), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4279) );
  AOI22_X1 U5306 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n3206), .B1(n3484), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U5307 ( .A1(n4415), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5308 ( .A1(n3678), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4276) );
  NAND4_X1 U5309 ( .A1(n4279), .A2(n4278), .A3(n4277), .A4(n4276), .ZN(n4285)
         );
  AOI22_X1 U5310 ( .A1(n4431), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4283) );
  AOI22_X1 U5311 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n3210), .B1(n4414), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4282) );
  AOI22_X1 U5312 ( .A1(n3561), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U5313 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n4299), .B1(n3446), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4280) );
  NAND4_X1 U5314 ( .A1(n4283), .A2(n4282), .A3(n4281), .A4(n4280), .ZN(n4284)
         );
  NOR2_X1 U5315 ( .A1(n4285), .A2(n4284), .ZN(n4292) );
  XOR2_X1 U5316 ( .A(n4291), .B(n4292), .Z(n4286) );
  NAND2_X1 U5317 ( .A1(n4455), .A2(n4286), .ZN(n4288) );
  AOI22_X1 U5318 ( .A1(EAX_REG_23__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6403), .ZN(n4287) );
  NAND3_X1 U5319 ( .A1(n4288), .A2(n4287), .A3(n4493), .ZN(n4289) );
  XNOR2_X1 U5320 ( .A(n4313), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5644)
         );
  NOR2_X1 U5321 ( .A1(n4292), .A2(n4291), .ZN(n4316) );
  AOI22_X1 U5322 ( .A1(n4431), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4298) );
  INV_X1 U5323 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4293) );
  INV_X1 U5324 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5111) );
  OAI22_X1 U5325 ( .A1(n4442), .A2(n4293), .B1(n4441), .B2(n5111), .ZN(n4294)
         );
  INV_X1 U5326 ( .A(n4294), .ZN(n4297) );
  AOI22_X1 U5327 ( .A1(n4407), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U5328 ( .A1(n4415), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4295) );
  NAND4_X1 U5329 ( .A1(n4298), .A2(n4297), .A3(n4296), .A4(n4295), .ZN(n4305)
         );
  AOI22_X1 U5330 ( .A1(n3484), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U5331 ( .A1(n3444), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4302) );
  AOI22_X1 U5332 ( .A1(n3209), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4301) );
  AOI22_X1 U5333 ( .A1(n3206), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4300) );
  NAND4_X1 U5334 ( .A1(n4303), .A2(n4302), .A3(n4301), .A4(n4300), .ZN(n4304)
         );
  OR2_X1 U5335 ( .A1(n4316), .A2(n4315), .ZN(n4310) );
  INV_X1 U5336 ( .A(n4455), .ZN(n4425) );
  AOI21_X1 U5337 ( .B1(n4316), .B2(n4315), .A(n4425), .ZN(n4309) );
  AOI22_X1 U5338 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n4459), .B1(n4306), 
        .B2(EAX_REG_24__SCAN_IN), .ZN(n4307) );
  INV_X1 U5339 ( .A(n4307), .ZN(n4308) );
  AOI21_X1 U5340 ( .B1(n4310), .B2(n4309), .A(n4308), .ZN(n4311) );
  NAND2_X1 U5341 ( .A1(n4312), .A2(n4311), .ZN(n4489) );
  NAND2_X1 U5342 ( .A1(n4486), .A2(n4489), .ZN(n4488) );
  INV_X1 U5343 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4484) );
  OAI21_X1 U5344 ( .B1(n4314), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n4333), 
        .ZN(n5730) );
  NAND2_X1 U5345 ( .A1(n4316), .A2(n4315), .ZN(n4334) );
  INV_X1 U5346 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4939) );
  NOR2_X1 U5347 ( .A1(n4441), .A2(n4939), .ZN(n4320) );
  OAI22_X1 U5348 ( .A1(n4343), .A2(n4318), .B1(n3203), .B2(n4317), .ZN(n4319)
         );
  AOI211_X1 U5349 ( .C1(INSTQUEUE_REG_8__2__SCAN_IN), .C2(n3208), .A(n4320), 
        .B(n4319), .ZN(n4323) );
  AOI22_X1 U5350 ( .A1(n4414), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U5351 ( .A1(n4299), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4321) );
  NAND3_X1 U5352 ( .A1(n4323), .A2(n4322), .A3(n4321), .ZN(n4329) );
  AOI22_X1 U5353 ( .A1(n4431), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U5354 ( .A1(n3444), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U5355 ( .A1(n3206), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U5356 ( .A1(n4407), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4324) );
  NAND4_X1 U5357 ( .A1(n4327), .A2(n4326), .A3(n4325), .A4(n4324), .ZN(n4328)
         );
  NOR2_X1 U5358 ( .A1(n4329), .A2(n4328), .ZN(n4335) );
  XNOR2_X1 U5359 ( .A(n4334), .B(n4335), .ZN(n4331) );
  AOI22_X1 U5360 ( .A1(EAX_REG_25__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6403), .ZN(n4330) );
  OAI21_X1 U5361 ( .B1(n4331), .B2(n4425), .A(n4330), .ZN(n4332) );
  AOI22_X1 U5362 ( .A1(n4458), .A2(n5730), .B1(n4332), .B2(n4493), .ZN(n5367)
         );
  NOR2_X2 U5363 ( .A1(n4488), .A2(n5367), .ZN(n5362) );
  INV_X1 U5364 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6913) );
  AOI21_X1 U5365 ( .B1(n6913), .B2(n4333), .A(n4354), .ZN(n5719) );
  NOR2_X1 U5366 ( .A1(n4335), .A2(n4334), .ZN(n4356) );
  AOI22_X1 U5367 ( .A1(n3484), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U5368 ( .A1(n3444), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U5369 ( .A1(n3206), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U5370 ( .A1(n3210), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4336) );
  NAND4_X1 U5371 ( .A1(n4339), .A2(n4338), .A3(n4337), .A4(n4336), .ZN(n4350)
         );
  INV_X1 U5372 ( .A(n4340), .ZN(n4343) );
  AOI22_X1 U5373 ( .A1(n4431), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U5374 ( .A1(n3202), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4341) );
  OAI211_X1 U5375 ( .C1(n4344), .C2(n4343), .A(n4342), .B(n4341), .ZN(n4349)
         );
  INV_X1 U5376 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4769) );
  INV_X1 U5377 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4345) );
  OAI22_X1 U5378 ( .A1(n3464), .A2(n4769), .B1(n3465), .B2(n4345), .ZN(n4348)
         );
  INV_X1 U5379 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4346) );
  INV_X1 U5380 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4830) );
  OAI22_X1 U5381 ( .A1(n4442), .A2(n4346), .B1(n4441), .B2(n4830), .ZN(n4347)
         );
  XOR2_X1 U5382 ( .A(n4356), .B(n4355), .Z(n4351) );
  AOI22_X1 U5383 ( .A1(n4455), .A2(n4351), .B1(n4306), .B2(EAX_REG_26__SCAN_IN), .ZN(n4353) );
  OAI21_X1 U5384 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n4392), .A(n6403), 
        .ZN(n4352) );
  NAND2_X1 U5385 ( .A1(n5362), .A2(n5364), .ZN(n5357) );
  OAI21_X1 U5386 ( .B1(n4354), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4402), 
        .ZN(n5627) );
  NAND2_X1 U5387 ( .A1(n4356), .A2(n4355), .ZN(n4372) );
  INV_X1 U5388 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4357) );
  INV_X1 U5389 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5006) );
  OAI22_X1 U5390 ( .A1(n4442), .A2(n4357), .B1(n4441), .B2(n5006), .ZN(n4358)
         );
  INV_X1 U5391 ( .A(n4358), .ZN(n4362) );
  AOI22_X1 U5392 ( .A1(n3444), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4361) );
  AOI22_X1 U5393 ( .A1(n4407), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U5394 ( .A1(n3561), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4359) );
  NAND4_X1 U5395 ( .A1(n4362), .A2(n4361), .A3(n4360), .A4(n4359), .ZN(n4368)
         );
  AOI22_X1 U5396 ( .A1(n4431), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4366) );
  AOI22_X1 U5397 ( .A1(n4414), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U5398 ( .A1(n3209), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U5399 ( .A1(n3206), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4363) );
  NAND4_X1 U5400 ( .A1(n4366), .A2(n4365), .A3(n4364), .A4(n4363), .ZN(n4367)
         );
  NOR2_X1 U5401 ( .A1(n4368), .A2(n4367), .ZN(n4373) );
  XNOR2_X1 U5402 ( .A(n4372), .B(n4373), .ZN(n4370) );
  AOI22_X1 U5403 ( .A1(EAX_REG_27__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6403), .ZN(n4369) );
  OAI21_X1 U5404 ( .B1(n4370), .B2(n4425), .A(n4369), .ZN(n4371) );
  AOI22_X1 U5405 ( .A1(n4458), .A2(n5627), .B1(n4371), .B2(n4493), .ZN(n5359)
         );
  NOR2_X2 U5406 ( .A1(n5357), .A2(n5359), .ZN(n5358) );
  XNOR2_X1 U5407 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(n4402), .ZN(n5614)
         );
  AOI22_X1 U5408 ( .A1(EAX_REG_28__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6403), .ZN(n4387) );
  NOR2_X1 U5409 ( .A1(n4373), .A2(n4372), .ZN(n4423) );
  INV_X1 U5410 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4374) );
  OAI22_X1 U5411 ( .A1(n4442), .A2(n4374), .B1(n4441), .B2(n4998), .ZN(n4376)
         );
  INV_X1 U5412 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5082) );
  NOR2_X1 U5413 ( .A1(n3464), .A2(n5082), .ZN(n4375) );
  AOI211_X1 U5414 ( .C1(INSTQUEUE_REG_12__5__SCAN_IN), .C2(n4439), .A(n4376), 
        .B(n4375), .ZN(n4384) );
  AOI22_X1 U5415 ( .A1(n4415), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U5416 ( .A1(n4431), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U5417 ( .A1(n3484), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4380) );
  AOI22_X1 U5418 ( .A1(n3444), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4379) );
  AOI22_X1 U5419 ( .A1(n3210), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4299), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U5420 ( .A1(n3206), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4377) );
  AND4_X1 U5421 ( .A1(n4380), .A2(n4379), .A3(n4378), .A4(n4377), .ZN(n4381)
         );
  NAND4_X1 U5422 ( .A1(n4384), .A2(n4383), .A3(n4382), .A4(n4381), .ZN(n4422)
         );
  XOR2_X1 U5423 ( .A(n4423), .B(n4422), .Z(n4385) );
  AOI21_X1 U5424 ( .B1(n4385), .B2(n4455), .A(n4458), .ZN(n4386) );
  AOI22_X1 U5425 ( .A1(n4458), .A2(n5614), .B1(n4387), .B2(n4386), .ZN(n4388)
         );
  INV_X1 U5426 ( .A(n4537), .ZN(n4390) );
  OR2_X1 U5427 ( .A1(n5358), .A2(n4388), .ZN(n4389) );
  NAND3_X1 U5428 ( .A1(n6523), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6536) );
  AOI21_X1 U5429 ( .B1(n6618), .B2(n6617), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n4391) );
  NAND2_X1 U5430 ( .A1(n6523), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4394) );
  INV_X1 U5431 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n4392) );
  NAND2_X1 U5432 ( .A1(n4392), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U5433 ( .A1(n4394), .A2(n4393), .ZN(n4639) );
  AOI22_X1 U5434 ( .A1(n6221), .A2(REIP_REG_28__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4395) );
  INV_X1 U5435 ( .A(n4395), .ZN(n4396) );
  NAND2_X1 U5436 ( .A1(n4400), .A2(n4399), .ZN(U2958) );
  INV_X1 U5437 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4401) );
  INV_X1 U5438 ( .A(n4403), .ZN(n4405) );
  INV_X1 U5439 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U5440 ( .A1(n4405), .A2(n4404), .ZN(n4406) );
  NAND2_X1 U5441 ( .A1(n4470), .A2(n4406), .ZN(n5608) );
  AOI22_X1 U5442 ( .A1(n3208), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4412) );
  AOI22_X1 U5443 ( .A1(n3206), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U5444 ( .A1(n3561), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4439), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U5445 ( .A1(n3444), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4409) );
  NAND4_X1 U5446 ( .A1(n4412), .A2(n4411), .A3(n4410), .A4(n4409), .ZN(n4421)
         );
  AOI22_X1 U5447 ( .A1(n4413), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4419) );
  AOI22_X1 U5448 ( .A1(n3484), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U5449 ( .A1(n4415), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4417) );
  AOI22_X1 U5450 ( .A1(n4299), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4416) );
  NAND4_X1 U5451 ( .A1(n4419), .A2(n4418), .A3(n4417), .A4(n4416), .ZN(n4420)
         );
  NOR2_X1 U5452 ( .A1(n4421), .A2(n4420), .ZN(n4430) );
  NAND2_X1 U5453 ( .A1(n4423), .A2(n4422), .ZN(n4429) );
  XNOR2_X1 U5454 ( .A(n4430), .B(n4429), .ZN(n4426) );
  AOI22_X1 U5455 ( .A1(EAX_REG_29__SCAN_IN), .A2(n4306), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6403), .ZN(n4424) );
  OAI211_X1 U5456 ( .C1(n4426), .C2(n4425), .A(n4424), .B(n4493), .ZN(n4427)
         );
  XNOR2_X1 U5457 ( .A(n4470), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5598)
         );
  NOR2_X1 U5458 ( .A1(n4430), .A2(n4429), .ZN(n4451) );
  AOI22_X1 U5459 ( .A1(n4431), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3561), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4435) );
  AOI22_X1 U5460 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n3484), .B1(n3209), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4434) );
  AOI22_X1 U5461 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n3444), .B1(n4408), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U5462 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n4299), .B1(n3446), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4432) );
  NAND4_X1 U5463 ( .A1(n4435), .A2(n4434), .A3(n4433), .A4(n4432), .ZN(n4449)
         );
  OAI22_X1 U5464 ( .A1(n4343), .A2(n4437), .B1(n3203), .B2(n4436), .ZN(n4447)
         );
  INV_X1 U5465 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4814) );
  INV_X1 U5466 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4784) );
  OAI22_X1 U5467 ( .A1(n4814), .A2(n3198), .B1(n4438), .B2(n4784), .ZN(n4446)
         );
  INV_X1 U5468 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4766) );
  INV_X1 U5469 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4440) );
  OAI22_X1 U5470 ( .A1(n3464), .A2(n4766), .B1(n3465), .B2(n4440), .ZN(n4445)
         );
  INV_X1 U5471 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4443) );
  INV_X1 U5472 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n7029) );
  OAI22_X1 U5473 ( .A1(n4443), .A2(n4442), .B1(n4441), .B2(n7029), .ZN(n4444)
         );
  OR4_X1 U5474 ( .A1(n4447), .A2(n4446), .A3(n4445), .A4(n4444), .ZN(n4448) );
  NOR2_X1 U5475 ( .A1(n4449), .A2(n4448), .ZN(n4450) );
  XNOR2_X1 U5476 ( .A(n4451), .B(n4450), .ZN(n4456) );
  INV_X1 U5477 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4453) );
  OAI21_X1 U5478 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n4392), .A(n6403), 
        .ZN(n4452) );
  OAI21_X1 U5479 ( .B1(n3298), .B2(n4453), .A(n4452), .ZN(n4454) );
  AOI21_X1 U5480 ( .B1(n4456), .B2(n4455), .A(n4454), .ZN(n4457) );
  AOI21_X1 U5481 ( .B1(n5598), .B2(n4458), .A(n4457), .ZN(n4557) );
  AOI22_X1 U5482 ( .A1(n4306), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4459), .ZN(n4460) );
  AND2_X1 U5483 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4462) );
  NAND2_X1 U5484 ( .A1(n4463), .A2(n4462), .ZN(n5452) );
  AND2_X1 U5485 ( .A1(n4464), .A2(n5481), .ZN(n5415) );
  NAND2_X1 U5486 ( .A1(n5415), .A2(n3302), .ZN(n4466) );
  OAI21_X1 U5487 ( .B1(n4467), .B2(n5452), .A(n4466), .ZN(n4468) );
  XNOR2_X1 U5488 ( .A(n4468), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5458)
         );
  INV_X1 U5489 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4469) );
  NOR2_X1 U5490 ( .A1(n6256), .A2(n4469), .ZN(n5450) );
  INV_X1 U5491 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5600) );
  INV_X1 U5492 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4471) );
  NOR2_X1 U5493 ( .A1(n5292), .A2(n6193), .ZN(n4473) );
  AOI211_X1 U5494 ( .C1(n6194), .C2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5450), 
        .B(n4473), .ZN(n4474) );
  NAND3_X1 U5495 ( .A1(n4476), .A2(n4475), .A3(n4474), .ZN(U2955) );
  NAND2_X1 U5496 ( .A1(n3725), .A2(n5541), .ZN(n4477) );
  XNOR2_X1 U5497 ( .A(n5756), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5431)
         );
  INV_X1 U5498 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4478) );
  XNOR2_X1 U5499 ( .A(n5754), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5514)
         );
  INV_X1 U5500 ( .A(n5513), .ZN(n4479) );
  NAND3_X1 U5501 ( .A1(n3725), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4480) );
  NOR2_X1 U5502 ( .A1(n3725), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5502)
         );
  NAND2_X1 U5503 ( .A1(n5513), .A2(n5502), .ZN(n5423) );
  XNOR2_X1 U5504 ( .A(n4482), .B(n4481), .ZN(n4542) );
  NAND2_X1 U5505 ( .A1(n5644), .A2(n6198), .ZN(n4483) );
  NAND2_X1 U5506 ( .A1(n6221), .A2(REIP_REG_24__SCAN_IN), .ZN(n4546) );
  OAI211_X1 U5507 ( .C1(n5741), .C2(n4484), .A(n4483), .B(n4546), .ZN(n4485)
         );
  AOI21_X1 U5508 ( .B1(n4542), .B2(n6199), .A(n4485), .ZN(n4491) );
  OAI21_X1 U5509 ( .B1(n4487), .B2(n4489), .A(n4488), .ZN(n5699) );
  NAND2_X1 U5510 ( .A1(n4491), .A2(n4490), .ZN(U2962) );
  NAND2_X1 U5511 ( .A1(n4492), .A2(n4565), .ZN(n4575) );
  NAND2_X1 U5512 ( .A1(n5334), .A2(n6403), .ZN(n6535) );
  NOR3_X1 U5513 ( .A1(n6523), .A2(n6605), .A3(n6535), .ZN(n6521) );
  NOR3_X1 U5514 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5334), .A3(n4493), .ZN(
        n6531) );
  INV_X1 U5515 ( .A(n6531), .ZN(n4494) );
  NAND2_X1 U5516 ( .A1(n6256), .A2(n4494), .ZN(n4495) );
  NOR2_X1 U5517 ( .A1(n6521), .A2(n4495), .ZN(n4496) );
  NAND2_X1 U5518 ( .A1(n5965), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5290) );
  INV_X1 U5519 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6597) );
  INV_X1 U5520 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6590) );
  NAND3_X1 U5521 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4509) );
  INV_X1 U5522 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6874) );
  INV_X1 U5523 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6579) );
  INV_X1 U5524 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U5525 ( .A1(n3834), .A2(n5596), .ZN(n4497) );
  NAND2_X1 U5526 ( .A1(n3821), .A2(n4392), .ZN(n5293) );
  AOI21_X1 U5527 ( .B1(n6075), .B2(n4497), .A(n5293), .ZN(n4498) );
  AND2_X2 U5528 ( .A1(n5299), .A2(n4498), .ZN(n5997) );
  INV_X1 U5529 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6572) );
  INV_X1 U5530 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6570) );
  INV_X1 U5531 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6568) );
  INV_X1 U5532 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6768) );
  INV_X1 U5533 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6563) );
  INV_X1 U5534 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6855) );
  INV_X1 U5535 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6559) );
  NAND3_X1 U5536 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5996) );
  NOR3_X1 U5537 ( .A1(n6855), .A2(n6559), .A3(n5996), .ZN(n5966) );
  NAND3_X1 U5538 ( .A1(n5966), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .ZN(n5954) );
  NOR2_X1 U5539 ( .A1(n6563), .A2(n5954), .ZN(n5937) );
  NAND2_X1 U5540 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5937), .ZN(n5933) );
  NOR2_X1 U5541 ( .A1(n6768), .A2(n5933), .ZN(n5930) );
  NAND2_X1 U5542 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5930), .ZN(n5906) );
  NOR2_X1 U5543 ( .A1(n6568), .A2(n5906), .ZN(n5909) );
  NAND2_X1 U5544 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5909), .ZN(n5898) );
  NOR2_X1 U5545 ( .A1(n6570), .A2(n5898), .ZN(n5880) );
  NAND2_X1 U5546 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5880), .ZN(n5879) );
  NOR2_X1 U5547 ( .A1(n6572), .A2(n5879), .ZN(n4505) );
  NAND2_X1 U5548 ( .A1(n5997), .A2(n4505), .ZN(n5872) );
  NAND3_X1 U5549 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        n5865), .ZN(n5669) );
  NAND2_X1 U5550 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5658), .ZN(n5660) );
  NAND2_X1 U5551 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5654), .ZN(n5639) );
  NOR2_X1 U5552 ( .A1(n4509), .A2(n5639), .ZN(n5623) );
  NAND2_X1 U5553 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5623), .ZN(n5617) );
  NOR2_X1 U5554 ( .A1(n6590), .A2(n5617), .ZN(n4510) );
  NAND2_X1 U5555 ( .A1(REIP_REG_29__SCAN_IN), .A2(n4510), .ZN(n4504) );
  NOR3_X1 U5556 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6597), .A3(n4504), .ZN(n4502) );
  NAND2_X1 U5557 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5299), .ZN(n4500) );
  INV_X1 U5558 ( .A(n5293), .ZN(n4499) );
  NAND2_X1 U5559 ( .A1(n5596), .A2(n4499), .ZN(n6520) );
  NAND2_X1 U5560 ( .A1(n4588), .A2(n6520), .ZN(n5294) );
  OAI22_X1 U5561 ( .A1(n4471), .A2(n6012), .B1(n4500), .B2(n5294), .ZN(n4501)
         );
  AOI21_X1 U5562 ( .B1(n4569), .B2(n5978), .A(n4503), .ZN(n4525) );
  NOR2_X1 U5563 ( .A1(REIP_REG_30__SCAN_IN), .A2(n4504), .ZN(n5602) );
  NAND2_X1 U5564 ( .A1(n5965), .A2(n5993), .ZN(n5676) );
  INV_X1 U5565 ( .A(n5676), .ZN(n4508) );
  INV_X1 U5566 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6583) );
  INV_X1 U5567 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6581) );
  NOR3_X1 U5568 ( .A1(n6583), .A2(n6874), .A3(n6581), .ZN(n4507) );
  NAND3_X1 U5569 ( .A1(REIP_REG_17__SCAN_IN), .A2(n4505), .A3(n5965), .ZN(
        n5675) );
  NAND3_X1 U5570 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4506) );
  OAI21_X1 U5571 ( .B1(n5675), .B2(n4506), .A(n5676), .ZN(n5668) );
  OAI21_X1 U5572 ( .B1(n4508), .B2(n4507), .A(n5668), .ZN(n5653) );
  AOI21_X1 U5573 ( .B1(n5676), .B2(n4509), .A(n5653), .ZN(n5629) );
  NAND2_X1 U5574 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5629), .ZN(n5624) );
  OAI21_X1 U5575 ( .B1(n6590), .B2(n5624), .A(n5676), .ZN(n5616) );
  INV_X1 U5576 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U5577 ( .A1(n4510), .A2(n5607), .ZN(n5612) );
  NAND2_X1 U5578 ( .A1(n5616), .A2(n5612), .ZN(n5603) );
  OAI21_X1 U5579 ( .B1(n5602), .B2(n5603), .A(REIP_REG_31__SCAN_IN), .ZN(n4524) );
  INV_X1 U5580 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4513) );
  MUX2_X1 U5581 ( .A(n4511), .B(n4513), .S(n3204), .Z(n4515) );
  NAND2_X1 U5582 ( .A1(n4513), .A2(n4512), .ZN(n4514) );
  NAND2_X1 U5583 ( .A1(n4515), .A2(n4514), .ZN(n4535) );
  NOR2_X1 U5584 ( .A1(n4536), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U5585 ( .A1(n4534), .A2(n4516), .ZN(n4518) );
  NAND2_X1 U5586 ( .A1(n4518), .A2(n4517), .ZN(n4520) );
  OAI22_X1 U5587 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n6075), .ZN(n4519) );
  INV_X1 U5588 ( .A(n6025), .ZN(n4522) );
  AND3_X1 U5589 ( .A1(n4530), .A2(EBX_REG_31__SCAN_IN), .A3(n5293), .ZN(n4521)
         );
  NAND3_X1 U5590 ( .A1(n4525), .A2(n4524), .A3(n4523), .ZN(U2796) );
  INV_X1 U5591 ( .A(n4606), .ZN(n4526) );
  NAND2_X1 U5592 ( .A1(n4623), .A2(n4526), .ZN(n4614) );
  NAND3_X1 U5593 ( .A1(n4527), .A2(n5328), .A3(n4999), .ZN(n4529) );
  OR2_X1 U5594 ( .A1(n4529), .A2(n4528), .ZN(n4564) );
  INV_X1 U5595 ( .A(n4564), .ZN(n4531) );
  NAND2_X1 U5596 ( .A1(n4531), .A2(n4530), .ZN(n4532) );
  NAND2_X1 U5597 ( .A1(n4614), .A2(n4532), .ZN(n4533) );
  INV_X1 U5598 ( .A(n6071), .ZN(n4541) );
  AOI21_X1 U5599 ( .B1(n4536), .B2(n4535), .A(n4534), .ZN(n5611) );
  INV_X1 U5600 ( .A(n5611), .ZN(n4540) );
  NOR2_X1 U5601 ( .A1(n4537), .A2(n4538), .ZN(n4539) );
  NAND2_X2 U5602 ( .A1(n6081), .A2(n4857), .ZN(n6083) );
  NAND2_X1 U5603 ( .A1(n4542), .A2(n3833), .ZN(n4552) );
  INV_X1 U5604 ( .A(n4543), .ZN(n5494) );
  INV_X1 U5605 ( .A(n4544), .ZN(n4545) );
  OAI21_X1 U5606 ( .B1(n5494), .B2(n4545), .A(n5638), .ZN(n5698) );
  OAI21_X1 U5607 ( .B1(n5698), .B2(n6258), .A(n4546), .ZN(n4550) );
  INV_X1 U5608 ( .A(n5531), .ZN(n4547) );
  NOR2_X1 U5609 ( .A1(n5543), .A2(n4547), .ZN(n5506) );
  NAND2_X1 U5610 ( .A1(n5506), .A2(n5507), .ZN(n5497) );
  AOI211_X1 U5611 ( .C1(n4481), .C2(n5497), .A(n4548), .B(n5779), .ZN(n4549)
         );
  NAND2_X1 U5612 ( .A1(n4552), .A2(n4551), .ZN(U2994) );
  NAND2_X1 U5613 ( .A1(n5598), .A2(n6198), .ZN(n4554) );
  OAI211_X1 U5614 ( .C1(n5600), .C2(n5741), .A(n4554), .B(n4553), .ZN(n4555)
         );
  AOI21_X1 U5615 ( .B1(n4556), .B2(n6199), .A(n4555), .ZN(n4560) );
  NAND2_X1 U5616 ( .A1(n4560), .A2(n4559), .ZN(U2956) );
  NAND2_X1 U5617 ( .A1(n4606), .A2(n4622), .ZN(n4563) );
  INV_X1 U5618 ( .A(n3829), .ZN(n5838) );
  NAND2_X1 U5619 ( .A1(n5838), .A2(n4561), .ZN(n4562) );
  NAND2_X1 U5620 ( .A1(n4563), .A2(n4562), .ZN(n4601) );
  INV_X1 U5621 ( .A(n3505), .ZN(n5289) );
  NOR2_X1 U5622 ( .A1(n4564), .A2(n5289), .ZN(n4566) );
  OAI21_X1 U5623 ( .B1(n4601), .B2(n4566), .A(n4565), .ZN(n4567) );
  NAND2_X1 U5624 ( .A1(n4569), .A2(n4568), .ZN(n4572) );
  AOI22_X1 U5625 ( .A1(EAX_REG_31__SCAN_IN), .A2(n6089), .B1(DATAI_31_), .B2(
        n6085), .ZN(n4571) );
  NAND2_X1 U5626 ( .A1(n4572), .A2(n4571), .ZN(U2860) );
  NOR2_X1 U5627 ( .A1(n6617), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5678) );
  INV_X1 U5628 ( .A(n4573), .ZN(n4574) );
  AOI211_X1 U5629 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4575), .A(n5678), .B(
        n4574), .ZN(n4576) );
  INV_X1 U5630 ( .A(n4576), .ZN(U2788) );
  NOR3_X1 U5631 ( .A1(n4583), .A2(n4577), .A3(n4622), .ZN(n4581) );
  INV_X1 U5632 ( .A(n4578), .ZN(n4579) );
  OAI22_X1 U5633 ( .A1(n4581), .A2(n4606), .B1(n4580), .B2(n4579), .ZN(n4582)
         );
  AOI21_X1 U5634 ( .B1(n4623), .B2(n4606), .A(n4582), .ZN(n6512) );
  INV_X1 U5635 ( .A(n4583), .ZN(n4603) );
  NAND2_X1 U5636 ( .A1(n4584), .A2(n4603), .ZN(n4586) );
  OR2_X1 U5637 ( .A1(n4606), .A2(n3505), .ZN(n4585) );
  NAND2_X1 U5638 ( .A1(n4586), .A2(n4585), .ZN(n5843) );
  INV_X1 U5639 ( .A(n4587), .ZN(n5298) );
  OR2_X1 U5640 ( .A1(n4588), .A2(n5298), .ZN(n4591) );
  AOI21_X1 U5641 ( .B1(n4591), .B2(n6543), .A(READY_N), .ZN(n6622) );
  NOR2_X1 U5642 ( .A1(n5843), .A2(n6622), .ZN(n6509) );
  OR2_X1 U5643 ( .A1(n6509), .A2(n6529), .ZN(n5848) );
  NAND2_X1 U5644 ( .A1(n5848), .A2(MORE_REG_SCAN_IN), .ZN(n4589) );
  OAI21_X1 U5645 ( .B1(n6512), .B2(n5848), .A(n4589), .ZN(U3471) );
  OAI21_X1 U5646 ( .B1(READREQUEST_REG_SCAN_IN), .B2(n5678), .A(n6616), .ZN(
        n4590) );
  OAI21_X1 U5647 ( .B1(n6616), .B2(n4591), .A(n4590), .ZN(U3474) );
  INV_X1 U5648 ( .A(DATAI_4_), .ZN(n5002) );
  OR2_X1 U5649 ( .A1(n4669), .A2(n5002), .ZN(n4681) );
  INV_X1 U5650 ( .A(n6519), .ZN(n5593) );
  NAND2_X1 U5651 ( .A1(n5597), .A2(n5593), .ZN(n6155) );
  AND2_X2 U5652 ( .A1(n4592), .A2(n6155), .ZN(n6152) );
  INV_X2 U5653 ( .A(n6155), .ZN(n6149) );
  AOI22_X1 U5654 ( .A1(n6152), .A2(UWORD_REG_4__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n4593) );
  NAND2_X1 U5655 ( .A1(n4681), .A2(n4593), .ZN(U2928) );
  AOI22_X1 U5656 ( .A1(n6152), .A2(UWORD_REG_3__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U5657 ( .A1(n6153), .A2(DATAI_3_), .ZN(n4673) );
  NAND2_X1 U5658 ( .A1(n4594), .A2(n4673), .ZN(U2927) );
  AOI22_X1 U5659 ( .A1(n6152), .A2(LWORD_REG_0__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U5660 ( .A1(n6153), .A2(DATAI_0_), .ZN(n4666) );
  NAND2_X1 U5661 ( .A1(n4595), .A2(n4666), .ZN(U2939) );
  AOI22_X1 U5662 ( .A1(n6152), .A2(LWORD_REG_9__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4596) );
  NAND2_X1 U5663 ( .A1(n6153), .A2(DATAI_9_), .ZN(n4662) );
  NAND2_X1 U5664 ( .A1(n4596), .A2(n4662), .ZN(U2948) );
  AOI22_X1 U5665 ( .A1(n6152), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6149), .ZN(n4597) );
  NAND2_X1 U5666 ( .A1(n6153), .A2(DATAI_2_), .ZN(n4688) );
  NAND2_X1 U5667 ( .A1(n4597), .A2(n4688), .ZN(U2926) );
  AOI22_X1 U5668 ( .A1(n6152), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6149), .ZN(n4598) );
  NAND2_X1 U5669 ( .A1(n6153), .A2(DATAI_5_), .ZN(n4686) );
  NAND2_X1 U5670 ( .A1(n4598), .A2(n4686), .ZN(U2929) );
  INV_X1 U5671 ( .A(n4600), .ZN(n4629) );
  INV_X1 U5672 ( .A(n4601), .ZN(n4612) );
  INV_X1 U5673 ( .A(n4602), .ZN(n4611) );
  NAND2_X1 U5674 ( .A1(n5594), .A2(n5596), .ZN(n4604) );
  NAND2_X1 U5675 ( .A1(n4604), .A2(n4603), .ZN(n4608) );
  INV_X1 U5676 ( .A(n4605), .ZN(n4607) );
  NAND3_X1 U5677 ( .A1(n4608), .A2(n4607), .A3(n4606), .ZN(n4609) );
  NAND2_X1 U5678 ( .A1(n4614), .A2(n4613), .ZN(n6498) );
  INV_X1 U5679 ( .A(n6498), .ZN(n4897) );
  NAND2_X1 U5680 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n5592) );
  OR2_X1 U5681 ( .A1(n6523), .A2(n5592), .ZN(n6603) );
  INV_X1 U5682 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5849) );
  OAI22_X1 U5683 ( .A1(n4897), .A2(n6529), .B1(n6603), .B2(n5849), .ZN(n5836)
         );
  NAND2_X1 U5684 ( .A1(n6523), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6604) );
  INV_X1 U5685 ( .A(n6604), .ZN(n4615) );
  AOI21_X1 U5686 ( .B1(n4629), .B2(n5343), .A(n5586), .ZN(n4633) );
  NAND4_X1 U5687 ( .A1(n3829), .A2(n4619), .A3(n4618), .A4(n3940), .ZN(n4620)
         );
  NOR2_X1 U5688 ( .A1(n4621), .A2(n4620), .ZN(n4655) );
  OR2_X1 U5689 ( .A1(n4623), .A2(n4622), .ZN(n4904) );
  XNOR2_X1 U5690 ( .A(n4600), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4626)
         );
  INV_X1 U5691 ( .A(n5594), .ZN(n5340) );
  XNOR2_X1 U5692 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4624) );
  OAI22_X1 U5693 ( .A1(n5340), .A2(n4624), .B1(n4909), .B2(n4626), .ZN(n4625)
         );
  AOI21_X1 U5694 ( .B1(n4904), .B2(n4626), .A(n4625), .ZN(n4627) );
  OAI21_X1 U5695 ( .B1(n4617), .B2(n4655), .A(n4627), .ZN(n4915) );
  INV_X1 U5696 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5697 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4628), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3536), .ZN(n5342) );
  NOR3_X1 U5698 ( .A1(n5334), .A2(n5562), .A3(n5342), .ZN(n4631) );
  NOR3_X1 U5699 ( .A1(n4629), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6524), 
        .ZN(n4630) );
  AOI211_X1 U5700 ( .C1(n4915), .C2(n5837), .A(n4631), .B(n4630), .ZN(n4632)
         );
  OAI22_X1 U5701 ( .A1(n4633), .A2(n3307), .B1(n5586), .B2(n4632), .ZN(U3459)
         );
  XNOR2_X1 U5702 ( .A(n4634), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4654)
         );
  NAND2_X1 U5703 ( .A1(n4636), .A2(n4635), .ZN(n4637) );
  NAND2_X1 U5704 ( .A1(n4638), .A2(n4637), .ZN(n6084) );
  INV_X1 U5705 ( .A(n6084), .ZN(n4643) );
  INV_X1 U5706 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6613) );
  NOR2_X1 U5707 ( .A1(n6256), .A2(n6613), .ZN(n4649) );
  INV_X1 U5708 ( .A(n4639), .ZN(n4641) );
  AOI21_X1 U5709 ( .B1(n5741), .B2(n4641), .A(n4640), .ZN(n4642) );
  AOI211_X1 U5710 ( .C1(n4643), .C2(n6189), .A(n4649), .B(n4642), .ZN(n4644)
         );
  OAI21_X1 U5711 ( .B1(n4654), .B2(n6179), .A(n4644), .ZN(U2986) );
  NOR2_X1 U5712 ( .A1(n4645), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4646)
         );
  OR2_X1 U5713 ( .A1(n4647), .A2(n4646), .ZN(n6080) );
  INV_X1 U5714 ( .A(n6080), .ZN(n4650) );
  AOI211_X1 U5715 ( .C1(n6245), .C2(n4650), .A(n4649), .B(n4648), .ZN(n4653)
         );
  OAI21_X1 U5716 ( .B1(n5828), .B2(n4651), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4652) );
  OAI211_X1 U5717 ( .C1(n4654), .C2(n6208), .A(n4653), .B(n4652), .ZN(U3018)
         );
  NAND2_X1 U5718 ( .A1(n5594), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6496) );
  INV_X1 U5719 ( .A(n5837), .ZN(n5584) );
  INV_X1 U5720 ( .A(n5586), .ZN(n5841) );
  OAI21_X1 U5721 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6524), .A(n5841), 
        .ZN(n5332) );
  INV_X1 U5722 ( .A(n4655), .ZN(n5335) );
  AOI22_X1 U5723 ( .A1(n6312), .A2(n5335), .B1(n5336), .B2(n4656), .ZN(n6497)
         );
  OAI22_X1 U5724 ( .A1(n6497), .A2(n5584), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5334), .ZN(n4657) );
  OAI22_X1 U5725 ( .A1(n5332), .A2(n4657), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5841), .ZN(n4658) );
  OAI21_X1 U5726 ( .B1(n6496), .B2(n5584), .A(n4658), .ZN(U3461) );
  AOI22_X1 U5727 ( .A1(n6152), .A2(UWORD_REG_1__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n4659) );
  NAND2_X1 U5728 ( .A1(n6153), .A2(DATAI_1_), .ZN(n4677) );
  NAND2_X1 U5729 ( .A1(n4659), .A2(n4677), .ZN(U2925) );
  AOI22_X1 U5730 ( .A1(n6152), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6149), .ZN(n4660) );
  NAND2_X1 U5731 ( .A1(n6153), .A2(DATAI_7_), .ZN(n4682) );
  NAND2_X1 U5732 ( .A1(n4660), .A2(n4682), .ZN(U2931) );
  AOI22_X1 U5733 ( .A1(n6152), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n6149), .ZN(n4661) );
  NAND2_X1 U5734 ( .A1(n6153), .A2(DATAI_12_), .ZN(n4675) );
  NAND2_X1 U5735 ( .A1(n4661), .A2(n4675), .ZN(U2936) );
  AOI22_X1 U5736 ( .A1(n6152), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6149), .ZN(n4663) );
  NAND2_X1 U5737 ( .A1(n4663), .A2(n4662), .ZN(U2933) );
  AOI22_X1 U5738 ( .A1(n6152), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6149), .ZN(n4664) );
  NAND2_X1 U5739 ( .A1(n6153), .A2(DATAI_14_), .ZN(n4684) );
  NAND2_X1 U5740 ( .A1(n4664), .A2(n4684), .ZN(U2938) );
  AOI22_X1 U5741 ( .A1(n6152), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6149), .ZN(n4665) );
  NAND2_X1 U5742 ( .A1(n6153), .A2(DATAI_8_), .ZN(n4690) );
  NAND2_X1 U5743 ( .A1(n4665), .A2(n4690), .ZN(U2932) );
  AOI22_X1 U5744 ( .A1(n6152), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6149), .ZN(n4667) );
  NAND2_X1 U5745 ( .A1(n4667), .A2(n4666), .ZN(U2924) );
  INV_X1 U5746 ( .A(DATAI_11_), .ZN(n5267) );
  OR2_X1 U5747 ( .A1(n4669), .A2(n5267), .ZN(n4671) );
  AOI22_X1 U5748 ( .A1(n6152), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n6149), .ZN(n4668) );
  NAND2_X1 U5749 ( .A1(n4671), .A2(n4668), .ZN(U2935) );
  INV_X1 U5750 ( .A(DATAI_13_), .ZN(n5326) );
  OR2_X1 U5751 ( .A1(n4669), .A2(n5326), .ZN(n4695) );
  AOI22_X1 U5752 ( .A1(n6152), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6149), .ZN(n4670) );
  NAND2_X1 U5753 ( .A1(n4695), .A2(n4670), .ZN(U2937) );
  AOI22_X1 U5754 ( .A1(n6152), .A2(LWORD_REG_11__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U5755 ( .A1(n4672), .A2(n4671), .ZN(U2950) );
  AOI22_X1 U5756 ( .A1(n6152), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6149), .ZN(n4674) );
  NAND2_X1 U5757 ( .A1(n4674), .A2(n4673), .ZN(U2942) );
  AOI22_X1 U5758 ( .A1(n6152), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6149), .ZN(n4676) );
  NAND2_X1 U5759 ( .A1(n4676), .A2(n4675), .ZN(U2951) );
  AOI22_X1 U5760 ( .A1(n6152), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6149), .ZN(n4678) );
  NAND2_X1 U5761 ( .A1(n4678), .A2(n4677), .ZN(U2940) );
  AOI22_X1 U5762 ( .A1(n6152), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6149), .ZN(n4679) );
  NAND2_X1 U5763 ( .A1(n6153), .A2(DATAI_6_), .ZN(n4692) );
  NAND2_X1 U5764 ( .A1(n4679), .A2(n4692), .ZN(U2930) );
  AOI22_X1 U5765 ( .A1(n6152), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6149), .ZN(n4680) );
  NAND2_X1 U5766 ( .A1(n4681), .A2(n4680), .ZN(U2943) );
  AOI22_X1 U5767 ( .A1(n6152), .A2(LWORD_REG_7__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U5768 ( .A1(n4683), .A2(n4682), .ZN(U2946) );
  AOI22_X1 U5769 ( .A1(n6152), .A2(LWORD_REG_14__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U5770 ( .A1(n4685), .A2(n4684), .ZN(U2953) );
  AOI22_X1 U5771 ( .A1(n6152), .A2(LWORD_REG_5__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4687) );
  NAND2_X1 U5772 ( .A1(n4687), .A2(n4686), .ZN(U2944) );
  AOI22_X1 U5773 ( .A1(n6152), .A2(LWORD_REG_2__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4689) );
  NAND2_X1 U5774 ( .A1(n4689), .A2(n4688), .ZN(U2941) );
  AOI22_X1 U5775 ( .A1(n6152), .A2(LWORD_REG_8__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4691) );
  NAND2_X1 U5776 ( .A1(n4691), .A2(n4690), .ZN(U2947) );
  AOI22_X1 U5777 ( .A1(n6152), .A2(LWORD_REG_6__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4693) );
  NAND2_X1 U5778 ( .A1(n4693), .A2(n4692), .ZN(U2945) );
  AOI22_X1 U5779 ( .A1(n6152), .A2(LWORD_REG_13__SCAN_IN), .B1(n6149), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n4694) );
  NAND2_X1 U5780 ( .A1(n4695), .A2(n4694), .ZN(U2952) );
  XOR2_X1 U5781 ( .A(n4697), .B(n4696), .Z(n5224) );
  INV_X1 U5782 ( .A(n5224), .ZN(n4707) );
  INV_X1 U5783 ( .A(n4698), .ZN(n4703) );
  INV_X1 U5784 ( .A(n4699), .ZN(n4702) );
  AOI21_X1 U5785 ( .B1(n4703), .B2(n4702), .A(n4701), .ZN(n6064) );
  AOI22_X1 U5786 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6221), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4704) );
  OAI21_X1 U5787 ( .B1(n6193), .B2(n6001), .A(n4704), .ZN(n4705) );
  AOI21_X1 U5788 ( .B1(n6064), .B2(n6189), .A(n4705), .ZN(n4706) );
  OAI21_X1 U5789 ( .B1(n4707), .B2(n6179), .A(n4706), .ZN(U2982) );
  XNOR2_X1 U5790 ( .A(n4709), .B(n4708), .ZN(n4888) );
  INV_X1 U5791 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6556) );
  NOR2_X1 U5792 ( .A1(n6256), .A2(n6556), .ZN(n4885) );
  NOR2_X1 U5793 ( .A1(n4710), .A2(n4711), .ZN(n4712) );
  OR2_X1 U5794 ( .A1(n4699), .A2(n4712), .ZN(n6070) );
  OAI22_X1 U5795 ( .A1(n6193), .A2(n6016), .B1(n6203), .B2(n6070), .ZN(n4713)
         );
  AOI211_X1 U5796 ( .C1(n6194), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4885), 
        .B(n4713), .ZN(n4714) );
  OAI21_X1 U5797 ( .B1(n4888), .B2(n6179), .A(n4714), .ZN(U2983) );
  NAND2_X1 U5798 ( .A1(n6189), .A2(DATAI_27_), .ZN(n6471) );
  OR2_X1 U5799 ( .A1(n6271), .A2(n4715), .ZN(n4757) );
  NOR2_X2 U5800 ( .A1(n5039), .A2(n4717), .ZN(n6467) );
  NAND2_X1 U5801 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4718) );
  NOR2_X2 U5802 ( .A1(n4724), .A2(n6308), .ZN(n5210) );
  INV_X1 U5803 ( .A(DATAI_19_), .ZN(n6963) );
  NOR2_X2 U5804 ( .A1(n6203), .A2(n6963), .ZN(n6468) );
  AOI22_X1 U5805 ( .A1(n6467), .A2(n3292), .B1(n5210), .B2(n6468), .ZN(n4731)
         );
  NAND2_X1 U5806 ( .A1(n5058), .A2(n6312), .ZN(n4968) );
  INV_X1 U5807 ( .A(n4968), .ZN(n4773) );
  INV_X1 U5808 ( .A(n4617), .ZN(n5302) );
  INV_X1 U5809 ( .A(n4721), .ZN(n4927) );
  NAND2_X1 U5810 ( .A1(n5302), .A2(n4927), .ZN(n6444) );
  INV_X1 U5811 ( .A(n6444), .ZN(n5054) );
  AOI21_X1 U5812 ( .B1(n4773), .B2(n5054), .A(n3292), .ZN(n4726) );
  NAND2_X1 U5813 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4722) );
  OAI22_X1 U5814 ( .A1(n4726), .A2(n6617), .B1(n4722), .B2(n6434), .ZN(n5205)
         );
  INV_X1 U5815 ( .A(DATAI_3_), .ZN(n5155) );
  NOR2_X2 U5816 ( .A1(n5155), .A2(n6353), .ZN(n6466) );
  INV_X1 U5817 ( .A(n4724), .ZN(n4725) );
  NAND2_X1 U5818 ( .A1(n4725), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5576) );
  NAND2_X1 U5819 ( .A1(n5576), .A2(n4726), .ZN(n4729) );
  NOR2_X1 U5820 ( .A1(n4948), .A2(n6434), .ZN(n4727) );
  OR2_X1 U5821 ( .A1(n6442), .A2(n4727), .ZN(n4728) );
  OAI21_X1 U5822 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6605), .A(n4867), 
        .ZN(n6400) );
  OAI211_X1 U5823 ( .C1(n4729), .C2(n6617), .A(n4728), .B(n6315), .ZN(n5116)
         );
  AOI22_X1 U5824 ( .A1(n5205), .A2(n6466), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n5116), .ZN(n4730) );
  OAI211_X1 U5825 ( .C1(n6471), .C2(n5212), .A(n4731), .B(n4730), .ZN(U3127)
         );
  NAND2_X1 U5826 ( .A1(n4738), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4733) );
  NAND2_X1 U5827 ( .A1(n4733), .A2(n6442), .ZN(n5061) );
  NOR2_X1 U5828 ( .A1(n6444), .A2(n4894), .ZN(n5062) );
  OR2_X1 U5829 ( .A1(n6434), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5059)
         );
  NOR2_X1 U5830 ( .A1(n6902), .A2(n5059), .ZN(n5196) );
  AOI21_X1 U5831 ( .B1(n5062), .B2(n6312), .A(n5196), .ZN(n4736) );
  OAI22_X1 U5832 ( .A1(n5061), .A2(n4736), .B1(n6403), .B2(n5059), .ZN(n4734)
         );
  INV_X1 U5833 ( .A(n6466), .ZN(n6288) );
  NAND2_X1 U5834 ( .A1(n4738), .A2(n4942), .ZN(n7024) );
  INV_X1 U5835 ( .A(n5061), .ZN(n4735) );
  AOI22_X1 U5836 ( .A1(n4736), .A2(n4735), .B1(n6617), .B2(n5059), .ZN(n4737)
         );
  NAND2_X1 U5837 ( .A1(n6315), .A2(n4737), .ZN(n5194) );
  AOI22_X1 U5838 ( .A1(n5195), .A2(n6468), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n5194), .ZN(n4741) );
  INV_X1 U5839 ( .A(n4738), .ZN(n4739) );
  INV_X1 U5840 ( .A(n6471), .ZN(n6414) );
  AOI22_X1 U5841 ( .A1(n5197), .A2(n6414), .B1(n6467), .B2(n5196), .ZN(n4740)
         );
  OAI211_X1 U5842 ( .C1(n5200), .C2(n6288), .A(n4741), .B(n4740), .ZN(U3063)
         );
  INV_X1 U5843 ( .A(DATAI_7_), .ZN(n6854) );
  NOR2_X2 U5844 ( .A1(n6854), .A2(n6353), .ZN(n7019) );
  INV_X1 U5845 ( .A(n7019), .ZN(n6306) );
  INV_X1 U5846 ( .A(DATAI_23_), .ZN(n4742) );
  NOR2_X2 U5847 ( .A1(n6203), .A2(n4742), .ZN(n7020) );
  AOI22_X1 U5848 ( .A1(n5195), .A2(n7020), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n5194), .ZN(n4745) );
  INV_X1 U5849 ( .A(DATAI_31_), .ZN(n4743) );
  NOR2_X1 U5850 ( .A1(n6203), .A2(n4743), .ZN(n6300) );
  NOR2_X2 U5851 ( .A1(n5039), .A2(n5328), .ZN(n7027) );
  AOI22_X1 U5852 ( .A1(n5197), .A2(n6300), .B1(n7027), .B2(n5196), .ZN(n4744)
         );
  OAI211_X1 U5853 ( .C1(n5200), .C2(n6306), .A(n4745), .B(n4744), .ZN(U3067)
         );
  XNOR2_X1 U5854 ( .A(n4746), .B(n4747), .ZN(n4856) );
  INV_X1 U5855 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4748) );
  NOR2_X1 U5856 ( .A1(n6256), .A2(n4748), .ZN(n4853) );
  NOR2_X1 U5857 ( .A1(n5741), .A2(n6921), .ZN(n4749) );
  AOI211_X1 U5858 ( .C1(n6198), .C2(n5979), .A(n4853), .B(n4749), .ZN(n4755)
         );
  AND2_X1 U5859 ( .A1(n4751), .A2(n4752), .ZN(n4753) );
  OR2_X1 U5860 ( .A1(n4750), .A2(n4753), .ZN(n6061) );
  INV_X1 U5861 ( .A(n6061), .ZN(n5977) );
  NAND2_X1 U5862 ( .A1(n5977), .A2(n6189), .ZN(n4754) );
  OAI211_X1 U5863 ( .C1(n4856), .C2(n6179), .A(n4755), .B(n4754), .ZN(U2980)
         );
  NOR2_X1 U5864 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4756), .ZN(n5120)
         );
  OAI21_X1 U5865 ( .B1(n6347), .B2(n6403), .A(n4867), .ZN(n4819) );
  OR2_X1 U5866 ( .A1(n4762), .A2(n6403), .ZN(n6448) );
  INV_X1 U5867 ( .A(n6448), .ZN(n5065) );
  NOR3_X1 U5868 ( .A1(n4819), .A2(n4948), .A3(n5065), .ZN(n4760) );
  OR2_X1 U5869 ( .A1(n4617), .A2(n4927), .ZN(n4820) );
  NOR2_X2 U5870 ( .A1(n4776), .A2(n4942), .ZN(n5126) );
  OAI21_X1 U5871 ( .B1(n5210), .B2(n5126), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4758) );
  NAND3_X1 U5872 ( .A1(n4820), .A2(n6442), .A3(n4758), .ZN(n4759) );
  OAI211_X1 U5873 ( .C1(n5120), .C2(n6605), .A(n4760), .B(n4759), .ZN(n4761)
         );
  INV_X1 U5874 ( .A(n4820), .ZN(n4772) );
  NAND2_X1 U5875 ( .A1(n4772), .A2(n6442), .ZN(n4826) );
  INV_X1 U5876 ( .A(n5058), .ZN(n6437) );
  AND2_X1 U5877 ( .A1(n4762), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5055) );
  NAND3_X1 U5878 ( .A1(n5055), .A2(n6347), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4763) );
  OAI21_X1 U5879 ( .B1(n4826), .B2(n6437), .A(n4763), .ZN(n5119) );
  AOI22_X1 U5880 ( .A1(n5210), .A2(n6300), .B1(n7019), .B2(n5119), .ZN(n4765)
         );
  AOI22_X1 U5881 ( .A1(n7027), .A2(n5120), .B1(n5126), .B2(n7020), .ZN(n4764)
         );
  OAI211_X1 U5882 ( .C1(n5124), .C2(n4766), .A(n4765), .B(n4764), .ZN(U3139)
         );
  AOI22_X1 U5883 ( .A1(n5210), .A2(n6414), .B1(n6466), .B2(n5119), .ZN(n4768)
         );
  AOI22_X1 U5884 ( .A1(n6467), .A2(n5120), .B1(n5126), .B2(n6468), .ZN(n4767)
         );
  OAI211_X1 U5885 ( .C1(n5124), .C2(n4769), .A(n4768), .B(n4767), .ZN(U3135)
         );
  INV_X1 U5886 ( .A(n4776), .ZN(n4770) );
  AND2_X1 U5887 ( .A1(n6442), .A2(n4392), .ZN(n4863) );
  INV_X1 U5888 ( .A(n4863), .ZN(n6351) );
  OAI21_X1 U5889 ( .B1(n4770), .B2(n6203), .A(n6351), .ZN(n4775) );
  INV_X1 U5890 ( .A(n4771), .ZN(n5127) );
  AOI21_X1 U5891 ( .B1(n4773), .B2(n4772), .A(n5127), .ZN(n4777) );
  OAI21_X1 U5892 ( .B1(n6442), .B2(n4779), .A(n6315), .ZN(n4774) );
  NOR2_X2 U5893 ( .A1(n4776), .A2(n6308), .ZN(n5241) );
  INV_X1 U5894 ( .A(n4777), .ZN(n4778) );
  NAND2_X1 U5895 ( .A1(n4778), .A2(n6442), .ZN(n4781) );
  NAND2_X1 U5896 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4779), .ZN(n4780) );
  NAND2_X1 U5897 ( .A1(n4781), .A2(n4780), .ZN(n5125) );
  AOI22_X1 U5898 ( .A1(n5241), .A2(n7020), .B1(n7019), .B2(n5125), .ZN(n4783)
         );
  AOI22_X1 U5899 ( .A1(n7027), .A2(n5127), .B1(n5126), .B2(n6300), .ZN(n4782)
         );
  OAI211_X1 U5900 ( .C1(n5131), .C2(n4784), .A(n4783), .B(n4782), .ZN(U3147)
         );
  INV_X1 U5901 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4787) );
  AOI22_X1 U5902 ( .A1(n5241), .A2(n6468), .B1(n6466), .B2(n5125), .ZN(n4786)
         );
  AOI22_X1 U5903 ( .A1(n6467), .A2(n5127), .B1(n5126), .B2(n6414), .ZN(n4785)
         );
  OAI211_X1 U5904 ( .C1(n5131), .C2(n4787), .A(n4786), .B(n4785), .ZN(U3143)
         );
  XNOR2_X1 U5905 ( .A(n4789), .B(n4788), .ZN(n6180) );
  NOR2_X1 U5906 ( .A1(n4849), .A2(n4848), .ZN(n4792) );
  NAND2_X1 U5907 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4791) );
  INV_X1 U5908 ( .A(n6262), .ZN(n4790) );
  AOI22_X1 U5909 ( .A1(n5558), .A2(n4791), .B1(n6243), .B2(n4790), .ZN(n6253)
         );
  OAI21_X1 U5910 ( .B1(n5804), .B2(n4792), .A(n6253), .ZN(n4852) );
  NOR2_X1 U5911 ( .A1(n3536), .A2(n4793), .ZN(n6250) );
  NAND2_X1 U5912 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6250), .ZN(n4850)
         );
  INV_X1 U5913 ( .A(n4794), .ZN(n4795) );
  OAI211_X1 U5914 ( .C1(n5220), .C2(n4850), .A(n4849), .B(n4795), .ZN(n4798)
         );
  OAI21_X1 U5915 ( .B1(n5215), .B2(n4796), .A(n5962), .ZN(n5982) );
  NOR2_X1 U5916 ( .A1(n5982), .A2(n6258), .ZN(n4797) );
  NOR2_X1 U5917 ( .A1(n6256), .A2(n6559), .ZN(n6182) );
  AOI211_X1 U5918 ( .C1(n4852), .C2(n4798), .A(n4797), .B(n6182), .ZN(n4799)
         );
  OAI21_X1 U5919 ( .B1(n6208), .B2(n6180), .A(n4799), .ZN(U3013) );
  NOR2_X1 U5920 ( .A1(n5055), .A2(n4819), .ZN(n4945) );
  INV_X1 U5921 ( .A(n6271), .ZN(n4800) );
  INV_X1 U5922 ( .A(n6396), .ZN(n4802) );
  AND2_X1 U5923 ( .A1(n6390), .A2(n6308), .ZN(n4801) );
  NAND2_X1 U5924 ( .A1(n5282), .A2(n6432), .ZN(n4803) );
  NAND2_X1 U5925 ( .A1(n4803), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4804) );
  NAND2_X1 U5926 ( .A1(n4804), .A2(n6442), .ZN(n4810) );
  AND2_X1 U5927 ( .A1(n4617), .A2(n4721), .ZN(n4943) );
  NAND2_X1 U5928 ( .A1(n4943), .A2(n5058), .ZN(n6397) );
  INV_X1 U5929 ( .A(n6397), .ZN(n4805) );
  NAND2_X1 U5930 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4940), .ZN(n6404) );
  NOR2_X1 U5931 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6404), .ZN(n5280)
         );
  OAI22_X1 U5932 ( .A1(n4810), .A2(n4805), .B1(n5280), .B2(n6605), .ZN(n4806)
         );
  INV_X1 U5933 ( .A(n4806), .ZN(n4807) );
  OAI211_X1 U5934 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6403), .A(n4945), .B(n4807), .ZN(n4808) );
  NAND3_X1 U5935 ( .A1(n5065), .A2(n6347), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4809) );
  OAI21_X1 U5936 ( .B1(n4810), .B2(n6397), .A(n4809), .ZN(n5284) );
  INV_X1 U5937 ( .A(n6300), .ZN(n7023) );
  AOI22_X1 U5938 ( .A1(n6421), .A2(n7020), .B1(n7027), .B2(n5280), .ZN(n4811)
         );
  OAI21_X1 U5939 ( .B1(n5282), .B2(n7023), .A(n4811), .ZN(n4812) );
  AOI21_X1 U5940 ( .B1(n5284), .B2(n7019), .A(n4812), .ZN(n4813) );
  OAI21_X1 U5941 ( .B1(n5287), .B2(n4814), .A(n4813), .ZN(U3107) );
  INV_X1 U5942 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4818) );
  AOI22_X1 U5943 ( .A1(n6421), .A2(n6468), .B1(n6467), .B2(n5280), .ZN(n4815)
         );
  OAI21_X1 U5944 ( .B1(n5282), .B2(n6471), .A(n4815), .ZN(n4816) );
  AOI21_X1 U5945 ( .B1(n5284), .B2(n6466), .A(n4816), .ZN(n4817) );
  OAI21_X1 U5946 ( .B1(n5287), .B2(n4818), .A(n4817), .ZN(U3103) );
  NOR2_X1 U5947 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6318), .ZN(n7026)
         );
  NOR3_X1 U5948 ( .A1(n4819), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5065), 
        .ZN(n4823) );
  AOI21_X1 U5949 ( .B1(n7024), .B2(n6343), .A(n4392), .ZN(n4821) );
  NOR2_X1 U5950 ( .A1(n4820), .A2(n4894), .ZN(n6313) );
  OR3_X1 U5951 ( .A1(n4821), .A2(n6313), .A3(n6617), .ZN(n4822) );
  OAI211_X1 U5952 ( .C1(n7026), .C2(n6605), .A(n4823), .B(n4822), .ZN(n4824)
         );
  NAND3_X1 U5953 ( .A1(n5055), .A2(n6347), .A3(n4948), .ZN(n4825) );
  OAI21_X1 U5954 ( .B1(n4826), .B2(n5058), .A(n4825), .ZN(n7018) );
  AOI22_X1 U5955 ( .A1(n7021), .A2(n6468), .B1(n6466), .B2(n7018), .ZN(n4827)
         );
  OAI21_X1 U5956 ( .B1(n7024), .B2(n6471), .A(n4827), .ZN(n4828) );
  AOI21_X1 U5957 ( .B1(n6467), .B2(n7026), .A(n4828), .ZN(n4829) );
  OAI21_X1 U5958 ( .B1(n7030), .B2(n4830), .A(n4829), .ZN(U3071) );
  INV_X1 U5959 ( .A(n7027), .ZN(n4976) );
  NAND3_X1 U5960 ( .A1(n4948), .A2(n6506), .A3(n6500), .ZN(n4865) );
  NOR2_X1 U5961 ( .A1(n6902), .A2(n4865), .ZN(n4831) );
  INV_X1 U5962 ( .A(n4831), .ZN(n5046) );
  NAND2_X1 U5963 ( .A1(n4617), .A2(n4927), .ZN(n6345) );
  OR2_X1 U5964 ( .A1(n6345), .A2(n5058), .ZN(n4872) );
  INV_X1 U5965 ( .A(n4872), .ZN(n4832) );
  AOI21_X1 U5966 ( .B1(n4832), .B2(n6312), .A(n4831), .ZN(n4837) );
  INV_X1 U5967 ( .A(n4941), .ZN(n4833) );
  INV_X1 U5968 ( .A(n4839), .ZN(n4834) );
  AOI21_X1 U5969 ( .B1(n4834), .B2(STATEBS16_REG_SCAN_IN), .A(n6617), .ZN(
        n4836) );
  AOI22_X1 U5970 ( .A1(n4837), .A2(n4836), .B1(n6617), .B2(n4865), .ZN(n4835)
         );
  NAND2_X1 U5971 ( .A1(n6315), .A2(n4835), .ZN(n5041) );
  INV_X1 U5972 ( .A(n4836), .ZN(n4838) );
  OAI22_X1 U5973 ( .A1(n4838), .A2(n4837), .B1(n6403), .B2(n4865), .ZN(n5040)
         );
  AOI22_X1 U5974 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5041), .B1(n7019), 
        .B2(n5040), .ZN(n4841) );
  NOR2_X2 U5975 ( .A1(n4839), .A2(n6308), .ZN(n5234) );
  AOI22_X1 U5976 ( .A1(n6300), .A2(n5243), .B1(n5234), .B2(n7020), .ZN(n4840)
         );
  OAI211_X1 U5977 ( .C1(n4976), .C2(n5046), .A(n4841), .B(n4840), .ZN(U3035)
         );
  INV_X1 U5978 ( .A(n6467), .ZN(n4979) );
  AOI22_X1 U5979 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5041), .B1(n6466), 
        .B2(n5040), .ZN(n4843) );
  AOI22_X1 U5980 ( .A1(n6414), .A2(n5243), .B1(n5234), .B2(n6468), .ZN(n4842)
         );
  OAI211_X1 U5981 ( .C1(n4979), .C2(n5046), .A(n4843), .B(n4842), .ZN(U3031)
         );
  INV_X1 U5982 ( .A(n5116), .ZN(n5208) );
  INV_X1 U5983 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4845) );
  AOI22_X1 U5984 ( .A1(n7027), .A2(n3292), .B1(n7019), .B2(n5205), .ZN(n4844)
         );
  OAI21_X1 U5985 ( .B1(n5208), .B2(n4845), .A(n4844), .ZN(n4846) );
  AOI21_X1 U5986 ( .B1(n5210), .B2(n7020), .A(n4846), .ZN(n4847) );
  OAI21_X1 U5987 ( .B1(n5212), .B2(n7023), .A(n4847), .ZN(U3131) );
  NOR3_X1 U5988 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4849), .A3(n4848), 
        .ZN(n4851) );
  NAND2_X1 U5989 ( .A1(n6243), .A2(n4850), .ZN(n4879) );
  AOI22_X1 U5990 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4852), .B1(n4851), 
        .B2(n4879), .ZN(n4855) );
  XOR2_X1 U5991 ( .A(n5961), .B(n5962), .Z(n6059) );
  AOI21_X1 U5992 ( .B1(n6059), .B2(n6245), .A(n4853), .ZN(n4854) );
  OAI211_X1 U5993 ( .C1(n6208), .C2(n4856), .A(n4855), .B(n4854), .ZN(U3012)
         );
  INV_X1 U5994 ( .A(n6064), .ZN(n4862) );
  NAND2_X1 U5995 ( .A1(n4858), .A2(n4857), .ZN(n4859) );
  INV_X1 U5996 ( .A(n4859), .ZN(n4860) );
  INV_X1 U5997 ( .A(n5406), .ZN(n5401) );
  AOI22_X1 U5998 ( .A1(n5401), .A2(DATAI_4_), .B1(n6089), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4861) );
  OAI21_X1 U5999 ( .B1(n4862), .B2(n5407), .A(n4861), .ZN(U2887) );
  NOR3_X1 U6000 ( .A1(n5243), .A2(n5241), .A3(n6617), .ZN(n4864) );
  OAI21_X1 U6001 ( .B1(n4864), .B2(n4863), .A(n4872), .ZN(n4870) );
  NOR2_X1 U6002 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4865), .ZN(n5242)
         );
  INV_X1 U6003 ( .A(n5242), .ZN(n4868) );
  INV_X1 U6004 ( .A(n6347), .ZN(n4866) );
  AND2_X1 U6005 ( .A1(n4866), .A2(n6346), .ZN(n5056) );
  OAI21_X1 U6006 ( .B1(n5056), .B2(n6403), .A(n4867), .ZN(n5063) );
  AOI211_X1 U6007 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4868), .A(n5055), .B(
        n5063), .ZN(n4869) );
  INV_X1 U6008 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U6009 ( .A1(n5056), .A2(n5065), .ZN(n4871) );
  OAI21_X1 U6010 ( .B1(n4872), .B2(n6617), .A(n4871), .ZN(n5240) );
  AOI22_X1 U6011 ( .A1(n5241), .A2(n6414), .B1(n6466), .B2(n5240), .ZN(n4874)
         );
  AOI22_X1 U6012 ( .A1(n5243), .A2(n6468), .B1(n6467), .B2(n5242), .ZN(n4873)
         );
  OAI211_X1 U6013 ( .C1(n5247), .C2(n4875), .A(n4874), .B(n4873), .ZN(U3023)
         );
  INV_X1 U6014 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4878) );
  AOI22_X1 U6015 ( .A1(n5241), .A2(n6300), .B1(n7019), .B2(n5240), .ZN(n4877)
         );
  AOI22_X1 U6016 ( .A1(n7020), .A2(n5243), .B1(n7027), .B2(n5242), .ZN(n4876)
         );
  OAI211_X1 U6017 ( .C1(n5247), .C2(n4878), .A(n4877), .B(n4876), .ZN(U3027)
         );
  OAI21_X1 U6018 ( .B1(n6243), .B2(n6239), .A(n6253), .ZN(n5217) );
  NAND2_X1 U6019 ( .A1(n6239), .A2(n4879), .ZN(n5102) );
  INV_X1 U6020 ( .A(n5102), .ZN(n5219) );
  AOI22_X1 U6021 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n5217), .B1(n5219), 
        .B2(n4880), .ZN(n4887) );
  INV_X1 U6022 ( .A(n5301), .ZN(n4882) );
  AOI21_X1 U6023 ( .B1(n4882), .B2(n5300), .A(n4881), .ZN(n4884) );
  INV_X1 U6024 ( .A(n5214), .ZN(n4883) );
  NOR2_X1 U6025 ( .A1(n4884), .A2(n4883), .ZN(n6067) );
  AOI21_X1 U6026 ( .B1(n6067), .B2(n6245), .A(n4885), .ZN(n4886) );
  OAI211_X1 U6027 ( .C1(n6208), .C2(n4888), .A(n4887), .B(n4886), .ZN(U3015)
         );
  NOR2_X2 U6028 ( .A1(n5039), .A2(n3438), .ZN(n6460) );
  INV_X1 U6029 ( .A(n6460), .ZN(n4893) );
  INV_X1 U6030 ( .A(DATAI_2_), .ZN(n5153) );
  NOR2_X2 U6031 ( .A1(n5153), .A2(n6353), .ZN(n6461) );
  AOI22_X1 U6032 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5041), .B1(n6461), 
        .B2(n5040), .ZN(n4892) );
  INV_X1 U6033 ( .A(DATAI_26_), .ZN(n4889) );
  NOR2_X1 U6034 ( .A1(n6203), .A2(n4889), .ZN(n6382) );
  INV_X1 U6035 ( .A(DATAI_18_), .ZN(n4890) );
  NOR2_X2 U6036 ( .A1(n6203), .A2(n4890), .ZN(n6462) );
  AOI22_X1 U6037 ( .A1(n6382), .A2(n5243), .B1(n5234), .B2(n6462), .ZN(n4891)
         );
  OAI211_X1 U6038 ( .C1(n4893), .C2(n5046), .A(n4892), .B(n4891), .ZN(U3030)
         );
  INV_X1 U6039 ( .A(n4894), .ZN(n6445) );
  NOR2_X1 U6040 ( .A1(n4895), .A2(n6445), .ZN(n4896) );
  XOR2_X1 U6041 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n4896), .Z(n6006) );
  AOI22_X1 U6042 ( .A1(n6006), .A2(n5838), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4897), .ZN(n4898) );
  NAND2_X1 U6043 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5849), .ZN(n4919) );
  OAI22_X1 U6044 ( .A1(n4898), .A2(STATE2_REG_1__SCAN_IN), .B1(n4919), .B2(
        n5840), .ZN(n4899) );
  INV_X1 U6045 ( .A(n4899), .ZN(n4922) );
  INV_X1 U6046 ( .A(n4900), .ZN(n4918) );
  MUX2_X1 U6047 ( .A(n4901), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4600), 
        .Z(n4902) );
  NOR2_X1 U6048 ( .A1(n4902), .A2(n4900), .ZN(n4903) );
  NAND2_X1 U6049 ( .A1(n4904), .A2(n4903), .ZN(n4913) );
  NAND2_X1 U6050 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4905) );
  XNOR2_X1 U6051 ( .A(n4905), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4911)
         );
  INV_X1 U6052 ( .A(n4906), .ZN(n4907) );
  OAI21_X1 U6053 ( .B1(n4600), .B2(n3750), .A(n4907), .ZN(n4908) );
  NOR2_X1 U6054 ( .A1(n4908), .A2(n3210), .ZN(n5583) );
  NOR2_X1 U6055 ( .A1(n4909), .A2(n5583), .ZN(n4910) );
  AOI21_X1 U6056 ( .B1(n5594), .B2(n4911), .A(n4910), .ZN(n4912) );
  NAND2_X1 U6057 ( .A1(n4913), .A2(n4912), .ZN(n4914) );
  AOI21_X1 U6058 ( .B1(n5058), .B2(n5335), .A(n4914), .ZN(n5585) );
  MUX2_X1 U6059 ( .A(n3750), .B(n5585), .S(n6498), .Z(n6507) );
  INV_X1 U6060 ( .A(n6507), .ZN(n4916) );
  MUX2_X1 U6061 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4915), .S(n6498), 
        .Z(n6505) );
  NAND3_X1 U6062 ( .A1(n4916), .A2(n6505), .A3(n5334), .ZN(n4917) );
  OAI211_X1 U6063 ( .C1(n4919), .C2(n4918), .A(n4922), .B(n4917), .ZN(n6514)
         );
  INV_X1 U6064 ( .A(n6514), .ZN(n4920) );
  AOI21_X1 U6065 ( .B1(n4922), .B2(n4921), .A(n4920), .ZN(n4924) );
  NOR2_X1 U6066 ( .A1(n4924), .A2(FLUSH_REG_SCAN_IN), .ZN(n4923) );
  NOR2_X1 U6067 ( .A1(n4924), .A2(n5592), .ZN(n6522) );
  AND2_X1 U6068 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6605), .ZN(n5580) );
  OAI22_X1 U6069 ( .A1(n6308), .A2(n6617), .B1(n3982), .B2(n5580), .ZN(n4925)
         );
  OAI21_X1 U6070 ( .B1(n6522), .B2(n4925), .A(n6264), .ZN(n4926) );
  OAI21_X1 U6071 ( .B1(n6264), .B2(n6902), .A(n4926), .ZN(U3465) );
  NAND2_X1 U6072 ( .A1(n6390), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6395) );
  INV_X1 U6073 ( .A(n6395), .ZN(n6272) );
  AOI211_X1 U6074 ( .C1(n6309), .C2(n4392), .A(n6617), .B(n6272), .ZN(n4929)
         );
  NOR2_X1 U6075 ( .A1(n4927), .A2(n5580), .ZN(n4928) );
  OAI21_X1 U6076 ( .B1(n4929), .B2(n4928), .A(n6264), .ZN(n4930) );
  OAI21_X1 U6077 ( .B1(n6264), .B2(n6500), .A(n4930), .ZN(U3464) );
  NOR2_X2 U6078 ( .A1(n5039), .A2(n6092), .ZN(n6440) );
  INV_X1 U6079 ( .A(n6440), .ZN(n4935) );
  INV_X1 U6080 ( .A(DATAI_0_), .ZN(n5154) );
  NOR2_X2 U6081 ( .A1(n5154), .A2(n6353), .ZN(n6439) );
  AOI22_X1 U6082 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5041), .B1(n6439), 
        .B2(n5040), .ZN(n4934) );
  INV_X1 U6083 ( .A(DATAI_24_), .ZN(n4931) );
  INV_X1 U6084 ( .A(DATAI_16_), .ZN(n4932) );
  NOR2_X2 U6085 ( .A1(n6203), .A2(n4932), .ZN(n6451) );
  AOI22_X1 U6086 ( .A1(n6394), .A2(n5243), .B1(n5234), .B2(n6451), .ZN(n4933)
         );
  OAI211_X1 U6087 ( .C1(n4935), .C2(n5046), .A(n4934), .B(n4933), .ZN(U3028)
         );
  INV_X1 U6088 ( .A(n6382), .ZN(n6465) );
  AOI22_X1 U6089 ( .A1(n7021), .A2(n6462), .B1(n6461), .B2(n7018), .ZN(n4936)
         );
  OAI21_X1 U6090 ( .B1(n7024), .B2(n6465), .A(n4936), .ZN(n4937) );
  AOI21_X1 U6091 ( .B1(n6460), .B2(n7026), .A(n4937), .ZN(n4938) );
  OAI21_X1 U6092 ( .B1(n7030), .B2(n4939), .A(n4938), .ZN(U3070) );
  NAND2_X1 U6093 ( .A1(n4940), .A2(n4948), .ZN(n6266) );
  NOR2_X1 U6094 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6266), .ZN(n5235)
         );
  NOR2_X2 U6095 ( .A1(n5060), .A2(n4942), .ZN(n6301) );
  OAI21_X1 U6096 ( .B1(n6301), .B2(n5234), .A(n6351), .ZN(n4944) );
  NAND2_X1 U6097 ( .A1(n6437), .A2(n4943), .ZN(n6267) );
  AOI21_X1 U6098 ( .B1(n4944), .B2(n6267), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4946) );
  OAI21_X1 U6099 ( .B1(n5235), .B2(n4946), .A(n4945), .ZN(n4947) );
  INV_X1 U6100 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4952) );
  NAND3_X1 U6101 ( .A1(n5065), .A2(n6347), .A3(n4948), .ZN(n4949) );
  OAI21_X1 U6102 ( .B1(n6267), .B2(n6617), .A(n4949), .ZN(n5233) );
  AOI22_X1 U6103 ( .A1(n5234), .A2(n6414), .B1(n6466), .B2(n5233), .ZN(n4951)
         );
  AOI22_X1 U6104 ( .A1(n6301), .A2(n6468), .B1(n6467), .B2(n5235), .ZN(n4950)
         );
  OAI211_X1 U6105 ( .C1(n5239), .C2(n4952), .A(n4951), .B(n4950), .ZN(U3039)
         );
  AOI22_X1 U6106 ( .A1(n5234), .A2(n6300), .B1(n7019), .B2(n5233), .ZN(n4954)
         );
  AOI22_X1 U6107 ( .A1(n6301), .A2(n7020), .B1(n7027), .B2(n5235), .ZN(n4953)
         );
  OAI211_X1 U6108 ( .C1(n5239), .C2(n4955), .A(n4954), .B(n4953), .ZN(U3043)
         );
  INV_X1 U6109 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4959) );
  INV_X1 U6110 ( .A(n6394), .ZN(n6454) );
  AOI22_X1 U6111 ( .A1(n7021), .A2(n6451), .B1(n6439), .B2(n7018), .ZN(n4956)
         );
  OAI21_X1 U6112 ( .B1(n7024), .B2(n6454), .A(n4956), .ZN(n4957) );
  AOI21_X1 U6113 ( .B1(n6440), .B2(n7026), .A(n4957), .ZN(n4958) );
  OAI21_X1 U6114 ( .B1(n7030), .B2(n4959), .A(n4958), .ZN(U3068) );
  INV_X1 U6115 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4962) );
  AOI22_X1 U6116 ( .A1(n5241), .A2(n6462), .B1(n6461), .B2(n5125), .ZN(n4961)
         );
  AOI22_X1 U6117 ( .A1(n6460), .A2(n5127), .B1(n5126), .B2(n6382), .ZN(n4960)
         );
  OAI211_X1 U6118 ( .C1(n5131), .C2(n4962), .A(n4961), .B(n4960), .ZN(U3142)
         );
  INV_X1 U6119 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U6120 ( .A1(n5210), .A2(n6382), .B1(n6461), .B2(n5119), .ZN(n4964)
         );
  AOI22_X1 U6121 ( .A1(n6460), .A2(n5120), .B1(n5126), .B2(n6462), .ZN(n4963)
         );
  OAI211_X1 U6122 ( .C1(n5124), .C2(n4965), .A(n4964), .B(n4963), .ZN(U3134)
         );
  NAND3_X1 U6123 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6506), .A3(n6500), .ZN(n6344) );
  NOR2_X1 U6124 ( .A1(n6902), .A2(n6344), .ZN(n6381) );
  INV_X1 U6125 ( .A(n6381), .ZN(n5024) );
  NOR2_X1 U6126 ( .A1(n6396), .A2(n6390), .ZN(n4966) );
  NAND2_X1 U6127 ( .A1(n4966), .A2(n6308), .ZN(n6349) );
  AOI22_X1 U6128 ( .A1(n6384), .A2(n7020), .B1(n6383), .B2(n6300), .ZN(n4975)
         );
  INV_X1 U6129 ( .A(n4966), .ZN(n4967) );
  OAI21_X1 U6130 ( .B1(n4967), .B2(n4392), .A(n6442), .ZN(n4973) );
  OR2_X1 U6131 ( .A1(n4968), .A2(n6345), .ZN(n4969) );
  NAND2_X1 U6132 ( .A1(n4969), .A2(n5024), .ZN(n4971) );
  OAI21_X1 U6133 ( .B1(n4973), .B2(n4971), .A(n6315), .ZN(n4970) );
  AOI21_X1 U6134 ( .B1(n6617), .B2(n6344), .A(n4970), .ZN(n6389) );
  INV_X1 U6135 ( .A(n6389), .ZN(n5021) );
  INV_X1 U6136 ( .A(n4971), .ZN(n4972) );
  OAI22_X1 U6137 ( .A1(n4973), .A2(n4972), .B1(n6344), .B2(n6403), .ZN(n6385)
         );
  AOI22_X1 U6138 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5021), .B1(n7019), 
        .B2(n6385), .ZN(n4974) );
  OAI211_X1 U6139 ( .C1(n4976), .C2(n5024), .A(n4975), .B(n4974), .ZN(U3099)
         );
  AOI22_X1 U6140 ( .A1(n6384), .A2(n6468), .B1(n6383), .B2(n6414), .ZN(n4978)
         );
  AOI22_X1 U6141 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5021), .B1(n6466), 
        .B2(n6385), .ZN(n4977) );
  OAI211_X1 U6142 ( .C1(n4979), .C2(n5024), .A(n4978), .B(n4977), .ZN(U3095)
         );
  INV_X1 U6143 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4982) );
  AOI22_X1 U6144 ( .A1(n5241), .A2(n6451), .B1(n6439), .B2(n5125), .ZN(n4981)
         );
  AOI22_X1 U6145 ( .A1(n6440), .A2(n5127), .B1(n5126), .B2(n6394), .ZN(n4980)
         );
  OAI211_X1 U6146 ( .C1(n5131), .C2(n4982), .A(n4981), .B(n4980), .ZN(U3140)
         );
  INV_X1 U6147 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4985) );
  AOI22_X1 U6148 ( .A1(n5210), .A2(n6394), .B1(n6439), .B2(n5119), .ZN(n4984)
         );
  AOI22_X1 U6149 ( .A1(n6440), .A2(n5120), .B1(n5126), .B2(n6451), .ZN(n4983)
         );
  OAI211_X1 U6150 ( .C1(n5124), .C2(n4985), .A(n4984), .B(n4983), .ZN(U3132)
         );
  INV_X1 U6151 ( .A(n6461), .ZN(n6285) );
  AOI22_X1 U6152 ( .A1(n5195), .A2(n6462), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n5194), .ZN(n4987) );
  AOI22_X1 U6153 ( .A1(n5197), .A2(n6382), .B1(n6460), .B2(n5196), .ZN(n4986)
         );
  OAI211_X1 U6154 ( .C1(n5200), .C2(n6285), .A(n4987), .B(n4986), .ZN(U3062)
         );
  INV_X1 U6155 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4992) );
  NOR2_X2 U6156 ( .A1(n5039), .A2(n4988), .ZN(n6484) );
  NAND2_X1 U6157 ( .A1(n6189), .A2(DATAI_30_), .ZN(n6488) );
  INV_X1 U6158 ( .A(DATAI_22_), .ZN(n6875) );
  NOR2_X2 U6159 ( .A1(n6203), .A2(n6875), .ZN(n6485) );
  INV_X1 U6160 ( .A(DATAI_6_), .ZN(n5149) );
  NOR2_X2 U6161 ( .A1(n5149), .A2(n6353), .ZN(n6483) );
  AOI22_X1 U6162 ( .A1(n7021), .A2(n6485), .B1(n6483), .B2(n7018), .ZN(n4989)
         );
  OAI21_X1 U6163 ( .B1(n7024), .B2(n6488), .A(n4989), .ZN(n4990) );
  AOI21_X1 U6164 ( .B1(n6484), .B2(n7026), .A(n4990), .ZN(n4991) );
  OAI21_X1 U6165 ( .B1(n7030), .B2(n4992), .A(n4991), .ZN(U3074) );
  NOR2_X2 U6166 ( .A1(n5039), .A2(n4993), .ZN(n6478) );
  NAND2_X1 U6167 ( .A1(n6189), .A2(DATAI_29_), .ZN(n6482) );
  INV_X1 U6168 ( .A(DATAI_21_), .ZN(n4994) );
  NOR2_X2 U6169 ( .A1(n6203), .A2(n4994), .ZN(n6479) );
  INV_X1 U6170 ( .A(DATAI_5_), .ZN(n5142) );
  NOR2_X2 U6171 ( .A1(n5142), .A2(n6353), .ZN(n6477) );
  AOI22_X1 U6172 ( .A1(n7021), .A2(n6479), .B1(n6477), .B2(n7018), .ZN(n4995)
         );
  OAI21_X1 U6173 ( .B1(n7024), .B2(n6482), .A(n4995), .ZN(n4996) );
  AOI21_X1 U6174 ( .B1(n6478), .B2(n7026), .A(n4996), .ZN(n4997) );
  OAI21_X1 U6175 ( .B1(n7030), .B2(n4998), .A(n4997), .ZN(U3073) );
  NOR2_X2 U6176 ( .A1(n5039), .A2(n4999), .ZN(n6473) );
  NAND2_X1 U6177 ( .A1(n6189), .A2(DATAI_28_), .ZN(n6476) );
  INV_X1 U6178 ( .A(DATAI_20_), .ZN(n5000) );
  NOR2_X2 U6179 ( .A1(n5002), .A2(n6353), .ZN(n6472) );
  AOI22_X1 U6180 ( .A1(n7021), .A2(n5001), .B1(n6472), .B2(n7018), .ZN(n5003)
         );
  OAI21_X1 U6181 ( .B1(n7024), .B2(n6476), .A(n5003), .ZN(n5004) );
  AOI21_X1 U6182 ( .B1(n6473), .B2(n7026), .A(n5004), .ZN(n5005) );
  OAI21_X1 U6183 ( .B1(n7030), .B2(n5006), .A(n5005), .ZN(U3072) );
  INV_X1 U6184 ( .A(n6439), .ZN(n6279) );
  AOI22_X1 U6185 ( .A1(n5195), .A2(n6451), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n5194), .ZN(n5008) );
  AOI22_X1 U6186 ( .A1(n5197), .A2(n6394), .B1(n6440), .B2(n5196), .ZN(n5007)
         );
  OAI211_X1 U6187 ( .C1(n5200), .C2(n6279), .A(n5008), .B(n5007), .ZN(U3060)
         );
  INV_X1 U6188 ( .A(n6473), .ZN(n5020) );
  AOI22_X1 U6189 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5041), .B1(n6472), 
        .B2(n5040), .ZN(n5010) );
  INV_X1 U6190 ( .A(n6476), .ZN(n6289) );
  AOI22_X1 U6191 ( .A1(n6289), .A2(n5243), .B1(n5234), .B2(n5001), .ZN(n5009)
         );
  OAI211_X1 U6192 ( .C1(n5020), .C2(n5046), .A(n5010), .B(n5009), .ZN(U3032)
         );
  INV_X1 U6193 ( .A(n6478), .ZN(n5017) );
  AOI22_X1 U6194 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5041), .B1(n6477), 
        .B2(n5040), .ZN(n5012) );
  INV_X1 U6195 ( .A(n6482), .ZN(n6420) );
  AOI22_X1 U6196 ( .A1(n6420), .A2(n5243), .B1(n5234), .B2(n6479), .ZN(n5011)
         );
  OAI211_X1 U6197 ( .C1(n5017), .C2(n5046), .A(n5012), .B(n5011), .ZN(U3033)
         );
  INV_X1 U6198 ( .A(n6484), .ZN(n5025) );
  AOI22_X1 U6199 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5041), .B1(n6483), 
        .B2(n5040), .ZN(n5014) );
  INV_X1 U6200 ( .A(n6488), .ZN(n6333) );
  AOI22_X1 U6201 ( .A1(n6333), .A2(n5243), .B1(n5234), .B2(n6485), .ZN(n5013)
         );
  OAI211_X1 U6202 ( .C1(n5025), .C2(n5046), .A(n5014), .B(n5013), .ZN(U3034)
         );
  AOI22_X1 U6203 ( .A1(n6384), .A2(n6479), .B1(n6383), .B2(n6420), .ZN(n5016)
         );
  AOI22_X1 U6204 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5021), .B1(n6477), 
        .B2(n6385), .ZN(n5015) );
  OAI211_X1 U6205 ( .C1(n5017), .C2(n5024), .A(n5016), .B(n5015), .ZN(U3097)
         );
  AOI22_X1 U6206 ( .A1(n6384), .A2(n5001), .B1(n6383), .B2(n6289), .ZN(n5019)
         );
  AOI22_X1 U6207 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5021), .B1(n6472), 
        .B2(n6385), .ZN(n5018) );
  OAI211_X1 U6208 ( .C1(n5020), .C2(n5024), .A(n5019), .B(n5018), .ZN(U3096)
         );
  AOI22_X1 U6209 ( .A1(n6384), .A2(n6485), .B1(n6383), .B2(n6333), .ZN(n5023)
         );
  AOI22_X1 U6210 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5021), .B1(n6483), 
        .B2(n6385), .ZN(n5022) );
  OAI211_X1 U6211 ( .C1(n5025), .C2(n5024), .A(n5023), .B(n5022), .ZN(U3098)
         );
  INV_X1 U6212 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5028) );
  AOI22_X1 U6213 ( .A1(n5234), .A2(n6382), .B1(n6461), .B2(n5233), .ZN(n5027)
         );
  AOI22_X1 U6214 ( .A1(n6301), .A2(n6462), .B1(n6460), .B2(n5235), .ZN(n5026)
         );
  OAI211_X1 U6215 ( .C1(n5239), .C2(n5028), .A(n5027), .B(n5026), .ZN(U3038)
         );
  INV_X1 U6216 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6217 ( .A1(n5241), .A2(n6382), .B1(n6461), .B2(n5240), .ZN(n5030)
         );
  AOI22_X1 U6218 ( .A1(n6462), .A2(n5243), .B1(n6460), .B2(n5242), .ZN(n5029)
         );
  OAI211_X1 U6219 ( .C1(n5247), .C2(n5031), .A(n5030), .B(n5029), .ZN(U3022)
         );
  INV_X1 U6220 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5034) );
  AOI22_X1 U6221 ( .A1(n5234), .A2(n6394), .B1(n6439), .B2(n5233), .ZN(n5033)
         );
  AOI22_X1 U6222 ( .A1(n6301), .A2(n6451), .B1(n6440), .B2(n5235), .ZN(n5032)
         );
  OAI211_X1 U6223 ( .C1(n5239), .C2(n5034), .A(n5033), .B(n5032), .ZN(U3036)
         );
  INV_X1 U6224 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5037) );
  AOI22_X1 U6225 ( .A1(n5241), .A2(n6394), .B1(n6439), .B2(n5240), .ZN(n5036)
         );
  AOI22_X1 U6226 ( .A1(n6451), .A2(n5243), .B1(n6440), .B2(n5242), .ZN(n5035)
         );
  OAI211_X1 U6227 ( .C1(n5247), .C2(n5037), .A(n5036), .B(n5035), .ZN(U3020)
         );
  NOR2_X2 U6228 ( .A1(n5039), .A2(n5038), .ZN(n6456) );
  INV_X1 U6229 ( .A(n6456), .ZN(n5047) );
  INV_X1 U6230 ( .A(DATAI_1_), .ZN(n5147) );
  NOR2_X2 U6231 ( .A1(n5147), .A2(n6353), .ZN(n6455) );
  AOI22_X1 U6232 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5041), .B1(n6455), 
        .B2(n5040), .ZN(n5045) );
  NAND2_X1 U6233 ( .A1(n6189), .A2(DATAI_25_), .ZN(n6459) );
  INV_X1 U6234 ( .A(n6459), .ZN(n6378) );
  INV_X1 U6235 ( .A(DATAI_17_), .ZN(n5042) );
  AOI22_X1 U6236 ( .A1(n6378), .A2(n5243), .B1(n5234), .B2(n5043), .ZN(n5044)
         );
  OAI211_X1 U6237 ( .C1(n5047), .C2(n5046), .A(n5045), .B(n5044), .ZN(U3029)
         );
  AOI22_X1 U6238 ( .A1(n6484), .A2(n3292), .B1(n5210), .B2(n6485), .ZN(n5049)
         );
  AOI22_X1 U6239 ( .A1(n5205), .A2(n6483), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n5116), .ZN(n5048) );
  OAI211_X1 U6240 ( .C1(n6488), .C2(n5212), .A(n5049), .B(n5048), .ZN(U3130)
         );
  AOI22_X1 U6241 ( .A1(n6473), .A2(n3292), .B1(n5210), .B2(n5001), .ZN(n5051)
         );
  AOI22_X1 U6242 ( .A1(n5205), .A2(n6472), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n5116), .ZN(n5050) );
  OAI211_X1 U6243 ( .C1(n6476), .C2(n5212), .A(n5051), .B(n5050), .ZN(U3128)
         );
  AOI22_X1 U6244 ( .A1(n6478), .A2(n3292), .B1(n5210), .B2(n6479), .ZN(n5053)
         );
  AOI22_X1 U6245 ( .A1(n5205), .A2(n6477), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n5116), .ZN(n5052) );
  OAI211_X1 U6246 ( .C1(n6482), .C2(n5212), .A(n5053), .B(n5052), .ZN(U3129)
         );
  INV_X1 U6247 ( .A(n6468), .ZN(n6417) );
  NAND2_X1 U6248 ( .A1(n5054), .A2(n6442), .ZN(n6438) );
  INV_X1 U6249 ( .A(n5055), .ZN(n6435) );
  INV_X1 U6250 ( .A(n5056), .ZN(n5057) );
  OAI22_X1 U6251 ( .A1(n6438), .A2(n5058), .B1(n6435), .B2(n5057), .ZN(n5227)
         );
  NOR2_X1 U6252 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5059), .ZN(n5228)
         );
  NOR2_X2 U6253 ( .A1(n5060), .A2(n6308), .ZN(n6302) );
  AOI211_X1 U6254 ( .C1(n6302), .C2(n6351), .A(n5062), .B(n5061), .ZN(n5064)
         );
  NOR3_X1 U6255 ( .A1(n5065), .A2(n5064), .A3(n5063), .ZN(n5066) );
  AOI22_X1 U6256 ( .A1(n5227), .A2(n6466), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5226), .ZN(n5068) );
  AOI22_X1 U6257 ( .A1(n6302), .A2(n6414), .B1(n6467), .B2(n5228), .ZN(n5067)
         );
  OAI211_X1 U6258 ( .C1(n5232), .C2(n6417), .A(n5068), .B(n5067), .ZN(U3055)
         );
  INV_X1 U6259 ( .A(n6451), .ZN(n6409) );
  AOI22_X1 U6260 ( .A1(n5227), .A2(n6439), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5226), .ZN(n5070) );
  AOI22_X1 U6261 ( .A1(n6302), .A2(n6394), .B1(n6440), .B2(n5228), .ZN(n5069)
         );
  OAI211_X1 U6262 ( .C1(n5232), .C2(n6409), .A(n5070), .B(n5069), .ZN(U3052)
         );
  INV_X1 U6263 ( .A(n6462), .ZN(n5073) );
  AOI22_X1 U6264 ( .A1(n5227), .A2(n6461), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5226), .ZN(n5072) );
  AOI22_X1 U6265 ( .A1(n6302), .A2(n6382), .B1(n6460), .B2(n5228), .ZN(n5071)
         );
  OAI211_X1 U6266 ( .C1(n5232), .C2(n5073), .A(n5072), .B(n5071), .ZN(U3054)
         );
  INV_X1 U6267 ( .A(n7020), .ZN(n5076) );
  AOI22_X1 U6268 ( .A1(n5227), .A2(n7019), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5226), .ZN(n5075) );
  AOI22_X1 U6269 ( .A1(n6302), .A2(n6300), .B1(n7027), .B2(n5228), .ZN(n5074)
         );
  OAI211_X1 U6270 ( .C1(n5232), .C2(n5076), .A(n5075), .B(n5074), .ZN(U3059)
         );
  INV_X1 U6271 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U6272 ( .A1(n5241), .A2(n6479), .B1(n6477), .B2(n5125), .ZN(n5078)
         );
  AOI22_X1 U6273 ( .A1(n6478), .A2(n5127), .B1(n5126), .B2(n6420), .ZN(n5077)
         );
  OAI211_X1 U6274 ( .C1(n5131), .C2(n5079), .A(n5078), .B(n5077), .ZN(U3145)
         );
  AOI22_X1 U6275 ( .A1(n5210), .A2(n6420), .B1(n6477), .B2(n5119), .ZN(n5081)
         );
  AOI22_X1 U6276 ( .A1(n6478), .A2(n5120), .B1(n5126), .B2(n6479), .ZN(n5080)
         );
  OAI211_X1 U6277 ( .C1(n5124), .C2(n5082), .A(n5081), .B(n5080), .ZN(U3137)
         );
  INV_X1 U6278 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5085) );
  AOI22_X1 U6279 ( .A1(n5210), .A2(n6289), .B1(n6472), .B2(n5119), .ZN(n5084)
         );
  AOI22_X1 U6280 ( .A1(n6473), .A2(n5120), .B1(n5126), .B2(n5001), .ZN(n5083)
         );
  OAI211_X1 U6281 ( .C1(n5124), .C2(n5085), .A(n5084), .B(n5083), .ZN(U3136)
         );
  INV_X1 U6282 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5088) );
  AOI22_X1 U6283 ( .A1(n5241), .A2(n6485), .B1(n6483), .B2(n5125), .ZN(n5087)
         );
  AOI22_X1 U6284 ( .A1(n6484), .A2(n5127), .B1(n5126), .B2(n6333), .ZN(n5086)
         );
  OAI211_X1 U6285 ( .C1(n5131), .C2(n5088), .A(n5087), .B(n5086), .ZN(U3146)
         );
  INV_X1 U6286 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5091) );
  AOI22_X1 U6287 ( .A1(n5241), .A2(n5001), .B1(n6472), .B2(n5125), .ZN(n5090)
         );
  AOI22_X1 U6288 ( .A1(n6473), .A2(n5127), .B1(n5126), .B2(n6289), .ZN(n5089)
         );
  OAI211_X1 U6289 ( .C1(n5131), .C2(n5091), .A(n5090), .B(n5089), .ZN(U3144)
         );
  INV_X1 U6290 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5094) );
  AOI22_X1 U6291 ( .A1(n5210), .A2(n6333), .B1(n6483), .B2(n5119), .ZN(n5093)
         );
  AOI22_X1 U6292 ( .A1(n6484), .A2(n5120), .B1(n5126), .B2(n6485), .ZN(n5092)
         );
  OAI211_X1 U6293 ( .C1(n5124), .C2(n5094), .A(n5093), .B(n5092), .ZN(U3138)
         );
  XNOR2_X1 U6294 ( .A(n3195), .B(n5096), .ZN(n5136) );
  INV_X1 U6295 ( .A(n5097), .ZN(n5099) );
  AOI22_X1 U6296 ( .A1(n5558), .A2(n5099), .B1(n5557), .B2(n5098), .ZN(n6238)
         );
  INV_X1 U6297 ( .A(n6238), .ZN(n5106) );
  AOI21_X1 U6298 ( .B1(n5100), .B2(n5963), .A(n5944), .ZN(n5101) );
  INV_X1 U6299 ( .A(n5101), .ZN(n6054) );
  OAI22_X1 U6300 ( .A1(n6054), .A2(n6258), .B1(n6563), .B2(n6256), .ZN(n5105)
         );
  INV_X1 U6301 ( .A(n5272), .ZN(n5271) );
  AOI211_X1 U6302 ( .C1(n6237), .C2(n6757), .A(n5271), .B(n6234), .ZN(n5104)
         );
  AOI211_X1 U6303 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n5106), .A(n5105), 
        .B(n5104), .ZN(n5107) );
  OAI21_X1 U6304 ( .B1(n6208), .B2(n5136), .A(n5107), .ZN(U3010) );
  AOI22_X1 U6305 ( .A1(n7021), .A2(n5043), .B1(n6455), .B2(n7018), .ZN(n5108)
         );
  OAI21_X1 U6306 ( .B1(n7024), .B2(n6459), .A(n5108), .ZN(n5109) );
  AOI21_X1 U6307 ( .B1(n6456), .B2(n7026), .A(n5109), .ZN(n5110) );
  OAI21_X1 U6308 ( .B1(n7030), .B2(n5111), .A(n5110), .ZN(U3069) );
  OAI21_X1 U6309 ( .B1(n5112), .B2(n5115), .A(n5114), .ZN(n6169) );
  INV_X1 U6310 ( .A(DATAI_9_), .ZN(n6936) );
  INV_X1 U6311 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6128) );
  OAI222_X1 U6312 ( .A1(n5398), .A2(n6169), .B1(n5406), .B2(n6936), .C1(n5405), 
        .C2(n6128), .ZN(U2882) );
  AOI22_X1 U6313 ( .A1(n6456), .A2(n3292), .B1(n5210), .B2(n5043), .ZN(n5118)
         );
  AOI22_X1 U6314 ( .A1(n5205), .A2(n6455), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n5116), .ZN(n5117) );
  OAI211_X1 U6315 ( .C1(n6459), .C2(n5212), .A(n5118), .B(n5117), .ZN(U3125)
         );
  INV_X1 U6316 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5123) );
  AOI22_X1 U6317 ( .A1(n5210), .A2(n6378), .B1(n6455), .B2(n5119), .ZN(n5122)
         );
  AOI22_X1 U6318 ( .A1(n6456), .A2(n5120), .B1(n5126), .B2(n5043), .ZN(n5121)
         );
  OAI211_X1 U6319 ( .C1(n5124), .C2(n5123), .A(n5122), .B(n5121), .ZN(U3133)
         );
  INV_X1 U6320 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5130) );
  AOI22_X1 U6321 ( .A1(n5241), .A2(n5043), .B1(n6455), .B2(n5125), .ZN(n5129)
         );
  AOI22_X1 U6322 ( .A1(n6456), .A2(n5127), .B1(n5126), .B2(n6378), .ZN(n5128)
         );
  OAI211_X1 U6323 ( .C1(n5131), .C2(n5130), .A(n5129), .B(n5128), .ZN(U3141)
         );
  NAND2_X1 U6324 ( .A1(n5132), .A2(n5133), .ZN(n5135) );
  INV_X1 U6325 ( .A(n5112), .ZN(n5134) );
  NAND2_X1 U6326 ( .A1(n5135), .A2(n5134), .ZN(n6056) );
  OR2_X1 U6327 ( .A1(n5136), .A2(n6179), .ZN(n5139) );
  OAI22_X1 U6328 ( .A1(n5741), .A2(n5952), .B1(n6256), .B2(n6563), .ZN(n5137)
         );
  AOI21_X1 U6329 ( .B1(n6198), .B2(n5957), .A(n5137), .ZN(n5138) );
  OAI211_X1 U6330 ( .C1(n6203), .C2(n6056), .A(n5139), .B(n5138), .ZN(U2978)
         );
  OR2_X1 U6331 ( .A1(n4701), .A2(n5140), .ZN(n5141) );
  NAND2_X1 U6332 ( .A1(n5141), .A2(n4751), .ZN(n6184) );
  INV_X1 U6333 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6867) );
  OAI222_X1 U6334 ( .A1(n6184), .A2(n5398), .B1(n5406), .B2(n5142), .C1(n5405), 
        .C2(n6867), .ZN(U2886) );
  OR2_X1 U6335 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  NAND2_X1 U6336 ( .A1(n5146), .A2(n5145), .ZN(n6202) );
  INV_X1 U6337 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6143) );
  OAI222_X1 U6338 ( .A1(n6202), .A2(n5398), .B1(n5406), .B2(n5147), .C1(n5405), 
        .C2(n6143), .ZN(U2890) );
  OAI21_X1 U6339 ( .B1(n4750), .B2(n5148), .A(n5132), .ZN(n6177) );
  INV_X1 U6340 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6132) );
  OAI222_X1 U6341 ( .A1(n6177), .A2(n5398), .B1(n5406), .B2(n6854), .C1(n5405), 
        .C2(n6132), .ZN(U2884) );
  INV_X1 U6342 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6134) );
  OAI222_X1 U6343 ( .A1(n6061), .A2(n5398), .B1(n5406), .B2(n5149), .C1(n5405), 
        .C2(n6134), .ZN(U2885) );
  NOR2_X1 U6344 ( .A1(n5150), .A2(n5151), .ZN(n5152) );
  NOR2_X1 U6345 ( .A1(n4710), .A2(n5152), .ZN(n6188) );
  INV_X1 U6346 ( .A(n6188), .ZN(n5310) );
  INV_X1 U6347 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6141) );
  OAI222_X1 U6348 ( .A1(n5310), .A2(n5398), .B1(n5406), .B2(n5153), .C1(n5405), 
        .C2(n6141), .ZN(U2889) );
  INV_X1 U6349 ( .A(DATAI_8_), .ZN(n6889) );
  INV_X1 U6350 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6130) );
  OAI222_X1 U6351 ( .A1(n6056), .A2(n5398), .B1(n5406), .B2(n6889), .C1(n5405), 
        .C2(n6130), .ZN(U2883) );
  INV_X1 U6352 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6147) );
  OAI222_X1 U6353 ( .A1(n6084), .A2(n5398), .B1(n5406), .B2(n5154), .C1(n5405), 
        .C2(n6147), .ZN(U2891) );
  INV_X1 U6354 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6139) );
  OAI222_X1 U6355 ( .A1(n6070), .A2(n5398), .B1(n5406), .B2(n5155), .C1(n5405), 
        .C2(n6139), .ZN(U2888) );
  INV_X1 U6356 ( .A(n6477), .ZN(n6295) );
  AOI22_X1 U6357 ( .A1(n5195), .A2(n6479), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n5194), .ZN(n5157) );
  AOI22_X1 U6358 ( .A1(n5197), .A2(n6420), .B1(n6478), .B2(n5196), .ZN(n5156)
         );
  OAI211_X1 U6359 ( .C1(n5200), .C2(n6295), .A(n5157), .B(n5156), .ZN(U3065)
         );
  INV_X1 U6360 ( .A(n6483), .ZN(n6298) );
  AOI22_X1 U6361 ( .A1(n5195), .A2(n6485), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n5194), .ZN(n5159) );
  AOI22_X1 U6362 ( .A1(n5197), .A2(n6333), .B1(n6484), .B2(n5196), .ZN(n5158)
         );
  OAI211_X1 U6363 ( .C1(n5200), .C2(n6298), .A(n5159), .B(n5158), .ZN(U3066)
         );
  INV_X1 U6364 ( .A(n6472), .ZN(n6292) );
  AOI22_X1 U6365 ( .A1(n5195), .A2(n5001), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n5194), .ZN(n5161) );
  AOI22_X1 U6366 ( .A1(n5197), .A2(n6289), .B1(n6473), .B2(n5196), .ZN(n5160)
         );
  OAI211_X1 U6367 ( .C1(n5200), .C2(n6292), .A(n5161), .B(n5160), .ZN(U3064)
         );
  INV_X1 U6368 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n5163) );
  AOI22_X1 U6369 ( .A1(n6440), .A2(n3292), .B1(n6439), .B2(n5205), .ZN(n5162)
         );
  OAI21_X1 U6370 ( .B1(n5208), .B2(n5163), .A(n5162), .ZN(n5164) );
  AOI21_X1 U6371 ( .B1(n5210), .B2(n6451), .A(n5164), .ZN(n5165) );
  OAI21_X1 U6372 ( .B1(n5212), .B2(n6454), .A(n5165), .ZN(U3124) );
  INV_X1 U6373 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5168) );
  AOI22_X1 U6374 ( .A1(n5241), .A2(n6420), .B1(n6477), .B2(n5240), .ZN(n5167)
         );
  AOI22_X1 U6375 ( .A1(n5243), .A2(n6479), .B1(n6478), .B2(n5242), .ZN(n5166)
         );
  OAI211_X1 U6376 ( .C1(n5247), .C2(n5168), .A(n5167), .B(n5166), .ZN(U3025)
         );
  INV_X1 U6377 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5171) );
  AOI22_X1 U6378 ( .A1(n5241), .A2(n6289), .B1(n6472), .B2(n5240), .ZN(n5170)
         );
  AOI22_X1 U6379 ( .A1(n5243), .A2(n5001), .B1(n6473), .B2(n5242), .ZN(n5169)
         );
  OAI211_X1 U6380 ( .C1(n5247), .C2(n5171), .A(n5170), .B(n5169), .ZN(U3024)
         );
  INV_X1 U6381 ( .A(n6485), .ZN(n6336) );
  AOI22_X1 U6382 ( .A1(n5227), .A2(n6483), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5226), .ZN(n5173) );
  AOI22_X1 U6383 ( .A1(n6302), .A2(n6333), .B1(n6484), .B2(n5228), .ZN(n5172)
         );
  OAI211_X1 U6384 ( .C1(n5232), .C2(n6336), .A(n5173), .B(n5172), .ZN(U3058)
         );
  AOI22_X1 U6385 ( .A1(n5234), .A2(n6333), .B1(n6483), .B2(n5233), .ZN(n5175)
         );
  AOI22_X1 U6386 ( .A1(n6301), .A2(n6485), .B1(n6484), .B2(n5235), .ZN(n5174)
         );
  OAI211_X1 U6387 ( .C1(n5239), .C2(n5176), .A(n5175), .B(n5174), .ZN(U3042)
         );
  INV_X1 U6388 ( .A(n6479), .ZN(n6424) );
  AOI22_X1 U6389 ( .A1(n5227), .A2(n6477), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5226), .ZN(n5178) );
  AOI22_X1 U6390 ( .A1(n6302), .A2(n6420), .B1(n6478), .B2(n5228), .ZN(n5177)
         );
  OAI211_X1 U6391 ( .C1(n5232), .C2(n6424), .A(n5178), .B(n5177), .ZN(U3057)
         );
  INV_X1 U6392 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5181) );
  AOI22_X1 U6393 ( .A1(n5234), .A2(n6420), .B1(n6477), .B2(n5233), .ZN(n5180)
         );
  AOI22_X1 U6394 ( .A1(n6301), .A2(n6479), .B1(n6478), .B2(n5235), .ZN(n5179)
         );
  OAI211_X1 U6395 ( .C1(n5239), .C2(n5181), .A(n5180), .B(n5179), .ZN(U3041)
         );
  AOI22_X1 U6396 ( .A1(n5234), .A2(n6289), .B1(n6472), .B2(n5233), .ZN(n5183)
         );
  AOI22_X1 U6397 ( .A1(n6301), .A2(n5001), .B1(n6473), .B2(n5235), .ZN(n5182)
         );
  OAI211_X1 U6398 ( .C1(n5239), .C2(n5184), .A(n5183), .B(n5182), .ZN(U3040)
         );
  INV_X1 U6399 ( .A(n5001), .ZN(n5187) );
  AOI22_X1 U6400 ( .A1(n5227), .A2(n6472), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5226), .ZN(n5186) );
  AOI22_X1 U6401 ( .A1(n6302), .A2(n6289), .B1(n6473), .B2(n5228), .ZN(n5185)
         );
  OAI211_X1 U6402 ( .C1(n5232), .C2(n5187), .A(n5186), .B(n5185), .ZN(U3056)
         );
  INV_X1 U6403 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6869) );
  AOI22_X1 U6404 ( .A1(n5241), .A2(n6333), .B1(n6483), .B2(n5240), .ZN(n5189)
         );
  AOI22_X1 U6405 ( .A1(n5243), .A2(n6485), .B1(n6484), .B2(n5242), .ZN(n5188)
         );
  OAI211_X1 U6406 ( .C1(n5247), .C2(n6869), .A(n5189), .B(n5188), .ZN(U3026)
         );
  INV_X1 U6407 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5193) );
  AOI22_X1 U6408 ( .A1(n6421), .A2(n6462), .B1(n6460), .B2(n5280), .ZN(n5190)
         );
  OAI21_X1 U6409 ( .B1(n5282), .B2(n6465), .A(n5190), .ZN(n5191) );
  AOI21_X1 U6410 ( .B1(n5284), .B2(n6461), .A(n5191), .ZN(n5192) );
  OAI21_X1 U6411 ( .B1(n5287), .B2(n5193), .A(n5192), .ZN(U3102) );
  INV_X1 U6412 ( .A(n6455), .ZN(n6282) );
  AOI22_X1 U6413 ( .A1(n5195), .A2(n5043), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n5194), .ZN(n5199) );
  AOI22_X1 U6414 ( .A1(n5197), .A2(n6378), .B1(n6456), .B2(n5196), .ZN(n5198)
         );
  OAI211_X1 U6415 ( .C1(n5200), .C2(n6282), .A(n5199), .B(n5198), .ZN(U3061)
         );
  INV_X1 U6416 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5204) );
  AOI22_X1 U6417 ( .A1(n6421), .A2(n6451), .B1(n6440), .B2(n5280), .ZN(n5201)
         );
  OAI21_X1 U6418 ( .B1(n5282), .B2(n6454), .A(n5201), .ZN(n5202) );
  AOI21_X1 U6419 ( .B1(n5284), .B2(n6439), .A(n5202), .ZN(n5203) );
  OAI21_X1 U6420 ( .B1(n5287), .B2(n5204), .A(n5203), .ZN(U3100) );
  INV_X1 U6421 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n5207) );
  AOI22_X1 U6422 ( .A1(n6461), .A2(n5205), .B1(n6460), .B2(n3292), .ZN(n5206)
         );
  OAI21_X1 U6423 ( .B1(n5208), .B2(n5207), .A(n5206), .ZN(n5209) );
  AOI21_X1 U6424 ( .B1(n5210), .B2(n6462), .A(n5209), .ZN(n5211) );
  OAI21_X1 U6425 ( .B1(n5212), .B2(n6465), .A(n5211), .ZN(U3126) );
  AND2_X1 U6426 ( .A1(n5214), .A2(n5213), .ZN(n5216) );
  OR2_X1 U6427 ( .A1(n5216), .A2(n5215), .ZN(n6066) );
  AOI22_X1 U6428 ( .A1(n6221), .A2(REIP_REG_4__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n5217), .ZN(n5218) );
  OAI21_X1 U6429 ( .B1(n6066), .B2(n6258), .A(n5218), .ZN(n5223) );
  OAI211_X1 U6430 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5220), .B(n5219), .ZN(n5221) );
  INV_X1 U6431 ( .A(n5221), .ZN(n5222) );
  AOI211_X1 U6432 ( .C1(n5224), .C2(n3833), .A(n5223), .B(n5222), .ZN(n5225)
         );
  INV_X1 U6433 ( .A(n5225), .ZN(U3014) );
  INV_X1 U6434 ( .A(n5043), .ZN(n5231) );
  AOI22_X1 U6435 ( .A1(n5227), .A2(n6455), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5226), .ZN(n5230) );
  AOI22_X1 U6436 ( .A1(n6302), .A2(n6378), .B1(n6456), .B2(n5228), .ZN(n5229)
         );
  OAI211_X1 U6437 ( .C1(n5232), .C2(n5231), .A(n5230), .B(n5229), .ZN(U3053)
         );
  AOI22_X1 U6438 ( .A1(n5234), .A2(n6378), .B1(n6455), .B2(n5233), .ZN(n5237)
         );
  AOI22_X1 U6439 ( .A1(n6301), .A2(n5043), .B1(n6456), .B2(n5235), .ZN(n5236)
         );
  OAI211_X1 U6440 ( .C1(n5239), .C2(n5238), .A(n5237), .B(n5236), .ZN(U3037)
         );
  INV_X1 U6441 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U6442 ( .A1(n5241), .A2(n6378), .B1(n6455), .B2(n5240), .ZN(n5245)
         );
  AOI22_X1 U6443 ( .A1(n5243), .A2(n5043), .B1(n6456), .B2(n5242), .ZN(n5244)
         );
  OAI211_X1 U6444 ( .C1(n5247), .C2(n5246), .A(n5245), .B(n5244), .ZN(U3021)
         );
  NAND2_X1 U6445 ( .A1(n5114), .A2(n5248), .ZN(n5252) );
  INV_X1 U6446 ( .A(n5250), .ZN(n5251) );
  AOI22_X1 U6447 ( .A1(n5401), .A2(DATAI_10_), .B1(n6089), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5253) );
  OAI21_X1 U6448 ( .B1(n6051), .B2(n5407), .A(n5253), .ZN(U2881) );
  INV_X1 U6449 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U6450 ( .A1(n6421), .A2(n5001), .B1(n6473), .B2(n5280), .ZN(n5254)
         );
  OAI21_X1 U6451 ( .B1(n5282), .B2(n6476), .A(n5254), .ZN(n5255) );
  AOI21_X1 U6452 ( .B1(n5284), .B2(n6472), .A(n5255), .ZN(n5256) );
  OAI21_X1 U6453 ( .B1(n5287), .B2(n6743), .A(n5256), .ZN(U3104) );
  INV_X1 U6454 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5260) );
  AOI22_X1 U6455 ( .A1(n6421), .A2(n6485), .B1(n6484), .B2(n5280), .ZN(n5257)
         );
  OAI21_X1 U6456 ( .B1(n5282), .B2(n6488), .A(n5257), .ZN(n5258) );
  AOI21_X1 U6457 ( .B1(n5284), .B2(n6483), .A(n5258), .ZN(n5259) );
  OAI21_X1 U6458 ( .B1(n5287), .B2(n5260), .A(n5259), .ZN(U3106) );
  INV_X1 U6459 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5264) );
  AOI22_X1 U6460 ( .A1(n6421), .A2(n6479), .B1(n6478), .B2(n5280), .ZN(n5261)
         );
  OAI21_X1 U6461 ( .B1(n5282), .B2(n6482), .A(n5261), .ZN(n5262) );
  AOI21_X1 U6462 ( .B1(n5284), .B2(n6477), .A(n5262), .ZN(n5263) );
  OAI21_X1 U6463 ( .B1(n5287), .B2(n5264), .A(n5263), .ZN(U3105) );
  OAI21_X1 U6464 ( .B1(n5250), .B2(n5266), .A(n5265), .ZN(n6163) );
  INV_X1 U6465 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6886) );
  OAI222_X1 U6466 ( .A1(n5398), .A2(n6163), .B1(n5406), .B2(n5267), .C1(n5405), 
        .C2(n6886), .ZN(U2880) );
  NAND2_X1 U6467 ( .A1(n3238), .A2(n5269), .ZN(n5270) );
  XNOR2_X1 U6468 ( .A(n5268), .B(n5270), .ZN(n5322) );
  OAI21_X1 U6469 ( .B1(n5271), .B2(n5804), .A(n6238), .ZN(n6220) );
  NOR2_X1 U6470 ( .A1(n5272), .A2(n6234), .ZN(n6224) );
  OAI211_X1 U6471 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6224), .B(n5273), .ZN(n5277) );
  NAND2_X1 U6472 ( .A1(n5945), .A2(n5274), .ZN(n5275) );
  AND2_X1 U6473 ( .A1(n5924), .A2(n5275), .ZN(n6048) );
  NAND2_X1 U6474 ( .A1(n6048), .A2(n6245), .ZN(n5276) );
  OAI211_X1 U6475 ( .C1(n6768), .C2(n6256), .A(n5277), .B(n5276), .ZN(n5278)
         );
  AOI21_X1 U6476 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6220), .A(n5278), 
        .ZN(n5279) );
  OAI21_X1 U6477 ( .B1(n6208), .B2(n5322), .A(n5279), .ZN(U3008) );
  INV_X1 U6478 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5286) );
  AOI22_X1 U6479 ( .A1(n6421), .A2(n5043), .B1(n6456), .B2(n5280), .ZN(n5281)
         );
  OAI21_X1 U6480 ( .B1(n5282), .B2(n6459), .A(n5281), .ZN(n5283) );
  AOI21_X1 U6481 ( .B1(n5284), .B2(n6455), .A(n5283), .ZN(n5285) );
  OAI21_X1 U6482 ( .B1(n5287), .B2(n5286), .A(n5285), .ZN(U3101) );
  INV_X1 U6483 ( .A(n5299), .ZN(n5288) );
  OAI21_X1 U6484 ( .B1(n5289), .B2(n5288), .A(n3197), .ZN(n6004) );
  INV_X1 U6485 ( .A(n6004), .ZN(n6018) );
  INV_X1 U6486 ( .A(n5290), .ZN(n5291) );
  INV_X1 U6487 ( .A(n6192), .ZN(n5308) );
  INV_X1 U6488 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6026) );
  NAND3_X1 U6489 ( .A1(n3834), .A2(n6026), .A3(n5293), .ZN(n5295) );
  NAND2_X1 U6490 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  AND2_X2 U6491 ( .A1(n5299), .A2(n5296), .ZN(n6021) );
  AOI22_X1 U6492 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6021), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6000), .ZN(n5297) );
  INV_X1 U6493 ( .A(n5297), .ZN(n5307) );
  AOI21_X1 U6494 ( .B1(n5997), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5305) );
  OAI211_X1 U6495 ( .C1(REIP_REG_1__SCAN_IN), .C2(n5993), .A(
        REIP_REG_2__SCAN_IN), .B(n5965), .ZN(n6023) );
  INV_X1 U6496 ( .A(n6023), .ZN(n5304) );
  AND2_X1 U6497 ( .A1(n5299), .A2(n5298), .ZN(n6005) );
  XNOR2_X1 U6498 ( .A(n5301), .B(n5300), .ZN(n6244) );
  AOI22_X1 U6499 ( .A1(n5302), .A2(n6005), .B1(n5983), .B2(n6244), .ZN(n5303)
         );
  OAI21_X1 U6500 ( .B1(n5305), .B2(n5304), .A(n5303), .ZN(n5306) );
  AOI211_X1 U6501 ( .C1(n6002), .C2(n5308), .A(n5307), .B(n5306), .ZN(n5309)
         );
  OAI21_X1 U6502 ( .B1(n6018), .B2(n5310), .A(n5309), .ZN(U2825) );
  AOI21_X1 U6503 ( .B1(n5265), .B2(n5312), .A(n5311), .ZN(n6045) );
  INV_X1 U6504 ( .A(n6045), .ZN(n5314) );
  AOI22_X1 U6505 ( .A1(n5401), .A2(DATAI_12_), .B1(n6089), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5313) );
  OAI21_X1 U6506 ( .B1(n5314), .B2(n5407), .A(n5313), .ZN(U2879) );
  INV_X1 U6507 ( .A(n6005), .ZN(n6013) );
  NOR2_X1 U6508 ( .A1(n6013), .A2(n3982), .ZN(n5316) );
  OAI22_X1 U6509 ( .A1(n6082), .A2(n5951), .B1(n6015), .B2(n6080), .ZN(n5315)
         );
  AOI211_X1 U6510 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5676), .A(n5316), .B(n5315), 
        .ZN(n5318) );
  OAI21_X1 U6511 ( .B1(n6002), .B2(n6000), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5317) );
  OAI211_X1 U6512 ( .C1(n6018), .C2(n6084), .A(n5318), .B(n5317), .ZN(U2827)
         );
  OAI22_X1 U6513 ( .A1(n5741), .A2(n6771), .B1(n6256), .B2(n6768), .ZN(n5320)
         );
  NOR2_X1 U6514 ( .A1(n6051), .A2(n6203), .ZN(n5319) );
  AOI211_X1 U6515 ( .C1(n6198), .C2(n5936), .A(n5320), .B(n5319), .ZN(n5321)
         );
  OAI21_X1 U6516 ( .B1(n6179), .B2(n5322), .A(n5321), .ZN(U2976) );
  INV_X1 U6517 ( .A(n5324), .ZN(n5325) );
  XNOR2_X1 U6518 ( .A(n5323), .B(n5325), .ZN(n5904) );
  OAI222_X1 U6519 ( .A1(n6044), .A2(n5398), .B1(n5406), .B2(n5326), .C1(n5405), 
        .C2(n6832), .ZN(U2878) );
  NOR3_X1 U6520 ( .A1(n6089), .A2(n5328), .A3(n5327), .ZN(n5329) );
  AOI22_X1 U6521 ( .A1(n6088), .A2(DATAI_12_), .B1(n6089), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6522 ( .A1(n6085), .A2(DATAI_28_), .ZN(n5330) );
  OAI211_X1 U6523 ( .C1(n5618), .C2(n5407), .A(n5331), .B(n5330), .ZN(U2863)
         );
  INV_X1 U6524 ( .A(n5332), .ZN(n5345) );
  NOR2_X1 U6525 ( .A1(n5334), .A2(n5562), .ZN(n5341) );
  NAND2_X1 U6526 ( .A1(n4721), .A2(n5335), .ZN(n5339) );
  OAI21_X1 U6527 ( .B1(n5333), .B2(n5337), .A(n5336), .ZN(n5338) );
  OAI211_X1 U6528 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n5340), .A(n5339), .B(n5338), .ZN(n6499) );
  AOI222_X1 U6529 ( .A1(n5343), .A2(n5333), .B1(n5342), .B2(n5341), .C1(n6499), 
        .C2(n5837), .ZN(n5344) );
  OAI22_X1 U6530 ( .A1(n5345), .A2(n6818), .B1(n5586), .B2(n5344), .ZN(U3460)
         );
  INV_X1 U6531 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6532 ( .A1(n6021), .A2(EBX_REG_1__SCAN_IN), .ZN(n5348) );
  INV_X1 U6533 ( .A(n5965), .ZN(n5995) );
  OAI22_X1 U6534 ( .A1(REIP_REG_1__SCAN_IN), .A2(n5993), .B1(n6076), .B2(n6015), .ZN(n5346) );
  AOI21_X1 U6535 ( .B1(n5995), .B2(REIP_REG_1__SCAN_IN), .A(n5346), .ZN(n5347)
         );
  OAI211_X1 U6536 ( .C1(n5349), .C2(n6012), .A(n5348), .B(n5347), .ZN(n5351)
         );
  NOR2_X1 U6537 ( .A1(n6017), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5350)
         );
  AOI211_X1 U6538 ( .C1(n6005), .C2(n4721), .A(n5351), .B(n5350), .ZN(n5352)
         );
  OAI21_X1 U6539 ( .B1(n6018), .B2(n6202), .A(n5352), .ZN(U2826) );
  AOI22_X1 U6540 ( .A1(n6088), .A2(DATAI_14_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6089), .ZN(n5354) );
  NAND2_X1 U6541 ( .A1(n6085), .A2(DATAI_30_), .ZN(n5353) );
  OAI211_X1 U6542 ( .C1(n5686), .C2(n5407), .A(n5354), .B(n5353), .ZN(U2861)
         );
  AOI22_X1 U6543 ( .A1(n6088), .A2(DATAI_13_), .B1(n6089), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6544 ( .A1(n6085), .A2(DATAI_29_), .ZN(n5355) );
  OAI211_X1 U6545 ( .C1(n3223), .C2(n5398), .A(n5356), .B(n5355), .ZN(U2862)
         );
  AOI21_X1 U6546 ( .B1(n5357), .B2(n5359), .A(n5358), .ZN(n5418) );
  AOI22_X1 U6547 ( .A1(n6088), .A2(DATAI_11_), .B1(n6085), .B2(DATAI_27_), 
        .ZN(n5361) );
  NAND2_X1 U6548 ( .A1(n6089), .A2(EAX_REG_27__SCAN_IN), .ZN(n5360) );
  OAI211_X1 U6549 ( .C1(n5691), .C2(n5407), .A(n5361), .B(n5360), .ZN(U2864)
         );
  OAI21_X1 U6551 ( .B1(n5363), .B2(n5364), .A(n5357), .ZN(n5723) );
  AOI22_X1 U6552 ( .A1(n6088), .A2(DATAI_10_), .B1(n6089), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6553 ( .A1(n6085), .A2(DATAI_26_), .ZN(n5365) );
  OAI211_X1 U6554 ( .C1(n5723), .C2(n5398), .A(n5366), .B(n5365), .ZN(U2865)
         );
  NAND2_X1 U6555 ( .A1(n4488), .A2(n5367), .ZN(n5369) );
  INV_X1 U6556 ( .A(n5363), .ZN(n5368) );
  AOI22_X1 U6557 ( .A1(n6088), .A2(DATAI_9_), .B1(n6089), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6558 ( .A1(n6085), .A2(DATAI_25_), .ZN(n5370) );
  OAI211_X1 U6559 ( .C1(n5697), .C2(n5398), .A(n5371), .B(n5370), .ZN(U2866)
         );
  AOI22_X1 U6560 ( .A1(n6088), .A2(DATAI_8_), .B1(n6089), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6561 ( .A1(n6085), .A2(DATAI_24_), .ZN(n5372) );
  OAI211_X1 U6562 ( .C1(n5699), .C2(n5398), .A(n5373), .B(n5372), .ZN(U2867)
         );
  NOR2_X1 U6563 ( .A1(n5374), .A2(n5375), .ZN(n5376) );
  NOR2_X1 U6564 ( .A1(n4487), .A2(n5376), .ZN(n5652) );
  INV_X1 U6565 ( .A(n5652), .ZN(n5702) );
  AOI22_X1 U6566 ( .A1(n6088), .A2(DATAI_7_), .B1(n6089), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6567 ( .A1(n6085), .A2(DATAI_23_), .ZN(n5377) );
  OAI211_X1 U6568 ( .C1(n5702), .C2(n5398), .A(n5378), .B(n5377), .ZN(U2868)
         );
  INV_X1 U6569 ( .A(n5374), .ZN(n5380) );
  OAI21_X1 U6570 ( .B1(n5381), .B2(n5379), .A(n5380), .ZN(n5734) );
  AOI22_X1 U6571 ( .A1(n6088), .A2(DATAI_6_), .B1(n6089), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6572 ( .A1(n6085), .A2(DATAI_22_), .ZN(n5382) );
  OAI211_X1 U6573 ( .C1(n5734), .C2(n5407), .A(n5383), .B(n5382), .ZN(U2869)
         );
  AOI21_X1 U6574 ( .B1(n3219), .B2(n5384), .A(n5379), .ZN(n5738) );
  INV_X1 U6575 ( .A(n5738), .ZN(n5706) );
  AOI22_X1 U6576 ( .A1(n6088), .A2(DATAI_5_), .B1(n6089), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6577 ( .A1(n6085), .A2(DATAI_21_), .ZN(n5385) );
  OAI211_X1 U6578 ( .C1(n5706), .C2(n5398), .A(n5386), .B(n5385), .ZN(U2870)
         );
  OAI21_X1 U6579 ( .B1(n5387), .B2(n5390), .A(n5389), .ZN(n6029) );
  AOI22_X1 U6580 ( .A1(n6088), .A2(DATAI_2_), .B1(n6089), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6581 ( .A1(n6085), .A2(DATAI_18_), .ZN(n5391) );
  OAI211_X1 U6582 ( .C1(n6029), .C2(n5407), .A(n5392), .B(n5391), .ZN(U2873)
         );
  OAI21_X1 U6583 ( .B1(n5393), .B2(n5395), .A(n5394), .ZN(n6034) );
  AOI22_X1 U6584 ( .A1(n6088), .A2(DATAI_0_), .B1(n6089), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6585 ( .A1(n6085), .A2(DATAI_16_), .ZN(n5396) );
  OAI211_X1 U6586 ( .C1(n6034), .C2(n5398), .A(n5397), .B(n5396), .ZN(U2875)
         );
  XNOR2_X1 U6587 ( .A(n5399), .B(n5400), .ZN(n6038) );
  AOI22_X1 U6588 ( .A1(n5401), .A2(DATAI_15_), .B1(n6089), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5402) );
  OAI21_X1 U6589 ( .B1(n6038), .B2(n5407), .A(n5402), .ZN(U2876) );
  OAI21_X1 U6590 ( .B1(n5403), .B2(n5404), .A(n5399), .ZN(n6041) );
  INV_X1 U6591 ( .A(DATAI_14_), .ZN(n6942) );
  INV_X1 U6592 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6121) );
  OAI222_X1 U6593 ( .A1(n5407), .A2(n6041), .B1(n5406), .B2(n6942), .C1(n5405), 
        .C2(n6121), .ZN(U2877) );
  INV_X1 U6594 ( .A(n5408), .ZN(n5410) );
  NAND2_X1 U6595 ( .A1(n5410), .A2(n5409), .ZN(n5411) );
  XNOR2_X1 U6596 ( .A(n5411), .B(n5461), .ZN(n5459) );
  NOR2_X1 U6597 ( .A1(n6256), .A2(n5607), .ZN(n5460) );
  AOI21_X1 U6598 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5460), 
        .ZN(n5412) );
  OAI21_X1 U6599 ( .B1(n5608), .B2(n6193), .A(n5412), .ZN(n5413) );
  AOI21_X1 U6600 ( .B1(n5459), .B2(n6199), .A(n5413), .ZN(n5414) );
  OAI21_X1 U6601 ( .B1(n3223), .B2(n6203), .A(n5414), .ZN(U2957) );
  NOR2_X1 U6602 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  XOR2_X1 U6603 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(n5417), .Z(n5478) );
  NAND2_X1 U6604 ( .A1(n5418), .A2(n6189), .ZN(n5422) );
  INV_X1 U6605 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5419) );
  NOR2_X1 U6606 ( .A1(n6256), .A2(n5419), .ZN(n5473) );
  NOR2_X1 U6607 ( .A1(n5627), .A2(n6193), .ZN(n5420) );
  AOI211_X1 U6608 ( .C1(n6194), .C2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5473), 
        .B(n5420), .ZN(n5421) );
  OAI211_X1 U6609 ( .C1(n5478), .C2(n6179), .A(n5422), .B(n5421), .ZN(U2959)
         );
  NAND3_X1 U6610 ( .A1(n3725), .A2(n5531), .A3(n5507), .ZN(n5424) );
  OAI21_X1 U6611 ( .B1(n5425), .B2(n5424), .A(n5423), .ZN(n5426) );
  XNOR2_X1 U6612 ( .A(n5426), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5501)
         );
  NOR2_X1 U6613 ( .A1(n6256), .A2(n6583), .ZN(n5495) );
  AOI21_X1 U6614 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5495), 
        .ZN(n5427) );
  OAI21_X1 U6615 ( .B1(n5650), .B2(n6193), .A(n5427), .ZN(n5428) );
  AOI21_X1 U6616 ( .B1(n5652), .B2(n6189), .A(n5428), .ZN(n5429) );
  OAI21_X1 U6617 ( .B1(n5501), .B2(n6179), .A(n5429), .ZN(U2963) );
  XOR2_X1 U6618 ( .A(n5431), .B(n5430), .Z(n5539) );
  XOR2_X1 U6619 ( .A(n5432), .B(n5433), .Z(n5714) );
  NAND2_X1 U6620 ( .A1(n5714), .A2(n6189), .ZN(n5436) );
  NAND2_X1 U6621 ( .A1(n6221), .A2(REIP_REG_20__SCAN_IN), .ZN(n5529) );
  OAI21_X1 U6622 ( .B1(n5741), .B2(n6780), .A(n5529), .ZN(n5434) );
  AOI21_X1 U6623 ( .B1(n5672), .B2(n6198), .A(n5434), .ZN(n5435) );
  OAI211_X1 U6624 ( .C1(n5539), .C2(n6179), .A(n5436), .B(n5435), .ZN(U2966)
         );
  NAND2_X1 U6625 ( .A1(n6221), .A2(REIP_REG_13__SCAN_IN), .ZN(n5830) );
  OAI21_X1 U6626 ( .B1(n5741), .B2(n4113), .A(n5830), .ZN(n5442) );
  INV_X1 U6627 ( .A(n5437), .ZN(n5438) );
  AOI21_X1 U6628 ( .B1(n5440), .B2(n5439), .A(n5438), .ZN(n5820) );
  NOR2_X1 U6629 ( .A1(n5820), .A2(n6179), .ZN(n5441) );
  AOI211_X1 U6630 ( .C1(n6198), .C2(n5905), .A(n5442), .B(n5441), .ZN(n5443)
         );
  OAI21_X1 U6631 ( .B1(n6044), .B2(n6203), .A(n5443), .ZN(U2973) );
  XNOR2_X1 U6632 ( .A(n3725), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5445)
         );
  XNOR2_X1 U6633 ( .A(n5444), .B(n5445), .ZN(n6209) );
  INV_X1 U6634 ( .A(n5918), .ZN(n5447) );
  AOI22_X1 U6635 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6221), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5446) );
  OAI21_X1 U6636 ( .B1(n6193), .B2(n5447), .A(n5446), .ZN(n5448) );
  AOI21_X1 U6637 ( .B1(n6045), .B2(n6189), .A(n5448), .ZN(n5449) );
  OAI21_X1 U6638 ( .B1(n6209), .B2(n6179), .A(n5449), .ZN(U2974) );
  INV_X1 U6639 ( .A(n5463), .ZN(n5474) );
  NOR2_X1 U6640 ( .A1(n5452), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5451)
         );
  AOI21_X1 U6641 ( .B1(n5474), .B2(n5451), .A(n5450), .ZN(n5457) );
  NAND2_X1 U6642 ( .A1(n6255), .A2(n5452), .ZN(n5453) );
  NAND2_X1 U6643 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  NAND2_X1 U6644 ( .A1(n5455), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5456) );
  INV_X1 U6645 ( .A(n5459), .ZN(n5468) );
  AOI21_X1 U6646 ( .B1(n5611), .B2(n6245), .A(n5460), .ZN(n5467) );
  OAI21_X1 U6647 ( .B1(n5463), .B2(n5462), .A(n5461), .ZN(n5464) );
  NAND2_X1 U6648 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  OAI211_X1 U6649 ( .C1(n5468), .C2(n6208), .A(n5467), .B(n5466), .ZN(U2989)
         );
  INV_X1 U6650 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6919) );
  INV_X1 U6651 ( .A(n5469), .ZN(n5470) );
  OAI21_X1 U6652 ( .B1(n5471), .B2(n5484), .A(n5470), .ZN(n5693) );
  NOR2_X1 U6653 ( .A1(n5693), .A2(n6258), .ZN(n5472) );
  AOI211_X1 U6654 ( .C1(n5474), .C2(n6919), .A(n5473), .B(n5472), .ZN(n5477)
         );
  NAND2_X1 U6655 ( .A1(n5475), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5476) );
  OAI211_X1 U6656 ( .C1(n5478), .C2(n6208), .A(n5477), .B(n5476), .ZN(U2991)
         );
  NOR2_X1 U6657 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  XNOR2_X1 U6658 ( .A(n5479), .B(n5482), .ZN(n5720) );
  NAND2_X1 U6659 ( .A1(n5720), .A2(n3833), .ZN(n5491) );
  AOI21_X1 U6660 ( .B1(n5492), .B2(n5778), .A(n5483), .ZN(n5489) );
  AOI21_X1 U6661 ( .B1(n5485), .B2(n5636), .A(n5484), .ZN(n5486) );
  INV_X1 U6662 ( .A(n5486), .ZN(n5695) );
  INV_X1 U6663 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5487) );
  OAI22_X1 U6664 ( .A1(n5695), .A2(n6258), .B1(n6256), .B2(n5487), .ZN(n5488)
         );
  AOI21_X1 U6665 ( .B1(n5773), .B2(n5489), .A(n5488), .ZN(n5490) );
  OAI211_X1 U6666 ( .C1(n5779), .C2(n5492), .A(n5491), .B(n5490), .ZN(U2992)
         );
  INV_X1 U6667 ( .A(n5493), .ZN(n5499) );
  AOI21_X1 U6668 ( .B1(n3239), .B2(n3228), .A(n5494), .ZN(n5700) );
  AOI21_X1 U6669 ( .B1(n5700), .B2(n6245), .A(n5495), .ZN(n5496) );
  OAI21_X1 U6670 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5497), .A(n5496), 
        .ZN(n5498) );
  AOI21_X1 U6671 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5499), .A(n5498), 
        .ZN(n5500) );
  OAI21_X1 U6672 ( .B1(n5501), .B2(n6208), .A(n5500), .ZN(U2995) );
  AOI21_X1 U6673 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3725), .A(n5502), 
        .ZN(n5504) );
  INV_X1 U6674 ( .A(n5732), .ZN(n5512) );
  INV_X1 U6675 ( .A(n5519), .ZN(n5505) );
  OAI21_X1 U6676 ( .B1(n5505), .B2(n3240), .A(n3228), .ZN(n5704) );
  OAI22_X1 U6677 ( .A1(n5704), .A2(n6258), .B1(n6256), .B2(n6874), .ZN(n5510)
         );
  INV_X1 U6678 ( .A(n5506), .ZN(n5521) );
  NOR3_X1 U6679 ( .A1(n5521), .A2(n5508), .A3(n5507), .ZN(n5509) );
  AOI211_X1 U6680 ( .C1(n5523), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5510), .B(n5509), .ZN(n5511) );
  OAI21_X1 U6681 ( .B1(n5512), .B2(n6208), .A(n5511), .ZN(U2996) );
  AOI21_X1 U6682 ( .B1(n5515), .B2(n5514), .A(n5513), .ZN(n5736) );
  NAND2_X1 U6683 ( .A1(n6221), .A2(REIP_REG_21__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U6684 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  AND2_X1 U6685 ( .A1(n5519), .A2(n5518), .ZN(n5705) );
  NAND2_X1 U6686 ( .A1(n5705), .A2(n6245), .ZN(n5520) );
  OAI211_X1 U6687 ( .C1(n5521), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5739), .B(n5520), .ZN(n5522) );
  AOI21_X1 U6688 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5523), .A(n5522), 
        .ZN(n5524) );
  OAI21_X1 U6689 ( .B1(n5736), .B2(n6208), .A(n5524), .ZN(U2997) );
  MUX2_X1 U6690 ( .A(n5526), .B(n5546), .S(n5525), .Z(n5528) );
  XNOR2_X1 U6691 ( .A(n5528), .B(n5527), .ZN(n5709) );
  INV_X1 U6692 ( .A(n5529), .ZN(n5533) );
  NOR3_X1 U6693 ( .A1(n5531), .A2(n5530), .A3(n5543), .ZN(n5532) );
  AOI211_X1 U6694 ( .C1(n5709), .C2(n6245), .A(n5533), .B(n5532), .ZN(n5538)
         );
  OAI21_X1 U6695 ( .B1(n5795), .B2(n5534), .A(n5557), .ZN(n5536) );
  NAND2_X1 U6696 ( .A1(n5536), .A2(n5535), .ZN(n5794) );
  AOI21_X1 U6697 ( .B1(n6205), .B2(n5795), .A(n5794), .ZN(n5788) );
  OAI21_X1 U6698 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5804), .A(n5788), 
        .ZN(n5551) );
  NAND2_X1 U6699 ( .A1(n5551), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5537) );
  OAI211_X1 U6700 ( .C1(n5539), .C2(n6208), .A(n5538), .B(n5537), .ZN(U2998)
         );
  XNOR2_X1 U6701 ( .A(n3725), .B(n5541), .ZN(n5542) );
  XNOR2_X1 U6702 ( .A(n5540), .B(n5542), .ZN(n5743) );
  INV_X1 U6703 ( .A(n5743), .ZN(n5553) );
  NOR2_X1 U6704 ( .A1(n5543), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5550)
         );
  INV_X1 U6705 ( .A(n5790), .ZN(n5783) );
  MUX2_X1 U6706 ( .A(n5546), .B(n5545), .S(n3204), .Z(n5782) );
  NOR2_X1 U6707 ( .A1(n5783), .A2(n5782), .ZN(n5781) );
  XNOR2_X1 U6708 ( .A(n5781), .B(n5547), .ZN(n5711) );
  INV_X1 U6709 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5548) );
  OAI22_X1 U6710 ( .A1(n5711), .A2(n6258), .B1(n6256), .B2(n5548), .ZN(n5549)
         );
  AOI211_X1 U6711 ( .C1(n5551), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5550), .B(n5549), .ZN(n5552) );
  OAI21_X1 U6712 ( .B1(n5553), .B2(n6208), .A(n5552), .ZN(U2999) );
  XNOR2_X1 U6713 ( .A(n3725), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5555)
         );
  XNOR2_X1 U6714 ( .A(n5554), .B(n5555), .ZN(n5770) );
  INV_X1 U6715 ( .A(n5770), .ZN(n5573) );
  AOI22_X1 U6716 ( .A1(n5558), .A2(n5825), .B1(n5557), .B2(n5556), .ZN(n6219)
         );
  OAI21_X1 U6717 ( .B1(n5566), .B2(n5559), .A(n6219), .ZN(n5560) );
  AOI21_X1 U6718 ( .B1(n6204), .B2(n5561), .A(n5560), .ZN(n5835) );
  NOR3_X1 U6719 ( .A1(n5563), .A2(n5825), .A3(n5562), .ZN(n5564) );
  NOR2_X1 U6720 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6204), .ZN(n5827)
         );
  OAI21_X1 U6721 ( .B1(n5565), .B2(n5564), .A(n5827), .ZN(n5833) );
  AOI21_X1 U6722 ( .B1(n5835), .B2(n5833), .A(n5567), .ZN(n5571) );
  INV_X1 U6723 ( .A(n5801), .ZN(n6215) );
  AND3_X1 U6724 ( .A1(n5567), .A2(n6215), .A3(n5566), .ZN(n5570) );
  OAI21_X1 U6725 ( .B1(n5822), .B2(n5568), .A(n3217), .ZN(n6039) );
  OAI22_X1 U6726 ( .A1(n6039), .A2(n6258), .B1(n6256), .B2(n6570), .ZN(n5569)
         );
  NOR3_X1 U6727 ( .A1(n5571), .A2(n5570), .A3(n5569), .ZN(n5572) );
  OAI21_X1 U6728 ( .B1(n5573), .B2(n6208), .A(n5572), .ZN(U3004) );
  XNOR2_X1 U6729 ( .A(n6271), .B(n6395), .ZN(n5574) );
  OAI22_X1 U6730 ( .A1(n5574), .A2(n6617), .B1(n4617), .B2(n5580), .ZN(n5575)
         );
  MUX2_X1 U6731 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5575), .S(n6264), 
        .Z(U3463) );
  INV_X1 U6732 ( .A(n5576), .ZN(n5579) );
  NOR2_X1 U6733 ( .A1(n6310), .A2(n6395), .ZN(n6311) );
  OAI21_X1 U6734 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5577), .A(n6396), .ZN(
        n5578) );
  NOR3_X1 U6735 ( .A1(n5579), .A2(n6311), .A3(n5578), .ZN(n5581) );
  OAI22_X1 U6736 ( .A1(n5581), .A2(n6617), .B1(n6437), .B2(n5580), .ZN(n5582)
         );
  MUX2_X1 U6737 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5582), .S(n6264), 
        .Z(U3462) );
  OAI22_X1 U6738 ( .A1(n5585), .A2(n5584), .B1(n5583), .B2(n6524), .ZN(n5587)
         );
  MUX2_X1 U6739 ( .A(n5587), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5586), 
        .Z(U3456) );
  AOI22_X1 U6740 ( .A1(n6221), .A2(REIP_REG_15__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U6741 ( .A(n5588), .B(n5589), .ZN(n5813) );
  AOI22_X1 U6742 ( .A1(n5813), .A2(n6199), .B1(n6198), .B2(n5890), .ZN(n5590)
         );
  OAI211_X1 U6743 ( .C1(n6203), .C2(n6038), .A(n5591), .B(n5590), .ZN(U2971)
         );
  AND2_X1 U6744 ( .A1(n6144), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6745 ( .A(n5598), .ZN(n5599) );
  OAI22_X1 U6746 ( .A1(n5600), .A2(n6012), .B1(n5599), .B2(n6017), .ZN(n5601)
         );
  AOI211_X1 U6747 ( .C1(EBX_REG_30__SCAN_IN), .C2(n6021), .A(n5602), .B(n5601), 
        .ZN(n5605) );
  AOI22_X1 U6748 ( .A1(n5687), .A2(n5983), .B1(REIP_REG_30__SCAN_IN), .B2(
        n5603), .ZN(n5604) );
  OAI211_X1 U6749 ( .C1(n5686), .C2(n3197), .A(n5605), .B(n5604), .ZN(U2797)
         );
  AOI22_X1 U6750 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6021), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6000), .ZN(n5606) );
  INV_X1 U6751 ( .A(n5606), .ZN(n5610) );
  OAI22_X1 U6752 ( .A1(n5608), .A2(n6017), .B1(n5607), .B2(n5616), .ZN(n5609)
         );
  AOI211_X1 U6753 ( .C1(n5611), .C2(n5983), .A(n5610), .B(n5609), .ZN(n5613)
         );
  OAI211_X1 U6754 ( .C1(n3223), .C2(n3197), .A(n5613), .B(n5612), .ZN(U2798)
         );
  AOI22_X1 U6755 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6000), .B1(n5614), 
        .B2(n6002), .ZN(n5615) );
  OAI21_X1 U6756 ( .B1(n6590), .B2(n5616), .A(n5615), .ZN(n5620) );
  OAI21_X1 U6757 ( .B1(n5618), .B2(n3197), .A(n3297), .ZN(n5619) );
  AOI211_X2 U6758 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6021), .A(n5620), .B(n5619), 
        .ZN(n5621) );
  OAI21_X1 U6759 ( .B1(n5690), .B2(n6015), .A(n5621), .ZN(U2799) );
  AOI22_X1 U6760 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6021), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6000), .ZN(n5626) );
  OAI22_X1 U6761 ( .A1(n5691), .A2(n3197), .B1(n5693), .B2(n6015), .ZN(n5622)
         );
  OAI211_X1 U6762 ( .C1(n5627), .C2(n6017), .A(n5626), .B(n5625), .ZN(U2800)
         );
  AOI22_X1 U6763 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6021), .B1(n5719), .B2(n6002), .ZN(n5633) );
  INV_X1 U6764 ( .A(n5723), .ZN(n5631) );
  INV_X1 U6765 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6585) );
  NOR2_X1 U6766 ( .A1(n6585), .A2(n5639), .ZN(n5634) );
  AOI21_X1 U6767 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5634), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5628) );
  OAI22_X1 U6768 ( .A1(n5629), .A2(n5628), .B1(n5695), .B2(n6015), .ZN(n5630)
         );
  AOI21_X1 U6769 ( .B1(n5631), .B2(n5978), .A(n5630), .ZN(n5632) );
  OAI211_X1 U6770 ( .C1(n6913), .C2(n6012), .A(n5633), .B(n5632), .ZN(U2801)
         );
  AOI22_X1 U6771 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6021), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6000), .ZN(n5643) );
  INV_X1 U6772 ( .A(n5730), .ZN(n5635) );
  INV_X1 U6773 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6755) );
  AOI22_X1 U6774 ( .A1(n5635), .A2(n6002), .B1(n5634), .B2(n6755), .ZN(n5642)
         );
  AOI21_X1 U6775 ( .B1(n5638), .B2(n5637), .A(n3253), .ZN(n5774) );
  AOI22_X1 U6776 ( .A1(n5983), .A2(n5774), .B1(n5978), .B2(n5727), .ZN(n5641)
         );
  NOR2_X1 U6777 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5639), .ZN(n5647) );
  OAI21_X1 U6778 ( .B1(n5647), .B2(n5653), .A(REIP_REG_25__SCAN_IN), .ZN(n5640) );
  NAND4_X1 U6779 ( .A1(n5643), .A2(n5642), .A3(n5641), .A4(n5640), .ZN(U2802)
         );
  AOI22_X1 U6780 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6021), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6000), .ZN(n5646) );
  AOI22_X1 U6781 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5653), .B1(n5644), .B2(
        n6002), .ZN(n5645) );
  OAI211_X1 U6782 ( .C1(n5699), .C2(n3197), .A(n5646), .B(n5645), .ZN(n5648)
         );
  NOR2_X1 U6783 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  OAI21_X1 U6784 ( .B1(n5698), .B2(n6015), .A(n5649), .ZN(U2803) );
  INV_X1 U6785 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6793) );
  OAI22_X1 U6786 ( .A1(n6793), .A2(n6012), .B1(n5650), .B2(n6017), .ZN(n5651)
         );
  AOI21_X1 U6787 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6021), .A(n5651), .ZN(n5657)
         );
  AOI22_X1 U6788 ( .A1(n5652), .A2(n5978), .B1(n5700), .B2(n5983), .ZN(n5656)
         );
  OAI21_X1 U6789 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5654), .A(n5653), .ZN(n5655) );
  NAND3_X1 U6790 ( .A1(n5657), .A2(n5656), .A3(n5655), .ZN(U2804) );
  NAND2_X1 U6791 ( .A1(n5658), .A2(n6581), .ZN(n5666) );
  AOI22_X1 U6792 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6000), .B1(n5731), 
        .B2(n6002), .ZN(n5659) );
  OAI21_X1 U6793 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5660), .A(n5659), .ZN(n5662) );
  OAI22_X1 U6794 ( .A1(n5734), .A2(n3197), .B1(n5704), .B2(n6015), .ZN(n5661)
         );
  AOI211_X1 U6795 ( .C1(EBX_REG_22__SCAN_IN), .C2(n6021), .A(n5662), .B(n5661), 
        .ZN(n5663) );
  OAI221_X1 U6796 ( .B1(n6874), .B2(n5668), .C1(n6874), .C2(n5666), .A(n5663), 
        .ZN(U2805) );
  INV_X1 U6797 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5742) );
  OAI22_X1 U6798 ( .A1(n5707), .A2(n5951), .B1(n5742), .B2(n6012), .ZN(n5665)
         );
  OAI22_X1 U6799 ( .A1(n5735), .A2(n6017), .B1(n6581), .B2(n5668), .ZN(n5664)
         );
  AOI211_X1 U6800 ( .C1(n5705), .C2(n5983), .A(n5665), .B(n5664), .ZN(n5667)
         );
  OAI211_X1 U6801 ( .C1(n3197), .C2(n5706), .A(n5667), .B(n5666), .ZN(U2806)
         );
  AOI21_X1 U6802 ( .B1(n6579), .B2(n5669), .A(n5668), .ZN(n5671) );
  OAI22_X1 U6803 ( .A1(n3890), .A2(n5951), .B1(n6780), .B2(n6012), .ZN(n5670)
         );
  AOI211_X1 U6804 ( .C1(n6002), .C2(n5672), .A(n5671), .B(n5670), .ZN(n5674)
         );
  AOI22_X1 U6805 ( .A1(n5983), .A2(n5709), .B1(n5978), .B2(n5714), .ZN(n5673)
         );
  NAND2_X1 U6806 ( .A1(n5674), .A2(n5673), .ZN(U2807) );
  AND2_X1 U6807 ( .A1(n5676), .A2(n5675), .ZN(n5875) );
  INV_X1 U6808 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U6809 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5677) );
  OAI211_X1 U6810 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5865), .B(n5677), .ZN(n5679) );
  NAND2_X1 U6811 ( .A1(n5678), .A2(n5965), .ZN(n5984) );
  OAI211_X1 U6812 ( .C1(n6012), .C2(n5680), .A(n5679), .B(n5984), .ZN(n5681)
         );
  AOI21_X1 U6813 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5875), .A(n5681), .ZN(n5685) );
  AOI21_X1 U6814 ( .B1(n5389), .B2(n5682), .A(n5432), .ZN(n5744) );
  OAI22_X1 U6815 ( .A1(n5711), .A2(n6015), .B1(n5747), .B2(n6017), .ZN(n5683)
         );
  AOI21_X1 U6816 ( .B1(n5978), .B2(n5744), .A(n5683), .ZN(n5684) );
  OAI211_X1 U6817 ( .C1(n5712), .C2(n5951), .A(n5685), .B(n5684), .ZN(U2808)
         );
  AOI22_X1 U6818 ( .A1(EBX_REG_30__SCAN_IN), .A2(n6068), .B1(n5687), .B2(n6071), .ZN(n5688) );
  OAI21_X1 U6819 ( .B1(n5686), .B2(n6083), .A(n5688), .ZN(U2829) );
  INV_X1 U6820 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5689) );
  OAI222_X1 U6821 ( .A1(n4541), .A2(n5690), .B1(n5689), .B2(n6081), .C1(n5618), 
        .C2(n6083), .ZN(U2831) );
  INV_X1 U6822 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5692) );
  OAI222_X1 U6823 ( .A1(n4541), .A2(n5693), .B1(n5692), .B2(n6081), .C1(n5691), 
        .C2(n6083), .ZN(U2832) );
  INV_X1 U6824 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5694) );
  OAI222_X1 U6825 ( .A1(n4541), .A2(n5695), .B1(n5694), .B2(n6081), .C1(n5723), 
        .C2(n6083), .ZN(U2833) );
  AOI22_X1 U6826 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6068), .B1(n6071), .B2(n5774), .ZN(n5696) );
  OAI21_X1 U6827 ( .B1(n6083), .B2(n5697), .A(n5696), .ZN(U2834) );
  INV_X1 U6828 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6837) );
  OAI222_X1 U6829 ( .A1(n6083), .A2(n5699), .B1(n6837), .B2(n6081), .C1(n5698), 
        .C2(n4541), .ZN(U2835) );
  AOI22_X1 U6830 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6068), .B1(n5700), .B2(n6071), .ZN(n5701) );
  OAI21_X1 U6831 ( .B1(n5702), .B2(n6083), .A(n5701), .ZN(U2836) );
  INV_X1 U6832 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5703) );
  OAI222_X1 U6833 ( .A1(n4541), .A2(n5704), .B1(n5703), .B2(n6081), .C1(n5734), 
        .C2(n6083), .ZN(U2837) );
  INV_X1 U6834 ( .A(n5705), .ZN(n5708) );
  OAI222_X1 U6835 ( .A1(n4541), .A2(n5708), .B1(n5707), .B2(n6081), .C1(n5706), 
        .C2(n6083), .ZN(U2838) );
  AOI22_X1 U6836 ( .A1(n6072), .A2(n5714), .B1(n6071), .B2(n5709), .ZN(n5710)
         );
  OAI21_X1 U6837 ( .B1(n6081), .B2(n3890), .A(n5710), .ZN(U2839) );
  INV_X1 U6838 ( .A(n5744), .ZN(n5713) );
  OAI222_X1 U6839 ( .A1(n5713), .A2(n6083), .B1(n5712), .B2(n6081), .C1(n4541), 
        .C2(n5711), .ZN(U2840) );
  AOI22_X1 U6840 ( .A1(n5714), .A2(n6086), .B1(n6085), .B2(DATAI_20_), .ZN(
        n5716) );
  AOI22_X1 U6841 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6089), .B1(n6088), .B2(
        DATAI_4_), .ZN(n5715) );
  NAND2_X1 U6842 ( .A1(n5716), .A2(n5715), .ZN(U2871) );
  AOI22_X1 U6843 ( .A1(n5744), .A2(n6086), .B1(n6085), .B2(DATAI_19_), .ZN(
        n5718) );
  AOI22_X1 U6844 ( .A1(EAX_REG_19__SCAN_IN), .A2(n6089), .B1(n6088), .B2(
        DATAI_3_), .ZN(n5717) );
  NAND2_X1 U6845 ( .A1(n5718), .A2(n5717), .ZN(U2872) );
  AOI22_X1 U6846 ( .A1(n6221), .A2(REIP_REG_26__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5722) );
  AOI22_X1 U6847 ( .A1(n5720), .A2(n6199), .B1(n6198), .B2(n5719), .ZN(n5721)
         );
  OAI211_X1 U6848 ( .C1(n6203), .C2(n5723), .A(n5722), .B(n5721), .ZN(U2960)
         );
  AOI22_X1 U6849 ( .A1(n6221), .A2(REIP_REG_25__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5729) );
  OAI21_X1 U6850 ( .B1(n5726), .B2(n5725), .A(n5724), .ZN(n5775) );
  AOI22_X1 U6851 ( .A1(n5727), .A2(n6189), .B1(n6199), .B2(n5775), .ZN(n5728)
         );
  OAI211_X1 U6852 ( .C1(n6193), .C2(n5730), .A(n5729), .B(n5728), .ZN(U2961)
         );
  AOI22_X1 U6853 ( .A1(n6221), .A2(REIP_REG_22__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5733) );
  OAI22_X1 U6854 ( .A1(n5736), .A2(n6179), .B1(n5735), .B2(n6193), .ZN(n5737)
         );
  OAI211_X1 U6855 ( .C1(n5742), .C2(n5741), .A(n5740), .B(n5739), .ZN(U2965)
         );
  AOI22_X1 U6856 ( .A1(n6221), .A2(REIP_REG_19__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5746) );
  AOI22_X1 U6857 ( .A1(n5744), .A2(n6189), .B1(n6199), .B2(n5743), .ZN(n5745)
         );
  OAI211_X1 U6858 ( .C1(n6193), .C2(n5747), .A(n5746), .B(n5745), .ZN(U2967)
         );
  AOI22_X1 U6859 ( .A1(n6221), .A2(REIP_REG_18__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5753) );
  INV_X1 U6860 ( .A(n5757), .ZN(n5748) );
  NOR3_X1 U6861 ( .A1(n5748), .A2(n5754), .A3(n5795), .ZN(n5760) );
  NOR3_X1 U6862 ( .A1(n5750), .A2(n3725), .A3(n5749), .ZN(n5758) );
  NOR2_X1 U6863 ( .A1(n5760), .A2(n5758), .ZN(n5751) );
  XNOR2_X1 U6864 ( .A(n5751), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5784)
         );
  AOI22_X1 U6865 ( .A1(n6199), .A2(n5784), .B1(n6198), .B2(n5869), .ZN(n5752)
         );
  OAI211_X1 U6866 ( .C1(n6203), .C2(n6029), .A(n5753), .B(n5752), .ZN(U2968)
         );
  AOI22_X1 U6867 ( .A1(n6221), .A2(REIP_REG_17__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5764) );
  NAND3_X1 U6868 ( .A1(n5748), .A2(n5754), .A3(n5805), .ZN(n5755) );
  AOI22_X1 U6869 ( .A1(n5757), .A2(n3725), .B1(n5755), .B2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5761) );
  INV_X1 U6870 ( .A(n5758), .ZN(n5759) );
  OAI21_X1 U6871 ( .B1(n5761), .B2(n5760), .A(n5759), .ZN(n5792) );
  AOI21_X1 U6872 ( .B1(n5394), .B2(n5762), .A(n5387), .ZN(n6087) );
  AOI22_X1 U6873 ( .A1(n6199), .A2(n5792), .B1(n6189), .B2(n6087), .ZN(n5763)
         );
  OAI211_X1 U6874 ( .C1(n6193), .C2(n5878), .A(n5764), .B(n5763), .ZN(U2969)
         );
  AOI22_X1 U6875 ( .A1(n6221), .A2(REIP_REG_16__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5769) );
  XNOR2_X1 U6876 ( .A(n3725), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5767)
         );
  XNOR2_X1 U6877 ( .A(n5766), .B(n5767), .ZN(n5800) );
  AOI22_X1 U6878 ( .A1(n5800), .A2(n6199), .B1(n6198), .B2(n5884), .ZN(n5768)
         );
  OAI211_X1 U6879 ( .C1(n6203), .C2(n6034), .A(n5769), .B(n5768), .ZN(U2970)
         );
  AOI22_X1 U6880 ( .A1(n6221), .A2(REIP_REG_14__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5772) );
  AOI22_X1 U6881 ( .A1(n5770), .A2(n6199), .B1(n6198), .B2(n5901), .ZN(n5771)
         );
  OAI211_X1 U6882 ( .C1(n6203), .C2(n6041), .A(n5772), .B(n5771), .ZN(U2972)
         );
  AOI22_X1 U6883 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6221), .B1(n5773), .B2(
        n5778), .ZN(n5777) );
  AOI22_X1 U6884 ( .A1(n5775), .A2(n3833), .B1(n5774), .B2(n6245), .ZN(n5776)
         );
  OAI211_X1 U6885 ( .C1(n5779), .C2(n5778), .A(n5777), .B(n5776), .ZN(U2993)
         );
  INV_X1 U6886 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5787) );
  NOR2_X1 U6887 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5795), .ZN(n5780)
         );
  AOI22_X1 U6888 ( .A1(n6221), .A2(REIP_REG_18__SCAN_IN), .B1(n5796), .B2(
        n5780), .ZN(n5786) );
  AOI21_X1 U6889 ( .B1(n5783), .B2(n5782), .A(n5781), .ZN(n6027) );
  AOI22_X1 U6890 ( .A1(n5784), .A2(n3833), .B1(n6245), .B2(n6027), .ZN(n5785)
         );
  OAI211_X1 U6891 ( .C1(n5788), .C2(n5787), .A(n5786), .B(n5785), .ZN(U3000)
         );
  AOI21_X1 U6892 ( .B1(n3249), .B2(n5799), .A(n5789), .ZN(n5791) );
  AOI22_X1 U6893 ( .A1(n5792), .A2(n3833), .B1(n6245), .B2(n3236), .ZN(n5798)
         );
  NOR2_X1 U6894 ( .A1(n6256), .A2(n6574), .ZN(n5793) );
  AOI221_X1 U6895 ( .B1(n5796), .B2(n5795), .C1(n5794), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5793), .ZN(n5797) );
  NAND2_X1 U6896 ( .A1(n5798), .A2(n5797), .ZN(U3001) );
  XNOR2_X1 U6897 ( .A(n5816), .B(n5799), .ZN(n6032) );
  AOI22_X1 U6898 ( .A1(n5800), .A2(n3833), .B1(n6245), .B2(n6032), .ZN(n5810)
         );
  NAND2_X1 U6899 ( .A1(n6221), .A2(REIP_REG_16__SCAN_IN), .ZN(n5809) );
  NOR3_X1 U6900 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5801), .A3(n5802), 
        .ZN(n5812) );
  INV_X1 U6901 ( .A(n5802), .ZN(n5803) );
  OAI21_X1 U6902 ( .B1(n5804), .B2(n5803), .A(n6219), .ZN(n5817) );
  OAI21_X1 U6903 ( .B1(n5812), .B2(n5817), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n5808) );
  NAND3_X1 U6904 ( .A1(n5806), .A2(n5805), .A3(n6215), .ZN(n5807) );
  NAND4_X1 U6905 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(U3002)
         );
  INV_X1 U6906 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6778) );
  NOR2_X1 U6907 ( .A1(n6256), .A2(n6778), .ZN(n5811) );
  AOI211_X1 U6908 ( .C1(n5813), .C2(n3833), .A(n5812), .B(n5811), .ZN(n5819)
         );
  NAND2_X1 U6909 ( .A1(n3217), .A2(n5814), .ZN(n5815) );
  AND2_X1 U6910 ( .A1(n5816), .A2(n5815), .ZN(n6035) );
  AOI22_X1 U6911 ( .A1(n5817), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .B1(n6245), .B2(n6035), .ZN(n5818) );
  NAND2_X1 U6912 ( .A1(n5819), .A2(n5818), .ZN(U3003) );
  INV_X1 U6913 ( .A(n5820), .ZN(n5832) );
  INV_X1 U6914 ( .A(n5923), .ZN(n5915) );
  OAI21_X1 U6915 ( .B1(n5915), .B2(n5914), .A(n5821), .ZN(n5824) );
  INV_X1 U6916 ( .A(n5822), .ZN(n5823) );
  NAND2_X1 U6917 ( .A1(n5824), .A2(n5823), .ZN(n6042) );
  INV_X1 U6918 ( .A(n5825), .ZN(n5826) );
  NAND3_X1 U6919 ( .A1(n5828), .A2(n5827), .A3(n5826), .ZN(n5829) );
  OAI211_X1 U6920 ( .C1(n6042), .C2(n6258), .A(n5830), .B(n5829), .ZN(n5831)
         );
  AOI21_X1 U6921 ( .B1(n5832), .B2(n3833), .A(n5831), .ZN(n5834) );
  OAI211_X1 U6922 ( .C1(n5835), .C2(n6752), .A(n5834), .B(n5833), .ZN(U3005)
         );
  NAND4_X1 U6923 ( .A1(n6006), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n5839)
         );
  OAI21_X1 U6924 ( .B1(n5841), .B2(n5840), .A(n5839), .ZN(U3455) );
  AOI21_X1 U6925 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6554), .A(n6545), .ZN(n5846) );
  INV_X1 U6926 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5842) );
  NOR2_X2 U6927 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6544), .ZN(n6631) );
  AOI21_X1 U6928 ( .B1(n5846), .B2(n5842), .A(n6631), .ZN(U2789) );
  OAI21_X1 U6929 ( .B1(n5843), .B2(n6529), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5844) );
  OAI21_X1 U6930 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6530), .A(n5844), .ZN(
        U2790) );
  NOR2_X1 U6931 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5847) );
  OAI21_X1 U6932 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5847), .A(n6629), .ZN(n5845)
         );
  OAI21_X1 U6933 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6629), .A(n5845), .ZN(
        U2791) );
  NOR2_X1 U6934 ( .A1(n6631), .A2(n5846), .ZN(n6602) );
  OAI21_X1 U6935 ( .B1(BS16_N), .B2(n5847), .A(n6602), .ZN(n6601) );
  OAI21_X1 U6936 ( .B1(n6602), .B2(n4392), .A(n6601), .ZN(U2792) );
  INV_X1 U6937 ( .A(n5848), .ZN(n5850) );
  OAI21_X1 U6938 ( .B1(n5850), .B2(n5849), .A(n6179), .ZN(U2793) );
  NOR4_X1 U6939 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5860) );
  NOR4_X1 U6940 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(
        n5859) );
  INV_X1 U6941 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6871) );
  INV_X1 U6942 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6794) );
  INV_X1 U6943 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6807) );
  INV_X1 U6944 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6895) );
  NAND4_X1 U6945 ( .A1(n6871), .A2(n6794), .A3(n6807), .A4(n6895), .ZN(n5857)
         );
  INV_X1 U6946 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6797) );
  INV_X1 U6947 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6852) );
  INV_X1 U6948 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6817) );
  INV_X1 U6949 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6823) );
  OAI211_X1 U6950 ( .C1(n6797), .C2(n6852), .A(n6817), .B(n6823), .ZN(n5856)
         );
  NOR4_X1 U6951 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5854) );
  NOR4_X1 U6952 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5853) );
  NOR4_X1 U6953 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5852) );
  NOR4_X1 U6954 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n5851) );
  NAND4_X1 U6955 ( .A1(n5854), .A2(n5853), .A3(n5852), .A4(n5851), .ZN(n5855)
         );
  NOR3_X1 U6956 ( .A1(n5857), .A2(n5856), .A3(n5855), .ZN(n5858) );
  NAND3_X1 U6957 ( .A1(n5860), .A2(n5859), .A3(n5858), .ZN(n6612) );
  NOR2_X1 U6958 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6612), .ZN(n6614) );
  INV_X1 U6959 ( .A(n6612), .ZN(n5861) );
  NOR2_X1 U6960 ( .A1(n5861), .A2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5862) );
  NAND4_X1 U6961 ( .A1(n5861), .A2(n6852), .A3(n6797), .A4(n6613), .ZN(n5863)
         );
  OAI21_X1 U6962 ( .B1(n6614), .B2(n5862), .A(n5863), .ZN(U2794) );
  AOI22_X1 U6963 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6612), .B1(n6614), 
        .B2(n6797), .ZN(n5864) );
  NAND2_X1 U6964 ( .A1(n5864), .A2(n5863), .ZN(U2795) );
  INV_X1 U6965 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6576) );
  AOI22_X1 U6966 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5875), .B1(n5865), .B2(
        n6576), .ZN(n5866) );
  OAI211_X1 U6967 ( .C1(n6012), .C2(n5867), .A(n5866), .B(n5984), .ZN(n5868)
         );
  AOI21_X1 U6968 ( .B1(EBX_REG_18__SCAN_IN), .B2(n6021), .A(n5868), .ZN(n5871)
         );
  AOI22_X1 U6969 ( .A1(n5869), .A2(n6002), .B1(n5983), .B2(n6027), .ZN(n5870)
         );
  OAI211_X1 U6970 ( .C1(n3197), .C2(n6029), .A(n5871), .B(n5870), .ZN(U2809)
         );
  NAND2_X1 U6971 ( .A1(n6574), .A2(n5872), .ZN(n5874) );
  INV_X1 U6972 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6782) );
  OAI22_X1 U6973 ( .A1(n6031), .A2(n5951), .B1(n6782), .B2(n6012), .ZN(n5873)
         );
  AOI211_X1 U6974 ( .C1(n5875), .C2(n5874), .A(n5999), .B(n5873), .ZN(n5877)
         );
  AOI22_X1 U6975 ( .A1(n5983), .A2(n3236), .B1(n5978), .B2(n6087), .ZN(n5876)
         );
  OAI211_X1 U6976 ( .C1(n5878), .C2(n6017), .A(n5877), .B(n5876), .ZN(U2810)
         );
  NOR3_X1 U6977 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5993), .A3(n5879), .ZN(n5883) );
  INV_X1 U6978 ( .A(n5880), .ZN(n5895) );
  NOR3_X1 U6979 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5993), .A3(n5895), .ZN(n5889) );
  OAI21_X1 U6980 ( .B1(n5880), .B2(n5993), .A(n5965), .ZN(n5893) );
  OAI21_X1 U6981 ( .B1(n5889), .B2(n5893), .A(REIP_REG_16__SCAN_IN), .ZN(n5881) );
  OAI211_X1 U6982 ( .C1(n6012), .C2(n6766), .A(n5984), .B(n5881), .ZN(n5882)
         );
  AOI211_X1 U6983 ( .C1(n6021), .C2(EBX_REG_16__SCAN_IN), .A(n5883), .B(n5882), 
        .ZN(n5886) );
  AOI22_X1 U6984 ( .A1(n5884), .A2(n6002), .B1(n5983), .B2(n6032), .ZN(n5885)
         );
  OAI211_X1 U6985 ( .C1(n3197), .C2(n6034), .A(n5886), .B(n5885), .ZN(U2811)
         );
  AOI22_X1 U6986 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6021), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5893), .ZN(n5887) );
  OAI211_X1 U6987 ( .C1(n6012), .C2(n6933), .A(n5887), .B(n5984), .ZN(n5888)
         );
  AOI211_X1 U6988 ( .C1(n6035), .C2(n5983), .A(n5889), .B(n5888), .ZN(n5892)
         );
  NAND2_X1 U6989 ( .A1(n5890), .A2(n6002), .ZN(n5891) );
  OAI211_X1 U6990 ( .C1(n6038), .C2(n3197), .A(n5892), .B(n5891), .ZN(U2812)
         );
  INV_X1 U6991 ( .A(n5893), .ZN(n5894) );
  OAI22_X1 U6992 ( .A1(n5894), .A2(n6570), .B1(n6015), .B2(n6039), .ZN(n5900)
         );
  NAND2_X1 U6993 ( .A1(n5997), .A2(n5895), .ZN(n5897) );
  AOI22_X1 U6994 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6021), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6000), .ZN(n5896) );
  OAI211_X1 U6995 ( .C1(n5898), .C2(n5897), .A(n5896), .B(n5984), .ZN(n5899)
         );
  AOI211_X1 U6996 ( .C1(n5901), .C2(n6002), .A(n5900), .B(n5899), .ZN(n5902)
         );
  OAI21_X1 U6997 ( .B1(n3197), .B2(n6041), .A(n5902), .ZN(U2813) );
  OAI22_X1 U6998 ( .A1(n6043), .A2(n5951), .B1(n6015), .B2(n6042), .ZN(n5903)
         );
  AOI211_X1 U6999 ( .C1(n6000), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5999), 
        .B(n5903), .ZN(n5913) );
  AOI22_X1 U7000 ( .A1(n5905), .A2(n6002), .B1(n5978), .B2(n5904), .ZN(n5912)
         );
  INV_X1 U7001 ( .A(n5906), .ZN(n5907) );
  OAI21_X1 U7002 ( .B1(n5907), .B2(n5993), .A(n5965), .ZN(n5929) );
  NAND3_X1 U7003 ( .A1(n6568), .A2(n5997), .A3(n5907), .ZN(n5920) );
  INV_X1 U7004 ( .A(n5920), .ZN(n5908) );
  OAI21_X1 U7005 ( .B1(n5929), .B2(n5908), .A(REIP_REG_13__SCAN_IN), .ZN(n5911) );
  INV_X1 U7006 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6951) );
  NAND3_X1 U7007 ( .A1(n5997), .A2(n5909), .A3(n6951), .ZN(n5910) );
  NAND4_X1 U7008 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(U2814)
         );
  AOI22_X1 U7009 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6021), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5929), .ZN(n5922) );
  XNOR2_X1 U7010 ( .A(n5915), .B(n5914), .ZN(n6207) );
  OAI22_X1 U7011 ( .A1(n5916), .A2(n6012), .B1(n6015), .B2(n6207), .ZN(n5917)
         );
  AOI211_X1 U7012 ( .C1(n5978), .C2(n6045), .A(n5999), .B(n5917), .ZN(n5921)
         );
  NAND2_X1 U7013 ( .A1(n5918), .A2(n6002), .ZN(n5919) );
  NAND4_X1 U7014 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(U2815)
         );
  AOI21_X1 U7015 ( .B1(n5925), .B2(n5924), .A(n5923), .ZN(n6214) );
  AOI22_X1 U7016 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6021), .B1(n5983), .B2(n6214), .ZN(n5926) );
  OAI211_X1 U7017 ( .C1(n6012), .C2(n5927), .A(n5926), .B(n5984), .ZN(n5928)
         );
  AOI21_X1 U7018 ( .B1(n6160), .B2(n6002), .A(n5928), .ZN(n5932) );
  OAI221_X1 U7019 ( .B1(REIP_REG_11__SCAN_IN), .B2(n5997), .C1(
        REIP_REG_11__SCAN_IN), .C2(n5930), .A(n5929), .ZN(n5931) );
  OAI211_X1 U7020 ( .C1(n6163), .C2(n3197), .A(n5932), .B(n5931), .ZN(U2816)
         );
  AOI22_X1 U7021 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6021), .B1(n5983), .B2(n6048), .ZN(n5941) );
  NOR3_X1 U7022 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5993), .A3(n5933), .ZN(n5934) );
  AOI211_X1 U7023 ( .C1(n6000), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5999), 
        .B(n5934), .ZN(n5940) );
  AOI22_X1 U7024 ( .A1(n5936), .A2(n6002), .B1(n5978), .B2(n5935), .ZN(n5939)
         );
  OAI21_X1 U7025 ( .B1(n5937), .B2(n5993), .A(n5965), .ZN(n5956) );
  INV_X1 U7026 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6783) );
  AND3_X1 U7027 ( .A1(n6783), .A2(n5997), .A3(n5937), .ZN(n5942) );
  OAI21_X1 U7028 ( .B1(n5956), .B2(n5942), .A(REIP_REG_10__SCAN_IN), .ZN(n5938) );
  NAND4_X1 U7029 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(U2817)
         );
  AOI21_X1 U7030 ( .B1(n5956), .B2(REIP_REG_9__SCAN_IN), .A(n5942), .ZN(n5950)
         );
  OR2_X1 U7031 ( .A1(n5944), .A2(n5943), .ZN(n5946) );
  AND2_X1 U7032 ( .A1(n5946), .A2(n5945), .ZN(n6222) );
  AOI22_X1 U7033 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6000), .B1(n5983), 
        .B2(n6222), .ZN(n5947) );
  OAI211_X1 U7034 ( .C1(n3197), .C2(n6169), .A(n5947), .B(n5984), .ZN(n5948)
         );
  AOI21_X1 U7035 ( .B1(n6166), .B2(n6002), .A(n5948), .ZN(n5949) );
  OAI211_X1 U7036 ( .C1(n6053), .C2(n5951), .A(n5950), .B(n5949), .ZN(U2818)
         );
  OAI22_X1 U7037 ( .A1(n5952), .A2(n6012), .B1(n6015), .B2(n6054), .ZN(n5953)
         );
  AOI211_X1 U7038 ( .C1(n6021), .C2(EBX_REG_8__SCAN_IN), .A(n5999), .B(n5953), 
        .ZN(n5959) );
  OAI21_X1 U7039 ( .B1(n5993), .B2(n5954), .A(n6563), .ZN(n5955) );
  AOI22_X1 U7040 ( .A1(n5957), .A2(n6002), .B1(n5956), .B2(n5955), .ZN(n5958)
         );
  OAI211_X1 U7041 ( .C1(n3197), .C2(n6056), .A(n5959), .B(n5958), .ZN(U2819)
         );
  INV_X1 U7042 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5968) );
  OAI21_X1 U7043 ( .B1(n5962), .B2(n5961), .A(n5960), .ZN(n5964) );
  AND2_X1 U7044 ( .A1(n5964), .A2(n5963), .ZN(n6230) );
  OAI21_X1 U7045 ( .B1(n5966), .B2(n5993), .A(n5965), .ZN(n5989) );
  AOI22_X1 U7046 ( .A1(n5983), .A2(n6230), .B1(REIP_REG_7__SCAN_IN), .B2(n5989), .ZN(n5967) );
  OAI211_X1 U7047 ( .C1(n6012), .C2(n5968), .A(n5967), .B(n5984), .ZN(n5971)
         );
  OAI22_X1 U7048 ( .A1(n6173), .A2(n6017), .B1(n3197), .B2(n6177), .ZN(n5970)
         );
  AOI211_X1 U7049 ( .C1(EBX_REG_7__SCAN_IN), .C2(n6021), .A(n5971), .B(n5970), 
        .ZN(n5973) );
  INV_X1 U7050 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6561) );
  NOR4_X1 U7051 ( .A1(n5993), .A2(n6855), .A3(n6559), .A4(n5996), .ZN(n5976)
         );
  OAI221_X1 U7052 ( .B1(REIP_REG_6__SCAN_IN), .B2(REIP_REG_7__SCAN_IN), .C1(
        n4748), .C2(n6561), .A(n5976), .ZN(n5972) );
  NAND2_X1 U7053 ( .A1(n5973), .A2(n5972), .ZN(U2820) );
  AOI22_X1 U7054 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6021), .B1(n5983), .B2(n6059), 
        .ZN(n5974) );
  OAI211_X1 U7055 ( .C1(n6012), .C2(n6921), .A(n5974), .B(n5984), .ZN(n5975)
         );
  AOI221_X1 U7056 ( .B1(n5976), .B2(n4748), .C1(n5989), .C2(
        REIP_REG_6__SCAN_IN), .A(n5975), .ZN(n5981) );
  AOI22_X1 U7057 ( .A1(n5979), .A2(n6002), .B1(n5978), .B2(n5977), .ZN(n5980)
         );
  NAND2_X1 U7058 ( .A1(n5981), .A2(n5980), .ZN(U2821) );
  INV_X1 U7059 ( .A(n6184), .ZN(n5988) );
  INV_X1 U7060 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5986) );
  INV_X1 U7061 ( .A(n5982), .ZN(n6062) );
  AOI22_X1 U7062 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6021), .B1(n5983), .B2(n6062), 
        .ZN(n5985) );
  OAI211_X1 U7063 ( .C1(n6012), .C2(n5986), .A(n5985), .B(n5984), .ZN(n5987)
         );
  AOI21_X1 U7064 ( .B1(n6004), .B2(n5988), .A(n5987), .ZN(n5992) );
  NOR3_X1 U7065 ( .A1(n5993), .A2(n6855), .A3(n5996), .ZN(n5990) );
  OAI21_X1 U7066 ( .B1(REIP_REG_5__SCAN_IN), .B2(n5990), .A(n5989), .ZN(n5991)
         );
  OAI211_X1 U7067 ( .C1(n6017), .C2(n6178), .A(n5992), .B(n5991), .ZN(U2822)
         );
  NOR2_X1 U7068 ( .A1(n5993), .A2(n5996), .ZN(n5994) );
  AOI22_X1 U7069 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6021), .B1(n5994), .B2(n6855), 
        .ZN(n6010) );
  AOI21_X1 U7070 ( .B1(n5997), .B2(n5996), .A(n5995), .ZN(n6024) );
  OAI22_X1 U7071 ( .A1(n6024), .A2(n6855), .B1(n6015), .B2(n6066), .ZN(n5998)
         );
  AOI211_X1 U7072 ( .C1(n6000), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5999), 
        .B(n5998), .ZN(n6009) );
  INV_X1 U7073 ( .A(n6001), .ZN(n6003) );
  AOI22_X1 U7074 ( .A1(n6004), .A2(n6064), .B1(n6003), .B2(n6002), .ZN(n6008)
         );
  NAND2_X1 U7075 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  NAND4_X1 U7076 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(U2823)
         );
  INV_X1 U7077 ( .A(n6067), .ZN(n6014) );
  OAI222_X1 U7078 ( .A1(n6015), .A2(n6014), .B1(n6013), .B2(n6437), .C1(n6012), 
        .C2(n6011), .ZN(n6020) );
  OAI22_X1 U7079 ( .A1(n6018), .A2(n6070), .B1(n6017), .B2(n6016), .ZN(n6019)
         );
  AOI211_X1 U7080 ( .C1(EBX_REG_3__SCAN_IN), .C2(n6021), .A(n6020), .B(n6019), 
        .ZN(n6022) );
  OAI221_X1 U7081 ( .B1(n6024), .B2(n6556), .C1(n6024), .C2(n6023), .A(n6022), 
        .ZN(U2824) );
  OAI22_X1 U7082 ( .A1(n6081), .A2(n6026), .B1(n6025), .B2(n4541), .ZN(U2828)
         );
  AOI22_X1 U7083 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6068), .B1(n6071), .B2(n6027), .ZN(n6028) );
  OAI21_X1 U7084 ( .B1(n6083), .B2(n6029), .A(n6028), .ZN(U2841) );
  AOI22_X1 U7085 ( .A1(n6072), .A2(n6087), .B1(n6071), .B2(n3236), .ZN(n6030)
         );
  OAI21_X1 U7086 ( .B1(n6081), .B2(n6031), .A(n6030), .ZN(U2842) );
  AOI22_X1 U7087 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6068), .B1(n6071), .B2(n6032), .ZN(n6033) );
  OAI21_X1 U7088 ( .B1(n6083), .B2(n6034), .A(n6033), .ZN(U2843) );
  INV_X1 U7089 ( .A(n6035), .ZN(n6036) );
  OAI222_X1 U7090 ( .A1(n6038), .A2(n6083), .B1(n6037), .B2(n6081), .C1(n4541), 
        .C2(n6036), .ZN(U2844) );
  INV_X1 U7091 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6040) );
  OAI222_X1 U7092 ( .A1(n6041), .A2(n6083), .B1(n6040), .B2(n6081), .C1(n4541), 
        .C2(n6039), .ZN(U2845) );
  OAI222_X1 U7093 ( .A1(n6044), .A2(n6083), .B1(n6043), .B2(n6081), .C1(n4541), 
        .C2(n6042), .ZN(U2846) );
  AOI22_X1 U7094 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6068), .B1(n6072), .B2(n6045), .ZN(n6046) );
  OAI21_X1 U7095 ( .B1(n4541), .B2(n6207), .A(n6046), .ZN(U2847) );
  AOI22_X1 U7096 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6068), .B1(n6071), .B2(n6214), .ZN(n6047) );
  OAI21_X1 U7097 ( .B1(n6083), .B2(n6163), .A(n6047), .ZN(U2848) );
  INV_X1 U7098 ( .A(n6048), .ZN(n6049) );
  OAI222_X1 U7099 ( .A1(n6051), .A2(n6083), .B1(n6050), .B2(n6081), .C1(n4541), 
        .C2(n6049), .ZN(U2849) );
  INV_X1 U7100 ( .A(n6222), .ZN(n6052) );
  OAI222_X1 U7101 ( .A1(n6169), .A2(n6083), .B1(n6053), .B2(n6081), .C1(n4541), 
        .C2(n6052), .ZN(U2850) );
  INV_X1 U7102 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6055) );
  OAI222_X1 U7103 ( .A1(n6056), .A2(n6083), .B1(n6055), .B2(n6081), .C1(n4541), 
        .C2(n6054), .ZN(U2851) );
  INV_X1 U7104 ( .A(n6230), .ZN(n6057) );
  OAI222_X1 U7105 ( .A1(n6177), .A2(n6083), .B1(n6058), .B2(n6081), .C1(n4541), 
        .C2(n6057), .ZN(U2852) );
  AOI22_X1 U7106 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6068), .B1(n6071), .B2(n6059), 
        .ZN(n6060) );
  OAI21_X1 U7107 ( .B1(n6083), .B2(n6061), .A(n6060), .ZN(U2853) );
  AOI22_X1 U7108 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6068), .B1(n6071), .B2(n6062), 
        .ZN(n6063) );
  OAI21_X1 U7109 ( .B1(n6083), .B2(n6184), .A(n6063), .ZN(U2854) );
  AOI22_X1 U7110 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6068), .B1(n6072), .B2(n6064), 
        .ZN(n6065) );
  OAI21_X1 U7111 ( .B1(n4541), .B2(n6066), .A(n6065), .ZN(U2855) );
  AOI22_X1 U7112 ( .A1(EBX_REG_3__SCAN_IN), .A2(n6068), .B1(n6071), .B2(n6067), 
        .ZN(n6069) );
  OAI21_X1 U7113 ( .B1(n6083), .B2(n6070), .A(n6069), .ZN(U2856) );
  AOI22_X1 U7114 ( .A1(n6072), .A2(n6188), .B1(n6071), .B2(n6244), .ZN(n6073)
         );
  OAI21_X1 U7115 ( .B1(n6081), .B2(n6074), .A(n6073), .ZN(U2857) );
  INV_X1 U7116 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7117 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  AND2_X1 U7118 ( .A1(n6078), .A2(n6077), .ZN(n6257) );
  OAI222_X1 U7119 ( .A1(n6202), .A2(n6083), .B1(n6079), .B2(n6081), .C1(n4541), 
        .C2(n6257), .ZN(U2858) );
  OAI222_X1 U7120 ( .A1(n6084), .A2(n6083), .B1(n6082), .B2(n6081), .C1(n4541), 
        .C2(n6080), .ZN(U2859) );
  AOI22_X1 U7121 ( .A1(n6087), .A2(n6086), .B1(n6085), .B2(DATAI_17_), .ZN(
        n6091) );
  AOI22_X1 U7122 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6089), .B1(n6088), .B2(
        DATAI_1_), .ZN(n6090) );
  NAND2_X1 U7123 ( .A1(n6091), .A2(n6090), .ZN(U2874) );
  INV_X1 U7124 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n6094) );
  AOI22_X1 U7125 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6110), .B1(n6144), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U7126 ( .B1(n6619), .B2(n6094), .A(n6093), .ZN(U2893) );
  INV_X1 U7127 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6096) );
  AOI22_X1 U7128 ( .A1(n3193), .A2(UWORD_REG_13__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7129 ( .B1(n6096), .B2(n6117), .A(n6095), .ZN(U2894) );
  INV_X1 U7130 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6098) );
  AOI22_X1 U7131 ( .A1(n3193), .A2(UWORD_REG_12__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7132 ( .B1(n6098), .B2(n6117), .A(n6097), .ZN(U2895) );
  INV_X1 U7133 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6100) );
  AOI22_X1 U7134 ( .A1(n3193), .A2(UWORD_REG_11__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n6099) );
  OAI21_X1 U7135 ( .B1(n6100), .B2(n6117), .A(n6099), .ZN(U2896) );
  INV_X1 U7136 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6882) );
  AOI22_X1 U7137 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6110), .B1(n3193), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6101) );
  OAI21_X1 U7138 ( .B1(n6882), .B2(n6126), .A(n6101), .ZN(U2897) );
  INV_X1 U7139 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6103) );
  AOI22_X1 U7140 ( .A1(n3193), .A2(UWORD_REG_9__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n6102) );
  OAI21_X1 U7141 ( .B1(n6103), .B2(n6117), .A(n6102), .ZN(U2898) );
  INV_X1 U7142 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n6916) );
  AOI22_X1 U7143 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6110), .B1(n3193), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7144 ( .B1(n6916), .B2(n6126), .A(n6104), .ZN(U2899) );
  INV_X1 U7145 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n6872) );
  INV_X1 U7146 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6958) );
  INV_X1 U7147 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6105) );
  OAI222_X1 U7148 ( .A1(n6126), .A2(n6872), .B1(n6117), .B2(n6958), .C1(n6619), 
        .C2(n6105), .ZN(U2900) );
  INV_X1 U7149 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6107) );
  AOI22_X1 U7150 ( .A1(n3193), .A2(UWORD_REG_6__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n6106) );
  OAI21_X1 U7151 ( .B1(n6107), .B2(n6117), .A(n6106), .ZN(U2901) );
  AOI22_X1 U7152 ( .A1(n3193), .A2(UWORD_REG_5__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n6108) );
  OAI21_X1 U7153 ( .B1(n6109), .B2(n6117), .A(n6108), .ZN(U2902) );
  INV_X1 U7154 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6946) );
  AOI22_X1 U7155 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6110), .B1(n3193), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7156 ( .B1(n6946), .B2(n6126), .A(n6111), .ZN(U2903) );
  INV_X1 U7157 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U7158 ( .A1(n3193), .A2(UWORD_REG_3__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7159 ( .B1(n6866), .B2(n6117), .A(n6112), .ZN(U2904) );
  INV_X1 U7160 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6114) );
  AOI22_X1 U7161 ( .A1(n3193), .A2(UWORD_REG_2__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7162 ( .B1(n6114), .B2(n6117), .A(n6113), .ZN(U2905) );
  INV_X1 U7163 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n6901) );
  INV_X1 U7164 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6115) );
  INV_X1 U7165 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6769) );
  OAI222_X1 U7166 ( .A1(n6126), .A2(n6901), .B1(n6117), .B2(n6115), .C1(n6619), 
        .C2(n6769), .ZN(U2906) );
  INV_X1 U7167 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6118) );
  AOI22_X1 U7168 ( .A1(n3193), .A2(UWORD_REG_0__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U7169 ( .B1(n6118), .B2(n6117), .A(n6116), .ZN(U2907) );
  INV_X1 U7170 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6961) );
  AOI22_X1 U7171 ( .A1(n3193), .A2(LWORD_REG_15__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6119) );
  OAI21_X1 U7172 ( .B1(n6961), .B2(n6146), .A(n6119), .ZN(U2908) );
  AOI22_X1 U7173 ( .A1(n3193), .A2(LWORD_REG_14__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7174 ( .B1(n6121), .B2(n6146), .A(n6120), .ZN(U2909) );
  AOI22_X1 U7175 ( .A1(n3193), .A2(LWORD_REG_13__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6122) );
  OAI21_X1 U7176 ( .B1(n6832), .B2(n6146), .A(n6122), .ZN(U2910) );
  INV_X1 U7177 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6948) );
  AOI22_X1 U7178 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6136), .B1(n6144), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7179 ( .B1(n6619), .B2(n6948), .A(n6123), .ZN(U2911) );
  INV_X1 U7180 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6836) );
  INV_X1 U7181 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6124) );
  OAI222_X1 U7182 ( .A1(n6126), .A2(n6836), .B1(n6146), .B2(n6886), .C1(n6619), 
        .C2(n6124), .ZN(U2912) );
  INV_X1 U7183 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6858) );
  AOI22_X1 U7184 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6136), .B1(n3193), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U7185 ( .B1(n6858), .B2(n6126), .A(n6125), .ZN(U2913) );
  AOI22_X1 U7186 ( .A1(n3193), .A2(LWORD_REG_9__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6127) );
  OAI21_X1 U7187 ( .B1(n6128), .B2(n6146), .A(n6127), .ZN(U2914) );
  AOI22_X1 U7188 ( .A1(n3193), .A2(LWORD_REG_8__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6129) );
  OAI21_X1 U7189 ( .B1(n6130), .B2(n6146), .A(n6129), .ZN(U2915) );
  AOI22_X1 U7190 ( .A1(n3193), .A2(LWORD_REG_7__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6131) );
  OAI21_X1 U7191 ( .B1(n6132), .B2(n6146), .A(n6131), .ZN(U2916) );
  AOI22_X1 U7192 ( .A1(n3193), .A2(LWORD_REG_6__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6133) );
  OAI21_X1 U7193 ( .B1(n6134), .B2(n6146), .A(n6133), .ZN(U2917) );
  AOI22_X1 U7194 ( .A1(n3193), .A2(LWORD_REG_5__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6135) );
  OAI21_X1 U7195 ( .B1(n6867), .B2(n6146), .A(n6135), .ZN(U2918) );
  AOI222_X1 U7196 ( .A1(n3193), .A2(LWORD_REG_4__SCAN_IN), .B1(n6136), .B2(
        EAX_REG_4__SCAN_IN), .C1(DATAO_REG_4__SCAN_IN), .C2(n6144), .ZN(n6137)
         );
  INV_X1 U7197 ( .A(n6137), .ZN(U2919) );
  AOI22_X1 U7198 ( .A1(n3193), .A2(LWORD_REG_3__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7199 ( .B1(n6139), .B2(n6146), .A(n6138), .ZN(U2920) );
  AOI22_X1 U7200 ( .A1(n3193), .A2(LWORD_REG_2__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7201 ( .B1(n6141), .B2(n6146), .A(n6140), .ZN(U2921) );
  AOI22_X1 U7202 ( .A1(n3193), .A2(LWORD_REG_1__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7203 ( .B1(n6143), .B2(n6146), .A(n6142), .ZN(U2922) );
  AOI22_X1 U7204 ( .A1(n3193), .A2(LWORD_REG_0__SCAN_IN), .B1(n6144), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6145) );
  OAI21_X1 U7205 ( .B1(n6147), .B2(n6146), .A(n6145), .ZN(U2923) );
  AOI22_X1 U7206 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6149), .B1(n6152), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7207 ( .A1(n6153), .A2(DATAI_10_), .ZN(n6150) );
  NAND2_X1 U7208 ( .A1(n6148), .A2(n6150), .ZN(U2934) );
  AOI22_X1 U7209 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6149), .B1(n6152), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7210 ( .A1(n6151), .A2(n6150), .ZN(U2949) );
  AOI22_X1 U7211 ( .A1(n6153), .A2(DATAI_15_), .B1(n6152), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6154) );
  OAI21_X1 U7212 ( .B1(n6961), .B2(n6155), .A(n6154), .ZN(U2954) );
  AOI22_X1 U7213 ( .A1(n6221), .A2(REIP_REG_11__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7214 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  XNOR2_X1 U7215 ( .A(n6156), .B(n6159), .ZN(n6216) );
  AOI22_X1 U7216 ( .A1(n6199), .A2(n6216), .B1(n6198), .B2(n6160), .ZN(n6161)
         );
  OAI211_X1 U7217 ( .C1(n6203), .C2(n6163), .A(n6162), .B(n6161), .ZN(U2975)
         );
  AOI22_X1 U7218 ( .A1(n6221), .A2(REIP_REG_9__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6168) );
  XNOR2_X1 U7219 ( .A(n3725), .B(n6227), .ZN(n6165) );
  XNOR2_X1 U7220 ( .A(n6164), .B(n6165), .ZN(n6223) );
  AOI22_X1 U7221 ( .A1(n6223), .A2(n6199), .B1(n6198), .B2(n6166), .ZN(n6167)
         );
  OAI211_X1 U7222 ( .C1(n6203), .C2(n6169), .A(n6168), .B(n6167), .ZN(U2977)
         );
  NOR2_X1 U7223 ( .A1(n6256), .A2(n6561), .ZN(n6229) );
  INV_X1 U7224 ( .A(n6171), .ZN(n6172) );
  XNOR2_X1 U7225 ( .A(n3194), .B(n6172), .ZN(n6231) );
  INV_X1 U7226 ( .A(n6231), .ZN(n6174) );
  OAI22_X1 U7227 ( .A1(n6174), .A2(n6179), .B1(n6173), .B2(n6193), .ZN(n6175)
         );
  AOI211_X1 U7228 ( .C1(PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n6194), .A(n6229), 
        .B(n6175), .ZN(n6176) );
  OAI21_X1 U7229 ( .B1(n6203), .B2(n6177), .A(n6176), .ZN(U2979) );
  OAI22_X1 U7230 ( .A1(n6180), .A2(n6179), .B1(n6178), .B2(n6193), .ZN(n6181)
         );
  AOI211_X1 U7231 ( .C1(PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n6194), .A(n6182), 
        .B(n6181), .ZN(n6183) );
  OAI21_X1 U7232 ( .B1(n6203), .B2(n6184), .A(n6183), .ZN(U2981) );
  AOI22_X1 U7233 ( .A1(n6221), .A2(REIP_REG_2__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6191) );
  XNOR2_X1 U7234 ( .A(n6185), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6186)
         );
  XNOR2_X1 U7235 ( .A(n6187), .B(n6186), .ZN(n6249) );
  AOI22_X1 U7236 ( .A1(n6189), .A2(n6188), .B1(n6249), .B2(n6199), .ZN(n6190)
         );
  OAI211_X1 U7237 ( .C1(n6193), .C2(n6192), .A(n6191), .B(n6190), .ZN(U2984)
         );
  AOI22_X1 U7238 ( .A1(n6221), .A2(REIP_REG_1__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6201) );
  INV_X1 U7239 ( .A(n6197), .ZN(n6260) );
  AOI22_X1 U7240 ( .A1(n6260), .A2(n6199), .B1(n6198), .B2(n5349), .ZN(n6200)
         );
  OAI211_X1 U7241 ( .C1(n6203), .C2(n6202), .A(n6201), .B(n6200), .ZN(U2985)
         );
  AOI21_X1 U7242 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6215), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6213) );
  INV_X1 U7243 ( .A(n6243), .ZN(n6206) );
  OAI21_X1 U7244 ( .B1(n6206), .B2(n6205), .A(n6204), .ZN(n6212) );
  OAI22_X1 U7245 ( .A1(n6209), .A2(n6208), .B1(n6207), .B2(n6258), .ZN(n6210)
         );
  AOI21_X1 U7246 ( .B1(n6221), .B2(REIP_REG_12__SCAN_IN), .A(n6210), .ZN(n6211) );
  OAI221_X1 U7247 ( .B1(n6213), .B2(n6219), .C1(n6213), .C2(n6212), .A(n6211), 
        .ZN(U3006) );
  AOI22_X1 U7248 ( .A1(n6214), .A2(n6245), .B1(n6221), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6218) );
  AOI22_X1 U7249 ( .A1(n6216), .A2(n3833), .B1(n6215), .B2(n6765), .ZN(n6217)
         );
  OAI211_X1 U7250 ( .C1(n6219), .C2(n6765), .A(n6218), .B(n6217), .ZN(U3007)
         );
  INV_X1 U7251 ( .A(n6220), .ZN(n6228) );
  AOI22_X1 U7252 ( .A1(n6222), .A2(n6245), .B1(n6221), .B2(REIP_REG_9__SCAN_IN), .ZN(n6226) );
  AOI22_X1 U7253 ( .A1(n6224), .A2(n6227), .B1(n6223), .B2(n3833), .ZN(n6225)
         );
  OAI211_X1 U7254 ( .C1(n6228), .C2(n6227), .A(n6226), .B(n6225), .ZN(U3009)
         );
  AOI21_X1 U7255 ( .B1(n6230), .B2(n6245), .A(n6229), .ZN(n6233) );
  NAND2_X1 U7256 ( .A1(n6231), .A2(n3833), .ZN(n6232) );
  OAI211_X1 U7257 ( .C1(n6234), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6233), 
        .B(n6232), .ZN(n6235) );
  INV_X1 U7258 ( .A(n6235), .ZN(n6236) );
  OAI21_X1 U7259 ( .B1(n6238), .B2(n6237), .A(n6236), .ZN(U3011) );
  INV_X1 U7260 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6555) );
  OAI21_X1 U7261 ( .B1(n6240), .B2(n3844), .A(n6239), .ZN(n6241) );
  INV_X1 U7262 ( .A(n6241), .ZN(n6242) );
  OR2_X1 U7263 ( .A1(n6243), .A2(n6242), .ZN(n6247) );
  NAND2_X1 U7264 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  OAI211_X1 U7265 ( .C1(n6555), .C2(n6256), .A(n6247), .B(n6246), .ZN(n6248)
         );
  INV_X1 U7266 ( .A(n6248), .ZN(n6252) );
  AOI22_X1 U7267 ( .A1(n6250), .A2(n3844), .B1(n3833), .B2(n6249), .ZN(n6251)
         );
  OAI211_X1 U7268 ( .C1(n6253), .C2(n3844), .A(n6252), .B(n6251), .ZN(U3016)
         );
  NAND2_X1 U7269 ( .A1(n6255), .A2(n6254), .ZN(n6263) );
  INV_X1 U7270 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6607) );
  OAI22_X1 U7271 ( .A1(n6258), .A2(n6257), .B1(n6607), .B2(n6256), .ZN(n6259)
         );
  AOI21_X1 U7272 ( .B1(n6260), .B2(n3833), .A(n6259), .ZN(n6261) );
  OAI221_X1 U7273 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6263), .C1(n3536), .C2(n6262), .A(n6261), .ZN(U3017) );
  NOR2_X1 U7274 ( .A1(n6265), .A2(n6264), .ZN(U3019) );
  INV_X1 U7275 ( .A(n6266), .ZN(n6276) );
  OR2_X1 U7276 ( .A1(n6267), .A2(n3982), .ZN(n6269) );
  NOR2_X1 U7277 ( .A1(n6392), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6299)
         );
  INV_X1 U7278 ( .A(n6299), .ZN(n6268) );
  AND2_X1 U7279 ( .A1(n6269), .A2(n6268), .ZN(n6273) );
  NOR2_X1 U7280 ( .A1(n6273), .A2(n6617), .ZN(n6270) );
  AOI21_X1 U7281 ( .B1(n6276), .B2(STATE2_REG_2__SCAN_IN), .A(n6270), .ZN(
        n6307) );
  AOI22_X1 U7282 ( .A1(n6394), .A2(n6301), .B1(n6440), .B2(n6299), .ZN(n6278)
         );
  NAND3_X1 U7283 ( .A1(n6396), .A2(n6272), .A3(n6271), .ZN(n6274) );
  NAND3_X1 U7284 ( .A1(n6274), .A2(n6442), .A3(n6273), .ZN(n6275) );
  OAI211_X1 U7285 ( .C1(n6442), .C2(n6276), .A(n6315), .B(n6275), .ZN(n6303)
         );
  AOI22_X1 U7286 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6303), .B1(n6451), 
        .B2(n6302), .ZN(n6277) );
  OAI211_X1 U7287 ( .C1(n6307), .C2(n6279), .A(n6278), .B(n6277), .ZN(U3044)
         );
  AOI22_X1 U7288 ( .A1(n6301), .A2(n6378), .B1(n6456), .B2(n6299), .ZN(n6281)
         );
  AOI22_X1 U7289 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6303), .B1(n5043), 
        .B2(n6302), .ZN(n6280) );
  OAI211_X1 U7290 ( .C1(n6307), .C2(n6282), .A(n6281), .B(n6280), .ZN(U3045)
         );
  AOI22_X1 U7291 ( .A1(n6301), .A2(n6382), .B1(n6460), .B2(n6299), .ZN(n6284)
         );
  AOI22_X1 U7292 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6303), .B1(n6462), 
        .B2(n6302), .ZN(n6283) );
  OAI211_X1 U7293 ( .C1(n6307), .C2(n6285), .A(n6284), .B(n6283), .ZN(U3046)
         );
  AOI22_X1 U7294 ( .A1(n6301), .A2(n6414), .B1(n6467), .B2(n6299), .ZN(n6287)
         );
  AOI22_X1 U7295 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6303), .B1(n6468), 
        .B2(n6302), .ZN(n6286) );
  OAI211_X1 U7296 ( .C1(n6307), .C2(n6288), .A(n6287), .B(n6286), .ZN(U3047)
         );
  AOI22_X1 U7297 ( .A1(n6301), .A2(n6289), .B1(n6473), .B2(n6299), .ZN(n6291)
         );
  AOI22_X1 U7298 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6303), .B1(n5001), 
        .B2(n6302), .ZN(n6290) );
  OAI211_X1 U7299 ( .C1(n6307), .C2(n6292), .A(n6291), .B(n6290), .ZN(U3048)
         );
  AOI22_X1 U7300 ( .A1(n6301), .A2(n6420), .B1(n6478), .B2(n6299), .ZN(n6294)
         );
  AOI22_X1 U7301 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6303), .B1(n6479), 
        .B2(n6302), .ZN(n6293) );
  OAI211_X1 U7302 ( .C1(n6307), .C2(n6295), .A(n6294), .B(n6293), .ZN(U3049)
         );
  AOI22_X1 U7303 ( .A1(n6301), .A2(n6333), .B1(n6484), .B2(n6299), .ZN(n6297)
         );
  AOI22_X1 U7304 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6303), .B1(n6485), 
        .B2(n6302), .ZN(n6296) );
  OAI211_X1 U7305 ( .C1(n6307), .C2(n6298), .A(n6297), .B(n6296), .ZN(U3050)
         );
  AOI22_X1 U7306 ( .A1(n6301), .A2(n6300), .B1(n7027), .B2(n6299), .ZN(n6305)
         );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6303), .B1(n7020), 
        .B2(n6302), .ZN(n6304) );
  OAI211_X1 U7308 ( .C1(n6307), .C2(n6306), .A(n6305), .B(n6304), .ZN(U3051)
         );
  AOI22_X1 U7309 ( .A1(n6338), .A2(n6440), .B1(n6394), .B2(n7021), .ZN(n6322)
         );
  NOR2_X1 U7310 ( .A1(n6311), .A2(n6617), .ZN(n6317) );
  AOI21_X1 U7311 ( .B1(n6313), .B2(n6312), .A(n6338), .ZN(n6319) );
  NAND2_X1 U7312 ( .A1(n6317), .A2(n6319), .ZN(n6314) );
  OAI211_X1 U7313 ( .C1(n6442), .C2(n6316), .A(n6315), .B(n6314), .ZN(n6340)
         );
  INV_X1 U7314 ( .A(n6317), .ZN(n6320) );
  OAI22_X1 U7315 ( .A1(n6320), .A2(n6319), .B1(n6318), .B2(n6403), .ZN(n6339)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6340), .B1(n6439), 
        .B2(n6339), .ZN(n6321) );
  OAI211_X1 U7317 ( .C1(n6409), .C2(n6375), .A(n6322), .B(n6321), .ZN(U3076)
         );
  INV_X1 U7318 ( .A(n6375), .ZN(n6337) );
  AOI22_X1 U7319 ( .A1(n6456), .A2(n6338), .B1(n5043), .B2(n6337), .ZN(n6324)
         );
  AOI22_X1 U7320 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6340), .B1(n6455), 
        .B2(n6339), .ZN(n6323) );
  OAI211_X1 U7321 ( .C1(n6459), .C2(n6343), .A(n6324), .B(n6323), .ZN(U3077)
         );
  AOI22_X1 U7322 ( .A1(n6338), .A2(n6460), .B1(n6462), .B2(n6337), .ZN(n6326)
         );
  AOI22_X1 U7323 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6340), .B1(n6461), 
        .B2(n6339), .ZN(n6325) );
  OAI211_X1 U7324 ( .C1(n6465), .C2(n6343), .A(n6326), .B(n6325), .ZN(U3078)
         );
  AOI22_X1 U7325 ( .A1(n6467), .A2(n6338), .B1(n6468), .B2(n6337), .ZN(n6328)
         );
  AOI22_X1 U7326 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6340), .B1(n6466), 
        .B2(n6339), .ZN(n6327) );
  OAI211_X1 U7327 ( .C1(n6471), .C2(n6343), .A(n6328), .B(n6327), .ZN(U3079)
         );
  AOI22_X1 U7328 ( .A1(n6473), .A2(n6338), .B1(n5001), .B2(n6337), .ZN(n6330)
         );
  AOI22_X1 U7329 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6340), .B1(n6472), 
        .B2(n6339), .ZN(n6329) );
  OAI211_X1 U7330 ( .C1(n6476), .C2(n6343), .A(n6330), .B(n6329), .ZN(U3080)
         );
  AOI22_X1 U7331 ( .A1(n6478), .A2(n6338), .B1(n6420), .B2(n7021), .ZN(n6332)
         );
  AOI22_X1 U7332 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6340), .B1(n6477), 
        .B2(n6339), .ZN(n6331) );
  OAI211_X1 U7333 ( .C1(n6424), .C2(n6375), .A(n6332), .B(n6331), .ZN(U3081)
         );
  AOI22_X1 U7334 ( .A1(n6484), .A2(n6338), .B1(n6333), .B2(n7021), .ZN(n6335)
         );
  AOI22_X1 U7335 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6340), .B1(n6483), 
        .B2(n6339), .ZN(n6334) );
  OAI211_X1 U7336 ( .C1(n6336), .C2(n6375), .A(n6335), .B(n6334), .ZN(U3082)
         );
  AOI22_X1 U7337 ( .A1(n6338), .A2(n7027), .B1(n7020), .B2(n6337), .ZN(n6342)
         );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6340), .B1(n7019), 
        .B2(n6339), .ZN(n6341) );
  OAI211_X1 U7339 ( .C1(n7023), .C2(n6343), .A(n6342), .B(n6341), .ZN(U3083)
         );
  NOR2_X1 U7340 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6344), .ZN(n6371)
         );
  NOR2_X1 U7341 ( .A1(n6437), .A2(n6345), .ZN(n6350) );
  INV_X1 U7342 ( .A(n6350), .ZN(n6348) );
  OR2_X1 U7343 ( .A1(n6347), .A2(n6346), .ZN(n6436) );
  OAI22_X1 U7344 ( .A1(n6348), .A2(n6617), .B1(n6448), .B2(n6436), .ZN(n6370)
         );
  AOI22_X1 U7345 ( .A1(n6440), .A2(n6371), .B1(n6439), .B2(n6370), .ZN(n6357)
         );
  NAND3_X1 U7346 ( .A1(n6349), .A2(n6442), .A3(n6375), .ZN(n6352) );
  AOI21_X1 U7347 ( .B1(n6352), .B2(n6351), .A(n6350), .ZN(n6355) );
  AOI21_X1 U7348 ( .B1(n6436), .B2(STATE2_REG_2__SCAN_IN), .A(n6353), .ZN(
        n6449) );
  OAI211_X1 U7349 ( .C1(n6605), .C2(n6371), .A(n6435), .B(n6449), .ZN(n6354)
         );
  AOI22_X1 U7350 ( .A1(n6372), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6451), 
        .B2(n6383), .ZN(n6356) );
  OAI211_X1 U7351 ( .C1(n6454), .C2(n6375), .A(n6357), .B(n6356), .ZN(U3084)
         );
  AOI22_X1 U7352 ( .A1(n6456), .A2(n6371), .B1(n6455), .B2(n6370), .ZN(n6359)
         );
  AOI22_X1 U7353 ( .A1(n6372), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5043), 
        .B2(n6383), .ZN(n6358) );
  OAI211_X1 U7354 ( .C1(n6459), .C2(n6375), .A(n6359), .B(n6358), .ZN(U3085)
         );
  AOI22_X1 U7355 ( .A1(n6461), .A2(n6370), .B1(n6460), .B2(n6371), .ZN(n6361)
         );
  AOI22_X1 U7356 ( .A1(n6372), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6462), 
        .B2(n6383), .ZN(n6360) );
  OAI211_X1 U7357 ( .C1(n6465), .C2(n6375), .A(n6361), .B(n6360), .ZN(U3086)
         );
  AOI22_X1 U7358 ( .A1(n6467), .A2(n6371), .B1(n6466), .B2(n6370), .ZN(n6363)
         );
  AOI22_X1 U7359 ( .A1(n6372), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6468), 
        .B2(n6383), .ZN(n6362) );
  OAI211_X1 U7360 ( .C1(n6471), .C2(n6375), .A(n6363), .B(n6362), .ZN(U3087)
         );
  AOI22_X1 U7361 ( .A1(n6473), .A2(n6371), .B1(n6472), .B2(n6370), .ZN(n6365)
         );
  AOI22_X1 U7362 ( .A1(n6372), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5001), 
        .B2(n6383), .ZN(n6364) );
  OAI211_X1 U7363 ( .C1(n6476), .C2(n6375), .A(n6365), .B(n6364), .ZN(U3088)
         );
  AOI22_X1 U7364 ( .A1(n6478), .A2(n6371), .B1(n6477), .B2(n6370), .ZN(n6367)
         );
  AOI22_X1 U7365 ( .A1(n6372), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6479), 
        .B2(n6383), .ZN(n6366) );
  OAI211_X1 U7366 ( .C1(n6482), .C2(n6375), .A(n6367), .B(n6366), .ZN(U3089)
         );
  AOI22_X1 U7367 ( .A1(n6484), .A2(n6371), .B1(n6483), .B2(n6370), .ZN(n6369)
         );
  AOI22_X1 U7368 ( .A1(n6372), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6485), 
        .B2(n6383), .ZN(n6368) );
  OAI211_X1 U7369 ( .C1(n6488), .C2(n6375), .A(n6369), .B(n6368), .ZN(U3090)
         );
  AOI22_X1 U7370 ( .A1(n7027), .A2(n6371), .B1(n7019), .B2(n6370), .ZN(n6374)
         );
  AOI22_X1 U7371 ( .A1(n6372), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n7020), 
        .B2(n6383), .ZN(n6373) );
  OAI211_X1 U7372 ( .C1(n7023), .C2(n6375), .A(n6374), .B(n6373), .ZN(U3091)
         );
  INV_X1 U7373 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6949) );
  AOI22_X1 U7374 ( .A1(n6383), .A2(n6394), .B1(n6440), .B2(n6381), .ZN(n6377)
         );
  AOI22_X1 U7375 ( .A1(n6385), .A2(n6439), .B1(n6384), .B2(n6451), .ZN(n6376)
         );
  OAI211_X1 U7376 ( .C1(n6389), .C2(n6949), .A(n6377), .B(n6376), .ZN(U3092)
         );
  INV_X1 U7377 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U7378 ( .A1(n6384), .A2(n5043), .B1(n6456), .B2(n6381), .ZN(n6380)
         );
  AOI22_X1 U7379 ( .A1(n6385), .A2(n6455), .B1(n6378), .B2(n6383), .ZN(n6379)
         );
  OAI211_X1 U7380 ( .C1(n6389), .C2(n6763), .A(n6380), .B(n6379), .ZN(U3093)
         );
  INV_X1 U7381 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6388) );
  AOI22_X1 U7382 ( .A1(n6383), .A2(n6382), .B1(n6460), .B2(n6381), .ZN(n6387)
         );
  AOI22_X1 U7383 ( .A1(n6385), .A2(n6461), .B1(n6384), .B2(n6462), .ZN(n6386)
         );
  OAI211_X1 U7384 ( .C1(n6389), .C2(n6388), .A(n6387), .B(n6386), .ZN(U3094)
         );
  INV_X1 U7385 ( .A(n6392), .ZN(n6393) );
  AND2_X1 U7386 ( .A1(n6393), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6427)
         );
  AOI22_X1 U7387 ( .A1(n6394), .A2(n6421), .B1(n6440), .B2(n6427), .ZN(n6408)
         );
  OAI21_X1 U7388 ( .B1(n6396), .B2(n6395), .A(n6442), .ZN(n6406) );
  OR2_X1 U7389 ( .A1(n6397), .A2(n3982), .ZN(n6399) );
  INV_X1 U7390 ( .A(n6427), .ZN(n6398) );
  NAND2_X1 U7391 ( .A1(n6399), .A2(n6398), .ZN(n6402) );
  AOI21_X1 U7392 ( .B1(n6404), .B2(n6617), .A(n6400), .ZN(n6401) );
  OAI21_X1 U7393 ( .B1(n6406), .B2(n6402), .A(n6401), .ZN(n6429) );
  INV_X1 U7394 ( .A(n6402), .ZN(n6405) );
  OAI22_X1 U7395 ( .A1(n6406), .A2(n6405), .B1(n6404), .B2(n6403), .ZN(n6428)
         );
  AOI22_X1 U7396 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6429), .B1(n6439), 
        .B2(n6428), .ZN(n6407) );
  OAI211_X1 U7397 ( .C1(n6409), .C2(n6495), .A(n6408), .B(n6407), .ZN(U3108)
         );
  AOI22_X1 U7398 ( .A1(n6441), .A2(n5043), .B1(n6456), .B2(n6427), .ZN(n6411)
         );
  AOI22_X1 U7399 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6429), .B1(n6455), 
        .B2(n6428), .ZN(n6410) );
  OAI211_X1 U7400 ( .C1(n6459), .C2(n6432), .A(n6411), .B(n6410), .ZN(U3109)
         );
  AOI22_X1 U7401 ( .A1(n6462), .A2(n6441), .B1(n6460), .B2(n6427), .ZN(n6413)
         );
  AOI22_X1 U7402 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6429), .B1(n6461), 
        .B2(n6428), .ZN(n6412) );
  OAI211_X1 U7403 ( .C1(n6465), .C2(n6432), .A(n6413), .B(n6412), .ZN(U3110)
         );
  AOI22_X1 U7404 ( .A1(n6421), .A2(n6414), .B1(n6467), .B2(n6427), .ZN(n6416)
         );
  AOI22_X1 U7405 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6429), .B1(n6466), 
        .B2(n6428), .ZN(n6415) );
  OAI211_X1 U7406 ( .C1(n6417), .C2(n6495), .A(n6416), .B(n6415), .ZN(U3111)
         );
  AOI22_X1 U7407 ( .A1(n6441), .A2(n5001), .B1(n6473), .B2(n6427), .ZN(n6419)
         );
  AOI22_X1 U7408 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6429), .B1(n6472), 
        .B2(n6428), .ZN(n6418) );
  OAI211_X1 U7409 ( .C1(n6476), .C2(n6432), .A(n6419), .B(n6418), .ZN(U3112)
         );
  AOI22_X1 U7410 ( .A1(n6421), .A2(n6420), .B1(n6478), .B2(n6427), .ZN(n6423)
         );
  AOI22_X1 U7411 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6429), .B1(n6477), 
        .B2(n6428), .ZN(n6422) );
  OAI211_X1 U7412 ( .C1(n6424), .C2(n6495), .A(n6423), .B(n6422), .ZN(U3113)
         );
  AOI22_X1 U7413 ( .A1(n6441), .A2(n6485), .B1(n6484), .B2(n6427), .ZN(n6426)
         );
  AOI22_X1 U7414 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6429), .B1(n6483), 
        .B2(n6428), .ZN(n6425) );
  OAI211_X1 U7415 ( .C1(n6488), .C2(n6432), .A(n6426), .B(n6425), .ZN(U3114)
         );
  AOI22_X1 U7416 ( .A1(n7020), .A2(n6441), .B1(n7027), .B2(n6427), .ZN(n6431)
         );
  AOI22_X1 U7417 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6429), .B1(n7019), 
        .B2(n6428), .ZN(n6430) );
  OAI211_X1 U7418 ( .C1(n7023), .C2(n6432), .A(n6431), .B(n6430), .ZN(U3115)
         );
  NAND2_X1 U7419 ( .A1(n6902), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6433) );
  OR2_X1 U7420 ( .A1(n6434), .A2(n6433), .ZN(n6446) );
  INV_X1 U7421 ( .A(n6446), .ZN(n6490) );
  OAI22_X1 U7422 ( .A1(n6438), .A2(n6437), .B1(n6436), .B2(n6435), .ZN(n6489)
         );
  AOI22_X1 U7423 ( .A1(n6440), .A2(n6490), .B1(n6439), .B2(n6489), .ZN(n6453)
         );
  OAI21_X1 U7424 ( .B1(n6441), .B2(n6491), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6443) );
  OAI211_X1 U7425 ( .C1(n6445), .C2(n6444), .A(n6443), .B(n6442), .ZN(n6450)
         );
  NAND2_X1 U7426 ( .A1(n6446), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6447) );
  NAND4_X1 U7427 ( .A1(n6450), .A2(n6449), .A3(n6448), .A4(n6447), .ZN(n6492)
         );
  AOI22_X1 U7428 ( .A1(n6492), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6451), 
        .B2(n6491), .ZN(n6452) );
  OAI211_X1 U7429 ( .C1(n6454), .C2(n6495), .A(n6453), .B(n6452), .ZN(U3116)
         );
  AOI22_X1 U7430 ( .A1(n6456), .A2(n6490), .B1(n6455), .B2(n6489), .ZN(n6458)
         );
  AOI22_X1 U7431 ( .A1(n6492), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5043), 
        .B2(n6491), .ZN(n6457) );
  OAI211_X1 U7432 ( .C1(n6459), .C2(n6495), .A(n6458), .B(n6457), .ZN(U3117)
         );
  AOI22_X1 U7433 ( .A1(n6461), .A2(n6489), .B1(n6460), .B2(n6490), .ZN(n6464)
         );
  AOI22_X1 U7434 ( .A1(n6492), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6462), 
        .B2(n6491), .ZN(n6463) );
  OAI211_X1 U7435 ( .C1(n6465), .C2(n6495), .A(n6464), .B(n6463), .ZN(U3118)
         );
  AOI22_X1 U7436 ( .A1(n6467), .A2(n6490), .B1(n6466), .B2(n6489), .ZN(n6470)
         );
  AOI22_X1 U7437 ( .A1(n6492), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6468), 
        .B2(n6491), .ZN(n6469) );
  OAI211_X1 U7438 ( .C1(n6471), .C2(n6495), .A(n6470), .B(n6469), .ZN(U3119)
         );
  AOI22_X1 U7439 ( .A1(n6473), .A2(n6490), .B1(n6472), .B2(n6489), .ZN(n6475)
         );
  AOI22_X1 U7440 ( .A1(n6492), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5001), 
        .B2(n6491), .ZN(n6474) );
  OAI211_X1 U7441 ( .C1(n6476), .C2(n6495), .A(n6475), .B(n6474), .ZN(U3120)
         );
  AOI22_X1 U7442 ( .A1(n6478), .A2(n6490), .B1(n6477), .B2(n6489), .ZN(n6481)
         );
  AOI22_X1 U7443 ( .A1(n6492), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6479), 
        .B2(n6491), .ZN(n6480) );
  OAI211_X1 U7444 ( .C1(n6482), .C2(n6495), .A(n6481), .B(n6480), .ZN(U3121)
         );
  AOI22_X1 U7445 ( .A1(n6484), .A2(n6490), .B1(n6483), .B2(n6489), .ZN(n6487)
         );
  AOI22_X1 U7446 ( .A1(n6492), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6485), 
        .B2(n6491), .ZN(n6486) );
  OAI211_X1 U7447 ( .C1(n6488), .C2(n6495), .A(n6487), .B(n6486), .ZN(U3122)
         );
  AOI22_X1 U7448 ( .A1(n7027), .A2(n6490), .B1(n7019), .B2(n6489), .ZN(n6494)
         );
  AOI22_X1 U7449 ( .A1(n6492), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n7020), 
        .B2(n6491), .ZN(n6493) );
  OAI211_X1 U7450 ( .C1(n7023), .C2(n6495), .A(n6494), .B(n6493), .ZN(U3123)
         );
  AND3_X1 U7451 ( .A1(n6497), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6496), 
        .ZN(n6503) );
  INV_X1 U7452 ( .A(n6503), .ZN(n6501) );
  OAI211_X1 U7453 ( .C1(n6501), .C2(n6500), .A(n6499), .B(n6498), .ZN(n6502)
         );
  OAI21_X1 U7454 ( .B1(n6503), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6502), 
        .ZN(n6504) );
  AOI222_X1 U7455 ( .A1(n6506), .A2(n6505), .B1(n6506), .B2(n6504), .C1(n6505), 
        .C2(n6504), .ZN(n6508) );
  OAI21_X1 U7456 ( .B1(n6508), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6507), 
        .ZN(n6516) );
  AOI21_X1 U7457 ( .B1(n6508), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6515) );
  OAI21_X1 U7458 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6509), 
        .ZN(n6510) );
  NAND3_X1 U7459 ( .A1(n6512), .A2(n6511), .A3(n6510), .ZN(n6513) );
  AOI211_X1 U7460 ( .C1(n6516), .C2(n6515), .A(n6514), .B(n6513), .ZN(n6527)
         );
  INV_X1 U7461 ( .A(n6527), .ZN(n6517) );
  OAI22_X1 U7462 ( .A1(n6517), .A2(n6529), .B1(n3821), .B2(n6619), .ZN(n6518)
         );
  OAI21_X1 U7463 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(n6606) );
  OAI21_X1 U7464 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3821), .A(n6606), .ZN(
        n6528) );
  AOI221_X1 U7465 ( .B1(n6522), .B2(STATE2_REG_0__SCAN_IN), .C1(n6528), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6521), .ZN(n6526) );
  OAI211_X1 U7466 ( .C1(n6535), .C2(n6524), .A(n6523), .B(n6606), .ZN(n6525)
         );
  OAI211_X1 U7467 ( .C1(n6527), .C2(n6529), .A(n6526), .B(n6525), .ZN(U3148)
         );
  OAI211_X1 U7468 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6528), .ZN(n6534) );
  OAI21_X1 U7469 ( .B1(READY_N), .B2(n6530), .A(n6529), .ZN(n6532) );
  AOI21_X1 U7470 ( .B1(n6532), .B2(n6606), .A(n6531), .ZN(n6533) );
  NAND2_X1 U7471 ( .A1(n6534), .A2(n6533), .ZN(U3149) );
  INV_X1 U7472 ( .A(n6535), .ZN(n6624) );
  OAI221_X1 U7473 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n3821), .A(n6603), .ZN(n6537) );
  OAI21_X1 U7474 ( .B1(n6624), .B2(n6537), .A(n6536), .ZN(U3150) );
  AND2_X1 U7475 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6600), .ZN(U3151) );
  NOR2_X1 U7476 ( .A1(n6602), .A2(n6794), .ZN(U3152) );
  AND2_X1 U7477 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6600), .ZN(U3153) );
  NOR2_X1 U7478 ( .A1(n6602), .A2(n6817), .ZN(U3154) );
  AND2_X1 U7479 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6600), .ZN(U3155) );
  AND2_X1 U7480 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6600), .ZN(U3156) );
  NOR2_X1 U7481 ( .A1(n6602), .A2(n6823), .ZN(U3157) );
  AND2_X1 U7482 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6600), .ZN(U3158) );
  NOR2_X1 U7483 ( .A1(n6602), .A2(n6871), .ZN(U3159) );
  AND2_X1 U7484 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6600), .ZN(U3160) );
  AND2_X1 U7485 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6600), .ZN(U3161) );
  AND2_X1 U7486 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6600), .ZN(U3162) );
  AND2_X1 U7487 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6600), .ZN(U3163) );
  AND2_X1 U7488 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6600), .ZN(U3164) );
  AND2_X1 U7489 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6600), .ZN(U3165) );
  AND2_X1 U7490 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6600), .ZN(U3166) );
  AND2_X1 U7491 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6600), .ZN(U3167) );
  AND2_X1 U7492 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6600), .ZN(U3168) );
  AND2_X1 U7493 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6600), .ZN(U3169) );
  NOR2_X1 U7494 ( .A1(n6602), .A2(n6807), .ZN(U3170) );
  NOR2_X1 U7495 ( .A1(n6602), .A2(n6895), .ZN(U3171) );
  AND2_X1 U7496 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6600), .ZN(U3172) );
  AND2_X1 U7497 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6600), .ZN(U3173) );
  AND2_X1 U7498 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6600), .ZN(U3174) );
  AND2_X1 U7499 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6600), .ZN(U3175) );
  INV_X1 U7500 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6912) );
  NOR2_X1 U7501 ( .A1(n6602), .A2(n6912), .ZN(U3176) );
  AND2_X1 U7502 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6600), .ZN(U3177) );
  AND2_X1 U7503 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6600), .ZN(U3178) );
  AND2_X1 U7504 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6600), .ZN(U3179) );
  AND2_X1 U7505 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6600), .ZN(U3180) );
  AOI22_X1 U7506 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6551) );
  AND2_X1 U7507 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6541) );
  INV_X1 U7508 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6539) );
  INV_X1 U7509 ( .A(NA_N), .ZN(n6548) );
  AOI211_X1 U7510 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6548), .A(
        STATE_REG_0__SCAN_IN), .B(n6547), .ZN(n6553) );
  AOI221_X1 U7511 ( .B1(n6541), .B2(n6629), .C1(n6539), .C2(n6629), .A(n6553), 
        .ZN(n6538) );
  OAI21_X1 U7512 ( .B1(n6547), .B2(n6551), .A(n6538), .ZN(U3181) );
  NOR2_X1 U7513 ( .A1(n6545), .A2(n6539), .ZN(n6549) );
  NAND2_X1 U7514 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6540) );
  OAI21_X1 U7515 ( .B1(n6549), .B2(n6541), .A(n6540), .ZN(n6542) );
  OAI211_X1 U7516 ( .C1(n6544), .C2(n3821), .A(n6543), .B(n6542), .ZN(U3182)
         );
  AOI221_X1 U7517 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n3821), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6546) );
  AOI221_X1 U7518 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6546), .C2(HOLD), .A(n6545), .ZN(n6552) );
  AOI21_X1 U7519 ( .B1(n6549), .B2(n6548), .A(n6547), .ZN(n6550) );
  OAI22_X1 U7520 ( .A1(n6553), .A2(n6552), .B1(n6551), .B2(n6550), .ZN(U3183)
         );
  NAND2_X1 U7521 ( .A1(n6631), .A2(n6554), .ZN(n6593) );
  INV_X1 U7522 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U7523 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6631), .ZN(n6596) );
  INV_X1 U7524 ( .A(n6596), .ZN(n6591) );
  OAI222_X1 U7525 ( .A1(n6593), .A2(n6555), .B1(n6796), .B2(n6631), .C1(n6607), 
        .C2(n6587), .ZN(U3184) );
  INV_X1 U7526 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6960) );
  OAI222_X1 U7527 ( .A1(n6596), .A2(n6555), .B1(n6960), .B2(n6631), .C1(n6556), 
        .C2(n6593), .ZN(U3185) );
  INV_X1 U7528 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6930) );
  OAI222_X1 U7529 ( .A1(n6596), .A2(n6556), .B1(n6930), .B2(n6631), .C1(n6855), 
        .C2(n6593), .ZN(U3186) );
  INV_X1 U7530 ( .A(n6593), .ZN(n6594) );
  AOI22_X1 U7531 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6629), .ZN(n6557) );
  OAI21_X1 U7532 ( .B1(n6855), .B2(n6596), .A(n6557), .ZN(U3187) );
  AOI22_X1 U7533 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6629), .ZN(n6558) );
  OAI21_X1 U7534 ( .B1(n6559), .B2(n6596), .A(n6558), .ZN(U3188) );
  AOI22_X1 U7535 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6629), .ZN(n6560) );
  OAI21_X1 U7536 ( .B1(n4748), .B2(n6596), .A(n6560), .ZN(U3189) );
  INV_X1 U7537 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6915) );
  OAI222_X1 U7538 ( .A1(n6596), .A2(n6561), .B1(n6915), .B2(n6631), .C1(n6563), 
        .C2(n6593), .ZN(U3190) );
  AOI22_X1 U7539 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6629), .ZN(n6562) );
  OAI21_X1 U7540 ( .B1(n6563), .B2(n6596), .A(n6562), .ZN(U3191) );
  AOI22_X1 U7541 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6629), .ZN(n6564) );
  OAI21_X1 U7542 ( .B1(n6783), .B2(n6587), .A(n6564), .ZN(U3192) );
  AOI22_X1 U7543 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6629), .ZN(n6565) );
  OAI21_X1 U7544 ( .B1(n6768), .B2(n6587), .A(n6565), .ZN(U3193) );
  INV_X1 U7545 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6943) );
  AOI22_X1 U7546 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6629), .ZN(n6566) );
  OAI21_X1 U7547 ( .B1(n6943), .B2(n6587), .A(n6566), .ZN(U3194) );
  AOI22_X1 U7548 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6629), .ZN(n6567) );
  OAI21_X1 U7549 ( .B1(n6568), .B2(n6587), .A(n6567), .ZN(U3195) );
  INV_X1 U7550 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6887) );
  OAI222_X1 U7551 ( .A1(n6587), .A2(n6951), .B1(n6887), .B2(n6631), .C1(n6570), 
        .C2(n6593), .ZN(U3196) );
  AOI22_X1 U7552 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6629), .ZN(n6569) );
  OAI21_X1 U7553 ( .B1(n6570), .B2(n6587), .A(n6569), .ZN(U3197) );
  AOI22_X1 U7554 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6629), .ZN(n6571) );
  OAI21_X1 U7555 ( .B1(n6778), .B2(n6587), .A(n6571), .ZN(U3198) );
  INV_X1 U7556 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6945) );
  OAI222_X1 U7557 ( .A1(n6587), .A2(n6572), .B1(n6945), .B2(n6631), .C1(n6574), 
        .C2(n6593), .ZN(U3199) );
  AOI22_X1 U7558 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6629), .ZN(n6573) );
  OAI21_X1 U7559 ( .B1(n6574), .B2(n6587), .A(n6573), .ZN(U3200) );
  AOI22_X1 U7560 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6629), .ZN(n6575) );
  OAI21_X1 U7561 ( .B1(n6576), .B2(n6587), .A(n6575), .ZN(U3201) );
  AOI22_X1 U7562 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6591), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6629), .ZN(n6577) );
  OAI21_X1 U7563 ( .B1(n6579), .B2(n6593), .A(n6577), .ZN(U3202) );
  AOI22_X1 U7564 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6629), .ZN(n6578) );
  OAI21_X1 U7565 ( .B1(n6579), .B2(n6587), .A(n6578), .ZN(U3203) );
  AOI22_X1 U7566 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6629), .ZN(n6580) );
  OAI21_X1 U7567 ( .B1(n6581), .B2(n6587), .A(n6580), .ZN(U3204) );
  AOI22_X1 U7568 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6591), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6629), .ZN(n6582) );
  OAI21_X1 U7569 ( .B1(n6583), .B2(n6593), .A(n6582), .ZN(U3205) );
  INV_X1 U7570 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6834) );
  OAI222_X1 U7571 ( .A1(n6587), .A2(n6583), .B1(n6834), .B2(n6631), .C1(n6585), 
        .C2(n6593), .ZN(U3206) );
  AOI22_X1 U7572 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6629), .ZN(n6584) );
  OAI21_X1 U7573 ( .B1(n6585), .B2(n6587), .A(n6584), .ZN(U3207) );
  AOI22_X1 U7574 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6629), .ZN(n6586) );
  OAI21_X1 U7575 ( .B1(n6755), .B2(n6596), .A(n6586), .ZN(U3208) );
  INV_X1 U7576 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6857) );
  OAI222_X1 U7577 ( .A1(n6587), .A2(n5487), .B1(n6857), .B2(n6631), .C1(n5419), 
        .C2(n6593), .ZN(U3209) );
  AOI22_X1 U7578 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6629), .ZN(n6588) );
  OAI21_X1 U7579 ( .B1(n5419), .B2(n6596), .A(n6588), .ZN(U3210) );
  AOI22_X1 U7580 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6629), .ZN(n6589) );
  OAI21_X1 U7581 ( .B1(n6590), .B2(n6596), .A(n6589), .ZN(U3211) );
  AOI22_X1 U7582 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6591), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6629), .ZN(n6592) );
  OAI21_X1 U7583 ( .B1(n6597), .B2(n6593), .A(n6592), .ZN(U3212) );
  AOI22_X1 U7584 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6594), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6629), .ZN(n6595) );
  OAI21_X1 U7585 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(U3213) );
  INV_X1 U7586 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6598) );
  INV_X1 U7587 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6964) );
  AOI22_X1 U7588 ( .A1(n6631), .A2(n6598), .B1(n6964), .B2(n6629), .ZN(U3445)
         );
  MUX2_X1 U7589 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6631), .Z(U3446) );
  MUX2_X1 U7590 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6631), .Z(U3447) );
  INV_X1 U7591 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6611) );
  INV_X1 U7592 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6899) );
  AOI22_X1 U7593 ( .A1(n6631), .A2(n6611), .B1(n6899), .B2(n6629), .ZN(U3448)
         );
  INV_X1 U7594 ( .A(n6601), .ZN(n6599) );
  AOI21_X1 U7595 ( .B1(n6852), .B2(n6600), .A(n6599), .ZN(U3451) );
  OAI21_X1 U7596 ( .B1(n6602), .B2(n6797), .A(n6601), .ZN(U3452) );
  OAI211_X1 U7597 ( .C1(n6606), .C2(n6605), .A(n6604), .B(n6603), .ZN(U3453)
         );
  OAI211_X1 U7598 ( .C1(n6852), .C2(n6613), .A(n6797), .B(n6614), .ZN(n6610)
         );
  NOR2_X1 U7599 ( .A1(n6612), .A2(n6607), .ZN(n6608) );
  AOI22_X1 U7600 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(n6612), .B1(
        REIP_REG_0__SCAN_IN), .B2(n6608), .ZN(n6609) );
  NAND2_X1 U7601 ( .A1(n6610), .A2(n6609), .ZN(U3468) );
  AOI22_X1 U7602 ( .A1(n6614), .A2(n6613), .B1(n6612), .B2(n6611), .ZN(U3469)
         );
  NAND2_X1 U7603 ( .A1(n6629), .A2(W_R_N_REG_SCAN_IN), .ZN(n6615) );
  OAI21_X1 U7604 ( .B1(n6629), .B2(READREQUEST_REG_SCAN_IN), .A(n6615), .ZN(
        U3470) );
  INV_X1 U7605 ( .A(n6616), .ZN(n6621) );
  OAI211_X1 U7606 ( .C1(READY_N), .C2(n6619), .A(n6618), .B(n6617), .ZN(n6620)
         );
  NOR2_X1 U7607 ( .A1(n6621), .A2(n6620), .ZN(n6628) );
  OAI211_X1 U7608 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6623), .A(n6622), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6625) );
  AOI21_X1 U7609 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6625), .A(n6624), .ZN(
        n6627) );
  NAND2_X1 U7610 ( .A1(n6628), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6626) );
  OAI21_X1 U7611 ( .B1(n6628), .B2(n6627), .A(n6626), .ZN(U3472) );
  INV_X1 U7612 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6630) );
  INV_X1 U7613 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6918) );
  AOI22_X1 U7614 ( .A1(n6631), .A2(n6630), .B1(n6918), .B2(n6629), .ZN(U3473)
         );
  OAI22_X1 U7615 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(keyinput51), .B1(
        keyinput75), .B2(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6632) );
  AOI221_X1 U7616 ( .B1(INSTQUEUE_REG_5__3__SCAN_IN), .B2(keyinput51), .C1(
        DATAWIDTH_REG_12__SCAN_IN), .C2(keyinput75), .A(n6632), .ZN(n6639) );
  OAI22_X1 U7617 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput48), .B1(
        DATAI_5_), .B2(keyinput50), .ZN(n6633) );
  AOI221_X1 U7618 ( .B1(PHYADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput48), .C1(
        keyinput50), .C2(DATAI_5_), .A(n6633), .ZN(n6638) );
  OAI22_X1 U7619 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput106), .B1(
        LWORD_REG_6__SCAN_IN), .B2(keyinput62), .ZN(n6634) );
  AOI221_X1 U7620 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput106), 
        .C1(keyinput62), .C2(LWORD_REG_6__SCAN_IN), .A(n6634), .ZN(n6637) );
  OAI22_X1 U7621 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(keyinput19), .B1(
        INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput90), .ZN(n6635) );
  AOI221_X1 U7622 ( .B1(INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput19), .C1(
        keyinput90), .C2(INSTQUEUE_REG_5__2__SCAN_IN), .A(n6635), .ZN(n6636)
         );
  NAND4_X1 U7623 ( .A1(n6639), .A2(n6638), .A3(n6637), .A4(n6636), .ZN(n6667)
         );
  OAI22_X1 U7624 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(keyinput43), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput79), .ZN(n6640) );
  AOI221_X1 U7625 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput43), 
        .C1(keyinput79), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n6640), .ZN(
        n6647) );
  OAI22_X1 U7626 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(keyinput13), .B1(
        keyinput117), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6641) );
  AOI221_X1 U7627 ( .B1(INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput13), .C1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput117), .A(n6641), .ZN(
        n6646) );
  OAI22_X1 U7628 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput82), .B1(
        EAX_REG_13__SCAN_IN), .B2(keyinput108), .ZN(n6642) );
  AOI221_X1 U7629 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput82), .C1(
        keyinput108), .C2(EAX_REG_13__SCAN_IN), .A(n6642), .ZN(n6645) );
  OAI22_X1 U7630 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(keyinput103), .B1(
        EBX_REG_20__SCAN_IN), .B2(keyinput15), .ZN(n6643) );
  AOI221_X1 U7631 ( .B1(INSTQUEUE_REG_5__6__SCAN_IN), .B2(keyinput103), .C1(
        keyinput15), .C2(EBX_REG_20__SCAN_IN), .A(n6643), .ZN(n6644) );
  NAND4_X1 U7632 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6666)
         );
  OAI22_X1 U7633 ( .A1(EBX_REG_2__SCAN_IN), .A2(keyinput112), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(keyinput10), .ZN(n6648) );
  AOI221_X1 U7634 ( .B1(EBX_REG_2__SCAN_IN), .B2(keyinput112), .C1(keyinput10), 
        .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6648), .ZN(n6655) );
  OAI22_X1 U7635 ( .A1(NA_N), .A2(keyinput12), .B1(keyinput107), .B2(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6649) );
  AOI221_X1 U7636 ( .B1(NA_N), .B2(keyinput12), .C1(DATAWIDTH_REG_1__SCAN_IN), 
        .C2(keyinput107), .A(n6649), .ZN(n6654) );
  OAI22_X1 U7637 ( .A1(n6793), .A2(keyinput47), .B1(keyinput61), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6650) );
  AOI221_X1 U7638 ( .B1(n6793), .B2(keyinput47), .C1(EAX_REG_25__SCAN_IN), 
        .C2(keyinput61), .A(n6650), .ZN(n6653) );
  OAI22_X1 U7639 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(keyinput21), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput64), .ZN(n6651) );
  AOI221_X1 U7640 ( .B1(INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput21), .C1(
        keyinput64), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n6651), .ZN(n6652) );
  NAND4_X1 U7641 ( .A1(n6655), .A2(n6654), .A3(n6653), .A4(n6652), .ZN(n6665)
         );
  OAI22_X1 U7642 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(keyinput26), .B1(
        keyinput57), .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6656) );
  AOI221_X1 U7643 ( .B1(INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput26), .C1(
        INSTQUEUE_REG_6__6__SCAN_IN), .C2(keyinput57), .A(n6656), .ZN(n6663)
         );
  OAI22_X1 U7644 ( .A1(DATAI_20_), .A2(keyinput60), .B1(keyinput44), .B2(
        BYTEENABLE_REG_2__SCAN_IN), .ZN(n6657) );
  AOI221_X1 U7645 ( .B1(DATAI_20_), .B2(keyinput60), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput44), .A(n6657), .ZN(n6662) );
  OAI22_X1 U7646 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(keyinput27), .B1(
        keyinput70), .B2(ADDRESS_REG_22__SCAN_IN), .ZN(n6658) );
  AOI221_X1 U7647 ( .B1(PHYADDRPOINTER_REG_16__SCAN_IN), .B2(keyinput27), .C1(
        ADDRESS_REG_22__SCAN_IN), .C2(keyinput70), .A(n6658), .ZN(n6661) );
  OAI22_X1 U7648 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput91), .B1(
        DATAO_REG_4__SCAN_IN), .B2(keyinput5), .ZN(n6659) );
  AOI221_X1 U7649 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput91), .C1(keyinput5), 
        .C2(DATAO_REG_4__SCAN_IN), .A(n6659), .ZN(n6660) );
  NAND4_X1 U7650 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n6664)
         );
  NOR4_X1 U7651 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n7017)
         );
  AOI22_X1 U7652 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(keyinput167), 
        .B1(INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput180), .ZN(n6668) );
  OAI221_X1 U7653 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput167), 
        .C1(INSTQUEUE_REG_9__4__SCAN_IN), .C2(keyinput180), .A(n6668), .ZN(
        n6675) );
  AOI22_X1 U7654 ( .A1(EAX_REG_14__SCAN_IN), .A2(keyinput224), .B1(
        INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput149), .ZN(n6669) );
  OAI221_X1 U7655 ( .B1(EAX_REG_14__SCAN_IN), .B2(keyinput224), .C1(
        INSTQUEUE_REG_4__7__SCAN_IN), .C2(keyinput149), .A(n6669), .ZN(n6674)
         );
  AOI22_X1 U7656 ( .A1(DATAI_5_), .A2(keyinput178), .B1(
        INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput218), .ZN(n6670) );
  OAI221_X1 U7657 ( .B1(DATAI_5_), .B2(keyinput178), .C1(
        INSTQUEUE_REG_5__2__SCAN_IN), .C2(keyinput218), .A(n6670), .ZN(n6673)
         );
  AOI22_X1 U7658 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(keyinput216), .B1(
        INSTQUEUE_REG_2__1__SCAN_IN), .B2(keyinput186), .ZN(n6671) );
  OAI221_X1 U7659 ( .B1(INSTQUEUE_REG_8__2__SCAN_IN), .B2(keyinput216), .C1(
        INSTQUEUE_REG_2__1__SCAN_IN), .C2(keyinput186), .A(n6671), .ZN(n6672)
         );
  NOR4_X1 U7660 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n6703)
         );
  AOI22_X1 U7661 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(keyinput195), .B1(
        INSTQUEUE_REG_11__1__SCAN_IN), .B2(keyinput221), .ZN(n6676) );
  OAI221_X1 U7662 ( .B1(INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput195), .C1(
        INSTQUEUE_REG_11__1__SCAN_IN), .C2(keyinput221), .A(n6676), .ZN(n6683)
         );
  AOI22_X1 U7663 ( .A1(EAX_REG_31__SCAN_IN), .A2(keyinput128), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput176), .ZN(n6677) );
  OAI221_X1 U7664 ( .B1(EAX_REG_31__SCAN_IN), .B2(keyinput128), .C1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .C2(keyinput176), .A(n6677), .ZN(n6682) );
  AOI22_X1 U7665 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(keyinput163), .B1(
        UWORD_REG_14__SCAN_IN), .B2(keyinput233), .ZN(n6678) );
  OAI221_X1 U7666 ( .B1(ADDRESS_REG_6__SCAN_IN), .B2(keyinput163), .C1(
        UWORD_REG_14__SCAN_IN), .C2(keyinput233), .A(n6678), .ZN(n6681) );
  AOI22_X1 U7667 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(keyinput250), .B1(
        INSTQUEUE_REG_1__3__SCAN_IN), .B2(keyinput151), .ZN(n6679) );
  OAI221_X1 U7668 ( .B1(INSTQUEUE_REG_11__3__SCAN_IN), .B2(keyinput250), .C1(
        INSTQUEUE_REG_1__3__SCAN_IN), .C2(keyinput151), .A(n6679), .ZN(n6680)
         );
  NOR4_X1 U7669 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6702)
         );
  AOI22_X1 U7670 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput172), .B1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput193), .ZN(n6684) );
  OAI221_X1 U7671 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput172), .C1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput193), .A(n6684), .ZN(
        n6691) );
  AOI22_X1 U7672 ( .A1(DATAO_REG_26__SCAN_IN), .A2(keyinput253), .B1(
        INSTQUEUE_REG_12__7__SCAN_IN), .B2(keyinput136), .ZN(n6685) );
  OAI221_X1 U7673 ( .B1(DATAO_REG_26__SCAN_IN), .B2(keyinput253), .C1(
        INSTQUEUE_REG_12__7__SCAN_IN), .C2(keyinput136), .A(n6685), .ZN(n6690)
         );
  AOI22_X1 U7674 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(keyinput217), .B1(
        INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput162), .ZN(n6686) );
  OAI221_X1 U7675 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(keyinput217), 
        .C1(INSTQUEUE_REG_9__0__SCAN_IN), .C2(keyinput162), .A(n6686), .ZN(
        n6689) );
  AOI22_X1 U7676 ( .A1(EBX_REG_20__SCAN_IN), .A2(keyinput143), .B1(
        INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput228), .ZN(n6687) );
  OAI221_X1 U7677 ( .B1(EBX_REG_20__SCAN_IN), .B2(keyinput143), .C1(
        INSTQUEUE_REG_9__7__SCAN_IN), .C2(keyinput228), .A(n6687), .ZN(n6688)
         );
  NOR4_X1 U7678 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6701)
         );
  AOI22_X1 U7679 ( .A1(EBX_REG_0__SCAN_IN), .A2(keyinput183), .B1(
        INSTQUEUE_REG_13__7__SCAN_IN), .B2(keyinput158), .ZN(n6692) );
  OAI221_X1 U7680 ( .B1(EBX_REG_0__SCAN_IN), .B2(keyinput183), .C1(
        INSTQUEUE_REG_13__7__SCAN_IN), .C2(keyinput158), .A(n6692), .ZN(n6699)
         );
  AOI22_X1 U7681 ( .A1(BE_N_REG_3__SCAN_IN), .A2(keyinput159), .B1(DATAI_22_), 
        .B2(keyinput213), .ZN(n6693) );
  OAI221_X1 U7682 ( .B1(BE_N_REG_3__SCAN_IN), .B2(keyinput159), .C1(DATAI_22_), 
        .C2(keyinput213), .A(n6693), .ZN(n6698) );
  AOI22_X1 U7683 ( .A1(NA_N), .A2(keyinput140), .B1(
        INSTQUEUE_REG_5__3__SCAN_IN), .B2(keyinput179), .ZN(n6694) );
  OAI221_X1 U7684 ( .B1(NA_N), .B2(keyinput140), .C1(
        INSTQUEUE_REG_5__3__SCAN_IN), .C2(keyinput179), .A(n6694), .ZN(n6697)
         );
  AOI22_X1 U7685 ( .A1(BE_N_REG_0__SCAN_IN), .A2(keyinput230), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput142), .ZN(n6695) );
  OAI221_X1 U7686 ( .B1(BE_N_REG_0__SCAN_IN), .B2(keyinput230), .C1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .C2(keyinput142), .A(n6695), .ZN(
        n6696) );
  NOR4_X1 U7687 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n6700)
         );
  NAND4_X1 U7688 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6849)
         );
  AOI22_X1 U7689 ( .A1(DATAI_20_), .A2(keyinput188), .B1(REIP_REG_21__SCAN_IN), 
        .B2(keyinput239), .ZN(n6704) );
  OAI221_X1 U7690 ( .B1(DATAI_20_), .B2(keyinput188), .C1(REIP_REG_21__SCAN_IN), .C2(keyinput239), .A(n6704), .ZN(n6711) );
  AOI22_X1 U7691 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput208), .B1(
        EAX_REG_11__SCAN_IN), .B2(keyinput204), .ZN(n6705) );
  OAI221_X1 U7692 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput208), .C1(
        EAX_REG_11__SCAN_IN), .C2(keyinput204), .A(n6705), .ZN(n6710) );
  AOI22_X1 U7693 ( .A1(EAX_REG_25__SCAN_IN), .A2(keyinput189), .B1(
        INSTQUEUE_REG_7__6__SCAN_IN), .B2(keyinput196), .ZN(n6706) );
  OAI221_X1 U7694 ( .B1(EAX_REG_25__SCAN_IN), .B2(keyinput189), .C1(
        INSTQUEUE_REG_7__6__SCAN_IN), .C2(keyinput196), .A(n6706), .ZN(n6709)
         );
  AOI22_X1 U7695 ( .A1(DATAI_12_), .A2(keyinput177), .B1(EBX_REG_2__SCAN_IN), 
        .B2(keyinput240), .ZN(n6707) );
  OAI221_X1 U7696 ( .B1(DATAI_12_), .B2(keyinput177), .C1(EBX_REG_2__SCAN_IN), 
        .C2(keyinput240), .A(n6707), .ZN(n6708) );
  NOR4_X1 U7697 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n6739)
         );
  AOI22_X1 U7698 ( .A1(DATAI_19_), .A2(keyinput173), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput145), .ZN(n6712) );
  OAI221_X1 U7699 ( .B1(DATAI_19_), .B2(keyinput173), .C1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput145), .A(n6712), .ZN(n6719) );
  AOI22_X1 U7700 ( .A1(LWORD_REG_4__SCAN_IN), .A2(keyinput206), .B1(
        INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput134), .ZN(n6713) );
  OAI221_X1 U7701 ( .B1(LWORD_REG_4__SCAN_IN), .B2(keyinput206), .C1(
        INSTQUEUE_REG_15__7__SCAN_IN), .C2(keyinput134), .A(n6713), .ZN(n6718)
         );
  AOI22_X1 U7702 ( .A1(ADDRESS_REG_2__SCAN_IN), .A2(keyinput181), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput150), .ZN(n6714) );
  OAI221_X1 U7703 ( .B1(ADDRESS_REG_2__SCAN_IN), .B2(keyinput181), .C1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .C2(keyinput150), .A(n6714), .ZN(
        n6717) );
  AOI22_X1 U7704 ( .A1(REIP_REG_13__SCAN_IN), .A2(keyinput139), .B1(DATAI_31_), 
        .B2(keyinput255), .ZN(n6715) );
  OAI221_X1 U7705 ( .B1(REIP_REG_13__SCAN_IN), .B2(keyinput139), .C1(DATAI_31_), .C2(keyinput255), .A(n6715), .ZN(n6716) );
  NOR4_X1 U7706 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6738)
         );
  AOI22_X1 U7707 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput210), .B1(
        INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput147), .ZN(n6720) );
  OAI221_X1 U7708 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput210), 
        .C1(INSTQUEUE_REG_12__6__SCAN_IN), .C2(keyinput147), .A(n6720), .ZN(
        n6727) );
  AOI22_X1 U7709 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(keyinput197), .B1(
        REIP_REG_4__SCAN_IN), .B2(keyinput160), .ZN(n6721) );
  OAI221_X1 U7710 ( .B1(DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput197), .C1(
        REIP_REG_4__SCAN_IN), .C2(keyinput160), .A(n6721), .ZN(n6726) );
  AOI22_X1 U7711 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(keyinput205), 
        .B1(INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput194), .ZN(n6722) );
  OAI221_X1 U7712 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput205), 
        .C1(INSTQUEUE_REG_10__5__SCAN_IN), .C2(keyinput194), .A(n6722), .ZN(
        n6725) );
  AOI22_X1 U7713 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput130), .B1(BS16_N), .B2(keyinput166), .ZN(n6723) );
  OAI221_X1 U7714 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput130), .C1(
        BS16_N), .C2(keyinput166), .A(n6723), .ZN(n6724) );
  NOR4_X1 U7715 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(n6737)
         );
  AOI22_X1 U7716 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(keyinput207), .B1(
        INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput226), .ZN(n6728) );
  OAI221_X1 U7717 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput207), 
        .C1(INSTQUEUE_REG_3__3__SCAN_IN), .C2(keyinput226), .A(n6728), .ZN(
        n6735) );
  AOI22_X1 U7718 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput129), .B1(
        EAX_REG_9__SCAN_IN), .B2(keyinput191), .ZN(n6729) );
  OAI221_X1 U7719 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput129), .C1(
        EAX_REG_9__SCAN_IN), .C2(keyinput191), .A(n6729), .ZN(n6734) );
  AOI22_X1 U7720 ( .A1(EAX_REG_15__SCAN_IN), .A2(keyinput187), .B1(
        INSTQUEUE_REG_10__1__SCAN_IN), .B2(keyinput238), .ZN(n6730) );
  OAI221_X1 U7721 ( .B1(EAX_REG_15__SCAN_IN), .B2(keyinput187), .C1(
        INSTQUEUE_REG_10__1__SCAN_IN), .C2(keyinput238), .A(n6730), .ZN(n6733)
         );
  AOI22_X1 U7722 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput225), .B1(
        EAX_REG_23__SCAN_IN), .B2(keyinput157), .ZN(n6731) );
  OAI221_X1 U7723 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput225), .C1(
        EAX_REG_23__SCAN_IN), .C2(keyinput157), .A(n6731), .ZN(n6732) );
  NOR4_X1 U7724 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6736)
         );
  NAND4_X1 U7725 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6848)
         );
  AOI22_X1 U7726 ( .A1(n6948), .A2(keyinput222), .B1(n6869), .B2(keyinput184), 
        .ZN(n6740) );
  OAI221_X1 U7727 ( .B1(n6948), .B2(keyinput222), .C1(n6869), .C2(keyinput184), 
        .A(n6740), .ZN(n6750) );
  INV_X1 U7728 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U7729 ( .A1(n6967), .A2(keyinput144), .B1(keyinput209), .B2(n6901), 
        .ZN(n6741) );
  OAI221_X1 U7730 ( .B1(n6967), .B2(keyinput144), .C1(n6901), .C2(keyinput209), 
        .A(n6741), .ZN(n6749) );
  INV_X1 U7731 ( .A(MORE_REG_SCAN_IN), .ZN(n6744) );
  AOI22_X1 U7732 ( .A1(n6744), .A2(keyinput219), .B1(n6743), .B2(keyinput141), 
        .ZN(n6742) );
  OAI221_X1 U7733 ( .B1(n6744), .B2(keyinput219), .C1(n6743), .C2(keyinput141), 
        .A(n6742), .ZN(n6748) );
  INV_X1 U7734 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6746) );
  AOI22_X1 U7735 ( .A1(n6946), .A2(keyinput227), .B1(keyinput190), .B2(n6746), 
        .ZN(n6745) );
  OAI221_X1 U7736 ( .B1(n6946), .B2(keyinput227), .C1(n6746), .C2(keyinput190), 
        .A(n6745), .ZN(n6747) );
  NOR4_X1 U7737 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6791)
         );
  AOI22_X1 U7738 ( .A1(n6752), .A2(keyinput252), .B1(keyinput246), .B2(n6857), 
        .ZN(n6751) );
  OAI221_X1 U7739 ( .B1(n6752), .B2(keyinput252), .C1(n6857), .C2(keyinput246), 
        .A(n6751), .ZN(n6761) );
  AOI22_X1 U7740 ( .A1(n6866), .A2(keyinput131), .B1(keyinput244), .B2(n4748), 
        .ZN(n6753) );
  OAI221_X1 U7741 ( .B1(n6866), .B2(keyinput131), .C1(n4748), .C2(keyinput244), 
        .A(n6753), .ZN(n6760) );
  AOI22_X1 U7742 ( .A1(n6936), .A2(keyinput182), .B1(n6755), .B2(keyinput132), 
        .ZN(n6754) );
  OAI221_X1 U7743 ( .B1(n6936), .B2(keyinput182), .C1(n6755), .C2(keyinput132), 
        .A(n6754), .ZN(n6759) );
  AOI22_X1 U7744 ( .A1(n6757), .A2(keyinput234), .B1(keyinput223), .B2(n6854), 
        .ZN(n6756) );
  OAI221_X1 U7745 ( .B1(n6757), .B2(keyinput234), .C1(n6854), .C2(keyinput223), 
        .A(n6756), .ZN(n6758) );
  NOR4_X1 U7746 ( .A1(n6761), .A2(n6760), .A3(n6759), .A4(n6758), .ZN(n6790)
         );
  AOI22_X1 U7747 ( .A1(n6763), .A2(keyinput154), .B1(keyinput170), .B2(n6898), 
        .ZN(n6762) );
  OAI221_X1 U7748 ( .B1(n6763), .B2(keyinput154), .C1(n6898), .C2(keyinput170), 
        .A(n6762), .ZN(n6775) );
  AOI22_X1 U7749 ( .A1(n6769), .A2(keyinput243), .B1(n6768), .B2(keyinput211), 
        .ZN(n6767) );
  OAI221_X1 U7750 ( .B1(n6769), .B2(keyinput243), .C1(n6768), .C2(keyinput211), 
        .A(n6767), .ZN(n6773) );
  AOI22_X1 U7751 ( .A1(n6771), .A2(keyinput138), .B1(n6902), .B2(keyinput148), 
        .ZN(n6770) );
  OAI221_X1 U7752 ( .B1(n6771), .B2(keyinput138), .C1(n6902), .C2(keyinput148), 
        .A(n6770), .ZN(n6772) );
  NOR4_X1 U7753 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6789)
         );
  AOI22_X1 U7754 ( .A1(n4939), .A2(keyinput248), .B1(keyinput215), .B2(n6887), 
        .ZN(n6776) );
  OAI221_X1 U7755 ( .B1(n4939), .B2(keyinput248), .C1(n6887), .C2(keyinput215), 
        .A(n6776), .ZN(n6787) );
  AOI22_X1 U7756 ( .A1(n6778), .A2(keyinput201), .B1(keyinput214), .B2(n6945), 
        .ZN(n6777) );
  OAI221_X1 U7757 ( .B1(n6778), .B2(keyinput201), .C1(n6945), .C2(keyinput214), 
        .A(n6777), .ZN(n6786) );
  AOI22_X1 U7758 ( .A1(n6783), .A2(keyinput249), .B1(n6782), .B2(keyinput245), 
        .ZN(n6781) );
  OAI221_X1 U7759 ( .B1(n6783), .B2(keyinput249), .C1(n6782), .C2(keyinput245), 
        .A(n6781), .ZN(n6784) );
  NOR4_X1 U7760 ( .A1(n6787), .A2(n6786), .A3(n6785), .A4(n6784), .ZN(n6788)
         );
  NAND4_X1 U7761 ( .A1(n6791), .A2(n6790), .A3(n6789), .A4(n6788), .ZN(n6847)
         );
  AOI22_X1 U7762 ( .A1(n6794), .A2(keyinput242), .B1(n6793), .B2(keyinput175), 
        .ZN(n6792) );
  OAI221_X1 U7763 ( .B1(n6794), .B2(keyinput242), .C1(n6793), .C2(keyinput175), 
        .A(n6792), .ZN(n6805) );
  AOI22_X1 U7764 ( .A1(n6797), .A2(keyinput235), .B1(keyinput237), .B2(n6796), 
        .ZN(n6795) );
  OAI221_X1 U7765 ( .B1(n6797), .B2(keyinput235), .C1(n6796), .C2(keyinput237), 
        .A(n6795), .ZN(n6804) );
  INV_X1 U7766 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6799) );
  AOI22_X1 U7767 ( .A1(n4115), .A2(keyinput254), .B1(n6799), .B2(keyinput199), 
        .ZN(n6798) );
  OAI221_X1 U7768 ( .B1(n4115), .B2(keyinput254), .C1(n6799), .C2(keyinput199), 
        .A(n6798), .ZN(n6803) );
  INV_X1 U7769 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6932) );
  XOR2_X1 U7770 ( .A(n6932), .B(keyinput156), .Z(n6801) );
  XNOR2_X1 U7771 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput212), .ZN(
        n6800) );
  NAND2_X1 U7772 ( .A1(n6801), .A2(n6800), .ZN(n6802) );
  NOR4_X1 U7773 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6845)
         );
  AOI22_X1 U7774 ( .A1(n6858), .A2(keyinput229), .B1(keyinput203), .B2(n6807), 
        .ZN(n6806) );
  OAI221_X1 U7775 ( .B1(n6858), .B2(keyinput229), .C1(n6807), .C2(keyinput203), 
        .A(n6806), .ZN(n6815) );
  AOI22_X1 U7776 ( .A1(n6966), .A2(keyinput174), .B1(keyinput247), .B2(n6916), 
        .ZN(n6808) );
  OAI221_X1 U7777 ( .B1(n6966), .B2(keyinput174), .C1(n6916), .C2(keyinput247), 
        .A(n6808), .ZN(n6814) );
  AOI22_X1 U7778 ( .A1(n4640), .A2(keyinput241), .B1(n4992), .B2(keyinput185), 
        .ZN(n6809) );
  OAI221_X1 U7779 ( .B1(n4640), .B2(keyinput241), .C1(n4992), .C2(keyinput185), 
        .A(n6809), .ZN(n6813) );
  INV_X1 U7780 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6811) );
  AOI22_X1 U7781 ( .A1(n6942), .A2(keyinput146), .B1(keyinput133), .B2(n6811), 
        .ZN(n6810) );
  OAI221_X1 U7782 ( .B1(n6942), .B2(keyinput146), .C1(n6811), .C2(keyinput133), 
        .A(n6810), .ZN(n6812) );
  NOR4_X1 U7783 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6844)
         );
  AOI22_X1 U7784 ( .A1(n6817), .A2(keyinput137), .B1(n6889), .B2(keyinput220), 
        .ZN(n6816) );
  OAI221_X1 U7785 ( .B1(n6817), .B2(keyinput137), .C1(n6889), .C2(keyinput220), 
        .A(n6816), .ZN(n6821) );
  XNOR2_X1 U7786 ( .A(n6818), .B(keyinput169), .ZN(n6820) );
  XNOR2_X1 U7787 ( .A(n6895), .B(keyinput202), .ZN(n6819) );
  OR3_X1 U7788 ( .A1(n6821), .A2(n6820), .A3(n6819), .ZN(n6827) );
  AOI22_X1 U7789 ( .A1(n6823), .A2(keyinput153), .B1(n6867), .B2(keyinput200), 
        .ZN(n6822) );
  OAI221_X1 U7790 ( .B1(n6823), .B2(keyinput153), .C1(n6867), .C2(keyinput200), 
        .A(n6822), .ZN(n6826) );
  AOI22_X1 U7791 ( .A1(n6943), .A2(keyinput161), .B1(keyinput232), .B2(n6960), 
        .ZN(n6824) );
  OAI221_X1 U7792 ( .B1(n6943), .B2(keyinput161), .C1(n6960), .C2(keyinput232), 
        .A(n6824), .ZN(n6825) );
  NOR3_X1 U7793 ( .A1(n6827), .A2(n6826), .A3(n6825), .ZN(n6843) );
  INV_X1 U7794 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6829) );
  AOI22_X1 U7795 ( .A1(n6829), .A2(keyinput231), .B1(keyinput164), .B2(n4346), 
        .ZN(n6828) );
  OAI221_X1 U7796 ( .B1(n6829), .B2(keyinput231), .C1(n4346), .C2(keyinput164), 
        .A(n6828), .ZN(n6841) );
  AOI22_X1 U7797 ( .A1(n6832), .A2(keyinput236), .B1(n6831), .B2(keyinput152), 
        .ZN(n6830) );
  OAI221_X1 U7798 ( .B1(n6832), .B2(keyinput236), .C1(n6831), .C2(keyinput152), 
        .A(n6830), .ZN(n6840) );
  INV_X1 U7799 ( .A(DATAI_30_), .ZN(n6927) );
  AOI22_X1 U7800 ( .A1(n6834), .A2(keyinput198), .B1(n6927), .B2(keyinput168), 
        .ZN(n6833) );
  OAI221_X1 U7801 ( .B1(n6834), .B2(keyinput198), .C1(n6927), .C2(keyinput168), 
        .A(n6833), .ZN(n6839) );
  AOI22_X1 U7802 ( .A1(n6837), .A2(keyinput165), .B1(keyinput251), .B2(n6836), 
        .ZN(n6835) );
  OAI221_X1 U7803 ( .B1(n6837), .B2(keyinput165), .C1(n6836), .C2(keyinput251), 
        .A(n6835), .ZN(n6838) );
  NOR4_X1 U7804 ( .A1(n6841), .A2(n6840), .A3(n6839), .A4(n6838), .ZN(n6842)
         );
  NAND4_X1 U7805 ( .A1(n6845), .A2(n6844), .A3(n6843), .A4(n6842), .ZN(n6846)
         );
  NOR4_X1 U7806 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6978)
         );
  INV_X1 U7807 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6851) );
  AOI22_X1 U7808 ( .A1(n6852), .A2(keyinput2), .B1(n6851), .B2(keyinput122), 
        .ZN(n6850) );
  OAI221_X1 U7809 ( .B1(n6852), .B2(keyinput2), .C1(n6851), .C2(keyinput122), 
        .A(n6850), .ZN(n6864) );
  AOI22_X1 U7810 ( .A1(n6855), .A2(keyinput32), .B1(keyinput95), .B2(n6854), 
        .ZN(n6853) );
  OAI221_X1 U7811 ( .B1(n6855), .B2(keyinput32), .C1(n6854), .C2(keyinput95), 
        .A(n6853), .ZN(n6863) );
  AOI22_X1 U7812 ( .A1(n6858), .A2(keyinput101), .B1(n6857), .B2(keyinput118), 
        .ZN(n6856) );
  OAI221_X1 U7813 ( .B1(n6858), .B2(keyinput101), .C1(n6857), .C2(keyinput118), 
        .A(n6856), .ZN(n6862) );
  INV_X1 U7814 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7815 ( .A1(n4115), .A2(keyinput126), .B1(n6860), .B2(keyinput93), 
        .ZN(n6859) );
  OAI221_X1 U7816 ( .B1(n4115), .B2(keyinput126), .C1(n6860), .C2(keyinput93), 
        .A(n6859), .ZN(n6861) );
  NOR4_X1 U7817 ( .A1(n6864), .A2(n6863), .A3(n6862), .A4(n6861), .ZN(n6910)
         );
  AOI22_X1 U7818 ( .A1(n6867), .A2(keyinput72), .B1(keyinput3), .B2(n6866), 
        .ZN(n6865) );
  OAI221_X1 U7819 ( .B1(n6867), .B2(keyinput72), .C1(n6866), .C2(keyinput3), 
        .A(n6865), .ZN(n6879) );
  AOI22_X1 U7820 ( .A1(n6869), .A2(keyinput56), .B1(keyinput120), .B2(n4939), 
        .ZN(n6868) );
  OAI221_X1 U7821 ( .B1(n6869), .B2(keyinput56), .C1(n4939), .C2(keyinput120), 
        .A(n6868), .ZN(n6878) );
  AOI22_X1 U7822 ( .A1(n6872), .A2(keyinput7), .B1(n6871), .B2(keyinput1), 
        .ZN(n6870) );
  OAI221_X1 U7823 ( .B1(n6872), .B2(keyinput7), .C1(n6871), .C2(keyinput1), 
        .A(n6870), .ZN(n6877) );
  AOI22_X1 U7824 ( .A1(n6875), .A2(keyinput85), .B1(n6874), .B2(keyinput80), 
        .ZN(n6873) );
  OAI221_X1 U7825 ( .B1(n6875), .B2(keyinput85), .C1(n6874), .C2(keyinput80), 
        .A(n6873), .ZN(n6876) );
  NOR4_X1 U7826 ( .A1(n6879), .A2(n6878), .A3(n6877), .A4(n6876), .ZN(n6909)
         );
  INV_X1 U7827 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6881) );
  AOI22_X1 U7828 ( .A1(n6882), .A2(keyinput125), .B1(n6881), .B2(keyinput0), 
        .ZN(n6880) );
  OAI221_X1 U7829 ( .B1(n6882), .B2(keyinput125), .C1(n6881), .C2(keyinput0), 
        .A(n6880), .ZN(n6893) );
  INV_X1 U7830 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6884) );
  AOI22_X1 U7831 ( .A1(n6884), .A2(keyinput88), .B1(n4845), .B2(keyinput30), 
        .ZN(n6883) );
  OAI221_X1 U7832 ( .B1(n6884), .B2(keyinput88), .C1(n4845), .C2(keyinput30), 
        .A(n6883), .ZN(n6892) );
  AOI22_X1 U7833 ( .A1(n6887), .A2(keyinput87), .B1(n6886), .B2(keyinput76), 
        .ZN(n6885) );
  OAI221_X1 U7834 ( .B1(n6887), .B2(keyinput87), .C1(n6886), .C2(keyinput76), 
        .A(n6885), .ZN(n6891) );
  AOI22_X1 U7835 ( .A1(n6889), .A2(keyinput92), .B1(n5238), .B2(keyinput58), 
        .ZN(n6888) );
  OAI221_X1 U7836 ( .B1(n6889), .B2(keyinput92), .C1(n5238), .C2(keyinput58), 
        .A(n6888), .ZN(n6890) );
  NOR4_X1 U7837 ( .A1(n6893), .A2(n6892), .A3(n6891), .A4(n6890), .ZN(n6908)
         );
  AOI22_X1 U7838 ( .A1(n4743), .A2(keyinput127), .B1(keyinput74), .B2(n6895), 
        .ZN(n6894) );
  OAI221_X1 U7839 ( .B1(n4743), .B2(keyinput127), .C1(n6895), .C2(keyinput74), 
        .A(n6894), .ZN(n6906) );
  AOI22_X1 U7840 ( .A1(n4346), .A2(keyinput36), .B1(keyinput22), .B2(n4471), 
        .ZN(n6896) );
  OAI221_X1 U7841 ( .B1(n4346), .B2(keyinput36), .C1(n4471), .C2(keyinput22), 
        .A(n6896), .ZN(n6905) );
  AOI22_X1 U7842 ( .A1(n6899), .A2(keyinput102), .B1(n6898), .B2(keyinput42), 
        .ZN(n6897) );
  OAI221_X1 U7843 ( .B1(n6899), .B2(keyinput102), .C1(n6898), .C2(keyinput42), 
        .A(n6897), .ZN(n6904) );
  AOI22_X1 U7844 ( .A1(n6902), .A2(keyinput20), .B1(keyinput81), .B2(n6901), 
        .ZN(n6900) );
  OAI221_X1 U7845 ( .B1(n6902), .B2(keyinput20), .C1(n6901), .C2(keyinput81), 
        .A(n6900), .ZN(n6903) );
  NOR4_X1 U7846 ( .A1(n6906), .A2(n6905), .A3(n6904), .A4(n6903), .ZN(n6907)
         );
  NAND4_X1 U7847 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n6977)
         );
  AOI22_X1 U7848 ( .A1(n6916), .A2(keyinput119), .B1(n6915), .B2(keyinput35), 
        .ZN(n6914) );
  OAI221_X1 U7849 ( .B1(n6916), .B2(keyinput119), .C1(n6915), .C2(keyinput35), 
        .A(n6914), .ZN(n6924) );
  AOI22_X1 U7850 ( .A1(n6919), .A2(keyinput39), .B1(keyinput97), .B2(n6918), 
        .ZN(n6917) );
  OAI221_X1 U7851 ( .B1(n6919), .B2(keyinput39), .C1(n6918), .C2(keyinput97), 
        .A(n6917), .ZN(n6923) );
  AOI22_X1 U7852 ( .A1(n6921), .A2(keyinput17), .B1(n4440), .B2(keyinput8), 
        .ZN(n6920) );
  OAI221_X1 U7853 ( .B1(n6921), .B2(keyinput17), .C1(n4440), .C2(keyinput8), 
        .A(n6920), .ZN(n6922) );
  NOR4_X1 U7854 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n6975)
         );
  AOI22_X1 U7855 ( .A1(n4640), .A2(keyinput113), .B1(keyinput40), .B2(n6927), 
        .ZN(n6926) );
  OAI221_X1 U7856 ( .B1(n4640), .B2(keyinput113), .C1(n6927), .C2(keyinput40), 
        .A(n6926), .ZN(n6940) );
  INV_X1 U7857 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6929) );
  AOI22_X1 U7858 ( .A1(n6930), .A2(keyinput53), .B1(n6929), .B2(keyinput23), 
        .ZN(n6928) );
  OAI221_X1 U7859 ( .B1(n6930), .B2(keyinput53), .C1(n6929), .C2(keyinput23), 
        .A(n6928), .ZN(n6939) );
  AOI22_X1 U7860 ( .A1(n6933), .A2(keyinput65), .B1(n6932), .B2(keyinput28), 
        .ZN(n6931) );
  OAI221_X1 U7861 ( .B1(n6933), .B2(keyinput65), .C1(n6932), .C2(keyinput28), 
        .A(n6931), .ZN(n6938) );
  INV_X1 U7862 ( .A(DATAI_12_), .ZN(n6935) );
  AOI22_X1 U7863 ( .A1(n6936), .A2(keyinput54), .B1(n6935), .B2(keyinput49), 
        .ZN(n6934) );
  OAI221_X1 U7864 ( .B1(n6936), .B2(keyinput54), .C1(n6935), .C2(keyinput49), 
        .A(n6934), .ZN(n6937) );
  NOR4_X1 U7865 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6974)
         );
  AOI22_X1 U7866 ( .A1(n6943), .A2(keyinput33), .B1(keyinput18), .B2(n6942), 
        .ZN(n6941) );
  OAI221_X1 U7867 ( .B1(n6943), .B2(keyinput33), .C1(n6942), .C2(keyinput18), 
        .A(n6941), .ZN(n6956) );
  AOI22_X1 U7868 ( .A1(n6946), .A2(keyinput99), .B1(keyinput86), .B2(n6945), 
        .ZN(n6944) );
  OAI221_X1 U7869 ( .B1(n6946), .B2(keyinput99), .C1(n6945), .C2(keyinput86), 
        .A(n6944), .ZN(n6955) );
  AOI22_X1 U7870 ( .A1(n6949), .A2(keyinput34), .B1(keyinput94), .B2(n6948), 
        .ZN(n6947) );
  OAI221_X1 U7871 ( .B1(n6949), .B2(keyinput34), .C1(n6948), .C2(keyinput94), 
        .A(n6947), .ZN(n6954) );
  INV_X1 U7872 ( .A(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n6952) );
  AOI22_X1 U7873 ( .A1(n6952), .A2(keyinput68), .B1(keyinput11), .B2(n6951), 
        .ZN(n6950) );
  OAI221_X1 U7874 ( .B1(n6952), .B2(keyinput68), .C1(n6951), .C2(keyinput11), 
        .A(n6950), .ZN(n6953) );
  NOR4_X1 U7875 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n6973)
         );
  AOI22_X1 U7876 ( .A1(n6958), .A2(keyinput29), .B1(n4345), .B2(keyinput67), 
        .ZN(n6957) );
  OAI221_X1 U7877 ( .B1(n6958), .B2(keyinput29), .C1(n4345), .C2(keyinput67), 
        .A(n6957), .ZN(n6971) );
  AOI22_X1 U7878 ( .A1(n6961), .A2(keyinput59), .B1(keyinput104), .B2(n6960), 
        .ZN(n6959) );
  OAI221_X1 U7879 ( .B1(n6961), .B2(keyinput59), .C1(n6960), .C2(keyinput104), 
        .A(n6959), .ZN(n6970) );
  AOI22_X1 U7880 ( .A1(n6964), .A2(keyinput31), .B1(n6963), .B2(keyinput45), 
        .ZN(n6962) );
  OAI221_X1 U7881 ( .B1(n6964), .B2(keyinput31), .C1(n6963), .C2(keyinput45), 
        .A(n6962), .ZN(n6969) );
  AOI22_X1 U7882 ( .A1(n6967), .A2(keyinput16), .B1(keyinput46), .B2(n6966), 
        .ZN(n6965) );
  OAI221_X1 U7883 ( .B1(n6967), .B2(keyinput16), .C1(n6966), .C2(keyinput46), 
        .A(n6965), .ZN(n6968) );
  NOR4_X1 U7884 ( .A1(n6971), .A2(n6970), .A3(n6969), .A4(n6968), .ZN(n6972)
         );
  NAND4_X1 U7885 ( .A1(n6975), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n6976)
         );
  NOR3_X1 U7886 ( .A1(n6978), .A2(n6977), .A3(n6976), .ZN(n7016) );
  OAI22_X1 U7887 ( .A1(BS16_N), .A2(keyinput38), .B1(keyinput109), .B2(
        ADDRESS_REG_0__SCAN_IN), .ZN(n6979) );
  AOI221_X1 U7888 ( .B1(BS16_N), .B2(keyinput38), .C1(ADDRESS_REG_0__SCAN_IN), 
        .C2(keyinput109), .A(n6979), .ZN(n6986) );
  OAI22_X1 U7889 ( .A1(EBX_REG_0__SCAN_IN), .A2(keyinput55), .B1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput124), .ZN(n6980) );
  AOI221_X1 U7890 ( .B1(EBX_REG_0__SCAN_IN), .B2(keyinput55), .C1(keyinput124), 
        .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n6980), .ZN(n6985) );
  OAI22_X1 U7891 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(keyinput71), .B1(
        LWORD_REG_4__SCAN_IN), .B2(keyinput78), .ZN(n6981) );
  AOI221_X1 U7892 ( .B1(INSTQUEUE_REG_12__4__SCAN_IN), .B2(keyinput71), .C1(
        keyinput78), .C2(LWORD_REG_4__SCAN_IN), .A(n6981), .ZN(n6984) );
  OAI22_X1 U7893 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(keyinput41), .B1(
        EAX_REG_14__SCAN_IN), .B2(keyinput96), .ZN(n6982) );
  AOI221_X1 U7894 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(keyinput41), 
        .C1(keyinput96), .C2(EAX_REG_14__SCAN_IN), .A(n6982), .ZN(n6983) );
  NAND4_X1 U7895 ( .A1(n6986), .A2(n6985), .A3(n6984), .A4(n6983), .ZN(n7014)
         );
  OAI22_X1 U7896 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(keyinput24), .B1(
        keyinput111), .B2(REIP_REG_21__SCAN_IN), .ZN(n6987) );
  AOI221_X1 U7897 ( .B1(INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput24), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput111), .A(n6987), .ZN(n6994) );
  OAI22_X1 U7898 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(keyinput66), .B1(
        DATAWIDTH_REG_28__SCAN_IN), .B2(keyinput9), .ZN(n6988) );
  AOI221_X1 U7899 ( .B1(INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput66), .C1(
        keyinput9), .C2(DATAWIDTH_REG_28__SCAN_IN), .A(n6988), .ZN(n6993) );
  OAI22_X1 U7900 ( .A1(REIP_REG_15__SCAN_IN), .A2(keyinput73), .B1(keyinput25), 
        .B2(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6989) );
  AOI221_X1 U7901 ( .B1(REIP_REG_15__SCAN_IN), .B2(keyinput73), .C1(
        DATAWIDTH_REG_25__SCAN_IN), .C2(keyinput25), .A(n6989), .ZN(n6992) );
  OAI22_X1 U7902 ( .A1(EAX_REG_9__SCAN_IN), .A2(keyinput63), .B1(keyinput105), 
        .B2(UWORD_REG_14__SCAN_IN), .ZN(n6990) );
  AOI221_X1 U7903 ( .B1(EAX_REG_9__SCAN_IN), .B2(keyinput63), .C1(
        UWORD_REG_14__SCAN_IN), .C2(keyinput105), .A(n6990), .ZN(n6991) );
  NAND4_X1 U7904 ( .A1(n6994), .A2(n6993), .A3(n6992), .A4(n6991), .ZN(n7013)
         );
  OAI22_X1 U7905 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(keyinput98), .B1(
        keyinput4), .B2(REIP_REG_25__SCAN_IN), .ZN(n6995) );
  AOI221_X1 U7906 ( .B1(INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput98), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput4), .A(n6995), .ZN(n7002) );
  OAI22_X1 U7907 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(keyinput110), .B1(
        DATAWIDTH_REG_30__SCAN_IN), .B2(keyinput114), .ZN(n6996) );
  AOI221_X1 U7908 ( .B1(INSTQUEUE_REG_10__1__SCAN_IN), .B2(keyinput110), .C1(
        keyinput114), .C2(DATAWIDTH_REG_30__SCAN_IN), .A(n6996), .ZN(n7001) );
  OAI22_X1 U7909 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(keyinput84), .B1(
        keyinput83), .B2(REIP_REG_10__SCAN_IN), .ZN(n6997) );
  AOI221_X1 U7910 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(keyinput84), 
        .C1(REIP_REG_10__SCAN_IN), .C2(keyinput83), .A(n6997), .ZN(n7000) );
  OAI22_X1 U7911 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(keyinput6), .B1(
        keyinput123), .B2(DATAO_REG_11__SCAN_IN), .ZN(n6998) );
  AOI221_X1 U7912 ( .B1(INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput6), .C1(
        DATAO_REG_11__SCAN_IN), .C2(keyinput123), .A(n6998), .ZN(n6999) );
  NAND4_X1 U7913 ( .A1(n7002), .A2(n7001), .A3(n7000), .A4(n6999), .ZN(n7012)
         );
  OAI22_X1 U7914 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(keyinput77), .B1(
        keyinput14), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7003) );
  AOI221_X1 U7915 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput77), 
        .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(keyinput14), .A(n7003), .ZN(
        n7010) );
  OAI22_X1 U7916 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(keyinput52), .B1(
        UWORD_REG_1__SCAN_IN), .B2(keyinput115), .ZN(n7004) );
  AOI221_X1 U7917 ( .B1(INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput52), .C1(
        keyinput115), .C2(UWORD_REG_1__SCAN_IN), .A(n7004), .ZN(n7009) );
  OAI22_X1 U7918 ( .A1(REIP_REG_9__SCAN_IN), .A2(keyinput121), .B1(keyinput116), .B2(REIP_REG_6__SCAN_IN), .ZN(n7005) );
  AOI221_X1 U7919 ( .B1(REIP_REG_9__SCAN_IN), .B2(keyinput121), .C1(
        REIP_REG_6__SCAN_IN), .C2(keyinput116), .A(n7005), .ZN(n7008) );
  OAI22_X1 U7920 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(keyinput100), .B1(
        keyinput37), .B2(EBX_REG_24__SCAN_IN), .ZN(n7006) );
  AOI221_X1 U7921 ( .B1(INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput100), .C1(
        EBX_REG_24__SCAN_IN), .C2(keyinput37), .A(n7006), .ZN(n7007) );
  NAND4_X1 U7922 ( .A1(n7010), .A2(n7009), .A3(n7008), .A4(n7007), .ZN(n7011)
         );
  NOR4_X1 U7923 ( .A1(n7014), .A2(n7013), .A3(n7012), .A4(n7011), .ZN(n7015)
         );
  NAND3_X1 U7924 ( .A1(n7017), .A2(n7016), .A3(n7015), .ZN(n7032) );
  AOI22_X1 U7925 ( .A1(n7021), .A2(n7020), .B1(n7019), .B2(n7018), .ZN(n7022)
         );
  OAI21_X1 U7926 ( .B1(n7024), .B2(n7023), .A(n7022), .ZN(n7025) );
  AOI21_X1 U7927 ( .B1(n7027), .B2(n7026), .A(n7025), .ZN(n7028) );
  OAI21_X1 U7928 ( .B1(n7030), .B2(n7029), .A(n7028), .ZN(n7031) );
  XNOR2_X1 U7929 ( .A(n7032), .B(n7031), .ZN(U3075) );
  INV_X1 U3647 ( .A(n4441), .ZN(n4413) );
  NOR2_X2 U3781 ( .A1(n3834), .A2(n3827), .ZN(n3505) );
  CLKBUF_X1 U3649 ( .A(n3348), .Z(n4442) );
  CLKBUF_X1 U3658 ( .A(n3419), .Z(n3801) );
  CLKBUF_X1 U3662 ( .A(n5544), .Z(n3204) );
  CLKBUF_X1 U3689 ( .A(n3418), .Z(n4858) );
  CLKBUF_X1 U3733 ( .A(n4128), .Z(n5311) );
  CLKBUF_X2 U3765 ( .A(n3472), .Z(n6092) );
  CLKBUF_X1 U3798 ( .A(n5362), .Z(n5363) );
endmodule

