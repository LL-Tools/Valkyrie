

module b21_C_SARLock_k_128_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229;

  OR2_X1 U4895 ( .A1(n7854), .A2(n8884), .ZN(n8791) );
  INV_X2 U4896 ( .A(n5121), .ZN(n5306) );
  NAND2_X2 U4897 ( .A1(n7383), .A2(n7314), .ZN(n8001) );
  AND2_X4 U4898 ( .A1(n5818), .A2(n8479), .ZN(n5895) );
  CLKBUF_X2 U4899 ( .A(n5096), .Z(n5732) );
  AND4_X1 U4900 ( .A1(n5823), .A2(n5822), .A3(n5821), .A4(n5820), .ZN(n7286)
         );
  INV_X1 U4901 ( .A(n8172), .ZN(n4641) );
  NAND2_X1 U4902 ( .A1(n6283), .A2(n8467), .ZN(n5860) );
  OAI21_X1 U4903 ( .B1(n4653), .B2(n4938), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4996) );
  INV_X2 U4904 ( .A(n5279), .ZN(n4655) );
  NOR2_X2 U4905 ( .A1(n5279), .A2(n4522), .ZN(n4994) );
  INV_X1 U4906 ( .A(n6186), .ZN(n6231) );
  AND2_X1 U4907 ( .A1(n8043), .A2(n8044), .ZN(n8135) );
  AND3_X1 U4908 ( .A1(n5867), .A2(n5803), .A3(n5804), .ZN(n4561) );
  AND2_X1 U4909 ( .A1(n7878), .A2(n6881), .ZN(n5743) );
  INV_X1 U4910 ( .A(n5167), .ZN(n5740) );
  NAND2_X1 U4911 ( .A1(n6308), .A2(n5497), .ZN(n5121) );
  NOR2_X1 U4912 ( .A1(n6888), .A2(n6891), .ZN(n6947) );
  INV_X1 U4913 ( .A(n6765), .ZN(n9786) );
  XNOR2_X1 U4914 ( .A(n7831), .B(n7830), .ZN(n7829) );
  INV_X1 U4915 ( .A(n7833), .ZN(n5846) );
  NAND2_X1 U4916 ( .A1(n6122), .A2(n6121), .ZN(n8878) );
  AND4_X1 U4917 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n6718)
         );
  XNOR2_X1 U4918 ( .A(n5633), .B(n5650), .ZN(n7235) );
  NAND4_X1 U4919 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n9023)
         );
  INV_X2 U4920 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U4921 ( .A1(n9459), .A2(n8557), .ZN(n4389) );
  NOR3_X2 U4923 ( .A1(n8791), .A2(n4634), .A3(n8863), .ZN(n4636) );
  OAI21_X2 U4924 ( .B1(n5364), .B2(n5363), .A(n5365), .ZN(n5388) );
  OAI21_X2 U4925 ( .B1(n5675), .B2(n4731), .A(n5679), .ZN(n5697) );
  NAND2_X2 U4926 ( .A1(n8744), .A2(n8457), .ZN(n8731) );
  XNOR2_X2 U4927 ( .A(n5304), .B(n4953), .ZN(n6382) );
  AOI211_X2 U4928 ( .C1(n8834), .C2(n8806), .A(n8473), .B(n8472), .ZN(n8474)
         );
  XNOR2_X2 U4929 ( .A(n4615), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6598) );
  XNOR2_X2 U4930 ( .A(n5831), .B(n5830), .ZN(n7970) );
  AND2_X4 U4931 ( .A1(n5819), .A2(n7933), .ZN(n5896) );
  AOI21_X2 U4932 ( .B1(n8504), .B2(n8734), .A(n8730), .ZN(n8713) );
  OR2_X1 U4933 ( .A1(n6278), .A2(n6269), .ZN(n6280) );
  AOI21_X1 U4934 ( .B1(n9211), .B2(n9085), .A(n9084), .ZN(n9198) );
  INV_X4 U4935 ( .A(n8748), .ZN(n8863) );
  NAND2_X1 U4936 ( .A1(n5323), .A2(n5322), .ZN(n7172) );
  NAND2_X1 U4937 ( .A1(n4813), .A2(n4811), .ZN(n4810) );
  AOI21_X1 U4938 ( .B1(n7186), .B2(n7182), .A(n7184), .ZN(n7271) );
  OR2_X1 U4939 ( .A1(n5622), .A2(n5621), .ZN(n5652) );
  NAND2_X1 U4940 ( .A1(n7121), .A2(n6010), .ZN(n7186) );
  NAND2_X1 U4941 ( .A1(n6086), .A2(n6085), .ZN(n8895) );
  OAI21_X1 U4942 ( .B1(n7313), .B2(n4851), .A(n4848), .ZN(n9751) );
  OR2_X1 U4943 ( .A1(n9741), .A2(n9732), .ZN(n9742) );
  NAND2_X1 U4944 ( .A1(n7434), .A2(n7367), .ZN(n8022) );
  NAND2_X1 U4945 ( .A1(n8276), .A2(n8240), .ZN(n6990) );
  NAND2_X1 U4946 ( .A1(n5988), .A2(n5987), .ZN(n7434) );
  NAND2_X1 U4947 ( .A1(n5216), .A2(n5215), .ZN(n7044) );
  NOR2_X1 U4948 ( .A1(n8541), .A2(n9763), .ZN(n8527) );
  AND2_X1 U4949 ( .A1(n6348), .A2(n5887), .ZN(n5892) );
  AND2_X1 U4950 ( .A1(n5129), .A2(n5128), .ZN(n9663) );
  AND2_X1 U4951 ( .A1(n5915), .A2(n5914), .ZN(n9799) );
  AND2_X1 U4952 ( .A1(n6759), .A2(n5854), .ZN(n6754) );
  NAND2_X1 U4953 ( .A1(n7988), .A2(n7987), .ZN(n7282) );
  NAND2_X1 U4954 ( .A1(n7984), .A2(n7986), .ZN(n6558) );
  NAND2_X2 U4955 ( .A1(n6955), .A2(n9274), .ZN(n9276) );
  INV_X1 U4956 ( .A(n6884), .ZN(n4643) );
  XNOR2_X1 U4957 ( .A(n9027), .B(n9640), .ZN(n6884) );
  NAND2_X1 U4958 ( .A1(n6557), .A2(n6708), .ZN(n7984) );
  NAND4_X1 U4959 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n6751)
         );
  BUF_X4 U4960 ( .A(n5871), .Z(n6186) );
  NAND2_X2 U4961 ( .A1(n5848), .A2(n4822), .ZN(n7241) );
  INV_X2 U4963 ( .A(n7969), .ZN(n6741) );
  AND2_X2 U4964 ( .A1(n6304), .A2(n6893), .ZN(n7878) );
  NAND4_X1 U4965 ( .A1(n5041), .A2(n5040), .A3(n5039), .A4(n5038), .ZN(n9025)
         );
  INV_X2 U4966 ( .A(n7960), .ZN(n7948) );
  NAND2_X1 U4967 ( .A1(n5815), .A2(n5816), .ZN(n7933) );
  XNOR2_X1 U4968 ( .A(n5186), .B(SI_6_), .ZN(n5183) );
  XNOR2_X1 U4969 ( .A(n5209), .B(SI_7_), .ZN(n5206) );
  XNOR2_X1 U4970 ( .A(n5817), .B(n7836), .ZN(n8479) );
  NAND2_X1 U4971 ( .A1(n5816), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5817) );
  XNOR2_X1 U4972 ( .A(n5117), .B(SI_4_), .ZN(n5142) );
  OR2_X1 U4973 ( .A1(n6096), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5835) );
  NAND3_X1 U4974 ( .A1(n4846), .A2(n4766), .A3(n4765), .ZN(n5845) );
  NAND2_X1 U4975 ( .A1(n5825), .A2(n5824), .ZN(n6096) );
  INV_X1 U4976 ( .A(n6066), .ZN(n4846) );
  INV_X2 U4977 ( .A(n7833), .ZN(n4390) );
  NAND2_X1 U4978 ( .A1(n4583), .A2(n4580), .ZN(n5279) );
  NAND2_X1 U4979 ( .A1(n4939), .A2(n4963), .ZN(n4522) );
  OAI21_X1 U4980 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n4733), .ZN(n4732) );
  AND2_X1 U4981 ( .A1(n5867), .A2(n5803), .ZN(n5910) );
  NOR2_X1 U4982 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4584) );
  NOR2_X1 U4983 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5803) );
  INV_X1 U4984 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4736) );
  INV_X4 U4985 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AOI22_X2 U4986 ( .A1(n7618), .A2(n7617), .B1(n6107), .B2(n6106), .ZN(n7726)
         );
  AND2_X1 U4987 ( .A1(n4557), .A2(n4556), .ZN(n4770) );
  NOR2_X1 U4988 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4557) );
  AND2_X1 U4989 ( .A1(n4559), .A2(n4558), .ZN(n4771) );
  NOR2_X1 U4990 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4559) );
  NOR2_X1 U4991 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4558) );
  AND2_X1 U4992 ( .A1(n5788), .A2(n5787), .ZN(n9092) );
  OR2_X1 U4993 ( .A1(n7888), .A2(n5783), .ZN(n5788) );
  AND2_X1 U4994 ( .A1(n8135), .A2(n8040), .ZN(n4555) );
  INV_X1 U4995 ( .A(n8081), .ZN(n4547) );
  NAND2_X1 U4996 ( .A1(n4542), .A2(n8720), .ZN(n4536) );
  AND2_X1 U4997 ( .A1(n8398), .A2(n9096), .ZN(n4481) );
  NOR2_X1 U4998 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5801) );
  OR2_X1 U4999 ( .A1(n9073), .A2(n8226), .ZN(n8268) );
  NOR2_X1 U5000 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  INV_X1 U5001 ( .A(n7933), .ZN(n5818) );
  OR2_X1 U5002 ( .A1(n8838), .A2(n8483), .ZN(n8094) );
  OR2_X1 U5003 ( .A1(n8854), .A2(n8538), .ZN(n8085) );
  OR2_X1 U5004 ( .A1(n8873), .A2(n8799), .ZN(n8071) );
  OR2_X1 U5005 ( .A1(n9459), .A2(n7642), .ZN(n8043) );
  OR2_X1 U5006 ( .A1(n7677), .A2(n7688), .ZN(n8048) );
  OR2_X1 U5007 ( .A1(n9732), .A2(n7464), .ZN(n8031) );
  OR2_X1 U5008 ( .A1(n8888), .A2(n7846), .ZN(n8063) );
  NOR2_X1 U5009 ( .A1(n5809), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U5010 ( .A1(n4412), .A2(n4500), .ZN(n4496) );
  NAND2_X1 U5011 ( .A1(n4955), .A2(n8427), .ZN(n8428) );
  NAND2_X1 U5012 ( .A1(n4738), .A2(n9069), .ZN(n8440) );
  NAND2_X1 U5013 ( .A1(n9144), .A2(n9157), .ZN(n9105) );
  OR2_X1 U5014 ( .A1(n9312), .A2(n9174), .ZN(n9090) );
  INV_X1 U5015 ( .A(n9172), .ZN(n4944) );
  OR2_X1 U5016 ( .A1(n9324), .A2(n9202), .ZN(n8395) );
  NOR2_X1 U5017 ( .A1(n9346), .A2(n9341), .ZN(n4607) );
  INV_X1 U5018 ( .A(n4923), .ZN(n4921) );
  OR2_X1 U5019 ( .A1(n9341), .A2(n9246), .ZN(n8398) );
  OR2_X1 U5020 ( .A1(n9356), .A2(n7800), .ZN(n8377) );
  OR2_X1 U5021 ( .A1(n9025), .A2(n9645), .ZN(n8193) );
  AND4_X1 U5022 ( .A1(n5473), .A2(n4962), .A3(n4961), .A4(n9938), .ZN(n4963)
         );
  AND3_X1 U5023 ( .A1(n4858), .A2(n4857), .A3(n4856), .ZN(n4939) );
  NOR2_X1 U5024 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4858) );
  NOR2_X1 U5025 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4856) );
  NOR2_X1 U5026 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4857) );
  OAI21_X1 U5027 ( .B1(n5492), .B2(n4730), .A(n5496), .ZN(n5514) );
  INV_X1 U5028 ( .A(n5493), .ZN(n4730) );
  XNOR2_X1 U5029 ( .A(n5330), .B(SI_11_), .ZN(n5329) );
  NAND2_X1 U5030 ( .A1(n5276), .A2(n5275), .ZN(n5305) );
  NAND2_X1 U5031 ( .A1(n5023), .A2(n4490), .ZN(n5044) );
  AOI21_X1 U5032 ( .B1(n7833), .B2(n4492), .A(n4491), .ZN(n4490) );
  NAND2_X1 U5033 ( .A1(n5860), .A2(n7826), .ZN(n5908) );
  OR2_X1 U5034 ( .A1(n6293), .A2(n9780), .ZN(n6282) );
  INV_X1 U5035 ( .A(n6552), .ZN(n8159) );
  NAND2_X1 U5036 ( .A1(n8647), .A2(n4637), .ZN(n8656) );
  INV_X1 U5037 ( .A(n8830), .ZN(n4637) );
  XNOR2_X1 U5038 ( .A(n8843), .B(n8550), .ZN(n8685) );
  OR2_X1 U5039 ( .A1(n8868), .A2(n8493), .ZN(n8749) );
  AND2_X1 U5040 ( .A1(n9737), .A2(n7461), .ZN(n7462) );
  AND2_X1 U5041 ( .A1(n7460), .A2(n9736), .ZN(n7461) );
  INV_X1 U5042 ( .A(n6068), .ZN(n5825) );
  AOI21_X1 U5043 ( .B1(n4875), .B2(n4505), .A(n4401), .ZN(n4504) );
  OR2_X1 U5044 ( .A1(n5608), .A2(n5607), .ZN(n5638) );
  INV_X1 U5045 ( .A(n8949), .ZN(n4892) );
  INV_X1 U5046 ( .A(n4997), .ZN(n4638) );
  NOR2_X1 U5047 ( .A1(n6503), .A2(n6502), .ZN(n6505) );
  AOI21_X1 U5048 ( .B1(n4904), .B2(n9145), .A(n4439), .ZN(n4902) );
  INV_X1 U5049 ( .A(n9157), .ZN(n9128) );
  NAND2_X1 U5050 ( .A1(n9107), .A2(n9108), .ZN(n9123) );
  AOI21_X1 U5051 ( .B1(n4408), .B2(n9103), .A(n4681), .ZN(n4680) );
  INV_X1 U5052 ( .A(n9104), .ZN(n4681) );
  NAND2_X1 U5053 ( .A1(n9324), .A2(n9202), .ZN(n9168) );
  NOR2_X1 U5054 ( .A1(n9200), .A2(n9199), .ZN(n9183) );
  NAND2_X1 U5055 ( .A1(n9228), .A2(n4948), .ZN(n9211) );
  NAND2_X1 U5056 ( .A1(n9095), .A2(n4411), .ZN(n4692) );
  NAND2_X1 U5057 ( .A1(n9299), .A2(n9443), .ZN(n4685) );
  OR2_X1 U5058 ( .A1(n7866), .A2(n4501), .ZN(n6304) );
  NAND2_X1 U5059 ( .A1(n5750), .A2(n4977), .ZN(n4501) );
  OR2_X1 U5060 ( .A1(n9509), .A2(n9508), .ZN(n4564) );
  MUX2_X1 U5061 ( .A(n8325), .B(n8324), .S(n8424), .Z(n8328) );
  AND2_X1 U5062 ( .A1(n8046), .A2(n8045), .ZN(n4554) );
  NAND2_X1 U5063 ( .A1(n4555), .A2(n8041), .ZN(n4553) );
  NOR2_X1 U5064 ( .A1(n4552), .A2(n4550), .ZN(n4549) );
  INV_X1 U5065 ( .A(n4555), .ZN(n4550) );
  INV_X1 U5066 ( .A(n8049), .ZN(n4552) );
  NAND2_X1 U5067 ( .A1(n8069), .A2(n8795), .ZN(n4532) );
  NOR2_X1 U5068 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  INV_X1 U5069 ( .A(n8060), .ZN(n4531) );
  OR2_X1 U5070 ( .A1(n4532), .A2(n4533), .ZN(n4529) );
  AND2_X1 U5071 ( .A1(n8066), .A2(n8063), .ZN(n4533) );
  AOI21_X1 U5072 ( .B1(n8075), .B2(n4537), .A(n4535), .ZN(n4534) );
  INV_X1 U5073 ( .A(n4540), .ZN(n4537) );
  NAND2_X1 U5074 ( .A1(n4443), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U5075 ( .A1(n8077), .A2(n4539), .ZN(n4538) );
  NAND2_X1 U5076 ( .A1(n4541), .A2(n4540), .ZN(n4539) );
  INV_X1 U5077 ( .A(n4542), .ZN(n4541) );
  AND2_X1 U5078 ( .A1(n8390), .A2(n4482), .ZN(n8394) );
  NOR2_X1 U5079 ( .A1(n9103), .A2(n4483), .ZN(n4482) );
  NAND2_X1 U5080 ( .A1(n4704), .A2(n4700), .ZN(n4699) );
  INV_X1 U5081 ( .A(n7824), .ZN(n4700) );
  NOR2_X1 U5082 ( .A1(n7326), .A2(n4754), .ZN(n4753) );
  INV_X1 U5083 ( .A(n8001), .ZN(n4754) );
  AND2_X1 U5084 ( .A1(n5148), .A2(n5143), .ZN(n4489) );
  OR2_X1 U5085 ( .A1(n5145), .A2(n5142), .ZN(n5148) );
  INV_X1 U5086 ( .A(n5152), .ZN(n5153) );
  NOR2_X1 U5087 ( .A1(n6082), .A2(n7668), .ZN(n4821) );
  NAND2_X1 U5088 ( .A1(n5840), .A2(n7200), .ZN(n5871) );
  NOR2_X1 U5089 ( .A1(n6718), .A2(n6741), .ZN(n5886) );
  OR2_X1 U5090 ( .A1(n8825), .A2(n7963), .ZN(n8111) );
  INV_X1 U5091 ( .A(n8094), .ZN(n4740) );
  OR2_X1 U5092 ( .A1(n8628), .A2(n4474), .ZN(n7905) );
  OR2_X1 U5093 ( .A1(n8833), .A2(n8670), .ZN(n8103) );
  NAND2_X1 U5094 ( .A1(n4396), .A2(n7940), .ZN(n4841) );
  NAND2_X1 U5095 ( .A1(n8763), .A2(n4635), .ZN(n4634) );
  OR2_X1 U5096 ( .A1(n8878), .A2(n8456), .ZN(n8067) );
  NAND2_X1 U5097 ( .A1(n8053), .A2(n4828), .ZN(n4826) );
  NAND2_X1 U5098 ( .A1(n7847), .A2(n7846), .ZN(n4827) );
  NOR2_X1 U5099 ( .A1(n7677), .A2(n9459), .ZN(n4627) );
  OR2_X1 U5100 ( .A1(n7434), .A2(n7367), .ZN(n8015) );
  INV_X1 U5101 ( .A(n4753), .ZN(n4752) );
  AOI21_X1 U5102 ( .B1(n4751), .B2(n4753), .A(n4750), .ZN(n4749) );
  INV_X1 U5103 ( .A(n8006), .ZN(n4750) );
  NOR2_X1 U5104 ( .A1(n7298), .A2(n8566), .ZN(n4832) );
  NAND2_X1 U5105 ( .A1(n7286), .A2(n7241), .ZN(n7986) );
  AND2_X1 U5106 ( .A1(n7973), .A2(n7972), .ZN(n4768) );
  AND2_X1 U5107 ( .A1(n4847), .A2(n5810), .ZN(n4766) );
  AND2_X1 U5108 ( .A1(n5802), .A2(n5801), .ZN(n4769) );
  NOR2_X1 U5109 ( .A1(n4516), .A2(n4510), .ZN(n4509) );
  INV_X1 U5110 ( .A(n7787), .ZN(n4510) );
  NOR2_X1 U5111 ( .A1(n5511), .A2(n8987), .ZN(n4516) );
  OAI21_X1 U5112 ( .B1(n4885), .B2(n4515), .A(n4514), .ZN(n4513) );
  INV_X1 U5113 ( .A(n8987), .ZN(n4515) );
  NAND2_X1 U5114 ( .A1(n5511), .A2(n4886), .ZN(n4514) );
  NOR2_X1 U5115 ( .A1(n5511), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U5116 ( .A1(n8269), .A2(n9287), .ZN(n8422) );
  OR2_X1 U5117 ( .A1(n9299), .A2(n9129), .ZN(n8418) );
  OR2_X1 U5118 ( .A1(n9312), .A2(n9089), .ZN(n8236) );
  INV_X1 U5119 ( .A(n9093), .ZN(n4696) );
  NAND2_X1 U5120 ( .A1(n7482), .A2(n7483), .ZN(n4651) );
  INV_X1 U5121 ( .A(n8206), .ZN(n4664) );
  NOR2_X1 U5122 ( .A1(n8326), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U5123 ( .A1(n7045), .A2(n4669), .ZN(n4668) );
  NOR2_X1 U5124 ( .A1(n4662), .A2(n4661), .ZN(n4660) );
  AND2_X1 U5125 ( .A1(n6949), .A2(n8307), .ZN(n4661) );
  INV_X1 U5126 ( .A(n8201), .ZN(n4662) );
  NAND2_X1 U5127 ( .A1(n4660), .A2(n4658), .ZN(n4657) );
  INV_X1 U5128 ( .A(n8307), .ZN(n4658) );
  OR2_X1 U5129 ( .A1(n9024), .A2(n6926), .ZN(n8270) );
  NOR2_X1 U5130 ( .A1(n7759), .A2(n9356), .ZN(n7801) );
  INV_X1 U5131 ( .A(n5676), .ZN(n4731) );
  AOI21_X1 U5132 ( .B1(n4725), .B2(n4727), .A(n4722), .ZN(n4721) );
  INV_X1 U5133 ( .A(n5575), .ZN(n4722) );
  NOR2_X1 U5134 ( .A1(n5545), .A2(n4729), .ZN(n4728) );
  INV_X1 U5135 ( .A(n5516), .ZN(n4729) );
  AOI21_X1 U5136 ( .B1(n4711), .B2(n4710), .A(n4436), .ZN(n4709) );
  NAND2_X1 U5137 ( .A1(n5365), .A2(n5339), .ZN(n5363) );
  NAND2_X1 U5138 ( .A1(n5274), .A2(n5273), .ZN(n5304) );
  AND2_X1 U5139 ( .A1(n5305), .A2(n5278), .ZN(n4953) );
  INV_X1 U5140 ( .A(n5183), .ZN(n5184) );
  OAI21_X1 U5141 ( .B1(n5846), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4484), .ZN(
        n5117) );
  NAND2_X1 U5142 ( .A1(n5846), .A2(n5095), .ZN(n4484) );
  INV_X1 U5143 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U5144 ( .A1(n6850), .A2(n4786), .ZN(n4784) );
  INV_X1 U5145 ( .A(n6871), .ZN(n4797) );
  NOR2_X1 U5146 ( .A1(n6871), .A2(n4799), .ZN(n4798) );
  NAND2_X1 U5147 ( .A1(n4802), .A2(n4801), .ZN(n4800) );
  INV_X1 U5148 ( .A(n6824), .ZN(n4801) );
  INV_X1 U5149 ( .A(n6826), .ZN(n4802) );
  AOI21_X1 U5150 ( .B1(n4774), .B2(n4777), .A(n4431), .ZN(n4772) );
  INV_X1 U5151 ( .A(n4774), .ZN(n4773) );
  OR2_X1 U5152 ( .A1(n6810), .A2(n6807), .ZN(n6811) );
  OR2_X1 U5153 ( .A1(n8501), .A2(n4795), .ZN(n4794) );
  INV_X1 U5154 ( .A(n8500), .ZN(n4795) );
  AND2_X1 U5155 ( .A1(n8111), .A2(n8107), .ZN(n8148) );
  NAND2_X2 U5156 ( .A1(n6266), .A2(n8707), .ZN(n7969) );
  OR2_X1 U5157 ( .A1(n5912), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U5158 ( .A1(n8573), .A2(n8574), .ZN(n8572) );
  OR2_X1 U5159 ( .A1(n6732), .A2(n6731), .ZN(n4614) );
  NOR2_X1 U5160 ( .A1(n8630), .A2(n8629), .ZN(n8628) );
  OAI21_X1 U5161 ( .B1(n5844), .B2(n4622), .A(n4620), .ZN(n8467) );
  NAND2_X1 U5162 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n4622) );
  NOR2_X1 U5163 ( .A1(n5812), .A2(n4621), .ZN(n4620) );
  NOR2_X1 U5164 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4621) );
  AND4_X1 U5165 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n8483)
         );
  NAND2_X1 U5166 ( .A1(n8696), .A2(n7946), .ZN(n8699) );
  NOR2_X1 U5167 ( .A1(n8746), .A2(n8858), .ZN(n8714) );
  NAND2_X1 U5168 ( .A1(n4760), .A2(n8076), .ZN(n4759) );
  NAND2_X1 U5169 ( .A1(n7944), .A2(n4763), .ZN(n4760) );
  NAND2_X1 U5170 ( .A1(n4834), .A2(n4838), .ZN(n8744) );
  AOI21_X1 U5171 ( .B1(n4843), .B2(n4841), .A(n4839), .ZN(n4838) );
  NAND2_X1 U5172 ( .A1(n8775), .A2(n4835), .ZN(n4834) );
  NOR2_X1 U5173 ( .A1(n4840), .A2(n4836), .ZN(n4835) );
  INV_X1 U5174 ( .A(n4841), .ZN(n4840) );
  NOR2_X1 U5175 ( .A1(n8873), .A2(n8878), .ZN(n4635) );
  OR2_X1 U5176 ( .A1(n8873), .A2(n8551), .ZN(n4844) );
  NAND2_X1 U5177 ( .A1(n8775), .A2(n4959), .ZN(n4845) );
  NAND2_X1 U5178 ( .A1(n7938), .A2(n7937), .ZN(n8796) );
  NAND2_X1 U5179 ( .A1(n7814), .A2(n8141), .ZN(n7938) );
  AND2_X1 U5180 ( .A1(n8899), .A2(n8555), .ZN(n7706) );
  NAND2_X1 U5181 ( .A1(n7709), .A2(n8139), .ZN(n7807) );
  AOI21_X1 U5182 ( .B1(n4854), .B2(n4853), .A(n4389), .ZN(n4852) );
  AND2_X1 U5183 ( .A1(n8135), .A2(n7496), .ZN(n4767) );
  AND4_X1 U5184 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(n7499)
         );
  AND4_X1 U5185 ( .A1(n6065), .A2(n6064), .A3(n6063), .A4(n6062), .ZN(n7688)
         );
  NAND2_X1 U5186 ( .A1(n7462), .A2(n8041), .ZN(n7503) );
  NAND2_X1 U5187 ( .A1(n4956), .A2(n4853), .ZN(n7497) );
  AND2_X1 U5188 ( .A1(n9728), .A2(n8031), .ZN(n4956) );
  AND2_X1 U5189 ( .A1(n4957), .A2(n7319), .ZN(n4833) );
  NAND2_X1 U5190 ( .A1(n6007), .A2(n6006), .ZN(n7456) );
  NAND2_X1 U5191 ( .A1(n7370), .A2(n8131), .ZN(n4478) );
  AND4_X1 U5192 ( .A1(n6003), .A2(n6002), .A3(n6001), .A4(n6000), .ZN(n7455)
         );
  AOI21_X1 U5193 ( .B1(n4850), .B2(n8820), .A(n4428), .ZN(n4848) );
  AND4_X1 U5195 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n9762)
         );
  AND2_X1 U5196 ( .A1(n8006), .A2(n8005), .ZN(n8128) );
  AND4_X1 U5197 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n5964), .ZN(n7384)
         );
  INV_X1 U5198 ( .A(n8128), .ZN(n7316) );
  AND2_X1 U5199 ( .A1(n7998), .A2(n8001), .ZN(n8820) );
  NAND2_X1 U5200 ( .A1(n8810), .A2(n8820), .ZN(n8809) );
  AND4_X1 U5201 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n7348)
         );
  NAND2_X1 U5202 ( .A1(n7353), .A2(n8125), .ZN(n7352) );
  NAND2_X1 U5203 ( .A1(n7285), .A2(n7987), .ZN(n6717) );
  AND4_X1 U5204 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n7297)
         );
  OAI21_X1 U5205 ( .B1(n7960), .B2(n6355), .A(n5849), .ZN(n4823) );
  NAND2_X1 U5206 ( .A1(n6193), .A2(n6192), .ZN(n8849) );
  NAND2_X1 U5207 ( .A1(n6147), .A2(n6146), .ZN(n8868) );
  NAND2_X1 U5208 ( .A1(n4809), .A2(n4808), .ZN(n4807) );
  NOR2_X1 U5209 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4808) );
  INV_X1 U5210 ( .A(n5835), .ZN(n5834) );
  INV_X1 U5211 ( .A(n5747), .ZN(n4894) );
  INV_X1 U5212 ( .A(n5362), .ZN(n4507) );
  AND2_X1 U5213 ( .A1(n8965), .A2(n5542), .ZN(n8931) );
  NAND2_X1 U5214 ( .A1(n5192), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U5215 ( .A1(n4878), .A2(n4876), .ZN(n7732) );
  NOR2_X1 U5216 ( .A1(n7734), .A2(n4877), .ZN(n4876) );
  INV_X1 U5217 ( .A(n4879), .ZN(n4877) );
  INV_X1 U5218 ( .A(n5205), .ZN(n4500) );
  NAND2_X1 U5219 ( .A1(n4499), .A2(n5205), .ZN(n4498) );
  INV_X1 U5220 ( .A(n5202), .ZN(n4499) );
  AOI21_X1 U5221 ( .B1(n5743), .B2(n6888), .A(n5010), .ZN(n6455) );
  NAND2_X1 U5222 ( .A1(n5478), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5502) );
  INV_X1 U5223 ( .A(n5480), .ZN(n5478) );
  NOR2_X1 U5224 ( .A1(n5161), .A2(n5160), .ZN(n5192) );
  NAND2_X1 U5225 ( .A1(n4435), .A2(n4891), .ZN(n4890) );
  NAND2_X1 U5226 ( .A1(n4892), .A2(n5674), .ZN(n4891) );
  NAND2_X1 U5227 ( .A1(n5428), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5454) );
  INV_X1 U5228 ( .A(n5430), .ZN(n5428) );
  NAND2_X1 U5229 ( .A1(n4591), .A2(n4589), .ZN(n5007) );
  NAND2_X1 U5230 ( .A1(n4590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U5231 ( .A1(n4592), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4591) );
  OR2_X1 U5232 ( .A1(n5104), .A2(n6451), .ZN(n5001) );
  NAND2_X1 U5233 ( .A1(n6408), .A2(n4563), .ZN(n6477) );
  NOR2_X1 U5234 ( .A1(n6331), .A2(n4562), .ZN(n4563) );
  INV_X1 U5235 ( .A(n6330), .ZN(n4562) );
  OR2_X1 U5236 ( .A1(n6473), .A2(n6472), .ZN(n6475) );
  OR2_X1 U5237 ( .A1(n6508), .A2(n6509), .ZN(n9513) );
  NOR2_X1 U5238 ( .A1(n6339), .A2(n6338), .ZN(n6624) );
  OR2_X1 U5239 ( .A1(n6627), .A2(n6626), .ZN(n4570) );
  OR2_X1 U5240 ( .A1(n9564), .A2(n4471), .ZN(n4574) );
  XNOR2_X1 U5241 ( .A(n9060), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9062) );
  XNOR2_X1 U5242 ( .A(n9041), .B(n4578), .ZN(n9063) );
  INV_X1 U5243 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n4578) );
  NOR2_X1 U5244 ( .A1(n9130), .A2(n9299), .ZN(n9115) );
  AOI21_X1 U5245 ( .B1(n4394), .B2(n4678), .A(n8298), .ZN(n4672) );
  NAND2_X1 U5246 ( .A1(n4902), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U5247 ( .A1(n4900), .A2(n4903), .ZN(n4899) );
  INV_X1 U5248 ( .A(n5707), .ZN(n5705) );
  OR2_X1 U5249 ( .A1(n9317), .A2(n9006), .ZN(n9153) );
  AOI21_X1 U5250 ( .B1(n4942), .B2(n4941), .A(n4437), .ZN(n4940) );
  INV_X1 U5251 ( .A(n9187), .ZN(n4941) );
  AND2_X1 U5252 ( .A1(n9153), .A2(n8299), .ZN(n9172) );
  NAND2_X1 U5253 ( .A1(n8395), .A2(n9168), .ZN(n9187) );
  AND2_X1 U5254 ( .A1(n5665), .A2(n5664), .ZN(n9202) );
  AND2_X1 U5255 ( .A1(n5614), .A2(n5613), .ZN(n9233) );
  AOI21_X1 U5256 ( .B1(n4411), .B2(n9094), .A(n4695), .ZN(n4694) );
  INV_X1 U5257 ( .A(n9096), .ZN(n4695) );
  OR2_X1 U5258 ( .A1(n5554), .A2(n5553), .ZN(n5580) );
  AND2_X1 U5259 ( .A1(n5587), .A2(n5586), .ZN(n9246) );
  NOR2_X1 U5260 ( .A1(n4423), .A2(n4924), .ZN(n4923) );
  NOR2_X1 U5261 ( .A1(n9079), .A2(n4925), .ZN(n4924) );
  INV_X1 U5262 ( .A(n4927), .ZN(n4925) );
  AND2_X1 U5263 ( .A1(n8378), .A2(n9096), .ZN(n9244) );
  INV_X1 U5264 ( .A(n9079), .ZN(n4926) );
  OR2_X1 U5265 ( .A1(n5502), .A2(n9982), .ZN(n5527) );
  AOI21_X1 U5266 ( .B1(n7798), .B2(n8372), .A(n7797), .ZN(n9095) );
  AND2_X1 U5267 ( .A1(n9356), .A2(n9011), .ZN(n4927) );
  AND2_X1 U5268 ( .A1(n8377), .A2(n8186), .ZN(n8259) );
  NOR2_X1 U5269 ( .A1(n7747), .A2(n8259), .ZN(n7795) );
  AOI22_X1 U5270 ( .A1(n7745), .A2(n7744), .B1(n9013), .B2(n7743), .ZN(n7758)
         );
  NAND2_X1 U5271 ( .A1(n7440), .A2(n4930), .ZN(n4929) );
  NOR2_X1 U5272 ( .A1(n4931), .A2(n4434), .ZN(n4930) );
  INV_X1 U5273 ( .A(n4947), .ZN(n4931) );
  AOI21_X1 U5274 ( .B1(n4649), .B2(n4647), .A(n4646), .ZN(n4645) );
  INV_X1 U5275 ( .A(n4649), .ZN(n4648) );
  INV_X1 U5276 ( .A(n8354), .ZN(n4646) );
  OR2_X1 U5277 ( .A1(n9371), .A2(n7529), .ZN(n4947) );
  INV_X1 U5278 ( .A(n4913), .ZN(n4912) );
  OAI21_X1 U5279 ( .B1(n8251), .B2(n4914), .A(n7438), .ZN(n4913) );
  INV_X1 U5280 ( .A(n7245), .ZN(n4918) );
  AND2_X1 U5281 ( .A1(n8343), .A2(n8342), .ZN(n8251) );
  OR2_X1 U5282 ( .A1(n5219), .A2(n5218), .ZN(n5245) );
  OAI21_X1 U5283 ( .B1(n7028), .B2(n4935), .A(n4932), .ZN(n7106) );
  AOI21_X1 U5284 ( .B1(n4934), .B2(n4933), .A(n4400), .ZN(n4932) );
  AND2_X1 U5285 ( .A1(n6941), .A2(n6939), .ZN(n4906) );
  NAND2_X1 U5286 ( .A1(n4909), .A2(n4907), .ZN(n7058) );
  NOR2_X1 U5287 ( .A1(n4951), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U5288 ( .A1(n4644), .A2(n6948), .ZN(n8197) );
  NAND2_X1 U5289 ( .A1(n5552), .A2(n5551), .ZN(n9346) );
  AND2_X1 U5290 ( .A1(n6439), .A2(n5767), .ZN(n9443) );
  AND3_X1 U5291 ( .A1(n5054), .A2(n5053), .A3(n5052), .ZN(n9645) );
  XNOR2_X1 U5292 ( .A(n4706), .B(n7835), .ZN(n8162) );
  OAI21_X1 U5293 ( .B1(n7829), .B2(n4707), .A(n7832), .ZN(n4706) );
  NAND2_X1 U5294 ( .A1(n7841), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4945) );
  XNOR2_X1 U5295 ( .A(n7829), .B(SI_30_), .ZN(n8165) );
  AND3_X1 U5296 ( .A1(n4967), .A2(n4966), .A3(n4965), .ZN(n4992) );
  AND2_X1 U5297 ( .A1(n4969), .A2(n5769), .ZN(n4965) );
  AND2_X1 U5298 ( .A1(n4991), .A2(n5005), .ZN(n4654) );
  INV_X1 U5299 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4995) );
  XNOR2_X1 U5300 ( .A(n7825), .B(n7704), .ZN(n8174) );
  OAI21_X1 U5301 ( .B1(n6219), .B2(n4704), .A(n4702), .ZN(n7825) );
  NAND2_X1 U5302 ( .A1(n4994), .A2(n4992), .ZN(n4972) );
  NOR2_X1 U5303 ( .A1(n4415), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4520) );
  INV_X1 U5304 ( .A(n4522), .ZN(n4521) );
  NAND2_X1 U5305 ( .A1(n5517), .A2(n5516), .ZN(n5546) );
  AND4_X1 U5306 ( .A1(n4588), .A2(n10058), .A3(n4582), .A4(n4581), .ZN(n4580)
         );
  AND4_X1 U5307 ( .A1(n4584), .A2(n4586), .A3(n4587), .A4(n4585), .ZN(n4583)
         );
  NOR2_X1 U5308 ( .A1(n5122), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5125) );
  OR2_X1 U5309 ( .A1(n5050), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U5310 ( .A1(n5047), .A2(n5046), .ZN(n5074) );
  XNOR2_X1 U5311 ( .A(n5075), .B(SI_2_), .ZN(n5073) );
  AND2_X1 U5312 ( .A1(n4588), .A2(n4587), .ZN(n5049) );
  NAND2_X1 U5313 ( .A1(n7842), .A2(n4586), .ZN(n4572) );
  INV_X1 U5314 ( .A(n6809), .ZN(n4805) );
  NAND2_X1 U5315 ( .A1(n6205), .A2(n6204), .ZN(n8843) );
  NAND2_X1 U5316 ( .A1(n7583), .A2(n7962), .ZN(n6205) );
  INV_X1 U5317 ( .A(n4782), .ZN(n4781) );
  OAI21_X1 U5318 ( .B1(n4783), .B2(n4785), .A(n6964), .ZN(n4782) );
  INV_X1 U5319 ( .A(n4784), .ZN(n4783) );
  NAND2_X1 U5320 ( .A1(n4780), .A2(n4784), .ZN(n6965) );
  NAND2_X1 U5321 ( .A1(n6848), .A2(n4785), .ZN(n4780) );
  INV_X1 U5322 ( .A(n6180), .ZN(n6181) );
  INV_X1 U5323 ( .A(n6179), .ZN(n6182) );
  NAND2_X1 U5324 ( .A1(n6028), .A2(n6027), .ZN(n8037) );
  OR2_X1 U5325 ( .A1(n6282), .A2(n6274), .ZN(n8522) );
  OR2_X1 U5326 ( .A1(n8156), .A2(n4525), .ZN(n4524) );
  AND2_X1 U5327 ( .A1(n8155), .A2(n8154), .ZN(n4525) );
  INV_X1 U5328 ( .A(n8160), .ZN(n4744) );
  NAND4_X1 U5329 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n8565)
         );
  INV_X1 U5330 ( .A(n8647), .ZN(n8654) );
  OR2_X1 U5331 ( .A1(n9780), .A2(n6543), .ZN(n8817) );
  AND2_X1 U5332 ( .A1(n7887), .A2(n9002), .ZN(n4518) );
  NAND2_X1 U5333 ( .A1(n7877), .A2(n7876), .ZN(n9303) );
  AND2_X1 U5334 ( .A1(n4895), .A2(n4449), .ZN(n7897) );
  XNOR2_X1 U5335 ( .A(n5029), .B(n7881), .ZN(n6520) );
  NAND2_X1 U5336 ( .A1(n7172), .A2(n5328), .ZN(n9441) );
  INV_X1 U5337 ( .A(n9324), .ZN(n9192) );
  NAND2_X1 U5338 ( .A1(n5373), .A2(n5372), .ZN(n7521) );
  OAI21_X1 U5339 ( .B1(n4720), .B2(n7020), .A(n4718), .ZN(n4717) );
  MUX2_X1 U5340 ( .A(n8435), .B(n8434), .S(n9275), .Z(n4720) );
  NOR2_X1 U5341 ( .A1(n4416), .A2(n4719), .ZN(n4718) );
  INV_X1 U5342 ( .A(n9092), .ZN(n9147) );
  NOR2_X1 U5343 ( .A1(n6505), .A2(n4425), .ZN(n9509) );
  NOR2_X1 U5344 ( .A1(n9566), .A2(n9565), .ZN(n9564) );
  XNOR2_X1 U5345 ( .A(n4574), .B(n9581), .ZN(n9583) );
  AND2_X1 U5346 ( .A1(n4488), .A2(n4486), .ZN(n4576) );
  NOR2_X1 U5347 ( .A1(n9621), .A2(n6909), .ZN(n4488) );
  OR2_X1 U5348 ( .A1(n9062), .A2(n4487), .ZN(n4486) );
  OR2_X1 U5349 ( .A1(n9063), .A2(n9575), .ZN(n4577) );
  NAND2_X1 U5350 ( .A1(n4673), .A2(n4675), .ZN(n9126) );
  OR2_X1 U5351 ( .A1(n9170), .A2(n4678), .ZN(n4673) );
  NAND2_X1 U5352 ( .A1(n4905), .A2(n4904), .ZN(n9122) );
  AND2_X1 U5353 ( .A1(n4905), .A2(n4419), .ZN(n9124) );
  NAND2_X1 U5354 ( .A1(n4686), .A2(n4683), .ZN(n9380) );
  INV_X1 U5355 ( .A(n9297), .ZN(n4686) );
  NOR2_X1 U5356 ( .A1(n9298), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U5357 ( .A1(n9300), .A2(n4685), .ZN(n4684) );
  NAND2_X1 U5358 ( .A1(n4409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5006) );
  AOI21_X1 U5359 ( .B1(n4438), .B2(n8049), .A(n8138), .ZN(n4551) );
  NOR2_X1 U5360 ( .A1(n8081), .A2(n8112), .ZN(n4545) );
  AND2_X1 U5361 ( .A1(n4546), .A2(n4543), .ZN(n4542) );
  NAND2_X1 U5362 ( .A1(n8079), .A2(n7943), .ZN(n4543) );
  AND2_X1 U5363 ( .A1(n4529), .A2(n4452), .ZN(n4528) );
  NAND2_X1 U5364 ( .A1(n4546), .A2(n8098), .ZN(n4540) );
  NOR2_X1 U5365 ( .A1(n8392), .A2(n8400), .ZN(n4483) );
  NAND2_X1 U5366 ( .A1(n4544), .A2(n8084), .ZN(n8088) );
  NAND2_X1 U5367 ( .A1(n4538), .A2(n4534), .ZN(n4544) );
  NAND2_X1 U5368 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  AOI21_X1 U5369 ( .B1(n6219), .B2(n4701), .A(n4698), .ZN(n4697) );
  NOR2_X1 U5370 ( .A1(n4703), .A2(n7824), .ZN(n4701) );
  OAI21_X1 U5371 ( .B1(n4703), .B2(n4699), .A(n7823), .ZN(n4698) );
  INV_X1 U5372 ( .A(n4726), .ZN(n4725) );
  OAI21_X1 U5373 ( .B1(n4728), .B2(n4727), .A(n5573), .ZN(n4726) );
  INV_X1 U5374 ( .A(n5544), .ZN(n4727) );
  INV_X1 U5375 ( .A(n5305), .ZN(n4712) );
  INV_X1 U5376 ( .A(n5329), .ZN(n5332) );
  INV_X1 U5377 ( .A(n4953), .ZN(n4710) );
  NAND2_X1 U5378 ( .A1(n5269), .A2(n5238), .ZN(n5265) );
  INV_X1 U5379 ( .A(n6849), .ZN(n4786) );
  AND2_X1 U5380 ( .A1(n7778), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U5381 ( .A1(n7769), .A2(n4776), .ZN(n4775) );
  OR2_X1 U5382 ( .A1(n8849), .A2(n8503), .ZN(n8087) );
  INV_X1 U5383 ( .A(n4959), .ZN(n4836) );
  AND2_X1 U5384 ( .A1(n4626), .A2(n4627), .ZN(n4625) );
  AND2_X1 U5385 ( .A1(n6060), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6072) );
  NOR2_X1 U5386 ( .A1(n9810), .A2(n7314), .ZN(n4630) );
  NAND2_X1 U5387 ( .A1(n8570), .A2(n9786), .ZN(n7988) );
  AND2_X1 U5388 ( .A1(n5826), .A2(n5832), .ZN(n4809) );
  AND2_X1 U5389 ( .A1(n5802), .A2(n5801), .ZN(n4560) );
  INV_X1 U5390 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5909) );
  INV_X1 U5391 ( .A(n8978), .ZN(n4869) );
  AOI21_X1 U5392 ( .B1(n4864), .B2(n4867), .A(n4458), .ZN(n4863) );
  INV_X1 U5393 ( .A(n4868), .ZN(n4864) );
  INV_X1 U5394 ( .A(n4867), .ZN(n4865) );
  INV_X1 U5395 ( .A(n5743), .ZN(n7884) );
  NAND2_X1 U5396 ( .A1(n4593), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5397 ( .A1(n4994), .A2(n4993), .ZN(n4593) );
  AND2_X1 U5398 ( .A1(n8440), .A2(n4446), .ZN(n4737) );
  AOI21_X1 U5399 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9552), .A(n9048), .ZN(
        n9050) );
  NAND2_X1 U5400 ( .A1(n9306), .A2(n9128), .ZN(n8411) );
  AND2_X1 U5401 ( .A1(n9215), .A2(n4607), .ZN(n4606) );
  AND2_X1 U5402 ( .A1(n9215), .A2(n9083), .ZN(n9100) );
  OR2_X1 U5403 ( .A1(n5454), .A2(n7737), .ZN(n5480) );
  OR2_X1 U5404 ( .A1(n9365), .A2(n9014), .ZN(n7630) );
  NOR2_X1 U5405 ( .A1(n7628), .A2(n9365), .ZN(n4603) );
  NOR2_X1 U5406 ( .A1(n8253), .A2(n4650), .ZN(n4649) );
  INV_X1 U5407 ( .A(n8210), .ZN(n4650) );
  NAND2_X1 U5408 ( .A1(n4916), .A2(n4918), .ZN(n4914) );
  NOR2_X1 U5409 ( .A1(n8251), .A2(n4917), .ZN(n4915) );
  NOR2_X1 U5410 ( .A1(n7128), .A2(n7103), .ZN(n4598) );
  NAND2_X1 U5411 ( .A1(n4611), .A2(n4610), .ZN(n9130) );
  INV_X1 U5412 ( .A(n9191), .ZN(n4610) );
  NOR2_X1 U5413 ( .A1(n4391), .A2(n4612), .ZN(n4611) );
  NAND2_X1 U5414 ( .A1(n9136), .A2(n9144), .ZN(n4612) );
  NAND2_X1 U5415 ( .A1(n9203), .A2(n9192), .ZN(n9191) );
  AND2_X1 U5416 ( .A1(n9248), .A2(n4604), .ZN(n9203) );
  NOR2_X1 U5417 ( .A1(n4605), .A2(n9331), .ZN(n4604) );
  INV_X1 U5418 ( .A(n4606), .ZN(n4605) );
  NAND2_X1 U5419 ( .A1(n9248), .A2(n9259), .ZN(n9249) );
  AND2_X1 U5420 ( .A1(n7801), .A2(n9078), .ZN(n9248) );
  NOR2_X1 U5421 ( .A1(n6938), .A2(n7084), .ZN(n9272) );
  NAND2_X1 U5422 ( .A1(n6926), .A2(n4594), .ZN(n7084) );
  INV_X1 U5423 ( .A(n7011), .ZN(n4594) );
  INV_X1 U5424 ( .A(SI_30_), .ZN(n4707) );
  INV_X1 U5425 ( .A(n7698), .ZN(n4704) );
  AND2_X1 U5426 ( .A1(n4992), .A2(n4991), .ZN(n4993) );
  OAI21_X1 U5427 ( .B1(n5697), .B2(n5696), .A(n5698), .ZN(n5721) );
  INV_X1 U5428 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5769) );
  INV_X1 U5429 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U5430 ( .A1(n4978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4982) );
  INV_X1 U5431 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5473) );
  INV_X1 U5432 ( .A(n5265), .ZN(n5272) );
  NAND2_X1 U5433 ( .A1(n5148), .A2(n4950), .ZN(n5149) );
  XNOR2_X1 U5434 ( .A(n5140), .B(SI_5_), .ZN(n5152) );
  INV_X1 U5435 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5048) );
  AOI21_X1 U5436 ( .B1(n4790), .B2(n4793), .A(n6203), .ZN(n4788) );
  INV_X1 U5437 ( .A(n7476), .ZN(n4819) );
  OR2_X1 U5438 ( .A1(n6850), .A2(n4786), .ZN(n4785) );
  AOI21_X1 U5439 ( .B1(n5862), .B2(n7969), .A(n5861), .ZN(n6753) );
  AND2_X1 U5440 ( .A1(n4821), .A2(n4819), .ZN(n4817) );
  NAND2_X1 U5441 ( .A1(n4818), .A2(n4821), .ZN(n4816) );
  NAND2_X1 U5442 ( .A1(n6083), .A2(n6054), .ZN(n4818) );
  OR2_X1 U5443 ( .A1(n7297), .A2(n6230), .ZN(n5906) );
  INV_X1 U5444 ( .A(n4817), .ZN(n4811) );
  AND2_X1 U5445 ( .A1(n4816), .A2(n4814), .ZN(n4813) );
  INV_X1 U5446 ( .A(n7572), .ZN(n4814) );
  NAND2_X1 U5447 ( .A1(n5940), .A2(n5941), .ZN(n6807) );
  AND2_X1 U5448 ( .A1(n8537), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U5449 ( .A1(n4455), .A2(n4792), .ZN(n4791) );
  INV_X1 U5450 ( .A(n4794), .ZN(n4792) );
  INV_X1 U5451 ( .A(n4455), .ZN(n4793) );
  OR3_X1 U5452 ( .A1(n6195), .A2(n6194), .A3(n8539), .ZN(n6208) );
  NAND2_X1 U5453 ( .A1(n4526), .A2(n7021), .ZN(n8155) );
  INV_X1 U5454 ( .A(n8118), .ZN(n4526) );
  OAI21_X1 U5455 ( .B1(n8673), .B2(n4741), .A(n4433), .ZN(n7957) );
  INV_X1 U5456 ( .A(n8104), .ZN(n4741) );
  NAND2_X1 U5457 ( .A1(n8104), .A2(n4740), .ZN(n4739) );
  AND2_X1 U5458 ( .A1(n4614), .A2(n4613), .ZN(n8585) );
  NAND2_X1 U5459 ( .A1(n6735), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4613) );
  NOR2_X1 U5460 ( .A1(n7226), .A2(n4462), .ZN(n7230) );
  NAND2_X1 U5461 ( .A1(n7230), .A2(n7229), .ZN(n7398) );
  NAND2_X1 U5462 ( .A1(n7398), .A2(n4616), .ZN(n7400) );
  OR2_X1 U5463 ( .A1(n7399), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U5464 ( .A1(n7400), .A2(n7401), .ZN(n7595) );
  NOR2_X1 U5465 ( .A1(n8612), .A2(n4617), .ZN(n8630) );
  AND2_X1 U5466 ( .A1(n7902), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4617) );
  INV_X1 U5467 ( .A(n7905), .ZN(n7904) );
  AND2_X1 U5468 ( .A1(n8663), .A2(n8462), .ZN(n8647) );
  INV_X1 U5469 ( .A(n8668), .ZN(n8661) );
  OAI22_X1 U5470 ( .A1(n8679), .A2(n8685), .B1(n8843), .B2(n8550), .ZN(n8662)
         );
  NAND2_X1 U5471 ( .A1(n8695), .A2(n8715), .ZN(n8703) );
  OR2_X1 U5472 ( .A1(n8843), .A2(n8703), .ZN(n8680) );
  INV_X1 U5473 ( .A(n8685), .ZN(n8678) );
  NAND2_X1 U5474 ( .A1(n8087), .A2(n8089), .ZN(n8697) );
  AOI21_X1 U5475 ( .B1(n4759), .B2(n4762), .A(n4757), .ZN(n4756) );
  INV_X1 U5476 ( .A(n4759), .ZN(n4755) );
  INV_X1 U5477 ( .A(n8736), .ZN(n4757) );
  AND2_X1 U5478 ( .A1(n8085), .A2(n8082), .ZN(n8721) );
  AND2_X1 U5479 ( .A1(n8719), .A2(n8714), .ZN(n8715) );
  NOR2_X1 U5480 ( .A1(n8731), .A2(n8736), .ZN(n8730) );
  NAND2_X1 U5481 ( .A1(n8765), .A2(n7941), .ZN(n8770) );
  OR2_X1 U5482 ( .A1(n8780), .A2(n8779), .ZN(n8765) );
  AND4_X1 U5483 ( .A1(n6142), .A2(n6141), .A3(n6140), .A4(n6139), .ZN(n8799)
         );
  NOR2_X1 U5484 ( .A1(n8791), .A2(n8878), .ZN(n8790) );
  NAND2_X1 U5485 ( .A1(n4827), .A2(n4828), .ZN(n4825) );
  INV_X1 U5486 ( .A(n4827), .ZN(n4824) );
  AND2_X1 U5487 ( .A1(n7507), .A2(n4623), .ZN(n7808) );
  NOR2_X1 U5488 ( .A1(n8895), .A2(n4624), .ZN(n4623) );
  INV_X1 U5489 ( .A(n4625), .ZN(n4624) );
  NAND2_X1 U5490 ( .A1(n7713), .A2(n7712), .ZN(n7813) );
  NAND2_X1 U5491 ( .A1(n7684), .A2(n8048), .ZN(n7686) );
  NAND2_X1 U5492 ( .A1(n7507), .A2(n7506), .ZN(n7610) );
  NAND2_X1 U5493 ( .A1(n7507), .A2(n4627), .ZN(n7692) );
  NOR2_X1 U5494 ( .A1(n9742), .A2(n8037), .ZN(n7507) );
  AND4_X1 U5495 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n7642)
         );
  AND2_X1 U5496 ( .A1(n8031), .A2(n8033), .ZN(n9722) );
  OR2_X1 U5497 ( .A1(n9722), .A2(n9734), .ZN(n9736) );
  NAND2_X1 U5498 ( .A1(n4478), .A2(n4477), .ZN(n9734) );
  INV_X1 U5499 ( .A(n7459), .ZN(n4477) );
  OR2_X1 U5500 ( .A1(n7431), .A2(n7456), .ZN(n9741) );
  NAND2_X1 U5501 ( .A1(n8015), .A2(n8022), .ZN(n8130) );
  AND3_X1 U5502 ( .A1(n7322), .A2(n8814), .A3(n4398), .ZN(n7429) );
  NAND2_X1 U5503 ( .A1(n4748), .A2(n4746), .ZN(n7327) );
  AND2_X1 U5504 ( .A1(n4747), .A2(n8011), .ZN(n4746) );
  AND2_X1 U5505 ( .A1(n8016), .A2(n8023), .ZN(n7414) );
  NAND2_X1 U5506 ( .A1(n7318), .A2(n7317), .ZN(n9753) );
  OAI21_X1 U5507 ( .B1(n8810), .B2(n4752), .A(n4749), .ZN(n9760) );
  NAND2_X1 U5508 ( .A1(n8814), .A2(n4630), .ZN(n9754) );
  NAND2_X1 U5509 ( .A1(n8814), .A2(n9806), .ZN(n8813) );
  NAND2_X1 U5510 ( .A1(n4830), .A2(n4831), .ZN(n8821) );
  AOI21_X1 U5511 ( .B1(n4440), .B2(n9799), .A(n4832), .ZN(n4831) );
  AND4_X1 U5512 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), .ZN(n9764)
         );
  AND2_X1 U5513 ( .A1(n7355), .A2(n9799), .ZN(n8814) );
  NOR2_X1 U5514 ( .A1(n7354), .A2(n7358), .ZN(n7355) );
  NAND2_X1 U5515 ( .A1(n7303), .A2(n7972), .ZN(n7346) );
  OAI211_X1 U5516 ( .C1(n6575), .C2(n6681), .A(n5882), .B(n5881), .ZN(n6713)
         );
  OR2_X1 U5517 ( .A1(n7960), .A2(n9968), .ZN(n5881) );
  NOR2_X1 U5518 ( .A1(n7241), .A2(n7208), .ZN(n7279) );
  NAND2_X1 U5519 ( .A1(n6558), .A2(n6559), .ZN(n6710) );
  BUF_X1 U5520 ( .A(n5860), .Z(n6575) );
  NAND2_X1 U5521 ( .A1(n7950), .A2(n7949), .ZN(n8833) );
  NAND2_X1 U5522 ( .A1(n6221), .A2(n6220), .ZN(n8838) );
  AND2_X1 U5523 ( .A1(n6265), .A2(n6281), .ZN(n9824) );
  INV_X1 U5524 ( .A(n6713), .ZN(n7336) );
  INV_X1 U5525 ( .A(n7241), .ZN(n6708) );
  INV_X1 U5526 ( .A(n9824), .ZN(n9850) );
  NOR2_X1 U5527 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4765) );
  INV_X1 U5528 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4764) );
  INV_X1 U5529 ( .A(n4809), .ZN(n4806) );
  INV_X1 U5530 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5953) );
  OR2_X1 U5531 ( .A1(n5956), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U5532 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4615) );
  OAI21_X1 U5533 ( .B1(n6616), .B2(n4883), .A(n4881), .ZN(n6859) );
  AOI21_X1 U5534 ( .B1(n4882), .B2(n4884), .A(n4430), .ZN(n4881) );
  INV_X1 U5535 ( .A(n4884), .ZN(n4883) );
  OR2_X1 U5536 ( .A1(n4870), .A2(n4869), .ZN(n4868) );
  NAND2_X1 U5537 ( .A1(n4869), .A2(n4870), .ZN(n4867) );
  OAI21_X1 U5538 ( .B1(n8940), .B2(n4865), .A(n4859), .ZN(n8923) );
  NOR2_X1 U5539 ( .A1(n4861), .A2(n4860), .ZN(n4859) );
  NOR2_X1 U5540 ( .A1(n4865), .A2(n5595), .ZN(n4861) );
  INV_X1 U5541 ( .A(n4863), .ZN(n4860) );
  INV_X1 U5542 ( .A(n4513), .ZN(n4512) );
  NAND2_X1 U5543 ( .A1(n4493), .A2(n5016), .ZN(n6519) );
  NAND2_X1 U5544 ( .A1(n7586), .A2(n7587), .ZN(n4879) );
  OR2_X1 U5545 ( .A1(n7586), .A2(n7587), .ZN(n4880) );
  AND2_X1 U5546 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5131) );
  AND2_X1 U5547 ( .A1(n6685), .A2(n5092), .ZN(n4884) );
  AND2_X1 U5548 ( .A1(n4872), .A2(n4496), .ZN(n4495) );
  AND2_X1 U5549 ( .A1(n5260), .A2(n5232), .ZN(n4872) );
  NAND2_X1 U5550 ( .A1(n7785), .A2(n7787), .ZN(n7786) );
  NAND2_X1 U5551 ( .A1(n7786), .A2(n4885), .ZN(n8988) );
  NAND2_X1 U5552 ( .A1(n5399), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5430) );
  AOI21_X1 U5553 ( .B1(n4504), .B2(n4506), .A(n4460), .ZN(n4502) );
  NOR2_X1 U5554 ( .A1(n8437), .A2(n8436), .ZN(n4719) );
  AND4_X1 U5555 ( .A1(n5197), .A2(n5196), .A3(n5195), .A4(n5194), .ZN(n6943)
         );
  OR2_X1 U5556 ( .A1(n5104), .A2(n7083), .ZN(n5105) );
  OR2_X1 U5557 ( .A1(n6428), .A2(n6429), .ZN(n6431) );
  NAND2_X1 U5558 ( .A1(n9513), .A2(n6319), .ZN(n9510) );
  NAND2_X1 U5559 ( .A1(n9524), .A2(n4463), .ZN(n9525) );
  NAND2_X1 U5560 ( .A1(n9510), .A2(n4485), .ZN(n9528) );
  OR2_X1 U5561 ( .A1(n9516), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4485) );
  AND2_X1 U5562 ( .A1(n9525), .A2(n4565), .ZN(n6339) );
  INV_X1 U5563 ( .A(n9533), .ZN(n4565) );
  NAND2_X1 U5564 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U5565 ( .A1(n6694), .A2(n5288), .ZN(n4569) );
  AOI21_X1 U5566 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6700), .A(n6699), .ZN(
        n6703) );
  NAND2_X1 U5567 ( .A1(n4410), .A2(n9545), .ZN(n9544) );
  NOR2_X1 U5568 ( .A1(n9054), .A2(n9577), .ZN(n9590) );
  AOI21_X1 U5569 ( .B1(n9601), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9602), .ZN(
        n9614) );
  NAND2_X1 U5570 ( .A1(n8167), .A2(n8166), .ZN(n9073) );
  OR3_X1 U5571 ( .A1(n5781), .A2(n5780), .A3(n5779), .ZN(n9116) );
  AOI21_X1 U5572 ( .B1(n4677), .B2(n4680), .A(n4676), .ZN(n4675) );
  INV_X1 U5573 ( .A(n9105), .ZN(n4676) );
  NOR2_X1 U5574 ( .A1(n9106), .A2(n4408), .ZN(n4677) );
  NAND2_X1 U5575 ( .A1(n4679), .A2(n4680), .ZN(n4678) );
  INV_X1 U5576 ( .A(n9106), .ZN(n4679) );
  NOR2_X1 U5577 ( .A1(n4609), .A2(n9191), .ZN(n9140) );
  OR2_X1 U5578 ( .A1(n4391), .A2(n9306), .ZN(n4609) );
  AND2_X1 U5579 ( .A1(n8236), .A2(n9104), .ZN(n9155) );
  AND2_X1 U5580 ( .A1(n5707), .A2(n5687), .ZN(n9176) );
  OR2_X1 U5581 ( .A1(n5658), .A2(n5657), .ZN(n5686) );
  AND2_X1 U5582 ( .A1(n9334), .A2(n9083), .ZN(n9084) );
  OR2_X1 U5583 ( .A1(n4399), .A2(n9099), .ZN(n4689) );
  AND2_X1 U5584 ( .A1(n4411), .A2(n9098), .ZN(n4690) );
  NAND2_X1 U5585 ( .A1(n9248), .A2(n4607), .ZN(n9235) );
  INV_X1 U5586 ( .A(n5580), .ZN(n5578) );
  NAND2_X1 U5587 ( .A1(n4920), .A2(n4919), .ZN(n9229) );
  NAND2_X1 U5588 ( .A1(n4444), .A2(n4397), .ZN(n4919) );
  NAND2_X1 U5589 ( .A1(n5525), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5554) );
  AOI21_X1 U5590 ( .B1(n7750), .B2(n8362), .A(n8366), .ZN(n7764) );
  NAND2_X1 U5591 ( .A1(n7489), .A2(n4602), .ZN(n7759) );
  AND2_X1 U5592 ( .A1(n4404), .A2(n7794), .ZN(n4602) );
  NAND2_X1 U5593 ( .A1(n7489), .A2(n4404), .ZN(n7761) );
  AND2_X1 U5594 ( .A1(n7489), .A2(n4603), .ZN(n7654) );
  AND4_X1 U5595 ( .A1(n5459), .A2(n5458), .A3(n5457), .A4(n5456), .ZN(n7649)
         );
  NAND2_X1 U5596 ( .A1(n4651), .A2(n4649), .ZN(n7624) );
  NOR2_X1 U5597 ( .A1(n7488), .A2(n7521), .ZN(n7489) );
  INV_X1 U5598 ( .A(n4666), .ZN(n4665) );
  AOI21_X1 U5599 ( .B1(n8336), .B2(n4666), .A(n4664), .ZN(n4663) );
  NAND2_X1 U5600 ( .A1(n4668), .A2(n4666), .ZN(n7442) );
  NAND2_X1 U5601 ( .A1(n5346), .A2(n5345), .ZN(n9444) );
  NAND2_X1 U5602 ( .A1(n7052), .A2(n4595), .ZN(n7488) );
  AND2_X1 U5603 ( .A1(n4403), .A2(n4596), .ZN(n4595) );
  INV_X1 U5604 ( .A(n9444), .ZN(n4596) );
  NAND2_X1 U5605 ( .A1(n7052), .A2(n4403), .ZN(n7255) );
  AND2_X1 U5606 ( .A1(n4668), .A2(n4670), .ZN(n7248) );
  NAND2_X1 U5607 ( .A1(n7052), .A2(n4598), .ZN(n7140) );
  AND2_X1 U5608 ( .A1(n7052), .A2(n9687), .ZN(n7114) );
  AND2_X1 U5609 ( .A1(n7045), .A2(n8208), .ZN(n7134) );
  OR2_X1 U5610 ( .A1(n7061), .A2(n7029), .ZN(n7034) );
  AND4_X1 U5611 ( .A1(n5224), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n7046)
         );
  INV_X1 U5612 ( .A(n4660), .ZN(n4659) );
  OR2_X1 U5613 ( .A1(n6952), .A2(n8239), .ZN(n7024) );
  NAND2_X1 U5614 ( .A1(n6880), .A2(n6893), .ZN(n6944) );
  AND2_X1 U5615 ( .A1(n9272), .A2(n9663), .ZN(n9270) );
  AND2_X1 U5616 ( .A1(n5766), .A2(n7020), .ZN(n6988) );
  NAND2_X1 U5617 ( .A1(n6940), .A2(n6939), .ZN(n9282) );
  AND4_X1 U5618 ( .A1(n5166), .A2(n5165), .A3(n5164), .A4(n5163), .ZN(n9268)
         );
  NAND2_X1 U5619 ( .A1(n8306), .A2(n8307), .ZN(n9263) );
  AND2_X1 U5620 ( .A1(n8270), .A2(n8199), .ZN(n8240) );
  INV_X1 U5621 ( .A(n6988), .ZN(n6893) );
  XNOR2_X1 U5622 ( .A(n7699), .B(n7698), .ZN(n7875) );
  NAND2_X1 U5623 ( .A1(n6219), .A2(n6218), .ZN(n7699) );
  NAND2_X1 U5624 ( .A1(n5730), .A2(n5729), .ZN(n6219) );
  XNOR2_X1 U5625 ( .A(n5721), .B(n5720), .ZN(n7536) );
  XNOR2_X1 U5626 ( .A(n5604), .B(n5623), .ZN(n7215) );
  NAND2_X1 U5627 ( .A1(n5599), .A2(n5624), .ZN(n5604) );
  NAND2_X1 U5628 ( .A1(n4724), .A2(n5544), .ZN(n5574) );
  NAND2_X1 U5629 ( .A1(n5517), .A2(n4728), .ZN(n4724) );
  NAND2_X1 U5630 ( .A1(n4519), .A2(n4655), .ZN(n4987) );
  NOR2_X1 U5631 ( .A1(n4522), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4519) );
  NAND2_X1 U5632 ( .A1(n5304), .A2(n4953), .ZN(n4713) );
  OR2_X1 U5633 ( .A1(n5156), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5213) );
  XNOR2_X1 U5634 ( .A(n5022), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U5635 ( .A1(n4735), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U5636 ( .A1(n4736), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4735) );
  NOR2_X1 U5637 ( .A1(n8768), .A2(n6230), .ZN(n8491) );
  NAND2_X1 U5638 ( .A1(n5951), .A2(n5952), .ZN(n4804) );
  NAND2_X1 U5639 ( .A1(n5942), .A2(n4797), .ZN(n4803) );
  NAND2_X1 U5640 ( .A1(n6185), .A2(n6184), .ZN(n8854) );
  NAND2_X1 U5641 ( .A1(n4800), .A2(n6823), .ZN(n6809) );
  NAND2_X1 U5642 ( .A1(n4815), .A2(n4816), .ZN(n7573) );
  NAND2_X1 U5643 ( .A1(n4820), .A2(n4817), .ZN(n4815) );
  NAND2_X1 U5644 ( .A1(n6171), .A2(n6170), .ZN(n8858) );
  XNOR2_X1 U5645 ( .A(n6154), .B(n6148), .ZN(n8526) );
  AOI21_X1 U5646 ( .B1(n4781), .B2(n4783), .A(n5995), .ZN(n4779) );
  AND4_X1 U5647 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n7367)
         );
  AND4_X1 U5648 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n7464)
         );
  OAI211_X1 U5649 ( .C1(n7960), .C2(n9907), .A(n5870), .B(n5869), .ZN(n6765)
         );
  NAND2_X1 U5650 ( .A1(n6099), .A2(n6098), .ZN(n8888) );
  NAND2_X1 U5651 ( .A1(n8499), .A2(n4794), .ZN(n4789) );
  OAI21_X1 U5652 ( .B1(n8499), .B2(n4793), .A(n4790), .ZN(n8536) );
  INV_X1 U5653 ( .A(n8543), .ZN(n8515) );
  NAND2_X1 U5654 ( .A1(n6059), .A2(n6058), .ZN(n7677) );
  INV_X1 U5655 ( .A(n8549), .ZN(n8567) );
  AND2_X1 U5656 ( .A1(n8572), .A2(n6607), .ZN(n6732) );
  INV_X1 U5657 ( .A(n4614), .ZN(n6730) );
  NAND2_X1 U5658 ( .A1(n4619), .A2(n6612), .ZN(n6769) );
  AND2_X1 U5659 ( .A1(n6769), .A2(n4618), .ZN(n6773) );
  NAND2_X1 U5660 ( .A1(n6770), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4618) );
  AOI21_X1 U5661 ( .B1(n8162), .B2(n7962), .A(n7961), .ZN(n8651) );
  XNOR2_X1 U5662 ( .A(n8656), .B(n8825), .ZN(n8827) );
  NAND2_X1 U5663 ( .A1(n7952), .A2(n7951), .ZN(n8830) );
  NAND2_X1 U5664 ( .A1(n8699), .A2(n8089), .ZN(n8686) );
  INV_X1 U5665 ( .A(n8849), .ZN(n8695) );
  NAND2_X1 U5666 ( .A1(n4758), .A2(n4759), .ZN(n8735) );
  NAND2_X1 U5667 ( .A1(n8780), .A2(n4761), .ZN(n4758) );
  INV_X1 U5668 ( .A(n4837), .ZN(n8745) );
  AOI21_X1 U5669 ( .B1(n4845), .B2(n4842), .A(n4840), .ZN(n4837) );
  INV_X1 U5670 ( .A(n4635), .ZN(n4633) );
  NAND2_X1 U5671 ( .A1(n4845), .A2(n4844), .ZN(n8759) );
  NAND2_X1 U5672 ( .A1(n6116), .A2(n6115), .ZN(n8884) );
  INV_X1 U5673 ( .A(n8888), .ZN(n7847) );
  NAND2_X1 U5674 ( .A1(n7807), .A2(n4828), .ZN(n7849) );
  NAND2_X1 U5675 ( .A1(n7497), .A2(n7496), .ZN(n7498) );
  NAND2_X1 U5676 ( .A1(n7503), .A2(n4854), .ZN(n7607) );
  NAND2_X1 U5677 ( .A1(n6017), .A2(n6016), .ZN(n9732) );
  INV_X1 U5678 ( .A(n4478), .ZN(n7458) );
  NAND2_X1 U5679 ( .A1(n8809), .A2(n8001), .ZN(n7381) );
  NAND2_X1 U5680 ( .A1(n9803), .A2(n4850), .ZN(n7385) );
  AND2_X1 U5681 ( .A1(n9803), .A2(n7315), .ZN(n4946) );
  NAND2_X1 U5682 ( .A1(n7313), .A2(n4751), .ZN(n9803) );
  NAND2_X1 U5683 ( .A1(n7352), .A2(n7298), .ZN(n7312) );
  OR2_X1 U5684 ( .A1(n9749), .A2(n7206), .ZN(n9775) );
  INV_X1 U5685 ( .A(n9775), .ZN(n9731) );
  AND2_X1 U5686 ( .A1(n6391), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9785) );
  OR2_X1 U5687 ( .A1(n6233), .A2(n6238), .ZN(n5828) );
  INV_X1 U5688 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9907) );
  INV_X1 U5689 ( .A(n4889), .ZN(n4888) );
  OAI21_X1 U5690 ( .B1(n4890), .B2(n4892), .A(n4894), .ZN(n4889) );
  OAI21_X1 U5691 ( .B1(n7172), .B2(n4506), .A(n4504), .ZN(n7527) );
  NAND2_X1 U5692 ( .A1(n4862), .A2(n4523), .ZN(n8958) );
  AND2_X1 U5693 ( .A1(n4867), .A2(n4458), .ZN(n4523) );
  NAND2_X1 U5694 ( .A1(n4871), .A2(n4868), .ZN(n4862) );
  NAND2_X1 U5695 ( .A1(n6616), .A2(n6617), .ZN(n6615) );
  NAND2_X1 U5696 ( .A1(n6791), .A2(n5202), .ZN(n4497) );
  NOR2_X1 U5697 ( .A1(n8950), .A2(n8949), .ZN(n9000) );
  NAND2_X1 U5698 ( .A1(n5685), .A2(n5684), .ZN(n9317) );
  AND3_X1 U5699 ( .A1(n5484), .A2(n5483), .A3(n5482), .ZN(n8992) );
  NAND2_X1 U5700 ( .A1(n4878), .A2(n4879), .ZN(n7735) );
  NAND2_X1 U5701 ( .A1(n5453), .A2(n5452), .ZN(n7743) );
  AND3_X1 U5702 ( .A1(n5506), .A2(n5505), .A3(n5504), .ZN(n7800) );
  AOI21_X1 U5703 ( .B1(n8958), .B2(n8921), .A(n8957), .ZN(n8960) );
  AND2_X1 U5704 ( .A1(n6615), .A2(n5092), .ZN(n6686) );
  NAND2_X1 U5705 ( .A1(n6615), .A2(n4884), .ZN(n6684) );
  OAI21_X1 U5706 ( .B1(n6791), .B2(n4500), .A(n4412), .ZN(n4873) );
  NAND2_X1 U5707 ( .A1(n9439), .A2(n5362), .ZN(n7515) );
  NAND2_X1 U5708 ( .A1(n4871), .A2(n4870), .ZN(n8977) );
  NAND2_X1 U5709 ( .A1(n4866), .A2(n5618), .ZN(n8976) );
  INV_X1 U5710 ( .A(n4871), .ZN(n4866) );
  NAND2_X1 U5711 ( .A1(n4511), .A2(n5511), .ZN(n8990) );
  NAND2_X1 U5712 ( .A1(n7786), .A2(n5491), .ZN(n4511) );
  OR2_X1 U5713 ( .A1(n5791), .A2(n5772), .ZN(n9446) );
  INV_X1 U5714 ( .A(n8444), .ZN(n4716) );
  NAND2_X1 U5715 ( .A1(n5739), .A2(n5738), .ZN(n9157) );
  INV_X1 U5716 ( .A(n9233), .ZN(n9083) );
  AND4_X1 U5717 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n7177)
         );
  NAND4_X1 U5718 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n9024)
         );
  NAND2_X1 U5719 ( .A1(n5017), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5072) );
  OR2_X1 U5720 ( .A1(n8172), .A2(n6323), .ZN(n5040) );
  NAND2_X1 U5721 ( .A1(n4641), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4640) );
  OR2_X1 U5722 ( .A1(n8172), .A2(n5011), .ZN(n5000) );
  AND2_X1 U5723 ( .A1(n6408), .A2(n6330), .ZN(n6479) );
  NAND2_X1 U5724 ( .A1(n6475), .A2(n6315), .ZN(n6425) );
  AND2_X1 U5725 ( .A1(n4564), .A2(n4459), .ZN(n9532) );
  AOI21_X1 U5726 ( .B1(n6631), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6630), .ZN(
        n6634) );
  INV_X1 U5727 ( .A(n4570), .ZN(n6693) );
  AND2_X1 U5728 ( .A1(n4568), .A2(n4567), .ZN(n9029) );
  INV_X1 U5729 ( .A(n6695), .ZN(n4567) );
  INV_X1 U5730 ( .A(n4568), .ZN(n6696) );
  NOR2_X1 U5731 ( .A1(n9029), .A2(n4566), .ZN(n9540) );
  NOR2_X1 U5732 ( .A1(n9042), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4566) );
  AOI21_X1 U5733 ( .B1(n9032), .B2(n9033), .A(n9560), .ZN(n9566) );
  INV_X1 U5734 ( .A(n4574), .ZN(n9034) );
  NAND2_X1 U5735 ( .A1(n8164), .A2(n8163), .ZN(n9287) );
  NAND2_X1 U5736 ( .A1(n4687), .A2(n9113), .ZN(n9297) );
  OR2_X1 U5737 ( .A1(n9114), .A2(n9265), .ZN(n4687) );
  NAND2_X1 U5738 ( .A1(n4904), .A2(n9109), .ZN(n4901) );
  OAI21_X1 U5739 ( .B1(n4902), .B2(n9109), .A(n4898), .ZN(n4897) );
  NAND2_X1 U5740 ( .A1(n8176), .A2(n8175), .ZN(n9299) );
  INV_X1 U5741 ( .A(n9303), .ZN(n9136) );
  NAND2_X1 U5742 ( .A1(n4674), .A2(n4680), .ZN(n9146) );
  NAND2_X1 U5743 ( .A1(n9322), .A2(n4949), .ZN(n9167) );
  NAND2_X1 U5744 ( .A1(n9188), .A2(n9187), .ZN(n9322) );
  NAND2_X1 U5745 ( .A1(n5656), .A2(n5655), .ZN(n9324) );
  NAND2_X1 U5746 ( .A1(n5577), .A2(n5576), .ZN(n9341) );
  NAND2_X1 U5747 ( .A1(n4692), .A2(n4694), .ZN(n9230) );
  NAND2_X1 U5748 ( .A1(n4693), .A2(n9093), .ZN(n9243) );
  OR2_X1 U5749 ( .A1(n9095), .A2(n9094), .ZN(n4693) );
  NAND2_X1 U5750 ( .A1(n4922), .A2(n4923), .ZN(n9242) );
  NAND2_X1 U5751 ( .A1(n7795), .A2(n4926), .ZN(n4922) );
  NAND2_X1 U5752 ( .A1(n5524), .A2(n5523), .ZN(n9351) );
  NOR2_X1 U5753 ( .A1(n7795), .A2(n4927), .ZN(n9080) );
  NAND2_X1 U5754 ( .A1(n5501), .A2(n5500), .ZN(n9356) );
  AND2_X1 U5755 ( .A1(n4929), .A2(n4421), .ZN(n7650) );
  NAND2_X1 U5756 ( .A1(n7440), .A2(n4947), .ZN(n7629) );
  OAI21_X1 U5757 ( .B1(n7130), .B2(n4918), .A(n4916), .ZN(n7439) );
  NAND2_X1 U5758 ( .A1(n7130), .A2(n7129), .ZN(n7246) );
  NAND2_X1 U5759 ( .A1(n4937), .A2(n7030), .ZN(n7031) );
  NAND2_X1 U5760 ( .A1(n7028), .A2(n8239), .ZN(n4937) );
  AND2_X1 U5761 ( .A1(n4909), .A2(n4910), .ZN(n7059) );
  INV_X1 U5762 ( .A(n9645), .ZN(n7015) );
  XNOR2_X1 U5763 ( .A(n9291), .B(n9287), .ZN(n9289) );
  AOI211_X1 U5764 ( .C1(n9443), .C2(n9303), .A(n9302), .B(n9301), .ZN(n9304)
         );
  NOR2_X1 U5765 ( .A1(n4938), .A2(n5279), .ZN(n4652) );
  NAND2_X1 U5766 ( .A1(n6219), .A2(n5731), .ZN(n7583) );
  OR2_X1 U5767 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  NAND2_X1 U5768 ( .A1(n4973), .A2(n4972), .ZN(n7866) );
  OR2_X1 U5769 ( .A1(n5127), .A2(n5126), .ZN(n6372) );
  NOR2_X1 U5770 ( .A1(n5051), .A2(n4571), .ZN(n6470) );
  OAI21_X1 U5771 ( .B1(n4573), .B2(n5049), .A(n4572), .ZN(n4571) );
  NAND2_X1 U5772 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4573) );
  AOI21_X1 U5773 ( .B1(n4805), .B2(n4393), .A(n5942), .ZN(n6872) );
  OAI21_X1 U5774 ( .B1(n6848), .B2(n4783), .A(n4781), .ZN(n6963) );
  XNOR2_X1 U5775 ( .A(n7967), .B(n7966), .ZN(n4743) );
  AOI21_X1 U5776 ( .B1(n4524), .B2(n4745), .A(n4476), .ZN(n4742) );
  OAI211_X1 U5777 ( .C1(n7897), .C2(n7896), .A(n4517), .B(n7895), .ZN(P1_U3218) );
  NAND2_X1 U5778 ( .A1(n7897), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U5779 ( .A1(n4715), .A2(n4714), .ZN(P1_U3240) );
  INV_X1 U5780 ( .A(n8449), .ZN(n4714) );
  INV_X1 U5781 ( .A(n4564), .ZN(n9507) );
  OAI21_X1 U5782 ( .B1(n4579), .B2(n9275), .A(n4575), .ZN(n9066) );
  INV_X1 U5783 ( .A(n9064), .ZN(n4579) );
  NAND2_X1 U5784 ( .A1(n4577), .A2(n4576), .ZN(n4575) );
  OAI21_X1 U5785 ( .B1(n9289), .B2(n4601), .A(n4599), .ZN(P1_U3522) );
  NAND2_X1 U5786 ( .A1(n9696), .A2(n9366), .ZN(n4601) );
  INV_X1 U5787 ( .A(n4600), .ZN(n4599) );
  OAI21_X1 U5788 ( .B1(n4395), .B2(n9694), .A(n4465), .ZN(n4600) );
  NAND2_X1 U5789 ( .A1(n4682), .A2(n4466), .ZN(P1_U3520) );
  NAND2_X1 U5790 ( .A1(n9380), .A2(n9696), .ZN(n4682) );
  OR2_X1 U5791 ( .A1(n9312), .A2(n9317), .ZN(n4391) );
  NAND2_X1 U5792 ( .A1(n4829), .A2(n7708), .ZN(n4828) );
  AND2_X1 U5793 ( .A1(n8423), .A2(n8268), .ZN(n4392) );
  AND3_X1 U5794 ( .A1(n5083), .A2(n5082), .A3(n5081), .ZN(n6926) );
  INV_X1 U5795 ( .A(n4506), .ZN(n4505) );
  OR2_X1 U5796 ( .A1(n5386), .A2(n4507), .ZN(n4506) );
  INV_X1 U5797 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4969) );
  INV_X1 U5798 ( .A(n9144), .ZN(n9306) );
  OR2_X1 U5799 ( .A1(n8858), .A2(n8504), .ZN(n8079) );
  NOR2_X1 U5800 ( .A1(n6808), .A2(n5931), .ZN(n4393) );
  AND2_X1 U5801 ( .A1(n4675), .A2(n9107), .ZN(n4394) );
  AND2_X1 U5802 ( .A1(n9288), .A2(n9292), .ZN(n4395) );
  NAND2_X1 U5803 ( .A1(n8763), .A2(n8493), .ZN(n4396) );
  OR2_X1 U5804 ( .A1(n9346), .A2(n9081), .ZN(n4397) );
  AND2_X1 U5805 ( .A1(n4630), .A2(n4629), .ZN(n4398) );
  NAND2_X1 U5806 ( .A1(n9105), .A2(n8411), .ZN(n9106) );
  INV_X1 U5807 ( .A(n9106), .ZN(n9145) );
  NAND2_X1 U5808 ( .A1(n8078), .A2(n8076), .ZN(n8750) );
  INV_X1 U5809 ( .A(n8750), .ZN(n4839) );
  INV_X1 U5810 ( .A(n4777), .ZN(n4776) );
  NOR2_X1 U5811 ( .A1(n6133), .A2(n6132), .ZN(n4777) );
  AND2_X1 U5812 ( .A1(n6135), .A2(n6134), .ZN(n8778) );
  INV_X1 U5813 ( .A(n8778), .ZN(n8873) );
  AND2_X1 U5814 ( .A1(n4694), .A2(n4691), .ZN(n4399) );
  AND2_X1 U5815 ( .A1(n7044), .A2(n9018), .ZN(n4400) );
  AND2_X1 U5816 ( .A1(n6157), .A2(n6156), .ZN(n8748) );
  NOR2_X1 U5817 ( .A1(n7513), .A2(n7512), .ZN(n4401) );
  INV_X1 U5818 ( .A(n5845), .ZN(n5812) );
  AND3_X1 U5819 ( .A1(n4654), .A2(n4995), .A3(n4992), .ZN(n4402) );
  NAND2_X1 U5820 ( .A1(n4789), .A2(n4455), .ZN(n8534) );
  XNOR2_X1 U5821 ( .A(n4982), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5766) );
  AND2_X1 U5822 ( .A1(n4598), .A2(n4597), .ZN(n4403) );
  AND2_X1 U5823 ( .A1(n9479), .A2(n4603), .ZN(n4404) );
  NAND2_X1 U5824 ( .A1(n5397), .A2(n5396), .ZN(n7628) );
  OR2_X1 U5825 ( .A1(n8791), .A2(n4633), .ZN(n4405) );
  INV_X1 U5826 ( .A(n8895), .ZN(n4829) );
  NAND2_X1 U5827 ( .A1(n4873), .A2(n5232), .ZN(n6970) );
  AND2_X1 U5828 ( .A1(n7969), .A2(n7968), .ZN(n4406) );
  OR2_X1 U5829 ( .A1(n4406), .A2(n8161), .ZN(n4407) );
  AND2_X1 U5830 ( .A1(n8236), .A2(n9153), .ZN(n4408) );
  INV_X1 U5831 ( .A(n5897), .ZN(n7956) );
  INV_X2 U5832 ( .A(n5860), .ZN(n5921) );
  NAND3_X1 U5833 ( .A1(n4993), .A2(n4656), .A3(n4655), .ZN(n4409) );
  AND2_X1 U5834 ( .A1(n9044), .A2(n9043), .ZN(n4410) );
  INV_X1 U5835 ( .A(n5100), .ZN(n5374) );
  NOR2_X1 U5836 ( .A1(n4696), .A2(n9097), .ZN(n4411) );
  AND2_X1 U5837 ( .A1(n4498), .A2(n5229), .ZN(n4412) );
  NAND2_X1 U5838 ( .A1(n5834), .A2(n5826), .ZN(n4413) );
  NOR2_X1 U5839 ( .A1(n9191), .A2(n9317), .ZN(n4414) );
  INV_X1 U5840 ( .A(n9006), .ZN(n9185) );
  AOI21_X1 U5841 ( .B1(n9176), .B2(n6983), .A(n5691), .ZN(n9006) );
  OR2_X1 U5842 ( .A1(n4970), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4415) );
  INV_X1 U5843 ( .A(n9160), .ZN(n9312) );
  AND2_X1 U5844 ( .A1(n8418), .A2(n8415), .ZN(n9109) );
  INV_X1 U5845 ( .A(n9109), .ZN(n4900) );
  INV_X1 U5846 ( .A(n5491), .ZN(n4886) );
  AND4_X1 U5847 ( .A1(n8443), .A2(n8442), .A3(n8441), .A4(n8440), .ZN(n4416)
         );
  NAND2_X1 U5848 ( .A1(n5049), .A2(n4586), .ZN(n5050) );
  INV_X1 U5849 ( .A(n8238), .ZN(n4908) );
  AND4_X1 U5850 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n6816)
         );
  OR3_X1 U5851 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4417) );
  NOR2_X1 U5852 ( .A1(n9170), .A2(n9103), .ZN(n4418) );
  NAND2_X1 U5853 ( .A1(n9144), .A2(n9128), .ZN(n4419) );
  INV_X1 U5854 ( .A(n5618), .ZN(n4870) );
  AND2_X1 U5855 ( .A1(n8010), .A2(n8011), .ZN(n9750) );
  NAND2_X1 U5856 ( .A1(n5635), .A2(n5634), .ZN(n9331) );
  INV_X1 U5857 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6238) );
  OR2_X1 U5858 ( .A1(n6816), .A2(n9799), .ZN(n4420) );
  OR2_X1 U5859 ( .A1(n7628), .A2(n9015), .ZN(n4421) );
  AND2_X1 U5860 ( .A1(n9346), .A2(n9081), .ZN(n4422) );
  NAND2_X1 U5861 ( .A1(n8398), .A2(n9098), .ZN(n9231) );
  INV_X1 U5862 ( .A(n9231), .ZN(n4691) );
  NOR2_X1 U5863 ( .A1(n9078), .A2(n9247), .ZN(n4423) );
  INV_X1 U5864 ( .A(n4762), .ZN(n4761) );
  NAND2_X1 U5865 ( .A1(n7941), .A2(n8076), .ZN(n4762) );
  AND2_X1 U5866 ( .A1(n5734), .A2(n5733), .ZN(n9144) );
  AND2_X1 U5867 ( .A1(n9322), .A2(n4942), .ZN(n4424) );
  OR2_X1 U5868 ( .A1(n9303), .A2(n9092), .ZN(n9107) );
  AND2_X1 U5869 ( .A1(n6510), .A2(n6335), .ZN(n4425) );
  INV_X1 U5870 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4586) );
  INV_X1 U5871 ( .A(n4917), .ZN(n4916) );
  OAI21_X1 U5872 ( .B1(n7129), .B2(n4918), .A(n7247), .ZN(n4917) );
  AND2_X1 U5873 ( .A1(n4893), .A2(n5746), .ZN(n4426) );
  AND2_X1 U5874 ( .A1(n4692), .A2(n4399), .ZN(n4427) );
  NOR2_X1 U5875 ( .A1(n9810), .A2(n8564), .ZN(n4428) );
  NOR2_X1 U5876 ( .A1(n5154), .A2(n5153), .ZN(n4429) );
  AND2_X1 U5877 ( .A1(n5115), .A2(n5114), .ZN(n4430) );
  AND2_X1 U5878 ( .A1(n6145), .A2(n6144), .ZN(n4431) );
  OR2_X1 U5879 ( .A1(n6095), .A2(n6094), .ZN(n4432) );
  INV_X1 U5880 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5804) );
  AND2_X1 U5881 ( .A1(n8103), .A2(n4739), .ZN(n4433) );
  AND2_X1 U5882 ( .A1(n7628), .A2(n9015), .ZN(n4434) );
  INV_X1 U5883 ( .A(n4855), .ZN(n4854) );
  NAND2_X1 U5884 ( .A1(n7504), .A2(n7502), .ZN(n4855) );
  NOR2_X1 U5885 ( .A1(n8998), .A2(n8999), .ZN(n4435) );
  INV_X1 U5886 ( .A(n4935), .ZN(n4934) );
  NAND2_X1 U5887 ( .A1(n4936), .A2(n7030), .ZN(n4935) );
  INV_X1 U5888 ( .A(n4851), .ZN(n4850) );
  NAND2_X1 U5889 ( .A1(n7316), .A2(n7315), .ZN(n4851) );
  AND2_X1 U5890 ( .A1(n5331), .A2(SI_11_), .ZN(n4436) );
  AND2_X1 U5891 ( .A1(n9088), .A2(n9006), .ZN(n4437) );
  NAND2_X1 U5892 ( .A1(n4554), .A2(n4553), .ZN(n4438) );
  AND2_X1 U5893 ( .A1(n8208), .A2(n8329), .ZN(n8245) );
  INV_X1 U5894 ( .A(n8245), .ZN(n4936) );
  INV_X1 U5895 ( .A(n4887), .ZN(n4895) );
  INV_X1 U5896 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7842) );
  NOR2_X1 U5897 ( .A1(n5332), .A2(n4712), .ZN(n4711) );
  INV_X1 U5898 ( .A(n4875), .ZN(n4874) );
  NAND2_X1 U5899 ( .A1(n5359), .A2(n5328), .ZN(n4875) );
  INV_X1 U5900 ( .A(n4843), .ZN(n4842) );
  NAND2_X1 U5901 ( .A1(n4396), .A2(n4844), .ZN(n4843) );
  NOR2_X1 U5902 ( .A1(n9136), .A2(n9092), .ZN(n4439) );
  NOR2_X1 U5903 ( .A1(n8080), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5904 ( .A1(n7298), .A2(n8566), .ZN(n4440) );
  INV_X1 U5905 ( .A(n4904), .ZN(n4903) );
  AND2_X1 U5906 ( .A1(n9123), .A2(n4419), .ZN(n4904) );
  NOR2_X1 U5907 ( .A1(n9191), .A2(n4391), .ZN(n4441) );
  AND2_X1 U5908 ( .A1(n8685), .A2(n8089), .ZN(n4442) );
  NOR2_X1 U5909 ( .A1(n8712), .A2(n4545), .ZN(n4443) );
  AND2_X1 U5910 ( .A1(n5837), .A2(n4413), .ZN(n7966) );
  INV_X1 U5911 ( .A(n7966), .ZN(n8707) );
  OR2_X1 U5912 ( .A1(n4921), .A2(n4422), .ZN(n4444) );
  NAND2_X1 U5913 ( .A1(n8749), .A2(n8073), .ZN(n8766) );
  AND2_X1 U5914 ( .A1(n4902), .A2(n4900), .ZN(n4445) );
  AND3_X1 U5915 ( .A1(n8265), .A2(n8266), .A3(n9109), .ZN(n4446) );
  AND2_X1 U5916 ( .A1(n8125), .A2(n4420), .ZN(n4447) );
  AND2_X1 U5917 ( .A1(n4711), .A2(n5273), .ZN(n4448) );
  NOR2_X1 U5918 ( .A1(n5746), .A2(n5747), .ZN(n4449) );
  INV_X1 U5919 ( .A(n9215), .ZN(n9334) );
  AND2_X1 U5920 ( .A1(n5606), .A2(n5605), .ZN(n9215) );
  AND2_X1 U5921 ( .A1(n7848), .A2(n4826), .ZN(n4450) );
  AND2_X1 U5922 ( .A1(n7685), .A2(n8048), .ZN(n4451) );
  AND2_X1 U5923 ( .A1(n8071), .A2(n8067), .ZN(n4452) );
  AND2_X1 U5924 ( .A1(n6950), .A2(n4657), .ZN(n4453) );
  AND2_X1 U5925 ( .A1(n4397), .A2(n4926), .ZN(n4454) );
  INV_X1 U5926 ( .A(n4943), .ZN(n4942) );
  NAND2_X1 U5927 ( .A1(n4944), .A2(n4949), .ZN(n4943) );
  INV_X1 U5928 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4590) );
  INV_X1 U5929 ( .A(n8041), .ZN(n4853) );
  NAND2_X1 U5930 ( .A1(n9753), .A2(n7319), .ZN(n7454) );
  OR2_X1 U5931 ( .A1(n6191), .A2(n8500), .ZN(n4455) );
  AND2_X1 U5932 ( .A1(n8988), .A2(n8987), .ZN(n4456) );
  INV_X1 U5933 ( .A(n7483), .ZN(n4647) );
  NAND2_X1 U5934 ( .A1(n7489), .A2(n9484), .ZN(n4457) );
  INV_X1 U5935 ( .A(n8239), .ZN(n4933) );
  XOR2_X1 U5936 ( .A(n5647), .B(n6944), .Z(n4458) );
  OR2_X1 U5937 ( .A1(n9516), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4459) );
  AND2_X1 U5938 ( .A1(n7525), .A2(n5410), .ZN(n4460) );
  NAND2_X1 U5939 ( .A1(n7172), .A2(n4874), .ZN(n9439) );
  AND2_X1 U5940 ( .A1(n4820), .A2(n4819), .ZN(n4461) );
  AND2_X1 U5941 ( .A1(n7227), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4462) );
  AND2_X1 U5942 ( .A1(n8334), .A2(n8208), .ZN(n4669) );
  NAND2_X1 U5943 ( .A1(n5242), .A2(n5241), .ZN(n7103) );
  NAND2_X1 U5944 ( .A1(n7507), .A2(n4625), .ZN(n4628) );
  NAND2_X1 U5945 ( .A1(n9248), .A2(n4606), .ZN(n4608) );
  NAND2_X1 U5946 ( .A1(n5426), .A2(n5425), .ZN(n9365) );
  NOR2_X1 U5947 ( .A1(n6096), .A2(n4807), .ZN(n6233) );
  INV_X1 U5948 ( .A(SI_0_), .ZN(n4491) );
  OR2_X1 U5949 ( .A1(n6377), .A2(n5217), .ZN(n4463) );
  INV_X1 U5950 ( .A(n4632), .ZN(n8760) );
  NOR2_X1 U5951 ( .A1(n8791), .A2(n4634), .ZN(n4632) );
  INV_X1 U5952 ( .A(n8341), .ZN(n4667) );
  AND2_X1 U5953 ( .A1(n8587), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4464) );
  INV_X1 U5954 ( .A(n7794), .ZN(n9359) );
  AND2_X1 U5955 ( .A1(n5477), .A2(n5476), .ZN(n7794) );
  AND2_X1 U5956 ( .A1(n7207), .A2(n8817), .ZN(n9773) );
  NAND2_X1 U5957 ( .A1(n4846), .A2(n4766), .ZN(n6240) );
  INV_X1 U5958 ( .A(n4703), .ZN(n4702) );
  OAI21_X1 U5959 ( .B1(n4704), .B2(n6218), .A(n7703), .ZN(n4703) );
  OR2_X1 U5960 ( .A1(n9696), .A2(n6417), .ZN(n4465) );
  XNOR2_X1 U5961 ( .A(n5828), .B(n5827), .ZN(n6552) );
  OR2_X1 U5962 ( .A1(n9696), .A2(n10107), .ZN(n4466) );
  NAND2_X1 U5963 ( .A1(n4497), .A2(n5205), .ZN(n6833) );
  NAND2_X1 U5964 ( .A1(n6071), .A2(n6070), .ZN(n8899) );
  INV_X1 U5965 ( .A(n8899), .ZN(n4626) );
  NOR2_X1 U5966 ( .A1(n7439), .A2(n8251), .ZN(n4467) );
  AND2_X1 U5967 ( .A1(n7503), .A2(n7502), .ZN(n4468) );
  NAND2_X1 U5968 ( .A1(n8814), .A2(n4398), .ZN(n4631) );
  AND2_X1 U5969 ( .A1(n4651), .A2(n8210), .ZN(n4469) );
  AND2_X1 U5970 ( .A1(n4937), .A2(n4934), .ZN(n4470) );
  OR2_X1 U5971 ( .A1(n8583), .A2(n4464), .ZN(n4619) );
  AND2_X1 U5972 ( .A1(n9049), .A2(n5398), .ZN(n4471) );
  INV_X1 U5973 ( .A(n4951), .ZN(n4910) );
  AND2_X1 U5974 ( .A1(n4846), .A2(n4847), .ZN(n4472) );
  OR2_X1 U5975 ( .A1(n6552), .A2(n8707), .ZN(n6550) );
  INV_X1 U5976 ( .A(n9770), .ZN(n4629) );
  NAND2_X1 U5977 ( .A1(n5310), .A2(n5309), .ZN(n7249) );
  INV_X1 U5978 ( .A(n7249), .ZN(n4597) );
  INV_X1 U5979 ( .A(n9499), .ZN(n4487) );
  OR3_X1 U5980 ( .A1(n8158), .A2(n9763), .A3(n8157), .ZN(n4473) );
  INV_X1 U5981 ( .A(n6823), .ZN(n4799) );
  AND2_X1 U5982 ( .A1(n7915), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4474) );
  NOR2_X1 U5983 ( .A1(n6349), .A2(n6350), .ZN(n4475) );
  AND2_X1 U5984 ( .A1(n4473), .A2(n4744), .ZN(n4476) );
  INV_X1 U5985 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4492) );
  INV_X1 U5986 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9938) );
  INV_X1 U5987 ( .A(n8161), .ZN(n4745) );
  INV_X1 U5988 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4733) );
  OR2_X1 U5989 ( .A1(n6282), .A2(n6281), .ZN(n8541) );
  OR2_X1 U5990 ( .A1(n5443), .A2(n5442), .ZN(n5445) );
  NAND2_X1 U5991 ( .A1(n5470), .A2(n5469), .ZN(n5492) );
  NAND2_X1 U5992 ( .A1(n5390), .A2(n5389), .ZN(n5419) );
  NAND2_X1 U5993 ( .A1(n4723), .A2(n4721), .ZN(n5622) );
  NAND2_X1 U5994 ( .A1(n5654), .A2(n5653), .ZN(n5675) );
  NOR2_X4 U5995 ( .A1(n7707), .A2(n7706), .ZN(n7709) );
  OAI21_X2 U5996 ( .B1(n7462), .B2(n4855), .A(n4852), .ZN(n7679) );
  NAND2_X1 U5997 ( .A1(n4713), .A2(n5305), .ZN(n5333) );
  OAI21_X1 U5998 ( .B1(n8455), .B2(n8800), .A(n8454), .ZN(n8789) );
  MUX2_X2 U5999 ( .A(n8306), .B(n8305), .S(n8424), .Z(n8314) );
  NAND2_X1 U6000 ( .A1(n4479), .A2(n8412), .ZN(n8413) );
  NAND3_X1 U6001 ( .A1(n8409), .A2(n8410), .A3(n9145), .ZN(n4479) );
  NAND2_X1 U6002 ( .A1(n4480), .A2(n8386), .ZN(n8388) );
  NAND2_X1 U6003 ( .A1(n8396), .A2(n4481), .ZN(n4480) );
  NAND2_X2 U6004 ( .A1(n6990), .A2(n8270), .ZN(n8304) );
  MUX2_X2 U6005 ( .A(n8339), .B(n8338), .S(n8424), .Z(n8350) );
  OAI21_X1 U6006 ( .B1(n8350), .B2(n8349), .A(n8348), .ZN(n8360) );
  NAND2_X1 U6007 ( .A1(n4717), .A2(n4716), .ZN(n4715) );
  NAND2_X1 U6008 ( .A1(n4705), .A2(n5187), .ZN(n5208) );
  NAND2_X1 U6009 ( .A1(n8453), .A2(n8452), .ZN(n8454) );
  NAND2_X1 U6010 ( .A1(n5144), .A2(n4489), .ZN(n5150) );
  NAND2_X2 U6011 ( .A1(n4734), .A2(n4732), .ZN(n7833) );
  NAND2_X1 U6012 ( .A1(n5185), .A2(n5184), .ZN(n4705) );
  OAI22_X1 U6013 ( .A1(n7709), .A2(n4825), .B1(n4450), .B2(n4824), .ZN(n8453)
         );
  AOI21_X1 U6014 ( .B1(n7679), .B2(n8137), .A(n7678), .ZN(n7681) );
  OAI21_X1 U6015 ( .B1(n6454), .B2(n6455), .A(n4493), .ZN(n6539) );
  NAND2_X1 U6016 ( .A1(n6455), .A2(n6454), .ZN(n4493) );
  NAND2_X1 U6017 ( .A1(n6791), .A2(n4412), .ZN(n4494) );
  NAND2_X1 U6018 ( .A1(n4495), .A2(n4494), .ZN(n6971) );
  AND2_X2 U6019 ( .A1(n6304), .A2(n6988), .ZN(n5167) );
  NAND2_X1 U6020 ( .A1(n7172), .A2(n4504), .ZN(n4503) );
  NAND2_X1 U6021 ( .A1(n4503), .A2(n4502), .ZN(n5413) );
  NAND2_X1 U6022 ( .A1(n4508), .A2(n4512), .ZN(n5543) );
  NAND2_X1 U6023 ( .A1(n7785), .A2(n4509), .ZN(n4508) );
  NAND3_X1 U6024 ( .A1(n4655), .A2(n4521), .A3(n4520), .ZN(n5768) );
  NAND2_X1 U6025 ( .A1(n8064), .A2(n4530), .ZN(n4527) );
  NAND2_X1 U6026 ( .A1(n4527), .A2(n4528), .ZN(n8061) );
  NAND2_X1 U6027 ( .A1(n8042), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U6028 ( .A1(n4548), .A2(n4551), .ZN(n8054) );
  NAND3_X1 U6029 ( .A1(n7966), .A2(n6552), .A3(n8152), .ZN(n8112) );
  NOR2_X1 U6030 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4556) );
  NOR2_X2 U6031 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5867) );
  INV_X1 U6032 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4587) );
  INV_X1 U6033 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4585) );
  INV_X1 U6034 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10058) );
  INV_X1 U6035 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4582) );
  INV_X1 U6036 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4581) );
  INV_X1 U6037 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4588) );
  OAI21_X1 U6038 ( .B1(n9289), .B2(n9688), .A(n4395), .ZN(n9378) );
  NAND2_X1 U6039 ( .A1(n9115), .A2(n9294), .ZN(n9291) );
  INV_X1 U6040 ( .A(n4608), .ZN(n9212) );
  MUX2_X1 U6041 ( .A(n6597), .B(P2_REG2_REG_1__SCAN_IN), .S(n6598), .Z(n9399)
         );
  INV_X1 U6042 ( .A(n4628), .ZN(n7717) );
  INV_X1 U6043 ( .A(n4631), .ZN(n9755) );
  INV_X1 U6044 ( .A(n4636), .ZN(n8746) );
  NAND2_X2 U6045 ( .A1(n4638), .A2(n4998), .ZN(n5783) );
  NAND3_X1 U6046 ( .A1(n4638), .A2(n4998), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n4642) );
  OR2_X4 U6047 ( .A1(n4998), .A2(n4997), .ZN(n8172) );
  NAND2_X2 U6048 ( .A1(n4640), .A2(n4639), .ZN(n9027) );
  AND3_X1 U6049 ( .A1(n4642), .A2(n5020), .A3(n5021), .ZN(n4639) );
  INV_X1 U6050 ( .A(n4998), .ZN(n7827) );
  NAND2_X1 U6051 ( .A1(n4643), .A2(n6947), .ZN(n4644) );
  NAND2_X1 U6052 ( .A1(n8197), .A2(n8241), .ZN(n7005) );
  OAI21_X1 U6053 ( .B1(n7482), .B2(n4648), .A(n4645), .ZN(n7647) );
  INV_X1 U6054 ( .A(n4938), .ZN(n4656) );
  NAND2_X1 U6055 ( .A1(n4402), .A2(n4652), .ZN(n7841) );
  NAND3_X1 U6056 ( .A1(n4655), .A2(n4992), .A3(n4654), .ZN(n4653) );
  OAI21_X1 U6057 ( .B1(n8304), .B2(n4659), .A(n4453), .ZN(n6952) );
  OR2_X2 U6058 ( .A1(n8304), .A2(n6949), .ZN(n8306) );
  OAI21_X1 U6059 ( .B1(n7045), .B2(n4665), .A(n4663), .ZN(n7443) );
  INV_X1 U6060 ( .A(n8326), .ZN(n4670) );
  NAND2_X1 U6061 ( .A1(n4671), .A2(n4672), .ZN(n9110) );
  NAND2_X1 U6062 ( .A1(n9170), .A2(n4394), .ZN(n4671) );
  NAND2_X1 U6063 ( .A1(n9170), .A2(n4408), .ZN(n4674) );
  NAND2_X1 U6064 ( .A1(n9095), .A2(n4690), .ZN(n4688) );
  NAND2_X1 U6065 ( .A1(n4688), .A2(n4689), .ZN(n9216) );
  INV_X1 U6066 ( .A(n4697), .ZN(n7831) );
  AOI21_X2 U6067 ( .B1(n5150), .B2(n5149), .A(n4429), .ZN(n5185) );
  NAND2_X1 U6068 ( .A1(n5274), .A2(n4448), .ZN(n4708) );
  NAND2_X1 U6069 ( .A1(n4708), .A2(n4709), .ZN(n5364) );
  NAND2_X1 U6070 ( .A1(n5517), .A2(n4725), .ZN(n4723) );
  AOI21_X1 U6071 ( .B1(n4392), .B2(n4737), .A(n5766), .ZN(n8432) );
  INV_X1 U6072 ( .A(n9287), .ZN(n4738) );
  NAND2_X1 U6073 ( .A1(n5445), .A2(n5444), .ZN(n5468) );
  OAI21_X2 U6074 ( .B1(n5419), .B2(n5418), .A(n5417), .ZN(n5443) );
  NAND2_X1 U6075 ( .A1(n5723), .A2(n5722), .ZN(n5730) );
  NAND3_X2 U6076 ( .A1(n5026), .A2(n5025), .A3(n5024), .ZN(n6932) );
  AOI21_X1 U6077 ( .B1(n9216), .B2(n9101), .A(n9100), .ZN(n9200) );
  NOR2_X1 U6078 ( .A1(n9183), .A2(n9102), .ZN(n9170) );
  NAND2_X1 U6079 ( .A1(n5141), .A2(n5151), .ZN(n5145) );
  NAND2_X1 U6080 ( .A1(n4390), .A2(n5003), .ZN(n5023) );
  NAND2_X1 U6081 ( .A1(n8667), .A2(n8661), .ZN(n8673) );
  NAND2_X1 U6082 ( .A1(n8673), .A2(n8094), .ZN(n8464) );
  OAI21_X1 U6083 ( .B1(n4743), .B2(n4407), .A(n4742), .ZN(P2_U3244) );
  INV_X1 U6084 ( .A(n8820), .ZN(n4751) );
  NAND3_X1 U6085 ( .A1(n9750), .A2(n4749), .A3(n4752), .ZN(n4747) );
  NAND3_X1 U6086 ( .A1(n8810), .A2(n4749), .A3(n9750), .ZN(n4748) );
  INV_X1 U6087 ( .A(n7282), .ZN(n8122) );
  INV_X1 U6088 ( .A(n6718), .ZN(n8570) );
  OAI21_X2 U6089 ( .B1(n8780), .B2(n4755), .A(n4756), .ZN(n8723) );
  NAND2_X1 U6090 ( .A1(n7941), .A2(n8779), .ZN(n4763) );
  AND3_X1 U6091 ( .A1(n4766), .A2(n4846), .A3(n4764), .ZN(n5844) );
  NAND2_X1 U6092 ( .A1(n7684), .A2(n4451), .ZN(n7713) );
  NAND2_X1 U6093 ( .A1(n8699), .A2(n4442), .ZN(n7947) );
  NAND2_X1 U6094 ( .A1(n7497), .A2(n4767), .ZN(n7608) );
  NAND2_X1 U6095 ( .A1(n7303), .A2(n4768), .ZN(n7324) );
  NAND2_X1 U6096 ( .A1(n6717), .A2(n7981), .ZN(n7303) );
  NAND4_X1 U6097 ( .A1(n4771), .A2(n5910), .A3(n4769), .A4(n4770), .ZN(n6066)
         );
  OAI21_X2 U6098 ( .B1(n7770), .B2(n4773), .A(n4772), .ZN(n6154) );
  OAI21_X1 U6099 ( .B1(n7770), .B2(n7769), .A(n4776), .ZN(n7777) );
  NAND2_X1 U6100 ( .A1(n6848), .A2(n4781), .ZN(n4778) );
  NAND2_X1 U6101 ( .A1(n4778), .A2(n4779), .ZN(n7123) );
  NAND2_X1 U6102 ( .A1(n8499), .A2(n4790), .ZN(n4787) );
  NAND2_X1 U6103 ( .A1(n4787), .A2(n4788), .ZN(n8482) );
  NAND3_X1 U6104 ( .A1(n4796), .A2(n4803), .A3(n4804), .ZN(n6801) );
  NAND3_X1 U6105 ( .A1(n4800), .A2(n4798), .A3(n4393), .ZN(n4796) );
  OR3_X1 U6106 ( .A1(n6096), .A2(n4806), .A3(P2_IR_REG_18__SCAN_IN), .ZN(n5829) );
  OAI211_X2 U6107 ( .C1(n4812), .C2(n4820), .A(n4432), .B(n4810), .ZN(n7618)
         );
  INV_X1 U6108 ( .A(n4813), .ZN(n4812) );
  NOR2_X1 U6109 ( .A1(n4461), .A2(n6055), .ZN(n7663) );
  INV_X1 U6110 ( .A(n7475), .ZN(n4820) );
  INV_X1 U6111 ( .A(n4823), .ZN(n4822) );
  XNOR2_X1 U6112 ( .A(n5871), .B(n7241), .ZN(n5852) );
  NAND2_X1 U6113 ( .A1(n7353), .A2(n4447), .ZN(n4830) );
  NAND2_X1 U6114 ( .A1(n9753), .A2(n4833), .ZN(n9737) );
  AND2_X1 U6115 ( .A1(n8940), .A2(n5595), .ZN(n4871) );
  NAND2_X1 U6116 ( .A1(n7589), .A2(n4880), .ZN(n4878) );
  INV_X1 U6117 ( .A(n6617), .ZN(n4882) );
  AOI21_X1 U6118 ( .B1(n8960), .B2(n4892), .A(n4890), .ZN(n4887) );
  NOR2_X1 U6119 ( .A1(n8960), .A2(n5674), .ZN(n8950) );
  OAI21_X1 U6120 ( .B1(n8960), .B2(n4890), .A(n4888), .ZN(n4893) );
  NAND2_X1 U6121 ( .A1(n9139), .A2(n9106), .ZN(n4905) );
  OAI211_X1 U6122 ( .C1(n9139), .C2(n4901), .A(n4897), .B(n4896), .ZN(n9296)
         );
  NAND2_X1 U6123 ( .A1(n9139), .A2(n4445), .ZN(n4896) );
  NAND2_X1 U6124 ( .A1(n6940), .A2(n4906), .ZN(n4909) );
  NAND2_X1 U6125 ( .A1(n7130), .A2(n4915), .ZN(n4911) );
  NAND2_X1 U6126 ( .A1(n4911), .A2(n4912), .ZN(n7484) );
  NAND2_X1 U6127 ( .A1(n7795), .A2(n4454), .ZN(n4920) );
  NAND2_X1 U6128 ( .A1(n4929), .A2(n4928), .ZN(n7632) );
  AND2_X1 U6129 ( .A1(n7630), .A2(n4421), .ZN(n4928) );
  NAND3_X1 U6130 ( .A1(n4939), .A2(n4963), .A3(n4590), .ZN(n4938) );
  OAI21_X1 U6131 ( .B1(n9188), .B2(n4943), .A(n4940), .ZN(n9152) );
  AND2_X2 U6132 ( .A1(n4997), .A2(n4998), .ZN(n5017) );
  XNOR2_X2 U6133 ( .A(n4945), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4998) );
  OAI222_X1 U6134 ( .A1(n9725), .A2(n8470), .B1(n8483), .B2(n9763), .C1(n7964), 
        .C2(n8469), .ZN(n8471) );
  NOR2_X1 U6135 ( .A1(n7286), .A2(n5838), .ZN(n5853) );
  NAND2_X1 U6136 ( .A1(n6710), .A2(n6709), .ZN(n7278) );
  INV_X1 U6137 ( .A(n7286), .ZN(n6557) );
  NAND2_X1 U6138 ( .A1(n7962), .A2(n5847), .ZN(n5848) );
  NAND2_X1 U6139 ( .A1(n9152), .A2(n4958), .ZN(n9091) );
  OR2_X1 U6140 ( .A1(n9082), .A2(n9246), .ZN(n4948) );
  OR2_X1 U6141 ( .A1(n9192), .A2(n9202), .ZN(n4949) );
  NAND2_X1 U6142 ( .A1(n5147), .A2(n5146), .ZN(n4950) );
  AND2_X1 U6143 ( .A1(n9022), .A2(n9279), .ZN(n4951) );
  OR2_X1 U6144 ( .A1(n7655), .A2(n7631), .ZN(n4952) );
  INV_X1 U6145 ( .A(n9317), .ZN(n9088) );
  NOR2_X1 U6146 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4954) );
  OR2_X1 U6147 ( .A1(n8422), .A2(n8424), .ZN(n4955) );
  INV_X1 U6148 ( .A(n7628), .ZN(n9484) );
  NOR2_X1 U6149 ( .A1(n9733), .A2(n9722), .ZN(n4957) );
  OR2_X1 U6150 ( .A1(n9160), .A2(n9089), .ZN(n4958) );
  OR2_X1 U6151 ( .A1(n8778), .A2(n8799), .ZN(n4959) );
  NAND2_X1 U6152 ( .A1(n8923), .A2(n8922), .ZN(n8921) );
  INV_X1 U6153 ( .A(n8138), .ZN(n7685) );
  INV_X1 U6154 ( .A(n9281), .ZN(n6941) );
  AND2_X1 U6155 ( .A1(n9633), .A2(n6901), .ZN(n4960) );
  INV_X1 U6156 ( .A(n8429), .ZN(n8425) );
  OR2_X1 U6157 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  MUX2_X1 U6158 ( .A(n8418), .B(n8417), .S(n8424), .Z(n8419) );
  NAND2_X1 U6159 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  INV_X1 U6160 ( .A(n9750), .ZN(n7317) );
  INV_X1 U6161 ( .A(n7283), .ZN(n6716) );
  INV_X1 U6162 ( .A(n6973), .ZN(n5260) );
  INV_X1 U6163 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5160) );
  INV_X1 U6164 ( .A(n5638), .ZN(n5636) );
  INV_X1 U6165 ( .A(n5400), .ZN(n5399) );
  INV_X1 U6166 ( .A(n5527), .ZN(n5525) );
  INV_X1 U6167 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5218) );
  INV_X2 U6168 ( .A(n7826), .ZN(n5497) );
  INV_X1 U6169 ( .A(n5268), .ZN(n5271) );
  INV_X1 U6170 ( .A(n5206), .ZN(n5207) );
  AND2_X1 U6171 ( .A1(n6760), .A2(n6759), .ZN(n5874) );
  INV_X1 U6172 ( .A(n6153), .ZN(n6148) );
  AND2_X1 U6173 ( .A1(n6045), .A2(n6044), .ZN(n6060) );
  NAND2_X1 U6174 ( .A1(n6716), .A2(n8122), .ZN(n7285) );
  AND2_X1 U6175 ( .A1(n5286), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5312) );
  INV_X1 U6176 ( .A(n9442), .ZN(n5359) );
  AND2_X1 U6177 ( .A1(n5616), .A2(n5615), .ZN(n5618) );
  OR2_X1 U6178 ( .A1(n5686), .A2(n8951), .ZN(n5707) );
  NAND2_X1 U6179 ( .A1(n5636), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5658) );
  OR2_X1 U6180 ( .A1(n5376), .A2(n5375), .ZN(n5400) );
  NAND2_X1 U6181 ( .A1(n7583), .A2(n5306), .ZN(n5734) );
  NAND2_X1 U6182 ( .A1(n5578), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5608) );
  NOR2_X1 U6183 ( .A1(n5245), .A2(n5244), .ZN(n5286) );
  NAND2_X1 U6184 ( .A1(n5131), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5161) );
  INV_X1 U6185 ( .A(n5414), .ZN(n5418) );
  NAND2_X1 U6186 ( .A1(n5337), .A2(n5336), .ZN(n5365) );
  AOI21_X1 U6187 ( .B1(n5272), .B2(n5271), .A(n5270), .ZN(n5273) );
  INV_X1 U6188 ( .A(n6275), .ZN(n6276) );
  NAND2_X1 U6189 ( .A1(n6008), .A2(n6009), .ZN(n6010) );
  AND3_X1 U6190 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5925) );
  AND2_X1 U6191 ( .A1(n6350), .A2(n5890), .ZN(n5891) );
  OR3_X1 U6192 ( .A1(n5998), .A2(n5997), .A3(n5996), .ZN(n6018) );
  INV_X1 U6193 ( .A(n6807), .ZN(n6815) );
  INV_X1 U6194 ( .A(n8838), .ZN(n8666) );
  INV_X1 U6195 ( .A(n8868), .ZN(n8763) );
  NOR2_X1 U6196 ( .A1(n6018), .A2(n7188), .ZN(n6045) );
  NAND2_X1 U6197 ( .A1(n7278), .A2(n7282), .ZN(n7277) );
  MUX2_X1 U6198 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5841), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5842) );
  NAND2_X1 U6199 ( .A1(n5705), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U6200 ( .A1(n5312), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5348) );
  AND2_X1 U6201 ( .A1(n5695), .A2(n5694), .ZN(n8999) );
  OR2_X1 U6202 ( .A1(n9159), .A2(n5783), .ZN(n5714) );
  INV_X1 U6203 ( .A(n5100), .ZN(n8168) );
  INV_X1 U6204 ( .A(n9331), .ZN(n9208) );
  AND2_X1 U6205 ( .A1(n8351), .A2(n8210), .ZN(n7483) );
  AND2_X1 U6206 ( .A1(n8441), .A2(n8267), .ZN(n6439) );
  NAND2_X1 U6207 ( .A1(n7632), .A2(n4952), .ZN(n7745) );
  INV_X1 U6208 ( .A(n6932), .ZN(n9640) );
  AND2_X1 U6209 ( .A1(n5575), .A2(n5550), .ZN(n5573) );
  AND2_X1 U6210 ( .A1(n5469), .A2(n5448), .ZN(n5467) );
  AND2_X1 U6211 ( .A1(n5389), .A2(n5370), .ZN(n5387) );
  NAND2_X1 U6212 ( .A1(n5043), .A2(n5042), .ZN(n5047) );
  INV_X1 U6213 ( .A(n6299), .ZN(n6300) );
  AND2_X1 U6214 ( .A1(n6298), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8543) );
  AND4_X1 U6215 ( .A1(n6200), .A2(n6199), .A3(n6198), .A4(n6197), .ZN(n8503)
         );
  AND4_X1 U6216 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n7680)
         );
  AND2_X1 U6217 ( .A1(n6611), .A2(n6610), .ZN(n9710) );
  INV_X1 U6218 ( .A(n8651), .ZN(n8825) );
  NAND2_X1 U6219 ( .A1(n8103), .A2(n8104), .ZN(n8463) );
  AND2_X1 U6220 ( .A1(n8079), .A2(n8081), .ZN(n8736) );
  OR2_X1 U6221 ( .A1(n8828), .A2(n9842), .ZN(n8832) );
  AND2_X1 U6222 ( .A1(n7816), .A2(n7815), .ZN(n8891) );
  AND2_X1 U6223 ( .A1(n6247), .A2(n6246), .ZN(n9779) );
  NAND2_X1 U6224 ( .A1(n5843), .A2(n5842), .ZN(n6283) );
  INV_X1 U6225 ( .A(n9010), .ZN(n5797) );
  AND2_X1 U6226 ( .A1(n5719), .A2(n5718), .ZN(n5747) );
  OR2_X1 U6227 ( .A1(n5348), .A2(n5347), .ZN(n5376) );
  AND2_X1 U6228 ( .A1(n5714), .A2(n5713), .ZN(n9089) );
  AND4_X1 U6229 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n7516)
         );
  OR2_X1 U6230 ( .A1(n8172), .A2(n5098), .ZN(n5108) );
  NOR2_X1 U6231 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  AND2_X1 U6232 ( .A1(n9276), .A2(n6901), .ZN(n9280) );
  INV_X1 U6233 ( .A(n9443), .ZN(n9686) );
  AND2_X1 U6234 ( .A1(n5157), .A2(n5213), .ZN(n6334) );
  OR3_X1 U6235 ( .A1(n7344), .A2(n7540), .A3(n7411), .ZN(n6571) );
  NOR2_X1 U6236 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  INV_X1 U6237 ( .A(n8520), .ZN(n8546) );
  AND4_X1 U6238 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(n8504)
         );
  INV_X1 U6239 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7930) );
  INV_X1 U6240 ( .A(n7202), .ZN(n9749) );
  OR2_X1 U6241 ( .A1(n9773), .A2(n7201), .ZN(n8808) );
  OR2_X1 U6242 ( .A1(n6567), .A2(n7199), .ZN(n9870) );
  OR2_X1 U6243 ( .A1(n6567), .A2(n6548), .ZN(n9855) );
  INV_X1 U6244 ( .A(n9781), .ZN(n9903) );
  XNOR2_X1 U6245 ( .A(n5833), .B(n5832), .ZN(n7021) );
  INV_X1 U6246 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U6247 ( .A1(n9306), .A2(n5797), .ZN(n5798) );
  INV_X1 U6248 ( .A(n9351), .ZN(n9078) );
  INV_X1 U6249 ( .A(n9346), .ZN(n9259) );
  INV_X1 U6250 ( .A(n9089), .ZN(n9174) );
  INV_X1 U6251 ( .A(n9073), .ZN(n9294) );
  OR2_X1 U6252 ( .A1(n6446), .A2(n6898), .ZN(n9705) );
  OR2_X1 U6253 ( .A1(n6446), .A2(n9395), .ZN(n9694) );
  INV_X1 U6254 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9985) );
  INV_X1 U6255 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4962) );
  INV_X1 U6256 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4961) );
  INV_X1 U6257 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6258 ( .A1(n4981), .A2(n4964), .ZN(n4970) );
  INV_X1 U6259 ( .A(n4970), .ZN(n4967) );
  NOR2_X1 U6260 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4966) );
  NAND2_X1 U6261 ( .A1(n4972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4974) );
  INV_X1 U6262 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6263 ( .A1(n4974), .A2(n4989), .ZN(n4976) );
  NAND2_X1 U6264 ( .A1(n4976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4968) );
  XNOR2_X1 U6265 ( .A(n4968), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5750) );
  OAI21_X1 U6266 ( .B1(n5768), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4971) );
  MUX2_X1 U6267 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4971), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n4973) );
  OR2_X1 U6268 ( .A1(n4974), .A2(n4989), .ZN(n4975) );
  NAND2_X1 U6269 ( .A1(n4976), .A2(n4975), .ZN(n7409) );
  INV_X1 U6270 ( .A(n7409), .ZN(n4977) );
  NAND2_X1 U6271 ( .A1(n4987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4980) );
  INV_X1 U6272 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4979) );
  NAND2_X1 U6273 ( .A1(n4980), .A2(n4979), .ZN(n4978) );
  XNOR2_X1 U6274 ( .A(n4980), .B(n4979), .ZN(n7020) );
  NAND2_X1 U6275 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  NAND2_X1 U6276 ( .A1(n4983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4984) );
  XNOR2_X1 U6277 ( .A(n4984), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8445) );
  INV_X1 U6278 ( .A(n8445), .ZN(n8441) );
  INV_X1 U6279 ( .A(n4994), .ZN(n4985) );
  NAND2_X1 U6280 ( .A1(n4985), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4986) );
  MUX2_X1 U6281 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4986), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n4988) );
  NAND2_X1 U6282 ( .A1(n4988), .A2(n4987), .ZN(n6909) );
  AND2_X1 U6283 ( .A1(n7020), .A2(n6909), .ZN(n5773) );
  NAND2_X1 U6284 ( .A1(n8441), .A2(n5773), .ZN(n6881) );
  INV_X1 U6285 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4990) );
  AND2_X1 U6286 ( .A1(n4990), .A2(n4989), .ZN(n4991) );
  INV_X1 U6287 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5005) );
  XNOR2_X2 U6288 ( .A(n4996), .B(n4995), .ZN(n4997) );
  NAND2_X1 U6289 ( .A1(n7827), .A2(n4997), .ZN(n5100) );
  NAND2_X1 U6290 ( .A1(n5374), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5002) );
  INV_X1 U6291 ( .A(n5017), .ZN(n5104) );
  INV_X1 U6292 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6451) );
  INV_X1 U6293 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5011) );
  INV_X1 U6294 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6542) );
  OR2_X1 U6295 ( .A1(n5783), .A2(n6542), .ZN(n4999) );
  NAND4_X2 U6296 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n6888)
         );
  NOR2_X1 U6297 ( .A1(n7826), .A2(n4491), .ZN(n5004) );
  INV_X1 U6298 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5003) );
  XNOR2_X1 U6299 ( .A(n5004), .B(n5003), .ZN(n9396) );
  XNOR2_X2 U6300 ( .A(n5006), .B(n5005), .ZN(n5777) );
  NAND2_X1 U6301 ( .A1(n5007), .A2(n4409), .ZN(n9067) );
  NAND2_X2 U6302 ( .A1(n5777), .A2(n9067), .ZN(n6308) );
  MUX2_X1 U6303 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9396), .S(n6308), .Z(n6904) );
  INV_X1 U6304 ( .A(n6304), .ZN(n5008) );
  AOI22_X1 U6305 ( .A1(n6904), .A2(n5167), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5008), .ZN(n5009) );
  INV_X1 U6306 ( .A(n5009), .ZN(n5010) );
  NAND2_X1 U6307 ( .A1(n6888), .A2(n5167), .ZN(n5014) );
  NOR2_X1 U6308 ( .A1(n6304), .A2(n5011), .ZN(n5012) );
  AOI21_X1 U6309 ( .B1(n6904), .B2(n7878), .A(n5012), .ZN(n5013) );
  NAND2_X1 U6310 ( .A1(n5014), .A2(n5013), .ZN(n6454) );
  INV_X1 U6311 ( .A(n6454), .ZN(n5015) );
  NAND2_X1 U6312 ( .A1(n8445), .A2(n6909), .ZN(n6880) );
  NAND2_X1 U6313 ( .A1(n5015), .A2(n6944), .ZN(n5016) );
  NAND2_X1 U6314 ( .A1(n5017), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5021) );
  INV_X1 U6315 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5018) );
  INV_X1 U6316 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6324) );
  INV_X1 U6317 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5019) );
  OR2_X1 U6318 ( .A1(n5100), .A2(n5019), .ZN(n5020) );
  NAND2_X1 U6319 ( .A1(n9027), .A2(n5167), .ZN(n5028) );
  INV_X4 U6320 ( .A(n6308), .ZN(n5522) );
  NAND2_X1 U6321 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5022) );
  NAND2_X1 U6322 ( .A1(n5522), .A2(n6364), .ZN(n5026) );
  AND2_X1 U6323 ( .A1(n6308), .A2(n7833), .ZN(n5096) );
  NAND2_X1 U6324 ( .A1(n5096), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5025) );
  XNOR2_X1 U6325 ( .A(n5044), .B(SI_1_), .ZN(n5043) );
  MUX2_X1 U6326 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5846), .Z(n5042) );
  XNOR2_X1 U6327 ( .A(n5043), .B(n5042), .ZN(n6366) );
  OR2_X1 U6328 ( .A1(n5121), .A2(n6366), .ZN(n5024) );
  NAND2_X1 U6329 ( .A1(n6932), .A2(n7878), .ZN(n5027) );
  NAND2_X1 U6330 ( .A1(n5028), .A2(n5027), .ZN(n5029) );
  NAND2_X1 U6331 ( .A1(n6519), .A2(n6520), .ZN(n5032) );
  NAND2_X1 U6332 ( .A1(n9027), .A2(n5743), .ZN(n5031) );
  NAND2_X1 U6333 ( .A1(n6932), .A2(n5167), .ZN(n5030) );
  NAND2_X1 U6334 ( .A1(n5031), .A2(n5030), .ZN(n6518) );
  NAND2_X1 U6335 ( .A1(n5032), .A2(n6518), .ZN(n5036) );
  INV_X1 U6336 ( .A(n6519), .ZN(n5034) );
  INV_X1 U6337 ( .A(n6520), .ZN(n5033) );
  NAND2_X1 U6338 ( .A1(n5034), .A2(n5033), .ZN(n5035) );
  NAND2_X1 U6339 ( .A1(n5036), .A2(n5035), .ZN(n6531) );
  INV_X1 U6340 ( .A(n6531), .ZN(n5066) );
  INV_X1 U6341 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7009) );
  OR2_X1 U6342 ( .A1(n5783), .A2(n7009), .ZN(n5041) );
  INV_X1 U6343 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U6344 ( .A1(n5017), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5039) );
  INV_X1 U6345 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5037) );
  OR2_X1 U6346 ( .A1(n5100), .A2(n5037), .ZN(n5038) );
  NAND2_X1 U6347 ( .A1(n9025), .A2(n5167), .ZN(n5056) );
  NAND2_X1 U6348 ( .A1(n5096), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5054) );
  INV_X1 U6349 ( .A(n5044), .ZN(n5045) );
  NAND2_X1 U6350 ( .A1(n5045), .A2(SI_1_), .ZN(n5046) );
  MUX2_X1 U6351 ( .A(n9907), .B(n5048), .S(n4390), .Z(n5075) );
  XNOR2_X1 U6352 ( .A(n5074), .B(n5073), .ZN(n6361) );
  OR2_X1 U6353 ( .A1(n5121), .A2(n6361), .ZN(n5053) );
  INV_X1 U6354 ( .A(n5050), .ZN(n5051) );
  NAND2_X1 U6355 ( .A1(n5522), .A2(n6470), .ZN(n5052) );
  NAND2_X1 U6356 ( .A1(n7015), .A2(n7878), .ZN(n5055) );
  NAND2_X1 U6357 ( .A1(n5056), .A2(n5055), .ZN(n5057) );
  INV_X2 U6358 ( .A(n6944), .ZN(n7881) );
  XNOR2_X1 U6359 ( .A(n5057), .B(n7881), .ZN(n5060) );
  NAND2_X1 U6360 ( .A1(n9025), .A2(n5743), .ZN(n5059) );
  NAND2_X1 U6361 ( .A1(n7015), .A2(n5167), .ZN(n5058) );
  AND2_X1 U6362 ( .A1(n5059), .A2(n5058), .ZN(n5061) );
  NAND2_X1 U6363 ( .A1(n5060), .A2(n5061), .ZN(n5067) );
  INV_X1 U6364 ( .A(n5060), .ZN(n5063) );
  INV_X1 U6365 ( .A(n5061), .ZN(n5062) );
  NAND2_X1 U6366 ( .A1(n5063), .A2(n5062), .ZN(n5064) );
  NAND2_X1 U6367 ( .A1(n5067), .A2(n5064), .ZN(n6534) );
  INV_X1 U6368 ( .A(n6534), .ZN(n5065) );
  NAND2_X1 U6369 ( .A1(n5066), .A2(n5065), .ZN(n6532) );
  NAND2_X1 U6370 ( .A1(n6532), .A2(n5067), .ZN(n6616) );
  OR2_X1 U6371 ( .A1(n5783), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5071) );
  INV_X1 U6372 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6327) );
  OR2_X1 U6373 ( .A1(n8172), .A2(n6327), .ZN(n5070) );
  INV_X1 U6374 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6375 ( .A1(n5100), .A2(n5068), .ZN(n5069) );
  NAND2_X1 U6376 ( .A1(n9024), .A2(n5167), .ZN(n5085) );
  NAND2_X1 U6377 ( .A1(n5074), .A2(n5073), .ZN(n5078) );
  INV_X1 U6378 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U6379 ( .A1(n5076), .A2(SI_2_), .ZN(n5077) );
  NAND2_X2 U6380 ( .A1(n5078), .A2(n5077), .ZN(n5144) );
  MUX2_X1 U6381 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4390), .Z(n5093) );
  INV_X1 U6382 ( .A(SI_3_), .ZN(n5079) );
  XNOR2_X1 U6383 ( .A(n5093), .B(n5079), .ZN(n5143) );
  XNOR2_X1 U6384 ( .A(n5144), .B(n5143), .ZN(n7869) );
  OR2_X1 U6385 ( .A1(n5121), .A2(n7869), .ZN(n5083) );
  NAND2_X1 U6386 ( .A1(n5732), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6387 ( .A1(n5050), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5080) );
  XNOR2_X1 U6388 ( .A(n5080), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U6389 ( .A1(n5522), .A2(n7867), .ZN(n5081) );
  INV_X1 U6390 ( .A(n6926), .ZN(n6927) );
  NAND2_X1 U6391 ( .A1(n6927), .A2(n7878), .ZN(n5084) );
  NAND2_X1 U6392 ( .A1(n5085), .A2(n5084), .ZN(n5086) );
  XNOR2_X1 U6393 ( .A(n5086), .B(n7881), .ZN(n5091) );
  NAND2_X1 U6394 ( .A1(n9024), .A2(n5743), .ZN(n5088) );
  NAND2_X1 U6395 ( .A1(n6927), .A2(n5167), .ZN(n5087) );
  NAND2_X1 U6396 ( .A1(n5088), .A2(n5087), .ZN(n5089) );
  XNOR2_X1 U6397 ( .A(n5091), .B(n5089), .ZN(n6617) );
  INV_X1 U6398 ( .A(n5089), .ZN(n5090) );
  NAND2_X1 U6399 ( .A1(n5091), .A2(n5090), .ZN(n5092) );
  NAND2_X1 U6400 ( .A1(n5144), .A2(n5143), .ZN(n5094) );
  NAND2_X1 U6401 ( .A1(n5093), .A2(SI_3_), .ZN(n5147) );
  NAND2_X1 U6402 ( .A1(n5094), .A2(n5147), .ZN(n5116) );
  XNOR2_X1 U6403 ( .A(n5116), .B(n5142), .ZN(n7874) );
  OR2_X1 U6404 ( .A1(n7874), .A2(n5121), .ZN(n6930) );
  NAND2_X1 U6405 ( .A1(n5732), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U6406 ( .A1(n5122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5097) );
  XNOR2_X1 U6407 ( .A(n5097), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U6408 ( .A1(n5522), .A2(n7871), .ZN(n6928) );
  NAND3_X1 U6409 ( .A1(n6930), .A2(n6929), .A3(n6928), .ZN(n6938) );
  NAND2_X1 U6410 ( .A1(n6938), .A2(n7878), .ZN(n5110) );
  INV_X1 U6411 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5098) );
  INV_X1 U6412 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5099) );
  OR2_X1 U6413 ( .A1(n5100), .A2(n5099), .ZN(n5107) );
  INV_X1 U6414 ( .A(n5131), .ZN(n5103) );
  INV_X1 U6415 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5101) );
  INV_X1 U6416 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U6417 ( .A1(n5101), .A2(n6618), .ZN(n5102) );
  NAND2_X1 U6418 ( .A1(n5103), .A2(n5102), .ZN(n7082) );
  OR2_X1 U6419 ( .A1(n5783), .A2(n7082), .ZN(n5106) );
  INV_X1 U6420 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U6421 ( .A1(n9023), .A2(n5167), .ZN(n5109) );
  NAND2_X1 U6422 ( .A1(n5110), .A2(n5109), .ZN(n5111) );
  XNOR2_X1 U6423 ( .A(n5111), .B(n7881), .ZN(n5113) );
  NAND2_X1 U6424 ( .A1(n9023), .A2(n5743), .ZN(n5112) );
  OAI21_X1 U6425 ( .B1(n6931), .B2(n5740), .A(n5112), .ZN(n5114) );
  XNOR2_X1 U6426 ( .A(n5113), .B(n5114), .ZN(n6685) );
  INV_X1 U6427 ( .A(n5113), .ZN(n5115) );
  NAND2_X1 U6428 ( .A1(n5116), .A2(n5142), .ZN(n5119) );
  INV_X1 U6429 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6430 ( .A1(n5118), .A2(SI_4_), .ZN(n5141) );
  NAND2_X1 U6431 ( .A1(n5119), .A2(n5141), .ZN(n5120) );
  MUX2_X1 U6432 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4390), .Z(n5140) );
  XNOR2_X1 U6433 ( .A(n5120), .B(n5152), .ZN(n5907) );
  NAND2_X1 U6434 ( .A1(n5907), .A2(n5306), .ZN(n5129) );
  NOR2_X1 U6435 ( .A1(n5125), .A2(n7842), .ZN(n5123) );
  MUX2_X1 U6436 ( .A(n7842), .B(n5123), .S(P1_IR_REG_5__SCAN_IN), .Z(n5127) );
  INV_X1 U6437 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6438 ( .A1(n5125), .A2(n5124), .ZN(n5156) );
  INV_X1 U6439 ( .A(n5156), .ZN(n5126) );
  INV_X1 U6440 ( .A(n6372), .ZN(n6427) );
  AOI22_X1 U6441 ( .A1(n5732), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5522), .B2(
        n6427), .ZN(n5128) );
  INV_X1 U6442 ( .A(n7878), .ZN(n5741) );
  NAND2_X1 U6443 ( .A1(n5374), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5135) );
  INV_X1 U6444 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5130) );
  OR2_X1 U6445 ( .A1(n8172), .A2(n5130), .ZN(n5134) );
  OAI21_X1 U6446 ( .B1(n5131), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5161), .ZN(
        n9273) );
  OR2_X1 U6447 ( .A1(n5783), .A2(n9273), .ZN(n5133) );
  INV_X1 U6448 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6316) );
  OR2_X1 U6449 ( .A1(n5104), .A2(n6316), .ZN(n5132) );
  NAND4_X1 U6450 ( .A1(n5135), .A2(n5134), .A3(n5133), .A4(n5132), .ZN(n9022)
         );
  NAND2_X1 U6451 ( .A1(n9022), .A2(n5167), .ZN(n5136) );
  OAI21_X1 U6452 ( .B1(n9663), .B2(n5741), .A(n5136), .ZN(n5137) );
  XNOR2_X1 U6453 ( .A(n5137), .B(n6944), .ZN(n5173) );
  OR2_X1 U6454 ( .A1(n9663), .A2(n5740), .ZN(n5139) );
  NAND2_X1 U6455 ( .A1(n9022), .A2(n5743), .ZN(n5138) );
  NAND2_X1 U6456 ( .A1(n5139), .A2(n5138), .ZN(n6863) );
  AND2_X1 U6457 ( .A1(n5173), .A2(n6863), .ZN(n5177) );
  NAND2_X1 U6458 ( .A1(n5140), .A2(SI_5_), .ZN(n5151) );
  INV_X1 U6459 ( .A(n5145), .ZN(n5146) );
  INV_X1 U6460 ( .A(n5151), .ZN(n5154) );
  MUX2_X1 U6461 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5334), .Z(n5186) );
  XNOR2_X1 U6462 ( .A(n5185), .B(n5183), .ZN(n6358) );
  NAND2_X1 U6463 ( .A1(n6358), .A2(n5306), .ZN(n5159) );
  NAND2_X1 U6464 ( .A1(n5156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5155) );
  MUX2_X1 U6465 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5155), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5157) );
  AOI22_X1 U6466 ( .A1(n5732), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5522), .B2(
        n6334), .ZN(n5158) );
  NAND2_X1 U6467 ( .A1(n5159), .A2(n5158), .ZN(n7064) );
  NAND2_X1 U6468 ( .A1(n7064), .A2(n7878), .ZN(n5169) );
  NAND2_X1 U6469 ( .A1(n5374), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5166) );
  INV_X1 U6470 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6335) );
  OR2_X1 U6471 ( .A1(n8172), .A2(n6335), .ZN(n5165) );
  AND2_X1 U6472 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  OR2_X1 U6473 ( .A1(n5162), .A2(n5192), .ZN(n7062) );
  OR2_X1 U6474 ( .A1(n5783), .A2(n7062), .ZN(n5164) );
  INV_X1 U6475 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6318) );
  OR2_X1 U6476 ( .A1(n5104), .A2(n6318), .ZN(n5163) );
  OR2_X1 U6477 ( .A1(n9268), .A2(n5740), .ZN(n5168) );
  NAND2_X1 U6478 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  XNOR2_X1 U6479 ( .A(n5170), .B(n7881), .ZN(n5178) );
  NAND2_X1 U6480 ( .A1(n7064), .A2(n5167), .ZN(n5172) );
  OR2_X1 U6481 ( .A1(n9268), .A2(n7884), .ZN(n5171) );
  AND2_X1 U6482 ( .A1(n5172), .A2(n5171), .ZN(n5179) );
  NAND2_X1 U6483 ( .A1(n5178), .A2(n5179), .ZN(n6912) );
  INV_X1 U6484 ( .A(n5173), .ZN(n6860) );
  INV_X1 U6485 ( .A(n6863), .ZN(n5174) );
  NAND2_X1 U6486 ( .A1(n6860), .A2(n5174), .ZN(n5175) );
  AND2_X1 U6487 ( .A1(n6912), .A2(n5175), .ZN(n5176) );
  OAI21_X1 U6488 ( .B1(n6859), .B2(n5177), .A(n5176), .ZN(n5182) );
  INV_X1 U6489 ( .A(n5178), .ZN(n5181) );
  INV_X1 U6490 ( .A(n5179), .ZN(n5180) );
  NAND2_X1 U6491 ( .A1(n5181), .A2(n5180), .ZN(n6913) );
  NAND2_X1 U6492 ( .A1(n5182), .A2(n6913), .ZN(n6791) );
  NAND2_X1 U6493 ( .A1(n5186), .A2(SI_6_), .ZN(n5187) );
  MUX2_X1 U6494 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5497), .Z(n5209) );
  XNOR2_X1 U6495 ( .A(n5208), .B(n5206), .ZN(n6367) );
  NAND2_X1 U6496 ( .A1(n6367), .A2(n5306), .ZN(n5190) );
  NAND2_X1 U6497 ( .A1(n5213), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5188) );
  XNOR2_X1 U6498 ( .A(n5188), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9516) );
  AOI22_X1 U6499 ( .A1(n5732), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5522), .B2(
        n9516), .ZN(n5189) );
  NAND2_X1 U6500 ( .A1(n5190), .A2(n5189), .ZN(n7029) );
  NAND2_X1 U6501 ( .A1(n7029), .A2(n7878), .ZN(n5199) );
  NAND2_X1 U6502 ( .A1(n5374), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5197) );
  INV_X1 U6503 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5191) );
  OR2_X1 U6504 ( .A1(n8172), .A2(n5191), .ZN(n5196) );
  OR2_X1 U6505 ( .A1(n5192), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6506 ( .A1(n5219), .A2(n5193), .ZN(n6956) );
  OR2_X1 U6507 ( .A1(n5783), .A2(n6956), .ZN(n5195) );
  INV_X1 U6508 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6957) );
  OR2_X1 U6509 ( .A1(n5104), .A2(n6957), .ZN(n5194) );
  OR2_X1 U6510 ( .A1(n6943), .A2(n5740), .ZN(n5198) );
  NAND2_X1 U6511 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  XNOR2_X1 U6512 ( .A(n5200), .B(n7881), .ZN(n6789) );
  NOR2_X1 U6513 ( .A1(n6943), .A2(n7884), .ZN(n5201) );
  AOI21_X1 U6514 ( .B1(n7029), .B2(n5167), .A(n5201), .ZN(n5203) );
  NAND2_X1 U6515 ( .A1(n6789), .A2(n5203), .ZN(n5202) );
  INV_X1 U6516 ( .A(n6789), .ZN(n5204) );
  INV_X1 U6517 ( .A(n5203), .ZN(n6788) );
  NAND2_X1 U6518 ( .A1(n5204), .A2(n6788), .ZN(n5205) );
  NAND2_X1 U6519 ( .A1(n5208), .A2(n5207), .ZN(n5267) );
  NAND2_X1 U6520 ( .A1(n5209), .A2(SI_7_), .ZN(n5263) );
  NAND2_X1 U6521 ( .A1(n5267), .A2(n5263), .ZN(n5234) );
  INV_X1 U6522 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9951) );
  INV_X1 U6523 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9973) );
  MUX2_X1 U6524 ( .A(n9951), .B(n9973), .S(n5334), .Z(n5211) );
  INV_X1 U6525 ( .A(SI_8_), .ZN(n5210) );
  NAND2_X1 U6526 ( .A1(n5211), .A2(n5210), .ZN(n5268) );
  INV_X1 U6527 ( .A(n5211), .ZN(n5212) );
  NAND2_X1 U6528 ( .A1(n5212), .A2(SI_8_), .ZN(n5262) );
  NAND2_X1 U6529 ( .A1(n5268), .A2(n5262), .ZN(n5233) );
  XNOR2_X1 U6530 ( .A(n5234), .B(n5233), .ZN(n6376) );
  NAND2_X1 U6531 ( .A1(n6376), .A2(n5306), .ZN(n5216) );
  OAI21_X1 U6532 ( .B1(n5213), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5214) );
  XNOR2_X1 U6533 ( .A(n5214), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9531) );
  AOI22_X1 U6534 ( .A1(n5732), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5522), .B2(
        n9531), .ZN(n5215) );
  NAND2_X1 U6535 ( .A1(n7044), .A2(n7878), .ZN(n5226) );
  NAND2_X1 U6536 ( .A1(n5374), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5224) );
  INV_X1 U6537 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5217) );
  OR2_X1 U6538 ( .A1(n8172), .A2(n5217), .ZN(n5223) );
  INV_X1 U6539 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7033) );
  OR2_X1 U6540 ( .A1(n5104), .A2(n7033), .ZN(n5222) );
  NAND2_X1 U6541 ( .A1(n5219), .A2(n5218), .ZN(n5220) );
  NAND2_X1 U6542 ( .A1(n5245), .A2(n5220), .ZN(n7032) );
  OR2_X1 U6543 ( .A1(n5783), .A2(n7032), .ZN(n5221) );
  OR2_X1 U6544 ( .A1(n7046), .A2(n5740), .ZN(n5225) );
  NAND2_X1 U6545 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  XNOR2_X1 U6546 ( .A(n5227), .B(n7881), .ZN(n6835) );
  NOR2_X1 U6547 ( .A1(n7046), .A2(n7884), .ZN(n5228) );
  AOI21_X1 U6548 ( .B1(n7044), .B2(n5167), .A(n5228), .ZN(n5230) );
  NAND2_X1 U6549 ( .A1(n6835), .A2(n5230), .ZN(n5229) );
  INV_X1 U6550 ( .A(n6835), .ZN(n5231) );
  INV_X1 U6551 ( .A(n5230), .ZN(n6834) );
  NAND2_X1 U6552 ( .A1(n5231), .A2(n6834), .ZN(n5232) );
  OAI21_X1 U6553 ( .B1(n5234), .B2(n5233), .A(n5268), .ZN(n5239) );
  INV_X1 U6554 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6384) );
  INV_X1 U6555 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5235) );
  MUX2_X1 U6556 ( .A(n6384), .B(n5235), .S(n5334), .Z(n5236) );
  INV_X1 U6557 ( .A(SI_9_), .ZN(n10092) );
  NAND2_X1 U6558 ( .A1(n5236), .A2(n10092), .ZN(n5269) );
  INV_X1 U6559 ( .A(n5236), .ZN(n5237) );
  NAND2_X1 U6560 ( .A1(n5237), .A2(SI_9_), .ZN(n5238) );
  XNOR2_X1 U6561 ( .A(n5239), .B(n5272), .ZN(n6380) );
  NAND2_X1 U6562 ( .A1(n6380), .A2(n5306), .ZN(n5242) );
  NAND2_X1 U6563 ( .A1(n5279), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5240) );
  XNOR2_X1 U6564 ( .A(n5240), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6631) );
  AOI22_X1 U6565 ( .A1(n5732), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5522), .B2(
        n6631), .ZN(n5241) );
  NAND2_X1 U6566 ( .A1(n7103), .A2(n7878), .ZN(n5252) );
  NAND2_X1 U6567 ( .A1(n5374), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5250) );
  INV_X1 U6568 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5243) );
  OR2_X1 U6569 ( .A1(n8172), .A2(n5243), .ZN(n5249) );
  INV_X1 U6570 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5244) );
  AND2_X1 U6571 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  OR2_X1 U6572 ( .A1(n5246), .A2(n5286), .ZN(n7050) );
  OR2_X1 U6573 ( .A1(n5783), .A2(n7050), .ZN(n5248) );
  INV_X1 U6574 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7051) );
  OR2_X1 U6575 ( .A1(n5104), .A2(n7051), .ZN(n5247) );
  NAND4_X1 U6576 ( .A1(n5250), .A2(n5249), .A3(n5248), .A4(n5247), .ZN(n9017)
         );
  NAND2_X1 U6577 ( .A1(n9017), .A2(n5167), .ZN(n5251) );
  NAND2_X1 U6578 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  XNOR2_X1 U6579 ( .A(n5253), .B(n7881), .ZN(n5255) );
  AND2_X1 U6580 ( .A1(n9017), .A2(n5743), .ZN(n5254) );
  AOI21_X1 U6581 ( .B1(n7103), .B2(n5167), .A(n5254), .ZN(n5256) );
  NAND2_X1 U6582 ( .A1(n5255), .A2(n5256), .ZN(n5261) );
  INV_X1 U6583 ( .A(n5255), .ZN(n5258) );
  INV_X1 U6584 ( .A(n5256), .ZN(n5257) );
  NAND2_X1 U6585 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  NAND2_X1 U6586 ( .A1(n5261), .A2(n5259), .ZN(n6973) );
  NAND2_X1 U6587 ( .A1(n6971), .A2(n5261), .ZN(n7092) );
  NAND2_X1 U6588 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  NAND2_X1 U6589 ( .A1(n5267), .A2(n5266), .ZN(n5274) );
  INV_X1 U6590 ( .A(n5269), .ZN(n5270) );
  INV_X1 U6591 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6500) );
  MUX2_X1 U6592 ( .A(n6500), .B(n9985), .S(n5334), .Z(n5276) );
  INV_X1 U6593 ( .A(SI_10_), .ZN(n5275) );
  INV_X1 U6594 ( .A(n5276), .ZN(n5277) );
  NAND2_X1 U6595 ( .A1(n5277), .A2(SI_10_), .ZN(n5278) );
  NAND2_X1 U6596 ( .A1(n6382), .A2(n5306), .ZN(n5285) );
  NOR2_X1 U6597 ( .A1(n5279), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5341) );
  OR2_X1 U6598 ( .A1(n5341), .A2(n7842), .ZN(n5282) );
  INV_X1 U6599 ( .A(n5282), .ZN(n5280) );
  NAND2_X1 U6600 ( .A1(n5280), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5283) );
  INV_X1 U6601 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6602 ( .A1(n5282), .A2(n5281), .ZN(n5307) );
  AND2_X1 U6603 ( .A1(n5283), .A2(n5307), .ZN(n6700) );
  AOI22_X1 U6604 ( .A1(n5732), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5522), .B2(
        n6700), .ZN(n5284) );
  NAND2_X1 U6605 ( .A1(n5285), .A2(n5284), .ZN(n7128) );
  NAND2_X1 U6606 ( .A1(n7128), .A2(n7878), .ZN(n5295) );
  NAND2_X1 U6607 ( .A1(n5017), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5293) );
  NOR2_X1 U6608 ( .A1(n5286), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5287) );
  OR2_X1 U6609 ( .A1(n5312), .A2(n5287), .ZN(n7115) );
  OR2_X1 U6610 ( .A1(n5783), .A2(n7115), .ZN(n5292) );
  INV_X1 U6611 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5288) );
  OR2_X1 U6612 ( .A1(n8172), .A2(n5288), .ZN(n5291) );
  INV_X1 U6613 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5289) );
  OR2_X1 U6614 ( .A1(n5100), .A2(n5289), .ZN(n5290) );
  OR2_X1 U6615 ( .A1(n7177), .A2(n5740), .ZN(n5294) );
  NAND2_X1 U6616 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  XNOR2_X1 U6617 ( .A(n5296), .B(n6944), .ZN(n5299) );
  NAND2_X1 U6618 ( .A1(n7128), .A2(n5167), .ZN(n5298) );
  OR2_X1 U6619 ( .A1(n7177), .A2(n7884), .ZN(n5297) );
  NAND2_X1 U6620 ( .A1(n5298), .A2(n5297), .ZN(n5300) );
  NAND2_X1 U6621 ( .A1(n5299), .A2(n5300), .ZN(n7094) );
  NAND2_X1 U6622 ( .A1(n7092), .A2(n7094), .ZN(n5303) );
  INV_X1 U6623 ( .A(n5299), .ZN(n5302) );
  INV_X1 U6624 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U6625 ( .A1(n5302), .A2(n5301), .ZN(n7093) );
  NAND2_X1 U6626 ( .A1(n5303), .A2(n7093), .ZN(n7171) );
  INV_X1 U6627 ( .A(n7171), .ZN(n5323) );
  INV_X1 U6628 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10104) );
  INV_X1 U6629 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6387) );
  MUX2_X1 U6630 ( .A(n10104), .B(n6387), .S(n5334), .Z(n5330) );
  XNOR2_X1 U6631 ( .A(n5333), .B(n5329), .ZN(n6386) );
  NAND2_X1 U6632 ( .A1(n6386), .A2(n5306), .ZN(n5310) );
  NAND2_X1 U6633 ( .A1(n5307), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5308) );
  XNOR2_X1 U6634 ( .A(n5308), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9042) );
  AOI22_X1 U6635 ( .A1(n5732), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5522), .B2(
        n9042), .ZN(n5309) );
  NAND2_X1 U6636 ( .A1(n7249), .A2(n7878), .ZN(n5319) );
  NAND2_X1 U6637 ( .A1(n5374), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5317) );
  INV_X1 U6638 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5311) );
  OR2_X1 U6639 ( .A1(n8172), .A2(n5311), .ZN(n5316) );
  OR2_X1 U6640 ( .A1(n5312), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6641 ( .A1(n5348), .A2(n5313), .ZN(n7174) );
  OR2_X1 U6642 ( .A1(n5783), .A2(n7174), .ZN(n5315) );
  INV_X1 U6643 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7142) );
  OR2_X1 U6644 ( .A1(n5104), .A2(n7142), .ZN(n5314) );
  NAND4_X1 U6645 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n9016)
         );
  NAND2_X1 U6646 ( .A1(n9016), .A2(n5167), .ZN(n5318) );
  NAND2_X1 U6647 ( .A1(n5319), .A2(n5318), .ZN(n5320) );
  XNOR2_X1 U6648 ( .A(n5320), .B(n7881), .ZN(n5324) );
  AND2_X1 U6649 ( .A1(n9016), .A2(n5743), .ZN(n5321) );
  AOI21_X1 U6650 ( .B1(n7249), .B2(n5167), .A(n5321), .ZN(n5325) );
  XNOR2_X1 U6651 ( .A(n5324), .B(n5325), .ZN(n7170) );
  INV_X1 U6652 ( .A(n7170), .ZN(n5322) );
  INV_X1 U6653 ( .A(n5324), .ZN(n5327) );
  INV_X1 U6654 ( .A(n5325), .ZN(n5326) );
  NAND2_X1 U6655 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  INV_X1 U6656 ( .A(n5330), .ZN(n5331) );
  INV_X1 U6657 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6498) );
  INV_X1 U6658 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5335) );
  INV_X1 U6659 ( .A(n7826), .ZN(n5334) );
  MUX2_X1 U6660 ( .A(n6498), .B(n5335), .S(n5334), .Z(n5337) );
  INV_X1 U6661 ( .A(SI_12_), .ZN(n5336) );
  INV_X1 U6662 ( .A(n5337), .ZN(n5338) );
  NAND2_X1 U6663 ( .A1(n5338), .A2(SI_12_), .ZN(n5339) );
  XNOR2_X1 U6664 ( .A(n5364), .B(n5363), .ZN(n6401) );
  NAND2_X1 U6665 ( .A1(n6401), .A2(n5306), .ZN(n5346) );
  NOR2_X1 U6666 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5340) );
  NAND2_X1 U6667 ( .A1(n5341), .A2(n5340), .ZN(n5343) );
  NAND2_X1 U6668 ( .A1(n5343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5342) );
  MUX2_X1 U6669 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5342), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5344) );
  OR2_X1 U6670 ( .A1(n5343), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5391) );
  AND2_X1 U6671 ( .A1(n5344), .A2(n5391), .ZN(n9543) );
  AOI22_X1 U6672 ( .A1(n5732), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5522), .B2(
        n9543), .ZN(n5345) );
  NAND2_X1 U6673 ( .A1(n9444), .A2(n7878), .ZN(n5356) );
  NAND2_X1 U6674 ( .A1(n5017), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5354) );
  INV_X1 U6675 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9028) );
  OR2_X1 U6676 ( .A1(n8172), .A2(n9028), .ZN(n5353) );
  INV_X1 U6677 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6678 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6679 ( .A1(n5376), .A2(n5349), .ZN(n9451) );
  OR2_X1 U6680 ( .A1(n5783), .A2(n9451), .ZN(n5352) );
  INV_X1 U6681 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5350) );
  OR2_X1 U6682 ( .A1(n5100), .A2(n5350), .ZN(n5351) );
  OR2_X1 U6683 ( .A1(n7516), .A2(n5740), .ZN(n5355) );
  NAND2_X1 U6684 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  XNOR2_X1 U6685 ( .A(n5357), .B(n7881), .ZN(n5361) );
  NOR2_X1 U6686 ( .A1(n7516), .A2(n7884), .ZN(n5358) );
  AOI21_X1 U6687 ( .B1(n9444), .B2(n5167), .A(n5358), .ZN(n5360) );
  XNOR2_X1 U6688 ( .A(n5361), .B(n5360), .ZN(n9442) );
  NAND2_X1 U6689 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  INV_X1 U6690 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6516) );
  INV_X1 U6691 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5366) );
  MUX2_X1 U6692 ( .A(n6516), .B(n5366), .S(n5334), .Z(n5368) );
  INV_X1 U6693 ( .A(SI_13_), .ZN(n5367) );
  NAND2_X1 U6694 ( .A1(n5368), .A2(n5367), .ZN(n5389) );
  INV_X1 U6695 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6696 ( .A1(n5369), .A2(SI_13_), .ZN(n5370) );
  XNOR2_X1 U6697 ( .A(n5388), .B(n5387), .ZN(n6449) );
  NAND2_X1 U6698 ( .A1(n6449), .A2(n5306), .ZN(n5373) );
  NAND2_X1 U6699 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U6700 ( .A(n5371), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U6701 ( .A1(n5732), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5522), .B2(
        n9552), .ZN(n5372) );
  NAND2_X1 U6702 ( .A1(n7521), .A2(n7878), .ZN(n5383) );
  NAND2_X1 U6703 ( .A1(n5374), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5381) );
  INV_X1 U6704 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9032) );
  OR2_X1 U6705 ( .A1(n8172), .A2(n9032), .ZN(n5380) );
  INV_X1 U6706 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6707 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  NAND2_X1 U6708 ( .A1(n5400), .A2(n5377), .ZN(n7519) );
  OR2_X1 U6709 ( .A1(n5783), .A2(n7519), .ZN(n5379) );
  INV_X1 U6710 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9047) );
  OR2_X1 U6711 ( .A1(n5104), .A2(n9047), .ZN(n5378) );
  NAND4_X1 U6712 ( .A1(n5381), .A2(n5380), .A3(n5379), .A4(n5378), .ZN(n9437)
         );
  NAND2_X1 U6713 ( .A1(n9437), .A2(n5167), .ZN(n5382) );
  NAND2_X1 U6714 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  XNOR2_X1 U6715 ( .A(n5384), .B(n7881), .ZN(n7513) );
  AND2_X1 U6716 ( .A1(n9437), .A2(n5743), .ZN(n5385) );
  AOI21_X1 U6717 ( .B1(n7521), .B2(n5167), .A(n5385), .ZN(n7512) );
  AND2_X1 U6718 ( .A1(n7513), .A2(n7512), .ZN(n5386) );
  NAND2_X1 U6719 ( .A1(n5388), .A2(n5387), .ZN(n5390) );
  INV_X1 U6720 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6530) );
  INV_X1 U6721 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6528) );
  MUX2_X1 U6722 ( .A(n6530), .B(n6528), .S(n5497), .Z(n5415) );
  XNOR2_X1 U6723 ( .A(n5415), .B(SI_14_), .ZN(n5414) );
  XNOR2_X1 U6724 ( .A(n5419), .B(n5414), .ZN(n6527) );
  NAND2_X1 U6725 ( .A1(n6527), .A2(n5306), .ZN(n5397) );
  NOR2_X1 U6726 ( .A1(n5391), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5450) );
  OR2_X1 U6727 ( .A1(n5450), .A2(n7842), .ZN(n5394) );
  INV_X1 U6728 ( .A(n5394), .ZN(n5392) );
  NAND2_X1 U6729 ( .A1(n5392), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5395) );
  INV_X1 U6730 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6731 ( .A1(n5394), .A2(n5393), .ZN(n5423) );
  AND2_X1 U6732 ( .A1(n5395), .A2(n5423), .ZN(n9568) );
  AOI22_X1 U6733 ( .A1(n5732), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5522), .B2(
        n9568), .ZN(n5396) );
  NAND2_X1 U6734 ( .A1(n7628), .A2(n7878), .ZN(n5407) );
  NAND2_X1 U6735 ( .A1(n8168), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5405) );
  INV_X1 U6736 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5398) );
  OR2_X1 U6737 ( .A1(n8172), .A2(n5398), .ZN(n5404) );
  INV_X1 U6738 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U6739 ( .A1(n5400), .A2(n7528), .ZN(n5401) );
  NAND2_X1 U6740 ( .A1(n5430), .A2(n5401), .ZN(n7532) );
  OR2_X1 U6741 ( .A1(n5783), .A2(n7532), .ZN(n5403) );
  INV_X1 U6742 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7447) );
  OR2_X1 U6743 ( .A1(n5104), .A2(n7447), .ZN(n5402) );
  NAND4_X1 U6744 ( .A1(n5405), .A2(n5404), .A3(n5403), .A4(n5402), .ZN(n9015)
         );
  NAND2_X1 U6745 ( .A1(n9015), .A2(n5167), .ZN(n5406) );
  NAND2_X1 U6746 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  XNOR2_X1 U6747 ( .A(n5408), .B(n7881), .ZN(n7525) );
  AND2_X1 U6748 ( .A1(n9015), .A2(n5743), .ZN(n5409) );
  AOI21_X1 U6749 ( .B1(n7628), .B2(n5167), .A(n5409), .ZN(n5410) );
  INV_X1 U6750 ( .A(n7525), .ZN(n5411) );
  INV_X1 U6751 ( .A(n5410), .ZN(n7524) );
  NAND2_X1 U6752 ( .A1(n5411), .A2(n7524), .ZN(n5412) );
  NAND2_X1 U6753 ( .A1(n5413), .A2(n5412), .ZN(n7589) );
  INV_X1 U6754 ( .A(n5415), .ZN(n5416) );
  NAND2_X1 U6755 ( .A1(n5416), .A2(SI_14_), .ZN(n5417) );
  INV_X1 U6756 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6644) );
  INV_X1 U6757 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6642) );
  MUX2_X1 U6758 ( .A(n6644), .B(n6642), .S(n5497), .Z(n5420) );
  NAND2_X1 U6759 ( .A1(n5420), .A2(n9990), .ZN(n5444) );
  INV_X1 U6760 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6761 ( .A1(n5421), .A2(SI_15_), .ZN(n5422) );
  NAND2_X1 U6762 ( .A1(n5444), .A2(n5422), .ZN(n5442) );
  XNOR2_X1 U6763 ( .A(n5443), .B(n5442), .ZN(n6641) );
  NAND2_X1 U6764 ( .A1(n6641), .A2(n5306), .ZN(n5426) );
  NAND2_X1 U6765 ( .A1(n5423), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5424) );
  XNOR2_X1 U6766 ( .A(n5424), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9581) );
  AOI22_X1 U6767 ( .A1(n5732), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5522), .B2(
        n9581), .ZN(n5425) );
  NAND2_X1 U6768 ( .A1(n9365), .A2(n5167), .ZN(n5438) );
  NAND2_X1 U6769 ( .A1(n8168), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5436) );
  INV_X1 U6770 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5427) );
  OR2_X1 U6771 ( .A1(n8172), .A2(n5427), .ZN(n5435) );
  INV_X1 U6772 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6773 ( .A1(n5430), .A2(n5429), .ZN(n5431) );
  NAND2_X1 U6774 ( .A1(n5454), .A2(n5431), .ZN(n7656) );
  OR2_X1 U6775 ( .A1(n5783), .A2(n7656), .ZN(n5434) );
  INV_X1 U6776 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5432) );
  OR2_X1 U6777 ( .A1(n5104), .A2(n5432), .ZN(n5433) );
  NAND4_X1 U6778 ( .A1(n5436), .A2(n5435), .A3(n5434), .A4(n5433), .ZN(n9014)
         );
  NAND2_X1 U6779 ( .A1(n9014), .A2(n5743), .ZN(n5437) );
  NAND2_X1 U6780 ( .A1(n5438), .A2(n5437), .ZN(n7587) );
  NAND2_X1 U6781 ( .A1(n9365), .A2(n7878), .ZN(n5440) );
  NAND2_X1 U6782 ( .A1(n9014), .A2(n5167), .ZN(n5439) );
  NAND2_X1 U6783 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  XNOR2_X1 U6784 ( .A(n5441), .B(n6944), .ZN(n7586) );
  INV_X1 U6785 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6738) );
  INV_X1 U6786 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6740) );
  MUX2_X1 U6787 ( .A(n6738), .B(n6740), .S(n5497), .Z(n5446) );
  INV_X1 U6788 ( .A(SI_16_), .ZN(n10081) );
  NAND2_X1 U6789 ( .A1(n5446), .A2(n10081), .ZN(n5469) );
  INV_X1 U6790 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6791 ( .A1(n5447), .A2(SI_16_), .ZN(n5448) );
  XNOR2_X1 U6792 ( .A(n5468), .B(n5467), .ZN(n6737) );
  NAND2_X1 U6793 ( .A1(n6737), .A2(n5306), .ZN(n5453) );
  NOR2_X1 U6794 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5449) );
  NAND2_X1 U6795 ( .A1(n5450), .A2(n5449), .ZN(n5471) );
  NAND2_X1 U6796 ( .A1(n5471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5451) );
  XNOR2_X1 U6797 ( .A(n5451), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9593) );
  AOI22_X1 U6798 ( .A1(n5732), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5522), .B2(
        n9593), .ZN(n5452) );
  INV_X1 U6799 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U6800 ( .A1(n5454), .A2(n7737), .ZN(n5455) );
  AND2_X1 U6801 ( .A1(n5480), .A2(n5455), .ZN(n7736) );
  INV_X1 U6802 ( .A(n5783), .ZN(n6983) );
  NAND2_X1 U6803 ( .A1(n7736), .A2(n6983), .ZN(n5459) );
  NAND2_X1 U6804 ( .A1(n8168), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6805 ( .A1(n4641), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U6806 ( .A1(n5017), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5456) );
  NOR2_X1 U6807 ( .A1(n7649), .A2(n5740), .ZN(n5460) );
  AOI21_X1 U6808 ( .B1(n7743), .B2(n7878), .A(n5460), .ZN(n5461) );
  XNOR2_X1 U6809 ( .A(n5461), .B(n6944), .ZN(n5464) );
  NOR2_X1 U6810 ( .A1(n7649), .A2(n7884), .ZN(n5462) );
  AOI21_X1 U6811 ( .B1(n7743), .B2(n5167), .A(n5462), .ZN(n5463) );
  OR2_X1 U6812 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U6813 ( .A1(n5464), .A2(n5463), .ZN(n5466) );
  NAND2_X1 U6814 ( .A1(n5465), .A2(n5466), .ZN(n7734) );
  NAND2_X1 U6815 ( .A1(n7732), .A2(n5466), .ZN(n7785) );
  NAND2_X1 U6816 ( .A1(n5468), .A2(n5467), .ZN(n5470) );
  INV_X1 U6817 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6787) );
  INV_X1 U6818 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10053) );
  MUX2_X1 U6819 ( .A(n6787), .B(n10053), .S(n5497), .Z(n5494) );
  XNOR2_X1 U6820 ( .A(n5494), .B(SI_17_), .ZN(n5493) );
  XNOR2_X1 U6821 ( .A(n5492), .B(n5493), .ZN(n6785) );
  NAND2_X1 U6822 ( .A1(n6785), .A2(n5306), .ZN(n5477) );
  OR2_X1 U6823 ( .A1(n5471), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6824 ( .A1(n5472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5474) );
  OR2_X1 U6825 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  NAND2_X1 U6826 ( .A1(n5474), .A2(n5473), .ZN(n5498) );
  AND2_X1 U6827 ( .A1(n5475), .A2(n5498), .ZN(n9601) );
  AOI22_X1 U6828 ( .A1(n5732), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5522), .B2(
        n9601), .ZN(n5476) );
  INV_X1 U6829 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6830 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  NAND2_X1 U6831 ( .A1(n5502), .A2(n5481), .ZN(n7762) );
  OR2_X1 U6832 ( .A1(n7762), .A2(n5783), .ZN(n5484) );
  AOI22_X1 U6833 ( .A1(n4641), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n8168), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U6834 ( .A1(n5017), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5482) );
  OAI22_X1 U6835 ( .A1(n7794), .A2(n5741), .B1(n8992), .B2(n5740), .ZN(n5485)
         );
  XNOR2_X1 U6836 ( .A(n5485), .B(n7881), .ZN(n5490) );
  OR2_X1 U6837 ( .A1(n7794), .A2(n5740), .ZN(n5487) );
  INV_X1 U6838 ( .A(n8992), .ZN(n9012) );
  NAND2_X1 U6839 ( .A1(n9012), .A2(n5743), .ZN(n5486) );
  NAND2_X1 U6840 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  XNOR2_X1 U6841 ( .A(n5490), .B(n5488), .ZN(n7787) );
  INV_X1 U6842 ( .A(n5488), .ZN(n5489) );
  NAND2_X1 U6843 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  INV_X1 U6844 ( .A(n5494), .ZN(n5495) );
  NAND2_X1 U6845 ( .A1(n5495), .A2(SI_17_), .ZN(n5496) );
  MUX2_X1 U6846 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5497), .Z(n5515) );
  XNOR2_X1 U6847 ( .A(n5515), .B(SI_18_), .ZN(n5512) );
  XNOR2_X1 U6848 ( .A(n5514), .B(n5512), .ZN(n6844) );
  NAND2_X1 U6849 ( .A1(n6844), .A2(n5306), .ZN(n5501) );
  NAND2_X1 U6850 ( .A1(n5498), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5499) );
  XNOR2_X1 U6851 ( .A(n5499), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U6852 ( .A1(n5522), .A2(n9620), .B1(n5732), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6853 ( .A1(n9356), .A2(n7878), .ZN(n5508) );
  INV_X1 U6854 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U6855 ( .A1(n5502), .A2(n9982), .ZN(n5503) );
  AND2_X1 U6856 ( .A1(n5527), .A2(n5503), .ZN(n8994) );
  NAND2_X1 U6857 ( .A1(n8994), .A2(n6983), .ZN(n5506) );
  AOI22_X1 U6858 ( .A1(n4641), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8168), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5505) );
  INV_X1 U6859 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9057) );
  OR2_X1 U6860 ( .A1(n5104), .A2(n9057), .ZN(n5504) );
  INV_X1 U6861 ( .A(n7800), .ZN(n9011) );
  NAND2_X1 U6862 ( .A1(n9011), .A2(n5167), .ZN(n5507) );
  NAND2_X1 U6863 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  XNOR2_X1 U6864 ( .A(n5509), .B(n7881), .ZN(n5511) );
  NOR2_X1 U6865 ( .A1(n7800), .A2(n7884), .ZN(n5510) );
  AOI21_X1 U6866 ( .B1(n9356), .B2(n5167), .A(n5510), .ZN(n8987) );
  INV_X1 U6867 ( .A(n5512), .ZN(n5513) );
  NAND2_X1 U6868 ( .A1(n5514), .A2(n5513), .ZN(n5517) );
  NAND2_X1 U6869 ( .A1(n5515), .A2(SI_18_), .ZN(n5516) );
  INV_X1 U6870 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9924) );
  INV_X1 U6871 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6910) );
  MUX2_X1 U6872 ( .A(n9924), .B(n6910), .S(n5497), .Z(n5519) );
  INV_X1 U6873 ( .A(SI_19_), .ZN(n5518) );
  NAND2_X1 U6874 ( .A1(n5519), .A2(n5518), .ZN(n5544) );
  INV_X1 U6875 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U6876 ( .A1(n5520), .A2(SI_19_), .ZN(n5521) );
  NAND2_X1 U6877 ( .A1(n5544), .A2(n5521), .ZN(n5545) );
  XNOR2_X1 U6878 ( .A(n5546), .B(n5545), .ZN(n6908) );
  NAND2_X1 U6879 ( .A1(n6908), .A2(n5306), .ZN(n5524) );
  INV_X1 U6880 ( .A(n6909), .ZN(n9275) );
  AOI22_X1 U6881 ( .A1(n5732), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9275), .B2(
        n5522), .ZN(n5523) );
  NAND2_X1 U6882 ( .A1(n9351), .A2(n7878), .ZN(n5535) );
  INV_X1 U6883 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6884 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  NAND2_X1 U6885 ( .A1(n5554), .A2(n5528), .ZN(n8935) );
  OR2_X1 U6886 ( .A1(n8935), .A2(n5783), .ZN(n5533) );
  INV_X1 U6887 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U6888 ( .A1(n4641), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U6889 ( .A1(n8168), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5529) );
  OAI211_X1 U6890 ( .C1(n5104), .C2(n9061), .A(n5530), .B(n5529), .ZN(n5531)
         );
  INV_X1 U6891 ( .A(n5531), .ZN(n5532) );
  NAND2_X1 U6892 ( .A1(n5533), .A2(n5532), .ZN(n9077) );
  NAND2_X1 U6893 ( .A1(n9077), .A2(n5167), .ZN(n5534) );
  NAND2_X1 U6894 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  XNOR2_X1 U6895 ( .A(n5536), .B(n7881), .ZN(n5538) );
  AND2_X1 U6896 ( .A1(n9077), .A2(n5743), .ZN(n5537) );
  AOI21_X1 U6897 ( .B1(n9351), .B2(n5167), .A(n5537), .ZN(n5539) );
  NAND2_X1 U6898 ( .A1(n5538), .A2(n5539), .ZN(n8965) );
  INV_X1 U6899 ( .A(n5538), .ZN(n5541) );
  INV_X1 U6900 ( .A(n5539), .ZN(n5540) );
  NAND2_X1 U6901 ( .A1(n5541), .A2(n5540), .ZN(n5542) );
  NAND2_X1 U6902 ( .A1(n5543), .A2(n8931), .ZN(n8933) );
  NAND2_X1 U6903 ( .A1(n8933), .A2(n8965), .ZN(n5571) );
  INV_X1 U6904 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9936) );
  INV_X1 U6905 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7019) );
  MUX2_X1 U6906 ( .A(n9936), .B(n7019), .S(n5497), .Z(n5548) );
  INV_X1 U6907 ( .A(SI_20_), .ZN(n5547) );
  NAND2_X1 U6908 ( .A1(n5548), .A2(n5547), .ZN(n5575) );
  INV_X1 U6909 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U6910 ( .A1(n5549), .A2(SI_20_), .ZN(n5550) );
  XNOR2_X1 U6911 ( .A(n5574), .B(n5573), .ZN(n7018) );
  NAND2_X1 U6912 ( .A1(n7018), .A2(n5306), .ZN(n5552) );
  NAND2_X1 U6913 ( .A1(n5732), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6914 ( .A1(n9346), .A2(n7878), .ZN(n5563) );
  INV_X1 U6915 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U6916 ( .A1(n5554), .A2(n5553), .ZN(n5555) );
  AND2_X1 U6917 ( .A1(n5580), .A2(n5555), .ZN(n9255) );
  NAND2_X1 U6918 ( .A1(n9255), .A2(n6983), .ZN(n5561) );
  INV_X1 U6919 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U6920 ( .A1(n5017), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U6921 ( .A1(n8168), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5556) );
  OAI211_X1 U6922 ( .C1(n8172), .C2(n5558), .A(n5557), .B(n5556), .ZN(n5559)
         );
  INV_X1 U6923 ( .A(n5559), .ZN(n5560) );
  NAND2_X1 U6924 ( .A1(n5561), .A2(n5560), .ZN(n9081) );
  NAND2_X1 U6925 ( .A1(n9081), .A2(n5167), .ZN(n5562) );
  NAND2_X1 U6926 ( .A1(n5563), .A2(n5562), .ZN(n5564) );
  XNOR2_X1 U6927 ( .A(n5564), .B(n7881), .ZN(n5566) );
  AND2_X1 U6928 ( .A1(n9081), .A2(n5743), .ZN(n5565) );
  AOI21_X1 U6929 ( .B1(n9346), .B2(n5167), .A(n5565), .ZN(n5567) );
  NAND2_X1 U6930 ( .A1(n5566), .A2(n5567), .ZN(n5572) );
  INV_X1 U6931 ( .A(n5566), .ZN(n5569) );
  INV_X1 U6932 ( .A(n5567), .ZN(n5568) );
  NAND2_X1 U6933 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  AND2_X1 U6934 ( .A1(n5572), .A2(n5570), .ZN(n8966) );
  NAND2_X1 U6935 ( .A1(n5571), .A2(n8966), .ZN(n8969) );
  NAND2_X1 U6936 ( .A1(n8969), .A2(n5572), .ZN(n8941) );
  INV_X1 U6937 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7148) );
  INV_X1 U6938 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10003) );
  MUX2_X1 U6939 ( .A(n7148), .B(n10003), .S(n5497), .Z(n5597) );
  XNOR2_X1 U6940 ( .A(n5597), .B(SI_21_), .ZN(n5596) );
  XNOR2_X1 U6941 ( .A(n5622), .B(n5596), .ZN(n7147) );
  NAND2_X1 U6942 ( .A1(n7147), .A2(n5306), .ZN(n5577) );
  NAND2_X1 U6943 ( .A1(n5732), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U6944 ( .A1(n9341), .A2(n7878), .ZN(n5589) );
  INV_X1 U6945 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U6946 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  NAND2_X1 U6947 ( .A1(n5608), .A2(n5581), .ZN(n9237) );
  OR2_X1 U6948 ( .A1(n9237), .A2(n5783), .ZN(n5587) );
  INV_X1 U6949 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U6950 ( .A1(n8168), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U6951 ( .A1(n5017), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5582) );
  OAI211_X1 U6952 ( .C1(n8172), .C2(n5584), .A(n5583), .B(n5582), .ZN(n5585)
         );
  INV_X1 U6953 ( .A(n5585), .ZN(n5586) );
  INV_X1 U6954 ( .A(n9246), .ZN(n9221) );
  NAND2_X1 U6955 ( .A1(n9221), .A2(n5167), .ZN(n5588) );
  NAND2_X1 U6956 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  XNOR2_X1 U6957 ( .A(n5590), .B(n6944), .ZN(n5592) );
  NOR2_X1 U6958 ( .A1(n9246), .A2(n7884), .ZN(n5591) );
  AOI21_X1 U6959 ( .B1(n9341), .B2(n5167), .A(n5591), .ZN(n5593) );
  XNOR2_X1 U6960 ( .A(n5592), .B(n5593), .ZN(n8942) );
  NAND2_X1 U6961 ( .A1(n8941), .A2(n8942), .ZN(n8940) );
  INV_X1 U6962 ( .A(n5592), .ZN(n5594) );
  NAND2_X1 U6963 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  INV_X1 U6964 ( .A(n5596), .ZN(n5620) );
  OR2_X1 U6965 ( .A1(n5622), .A2(n5620), .ZN(n5599) );
  INV_X1 U6966 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U6967 ( .A1(n5598), .A2(SI_21_), .ZN(n5624) );
  INV_X1 U6968 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8451) );
  INV_X1 U6969 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7216) );
  MUX2_X1 U6970 ( .A(n8451), .B(n7216), .S(n5497), .Z(n5601) );
  INV_X1 U6971 ( .A(SI_22_), .ZN(n5600) );
  NAND2_X1 U6972 ( .A1(n5601), .A2(n5600), .ZN(n5619) );
  INV_X1 U6973 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U6974 ( .A1(n5602), .A2(SI_22_), .ZN(n5603) );
  NAND2_X1 U6975 ( .A1(n5619), .A2(n5603), .ZN(n5623) );
  NAND2_X1 U6976 ( .A1(n7215), .A2(n5306), .ZN(n5606) );
  NAND2_X1 U6977 ( .A1(n5732), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5605) );
  OR2_X1 U6978 ( .A1(n9215), .A2(n5740), .ZN(n5616) );
  INV_X1 U6979 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U6980 ( .A1(n5608), .A2(n5607), .ZN(n5609) );
  AND2_X1 U6981 ( .A1(n5638), .A2(n5609), .ZN(n9213) );
  NAND2_X1 U6982 ( .A1(n9213), .A2(n6983), .ZN(n5614) );
  INV_X1 U6983 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10094) );
  NAND2_X1 U6984 ( .A1(n5017), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U6985 ( .A1(n8168), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U6986 ( .C1(n8172), .C2(n10094), .A(n5611), .B(n5610), .ZN(n5612)
         );
  INV_X1 U6987 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U6988 ( .A1(n9083), .A2(n5743), .ZN(n5615) );
  OAI22_X1 U6989 ( .A1(n9215), .A2(n5741), .B1(n9233), .B2(n5740), .ZN(n5617)
         );
  XNOR2_X1 U6990 ( .A(n5617), .B(n7881), .ZN(n8978) );
  INV_X1 U6991 ( .A(n5619), .ZN(n5627) );
  OR2_X1 U6992 ( .A1(n5620), .A2(n5627), .ZN(n5621) );
  INV_X1 U6993 ( .A(n5623), .ZN(n5625) );
  AND2_X1 U6994 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  OR2_X1 U6995 ( .A1(n5627), .A2(n5626), .ZN(n5649) );
  INV_X1 U6997 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9940) );
  INV_X1 U6998 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5628) );
  MUX2_X1 U6999 ( .A(n9940), .B(n5628), .S(n5497), .Z(n5630) );
  INV_X1 U7000 ( .A(SI_23_), .ZN(n5629) );
  NAND2_X1 U7001 ( .A1(n5630), .A2(n5629), .ZN(n5653) );
  INV_X1 U7002 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U7003 ( .A1(n5631), .A2(SI_23_), .ZN(n5632) );
  AND2_X1 U7004 ( .A1(n5653), .A2(n5632), .ZN(n5650) );
  NAND2_X1 U7005 ( .A1(n7235), .A2(n5306), .ZN(n5635) );
  NAND2_X1 U7006 ( .A1(n5732), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7007 ( .A1(n9331), .A2(n7878), .ZN(n5646) );
  INV_X1 U7008 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7009 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  NAND2_X1 U7010 ( .A1(n5658), .A2(n5639), .ZN(n9204) );
  OR2_X1 U7011 ( .A1(n9204), .A2(n5783), .ZN(n5644) );
  INV_X1 U7012 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U7013 ( .A1(n5017), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7014 ( .A1(n4641), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5640) );
  OAI211_X1 U7015 ( .C1(n5100), .C2(n10068), .A(n5641), .B(n5640), .ZN(n5642)
         );
  INV_X1 U7016 ( .A(n5642), .ZN(n5643) );
  NAND2_X1 U7017 ( .A1(n5644), .A2(n5643), .ZN(n9219) );
  NAND2_X1 U7018 ( .A1(n9219), .A2(n5167), .ZN(n5645) );
  NAND2_X1 U7019 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  AND2_X1 U7020 ( .A1(n9219), .A2(n5743), .ZN(n5648) );
  AOI21_X1 U7021 ( .B1(n9331), .B2(n5167), .A(n5648), .ZN(n8922) );
  AND2_X1 U7022 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  NAND2_X1 U7023 ( .A1(n5652), .A2(n5651), .ZN(n5654) );
  INV_X1 U7024 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7343) );
  INV_X1 U7025 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7864) );
  MUX2_X1 U7026 ( .A(n7343), .B(n7864), .S(n5497), .Z(n5677) );
  XNOR2_X1 U7027 ( .A(n5677), .B(SI_24_), .ZN(n5676) );
  XNOR2_X1 U7028 ( .A(n5675), .B(n5676), .ZN(n7342) );
  NAND2_X1 U7029 ( .A1(n7342), .A2(n5306), .ZN(n5656) );
  NAND2_X1 U7030 ( .A1(n5732), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7031 ( .A1(n9324), .A2(n7878), .ZN(n5667) );
  INV_X1 U7032 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7033 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  NAND2_X1 U7034 ( .A1(n5686), .A2(n5659), .ZN(n9190) );
  OR2_X1 U7035 ( .A1(n9190), .A2(n5783), .ZN(n5665) );
  INV_X1 U7036 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7037 ( .A1(n8168), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7038 ( .A1(n5017), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5660) );
  OAI211_X1 U7039 ( .C1(n8172), .C2(n5662), .A(n5661), .B(n5660), .ZN(n5663)
         );
  INV_X1 U7040 ( .A(n5663), .ZN(n5664) );
  INV_X1 U7041 ( .A(n9202), .ZN(n9173) );
  NAND2_X1 U7042 ( .A1(n9173), .A2(n5167), .ZN(n5666) );
  NAND2_X1 U7043 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  XNOR2_X1 U7044 ( .A(n5668), .B(n7881), .ZN(n5671) );
  NOR2_X1 U7045 ( .A1(n9202), .A2(n7884), .ZN(n5669) );
  AOI21_X1 U7046 ( .B1(n9324), .B2(n5167), .A(n5669), .ZN(n5670) );
  NAND2_X1 U7047 ( .A1(n5671), .A2(n5670), .ZN(n5673) );
  OR2_X1 U7048 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  NAND2_X1 U7049 ( .A1(n5673), .A2(n5672), .ZN(n8957) );
  INV_X1 U7050 ( .A(n5673), .ZN(n5674) );
  INV_X1 U7051 ( .A(n5677), .ZN(n5678) );
  NAND2_X1 U7052 ( .A1(n5678), .A2(SI_24_), .ZN(n5679) );
  INV_X1 U7053 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7413) );
  INV_X1 U7054 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7410) );
  MUX2_X1 U7055 ( .A(n7413), .B(n7410), .S(n5497), .Z(n5681) );
  INV_X1 U7056 ( .A(SI_25_), .ZN(n5680) );
  NAND2_X1 U7057 ( .A1(n5681), .A2(n5680), .ZN(n5698) );
  INV_X1 U7058 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U7059 ( .A1(n5682), .A2(SI_25_), .ZN(n5683) );
  NAND2_X1 U7060 ( .A1(n5698), .A2(n5683), .ZN(n5696) );
  XNOR2_X1 U7061 ( .A(n5697), .B(n5696), .ZN(n7408) );
  NAND2_X1 U7062 ( .A1(n7408), .A2(n5306), .ZN(n5685) );
  NAND2_X1 U7063 ( .A1(n5732), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5684) );
  INV_X1 U7064 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U7065 ( .A1(n5686), .A2(n8951), .ZN(n5687) );
  INV_X1 U7066 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U7067 ( .A1(n5017), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7068 ( .A1(n8168), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5688) );
  OAI211_X1 U7069 ( .C1(n8172), .C2(n5690), .A(n5689), .B(n5688), .ZN(n5691)
         );
  AOI22_X1 U7070 ( .A1(n9317), .A2(n7878), .B1(n5167), .B2(n9185), .ZN(n5692)
         );
  XNOR2_X1 U7071 ( .A(n5692), .B(n6944), .ZN(n5695) );
  NOR2_X1 U7072 ( .A1(n9006), .A2(n7884), .ZN(n5693) );
  AOI21_X1 U7073 ( .B1(n9317), .B2(n5167), .A(n5693), .ZN(n5694) );
  XNOR2_X1 U7074 ( .A(n5695), .B(n5694), .ZN(n8949) );
  INV_X1 U7075 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7538) );
  INV_X1 U7076 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9934) );
  MUX2_X1 U7077 ( .A(n7538), .B(n9934), .S(n5497), .Z(n5700) );
  INV_X1 U7078 ( .A(SI_26_), .ZN(n5699) );
  NAND2_X1 U7079 ( .A1(n5700), .A2(n5699), .ZN(n5722) );
  INV_X1 U7080 ( .A(n5700), .ZN(n5701) );
  NAND2_X1 U7081 ( .A1(n5701), .A2(SI_26_), .ZN(n5702) );
  AND2_X1 U7082 ( .A1(n5722), .A2(n5702), .ZN(n5720) );
  NAND2_X1 U7083 ( .A1(n7536), .A2(n5306), .ZN(n5704) );
  NAND2_X1 U7084 ( .A1(n5732), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5703) );
  AND2_X2 U7085 ( .A1(n5704), .A2(n5703), .ZN(n9160) );
  INV_X1 U7086 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7087 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  NAND2_X1 U7088 ( .A1(n5781), .A2(n5708), .ZN(n9159) );
  INV_X1 U7089 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7090 ( .A1(n8168), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7091 ( .A1(n5017), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5709) );
  OAI211_X1 U7092 ( .C1(n8172), .C2(n5711), .A(n5710), .B(n5709), .ZN(n5712)
         );
  INV_X1 U7093 ( .A(n5712), .ZN(n5713) );
  OAI22_X1 U7094 ( .A1(n9160), .A2(n5741), .B1(n9089), .B2(n5740), .ZN(n5715)
         );
  XNOR2_X1 U7095 ( .A(n5715), .B(n6944), .ZN(n5719) );
  OR2_X1 U7096 ( .A1(n9160), .A2(n5740), .ZN(n5717) );
  NAND2_X1 U7097 ( .A1(n9174), .A2(n5743), .ZN(n5716) );
  NAND2_X1 U7098 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  XNOR2_X1 U7099 ( .A(n5719), .B(n5718), .ZN(n8998) );
  NAND2_X1 U7100 ( .A1(n5721), .A2(n5720), .ZN(n5723) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5724) );
  INV_X1 U7102 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9923) );
  MUX2_X1 U7103 ( .A(n5724), .B(n9923), .S(n5497), .Z(n5726) );
  INV_X1 U7104 ( .A(SI_27_), .ZN(n5725) );
  NAND2_X1 U7105 ( .A1(n5726), .A2(n5725), .ZN(n6218) );
  INV_X1 U7106 ( .A(n5726), .ZN(n5727) );
  NAND2_X1 U7107 ( .A1(n5727), .A2(SI_27_), .ZN(n5728) );
  AND2_X1 U7108 ( .A1(n6218), .A2(n5728), .ZN(n5729) );
  NAND2_X1 U7109 ( .A1(n5732), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5733) );
  XNOR2_X1 U7110 ( .A(n5781), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U7111 ( .A1(n9142), .A2(n6983), .ZN(n5739) );
  INV_X1 U7112 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U7113 ( .A1(n4641), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7114 ( .A1(n8168), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5735) );
  OAI211_X1 U7115 ( .C1(n10063), .C2(n5104), .A(n5736), .B(n5735), .ZN(n5737)
         );
  INV_X1 U7116 ( .A(n5737), .ZN(n5738) );
  OAI22_X1 U7117 ( .A1(n9144), .A2(n5741), .B1(n9128), .B2(n5740), .ZN(n5742)
         );
  XOR2_X1 U7118 ( .A(n6944), .B(n5742), .Z(n5745) );
  AOI22_X1 U7119 ( .A1(n9306), .A2(n5167), .B1(n5743), .B2(n9157), .ZN(n5744)
         );
  NAND2_X1 U7120 ( .A1(n5745), .A2(n5744), .ZN(n7891) );
  OAI21_X1 U7121 ( .B1(n5745), .B2(n5744), .A(n7891), .ZN(n5746) );
  NAND2_X1 U7122 ( .A1(n7409), .A2(P1_B_REG_SCAN_IN), .ZN(n5748) );
  MUX2_X1 U7123 ( .A(P1_B_REG_SCAN_IN), .B(n5748), .S(n7866), .Z(n5749) );
  AND2_X1 U7124 ( .A1(n5749), .A2(n5750), .ZN(n9632) );
  INV_X1 U7125 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U7126 ( .A1(n9632), .A2(n10011), .ZN(n5752) );
  INV_X1 U7127 ( .A(n5750), .ZN(n7537) );
  NAND2_X1 U7128 ( .A1(n7537), .A2(n7409), .ZN(n5751) );
  NAND2_X1 U7129 ( .A1(n5752), .A2(n5751), .ZN(n6899) );
  INV_X1 U7130 ( .A(n6899), .ZN(n6356) );
  INV_X1 U7131 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7132 ( .A1(n9632), .A2(n5753), .ZN(n5755) );
  NAND2_X1 U7133 ( .A1(n7537), .A2(n7866), .ZN(n5754) );
  NAND2_X1 U7134 ( .A1(n5755), .A2(n5754), .ZN(n6898) );
  INV_X1 U7135 ( .A(n6898), .ZN(n9395) );
  NOR4_X1 U7136 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5764) );
  NOR4_X1 U7137 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5763) );
  INV_X1 U7138 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10105) );
  INV_X1 U7139 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9916) );
  INV_X1 U7140 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9914) );
  INV_X1 U7141 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9921) );
  NAND4_X1 U7142 ( .A1(n10105), .A2(n9916), .A3(n9914), .A4(n9921), .ZN(n5761)
         );
  NOR4_X1 U7143 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5759) );
  NOR4_X1 U7144 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5758) );
  NOR4_X1 U7145 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5757) );
  NOR4_X1 U7146 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5756) );
  NAND4_X1 U7147 ( .A1(n5759), .A2(n5758), .A3(n5757), .A4(n5756), .ZN(n5760)
         );
  NOR4_X1 U7148 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5761), .A4(n5760), .ZN(n5762) );
  NAND3_X1 U7149 ( .A1(n5764), .A2(n5763), .A3(n5762), .ZN(n5765) );
  NAND2_X1 U7150 ( .A1(n9632), .A2(n5765), .ZN(n6896) );
  NAND3_X1 U7151 ( .A1(n6356), .A2(n9395), .A3(n6896), .ZN(n5791) );
  INV_X1 U7152 ( .A(n5766), .ZN(n8267) );
  INV_X1 U7153 ( .A(n5773), .ZN(n5767) );
  NAND2_X1 U7154 ( .A1(n5768), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5770) );
  XNOR2_X1 U7155 ( .A(n5770), .B(n5769), .ZN(n7212) );
  AND2_X1 U7156 ( .A1(n7212), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5771) );
  AND2_X1 U7157 ( .A1(n6304), .A2(n5771), .ZN(n9633) );
  NAND2_X1 U7158 ( .A1(n8445), .A2(n5766), .ZN(n6887) );
  NAND3_X1 U7159 ( .A1(n9686), .A2(n9633), .A3(n6887), .ZN(n5772) );
  INV_X1 U7160 ( .A(n9446), .ZN(n9002) );
  OAI21_X1 U7161 ( .B1(n7897), .B2(n4426), .A(n9002), .ZN(n5800) );
  OR2_X1 U7162 ( .A1(n6887), .A2(n5773), .ZN(n5794) );
  AND3_X1 U7163 ( .A1(n5794), .A2(n7212), .A3(n6304), .ZN(n5774) );
  NAND2_X1 U7164 ( .A1(n5791), .A2(n9686), .ZN(n5795) );
  NAND2_X1 U7165 ( .A1(n5774), .A2(n5795), .ZN(n5775) );
  NAND2_X1 U7166 ( .A1(n5775), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5776) );
  INV_X1 U7167 ( .A(n7020), .ZN(n8436) );
  AND2_X1 U7168 ( .A1(n6439), .A2(n8436), .ZN(n6901) );
  NAND2_X1 U7169 ( .A1(n5791), .A2(n4960), .ZN(n5796) );
  AND2_X1 U7170 ( .A1(n5776), .A2(n5796), .ZN(n9452) );
  INV_X1 U7171 ( .A(n9452), .ZN(n9003) );
  OR2_X1 U7172 ( .A1(n6893), .A2(n6880), .ZN(n6945) );
  INV_X1 U7173 ( .A(n6945), .ZN(n6440) );
  NAND2_X1 U7174 ( .A1(n6440), .A2(n9633), .ZN(n5789) );
  NOR2_X1 U7175 ( .A1(n5789), .A2(n5777), .ZN(n8448) );
  INV_X1 U7176 ( .A(n8448), .ZN(n5778) );
  OR2_X1 U7177 ( .A1(n5791), .A2(n5778), .ZN(n9435) );
  INV_X1 U7178 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5780) );
  OAI22_X1 U7179 ( .A1(n9089), .A2(n9435), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5780), .ZN(n5793) );
  INV_X1 U7180 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5779) );
  OAI21_X1 U7181 ( .B1(n5781), .B2(n5780), .A(n5779), .ZN(n5782) );
  NAND2_X1 U7182 ( .A1(n5782), .A2(n9116), .ZN(n7888) );
  INV_X1 U7183 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U7184 ( .A1(n5017), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7185 ( .A1(n8168), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5784) );
  OAI211_X1 U7186 ( .C1(n8172), .C2(n9906), .A(n5785), .B(n5784), .ZN(n5786)
         );
  INV_X1 U7187 ( .A(n5786), .ZN(n5787) );
  INV_X1 U7188 ( .A(n5777), .ZN(n9500) );
  OR2_X1 U7189 ( .A1(n5789), .A2(n9500), .ZN(n5790) );
  OR2_X1 U7190 ( .A1(n5791), .A2(n5790), .ZN(n8983) );
  NOR2_X1 U7191 ( .A1(n9092), .A2(n8983), .ZN(n5792) );
  AOI211_X1 U7192 ( .C1(n9142), .C2(n9003), .A(n5793), .B(n5792), .ZN(n5799)
         );
  AND2_X1 U7193 ( .A1(n9633), .A2(n5794), .ZN(n6897) );
  NAND3_X1 U7194 ( .A1(n5796), .A2(n5795), .A3(n6897), .ZN(n9445) );
  OR2_X1 U7195 ( .A1(n9445), .A2(n9686), .ZN(n9010) );
  NAND3_X1 U7196 ( .A1(n5800), .A2(n5799), .A3(n5798), .ZN(P1_U3212) );
  NOR2_X1 U7197 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5802) );
  NOR2_X1 U7198 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5808) );
  NOR2_X1 U7199 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5807) );
  NOR2_X1 U7200 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5806) );
  NOR2_X1 U7201 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5805) );
  NAND4_X1 U7202 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), .ZN(n5809)
         );
  INV_X1 U7203 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5810) );
  INV_X1 U7204 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7205 ( .A1(n5812), .A2(n5811), .ZN(n5843) );
  NAND2_X1 U7206 ( .A1(n5843), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5813) );
  MUX2_X1 U7207 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5813), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5815) );
  INV_X1 U7208 ( .A(n5845), .ZN(n5814) );
  NAND2_X1 U7209 ( .A1(n5814), .A2(n4954), .ZN(n5816) );
  INV_X1 U7210 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U7211 ( .A1(n5895), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5823) );
  INV_X1 U7212 ( .A(n8479), .ZN(n5819) );
  AND2_X2 U7213 ( .A1(n5818), .A2(n5819), .ZN(n5893) );
  NAND2_X1 U7214 ( .A1(n5893), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7215 ( .A1(n5896), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5821) );
  AND2_X2 U7216 ( .A1(n7933), .A2(n8479), .ZN(n5897) );
  NAND2_X1 U7217 ( .A1(n5897), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5820) );
  INV_X1 U7218 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5824) );
  INV_X1 U7219 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5826) );
  INV_X1 U7220 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5832) );
  INV_X1 U7221 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U7222 ( .A1(n5829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5831) );
  INV_X1 U7223 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7224 ( .A1(n6552), .A2(n7970), .ZN(n5839) );
  INV_X1 U7225 ( .A(n5839), .ZN(n6265) );
  NAND2_X1 U7226 ( .A1(n4413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5833) );
  AND2_X2 U7227 ( .A1(n6265), .A2(n7021), .ZN(n6266) );
  NAND2_X1 U7228 ( .A1(n5835), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5836) );
  MUX2_X1 U7229 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5836), .S(
        P2_IR_REG_19__SCAN_IN), .Z(n5837) );
  INV_X1 U7230 ( .A(n7969), .ZN(n5838) );
  INV_X1 U7231 ( .A(n5853), .ZN(n5851) );
  NAND3_X1 U7232 ( .A1(n6550), .A2(n5839), .A3(n7970), .ZN(n5840) );
  INV_X1 U7233 ( .A(n7970), .ZN(n8152) );
  NAND2_X1 U7234 ( .A1(n8152), .A2(n7021), .ZN(n7200) );
  NAND2_X1 U7235 ( .A1(n5845), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5841) );
  INV_X1 U7236 ( .A(n5844), .ZN(n6244) );
  NAND2_X2 U7237 ( .A1(n5860), .A2(n5497), .ZN(n7960) );
  INV_X1 U7238 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U7239 ( .A1(n5921), .A2(n6598), .ZN(n5849) );
  INV_X1 U7240 ( .A(n5846), .ZN(n7826) );
  INV_X1 U7241 ( .A(n6366), .ZN(n5847) );
  INV_X1 U7242 ( .A(n5852), .ZN(n5850) );
  NAND2_X1 U7243 ( .A1(n5851), .A2(n5850), .ZN(n6759) );
  NAND2_X1 U7244 ( .A1(n5853), .A2(n5852), .ZN(n5854) );
  NAND2_X1 U7245 ( .A1(n5895), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7246 ( .A1(n5893), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7247 ( .A1(n5896), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7248 ( .A1(n5897), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7249 ( .A1(n7833), .A2(SI_0_), .ZN(n5859) );
  XNOR2_X1 U7250 ( .A(n5859), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8920) );
  MUX2_X1 U7251 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8920), .S(n6575), .Z(n7208) );
  NAND2_X1 U7252 ( .A1(n6751), .A2(n7208), .ZN(n6559) );
  INV_X1 U7253 ( .A(n6559), .ZN(n5862) );
  NOR2_X1 U7254 ( .A1(n6186), .A2(n7208), .ZN(n5861) );
  NAND2_X1 U7255 ( .A1(n6754), .A2(n6753), .ZN(n6752) );
  NAND2_X1 U7256 ( .A1(n5893), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7257 ( .A1(n5895), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U7258 ( .A1(n5896), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7259 ( .A1(n5897), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5863) );
  INV_X1 U7260 ( .A(n5886), .ZN(n5873) );
  OR2_X1 U7261 ( .A1(n5867), .A2(n6238), .ZN(n5868) );
  XNOR2_X2 U7262 ( .A(n5868), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U7263 ( .A1(n5921), .A2(n9419), .ZN(n5870) );
  OR2_X1 U7264 ( .A1(n5908), .A2(n6361), .ZN(n5869) );
  XNOR2_X1 U7265 ( .A(n5871), .B(n6765), .ZN(n5885) );
  INV_X1 U7266 ( .A(n5885), .ZN(n5872) );
  NAND2_X1 U7267 ( .A1(n5873), .A2(n5872), .ZN(n6760) );
  NAND2_X1 U7268 ( .A1(n6752), .A2(n5874), .ZN(n6348) );
  INV_X1 U7269 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7270 ( .A1(n5893), .A2(n5875), .ZN(n5879) );
  NAND2_X1 U7271 ( .A1(n5895), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7272 ( .A1(n5896), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7273 ( .A1(n5897), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5876) );
  OR2_X1 U7274 ( .A1(n7348), .A2(n6741), .ZN(n5888) );
  INV_X1 U7275 ( .A(n5888), .ZN(n5884) );
  NAND2_X1 U7276 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4417), .ZN(n5880) );
  XNOR2_X1 U7277 ( .A(n5880), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6601) );
  INV_X1 U7278 ( .A(n6601), .ZN(n6681) );
  OR2_X1 U7279 ( .A1(n5908), .A2(n7869), .ZN(n5882) );
  INV_X1 U7280 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9968) );
  XNOR2_X1 U7281 ( .A(n7336), .B(n6186), .ZN(n5889) );
  INV_X1 U7282 ( .A(n5889), .ZN(n5883) );
  NAND2_X1 U7283 ( .A1(n5884), .A2(n5883), .ZN(n5890) );
  NAND2_X1 U7284 ( .A1(n5886), .A2(n5885), .ZN(n6761) );
  AND2_X1 U7285 ( .A1(n5890), .A2(n6761), .ZN(n5887) );
  XNOR2_X1 U7286 ( .A(n5889), .B(n5888), .ZN(n6350) );
  NOR2_X2 U7287 ( .A1(n5892), .A2(n5891), .ZN(n6826) );
  BUF_X4 U7288 ( .A(n5893), .Z(n6285) );
  INV_X1 U7289 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5894) );
  XNOR2_X1 U7290 ( .A(n5894), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n7359) );
  NAND2_X1 U7291 ( .A1(n6285), .A2(n7359), .ZN(n5901) );
  NAND2_X1 U7292 ( .A1(n5895), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7293 ( .A1(n5896), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7294 ( .A1(n6286), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5898) );
  OR2_X1 U7295 ( .A1(n5910), .A2(n6238), .ZN(n5902) );
  XNOR2_X1 U7296 ( .A(n5902), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7297 ( .A1(n5921), .A2(n6603), .ZN(n5904) );
  OR2_X1 U7298 ( .A1(n5908), .A2(n7874), .ZN(n5903) );
  OAI211_X1 U7299 ( .C1(n7960), .C2(n6375), .A(n5904), .B(n5903), .ZN(n7358)
         );
  XNOR2_X1 U7300 ( .A(n6231), .B(n7358), .ZN(n5905) );
  NOR2_X1 U7301 ( .A1(n5906), .A2(n5905), .ZN(n6824) );
  NAND2_X1 U7302 ( .A1(n5906), .A2(n5905), .ZN(n6823) );
  INV_X4 U7303 ( .A(n5908), .ZN(n7962) );
  NAND2_X1 U7304 ( .A1(n5907), .A2(n7962), .ZN(n5915) );
  NAND2_X1 U7305 ( .A1(n5910), .A2(n5909), .ZN(n5912) );
  NAND2_X1 U7306 ( .A1(n5912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  MUX2_X1 U7307 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5911), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5913) );
  AND2_X1 U7308 ( .A1(n5913), .A2(n5943), .ZN(n6604) );
  AOI22_X1 U7309 ( .A1(n7948), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5921), .B2(
        n6604), .ZN(n5914) );
  XNOR2_X1 U7310 ( .A(n9799), .B(n6186), .ZN(n5933) );
  AOI21_X1 U7311 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5916) );
  NOR2_X1 U7312 ( .A1(n5916), .A2(n5925), .ZN(n7301) );
  NAND2_X1 U7313 ( .A1(n6285), .A2(n7301), .ZN(n5920) );
  NAND2_X1 U7314 ( .A1(n5895), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5919) );
  INV_X2 U7315 ( .A(n7956), .ZN(n6286) );
  NAND2_X1 U7316 ( .A1(n6286), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7317 ( .A1(n5896), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5917) );
  OR2_X1 U7318 ( .A1(n6816), .A2(n6741), .ZN(n5932) );
  XNOR2_X1 U7319 ( .A(n5933), .B(n5932), .ZN(n6808) );
  NAND2_X1 U7320 ( .A1(n6358), .A2(n7962), .ZN(n5924) );
  NAND2_X1 U7321 ( .A1(n5943), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7322 ( .A(n5922), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8571) );
  AOI22_X1 U7323 ( .A1(n7948), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5921), .B2(
        n8571), .ZN(n5923) );
  AND2_X2 U7324 ( .A1(n5924), .A2(n5923), .ZN(n9806) );
  XNOR2_X1 U7325 ( .A(n9806), .B(n6186), .ZN(n5936) );
  NAND2_X1 U7326 ( .A1(n5925), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5962) );
  OAI21_X1 U7327 ( .B1(n5925), .B2(P2_REG3_REG_6__SCAN_IN), .A(n5962), .ZN(
        n8816) );
  INV_X1 U7328 ( .A(n8816), .ZN(n5926) );
  NAND2_X1 U7329 ( .A1(n6285), .A2(n5926), .ZN(n5930) );
  NAND2_X1 U7330 ( .A1(n5895), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7331 ( .A1(n5897), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7332 ( .A1(n5896), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7333 ( .A1(n8565), .A2(n7969), .ZN(n5937) );
  NAND2_X1 U7334 ( .A1(n5936), .A2(n5937), .ZN(n5941) );
  INV_X1 U7335 ( .A(n5941), .ZN(n5931) );
  INV_X1 U7336 ( .A(n5932), .ZN(n5935) );
  INV_X1 U7337 ( .A(n5933), .ZN(n5934) );
  AND2_X1 U7338 ( .A1(n5935), .A2(n5934), .ZN(n6810) );
  INV_X1 U7339 ( .A(n5936), .ZN(n5939) );
  INV_X1 U7340 ( .A(n5937), .ZN(n5938) );
  NAND2_X1 U7341 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  AND2_X1 U7342 ( .A1(n5941), .A2(n6811), .ZN(n5942) );
  NAND2_X1 U7343 ( .A1(n6367), .A2(n7962), .ZN(n5946) );
  NOR2_X1 U7344 ( .A1(n5943), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5954) );
  OR2_X1 U7345 ( .A1(n5954), .A2(n6238), .ZN(n5944) );
  XNOR2_X1 U7346 ( .A(n5944), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6735) );
  AOI22_X1 U7347 ( .A1(n7948), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5921), .B2(
        n6735), .ZN(n5945) );
  NAND2_X1 U7348 ( .A1(n5946), .A2(n5945), .ZN(n9810) );
  XNOR2_X1 U7349 ( .A(n9810), .B(n6186), .ZN(n5951) );
  XNOR2_X1 U7350 ( .A(n5962), .B(P2_REG3_REG_7__SCAN_IN), .ZN(n7387) );
  NAND2_X1 U7351 ( .A1(n6285), .A2(n7387), .ZN(n5950) );
  NAND2_X1 U7352 ( .A1(n5895), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7353 ( .A1(n5896), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7354 ( .A1(n6286), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5947) );
  NOR2_X1 U7355 ( .A1(n9764), .A2(n6230), .ZN(n5952) );
  XNOR2_X1 U7356 ( .A(n5951), .B(n5952), .ZN(n6871) );
  NAND2_X1 U7357 ( .A1(n6376), .A2(n7962), .ZN(n5959) );
  NAND2_X1 U7358 ( .A1(n5954), .A2(n5953), .ZN(n5956) );
  NAND2_X1 U7359 ( .A1(n5956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5955) );
  MUX2_X1 U7360 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5955), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5957) );
  AND2_X1 U7361 ( .A1(n5957), .A2(n5982), .ZN(n8587) );
  AOI22_X1 U7362 ( .A1(n7948), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5921), .B2(
        n8587), .ZN(n5958) );
  NAND2_X1 U7363 ( .A1(n5959), .A2(n5958), .ZN(n9770) );
  XNOR2_X1 U7364 ( .A(n9770), .B(n6231), .ZN(n5968) );
  INV_X1 U7365 ( .A(n5962), .ZN(n5960) );
  AOI21_X1 U7366 ( .B1(n5960), .B2(P2_REG3_REG_7__SCAN_IN), .A(
        P2_REG3_REG_8__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7367 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n5961) );
  NOR2_X1 U7368 ( .A1(n5962), .A2(n5961), .ZN(n5976) );
  OR2_X1 U7369 ( .A1(n5963), .A2(n5976), .ZN(n6803) );
  INV_X1 U7370 ( .A(n6803), .ZN(n9772) );
  NAND2_X1 U7371 ( .A1(n6285), .A2(n9772), .ZN(n5967) );
  NAND2_X1 U7372 ( .A1(n5895), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7373 ( .A1(n5896), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7374 ( .A1(n6286), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5964) );
  NOR2_X1 U7375 ( .A1(n7384), .A2(n6230), .ZN(n5969) );
  XNOR2_X1 U7376 ( .A(n5968), .B(n5969), .ZN(n6800) );
  NAND2_X1 U7377 ( .A1(n6801), .A2(n6800), .ZN(n5972) );
  INV_X1 U7378 ( .A(n5968), .ZN(n5970) );
  NAND2_X1 U7379 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  NAND2_X1 U7380 ( .A1(n5972), .A2(n5971), .ZN(n6848) );
  NAND2_X1 U7381 ( .A1(n6380), .A2(n7962), .ZN(n5975) );
  NAND2_X1 U7382 ( .A1(n5982), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U7383 ( .A(n5973), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U7384 ( .A1(n7948), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5921), .B2(
        n6770), .ZN(n5974) );
  NAND2_X1 U7385 ( .A1(n5975), .A2(n5974), .ZN(n9823) );
  XNOR2_X1 U7386 ( .A(n9823), .B(n6186), .ZN(n6850) );
  NAND2_X1 U7387 ( .A1(n5976), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7388 ( .A1(n5976), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5977) );
  AND2_X1 U7389 ( .A1(n5998), .A2(n5977), .ZN(n7320) );
  NAND2_X1 U7390 ( .A1(n6285), .A2(n7320), .ZN(n5981) );
  NAND2_X1 U7391 ( .A1(n5895), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7392 ( .A1(n6286), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7393 ( .A1(n5896), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5978) );
  INV_X1 U7394 ( .A(n9762), .ZN(n8562) );
  NAND2_X1 U7395 ( .A1(n8562), .A2(n7969), .ZN(n6849) );
  NAND2_X1 U7396 ( .A1(n6382), .A2(n7962), .ZN(n5988) );
  NOR2_X1 U7397 ( .A1(n5982), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6012) );
  NOR2_X1 U7398 ( .A1(n6012), .A2(n6238), .ZN(n5983) );
  NAND2_X1 U7399 ( .A1(n5983), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5986) );
  INV_X1 U7400 ( .A(n5983), .ZN(n5985) );
  INV_X1 U7401 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7402 ( .A1(n5985), .A2(n5984), .ZN(n6004) );
  AND2_X1 U7403 ( .A1(n5986), .A2(n6004), .ZN(n7151) );
  AOI22_X1 U7404 ( .A1(n7948), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5921), .B2(
        n7151), .ZN(n5987) );
  XNOR2_X1 U7405 ( .A(n7434), .B(n6231), .ZN(n5994) );
  XNOR2_X1 U7406 ( .A(n5998), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n7427) );
  NAND2_X1 U7407 ( .A1(n6285), .A2(n7427), .ZN(n5992) );
  NAND2_X1 U7408 ( .A1(n5895), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7409 ( .A1(n6286), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7410 ( .A1(n5896), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7411 ( .A1(n7367), .A2(n6230), .ZN(n5993) );
  NOR2_X1 U7412 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  AOI21_X1 U7413 ( .B1(n5994), .B2(n5993), .A(n5995), .ZN(n6964) );
  INV_X1 U7414 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5997) );
  INV_X1 U7415 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5996) );
  OAI21_X1 U7416 ( .B1(n5998), .B2(n5997), .A(n5996), .ZN(n5999) );
  AND2_X1 U7417 ( .A1(n5999), .A2(n6018), .ZN(n7375) );
  NAND2_X1 U7418 ( .A1(n6285), .A2(n7375), .ZN(n6003) );
  NAND2_X1 U7419 ( .A1(n5895), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7420 ( .A1(n6286), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7421 ( .A1(n5896), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6000) );
  NOR2_X1 U7422 ( .A1(n7455), .A2(n6741), .ZN(n6009) );
  NAND2_X1 U7423 ( .A1(n6386), .A2(n7962), .ZN(n6007) );
  NAND2_X1 U7424 ( .A1(n6004), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6005) );
  XNOR2_X1 U7425 ( .A(n6005), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8596) );
  AOI22_X1 U7426 ( .A1(n7948), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5921), .B2(
        n8596), .ZN(n6006) );
  XNOR2_X1 U7427 ( .A(n7456), .B(n6186), .ZN(n6008) );
  XOR2_X1 U7428 ( .A(n6009), .B(n6008), .Z(n7122) );
  NAND2_X1 U7429 ( .A1(n7123), .A2(n7122), .ZN(n7121) );
  NAND2_X1 U7430 ( .A1(n6401), .A2(n7962), .ZN(n6017) );
  NOR2_X1 U7431 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6011) );
  NAND2_X1 U7432 ( .A1(n6012), .A2(n6011), .ZN(n6014) );
  NAND2_X1 U7433 ( .A1(n6014), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6013) );
  MUX2_X1 U7434 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6013), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n6015) );
  OR2_X1 U7435 ( .A1(n6014), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6037) );
  AND2_X1 U7436 ( .A1(n6015), .A2(n6037), .ZN(n7227) );
  AOI22_X1 U7437 ( .A1(n7948), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5921), .B2(
        n7227), .ZN(n6016) );
  XNOR2_X1 U7438 ( .A(n9732), .B(n6231), .ZN(n6025) );
  NAND2_X1 U7439 ( .A1(n5895), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6023) );
  INV_X1 U7440 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7188) );
  AND2_X1 U7441 ( .A1(n6018), .A2(n7188), .ZN(n6019) );
  NOR2_X1 U7442 ( .A1(n6045), .A2(n6019), .ZN(n9730) );
  NAND2_X1 U7443 ( .A1(n6285), .A2(n9730), .ZN(n6022) );
  NAND2_X1 U7444 ( .A1(n5896), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7445 ( .A1(n6286), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6020) );
  OR2_X1 U7446 ( .A1(n7464), .A2(n6741), .ZN(n6024) );
  NAND2_X1 U7447 ( .A1(n6025), .A2(n6024), .ZN(n7182) );
  NOR2_X1 U7448 ( .A1(n6025), .A2(n6024), .ZN(n7184) );
  NAND2_X1 U7449 ( .A1(n6449), .A2(n7962), .ZN(n6028) );
  NAND2_X1 U7450 ( .A1(n6037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6026) );
  XNOR2_X1 U7451 ( .A(n6026), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7399) );
  AOI22_X1 U7452 ( .A1(n7948), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7399), .B2(
        n5921), .ZN(n6027) );
  XNOR2_X1 U7453 ( .A(n8037), .B(n6186), .ZN(n6033) );
  INV_X1 U7454 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7217) );
  XNOR2_X1 U7455 ( .A(n6045), .B(n7217), .ZN(n7469) );
  NAND2_X1 U7456 ( .A1(n6285), .A2(n7469), .ZN(n6032) );
  NAND2_X1 U7457 ( .A1(n5895), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7458 ( .A1(n6286), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7459 ( .A1(n5896), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6029) );
  NOR2_X1 U7460 ( .A1(n7499), .A2(n6230), .ZN(n6034) );
  XNOR2_X1 U7461 ( .A(n6033), .B(n6034), .ZN(n7270) );
  INV_X1 U7462 ( .A(n6033), .ZN(n6036) );
  INV_X1 U7463 ( .A(n6034), .ZN(n6035) );
  OAI22_X2 U7464 ( .A1(n7271), .A2(n7270), .B1(n6036), .B2(n6035), .ZN(n7475)
         );
  NAND2_X1 U7465 ( .A1(n6527), .A2(n7962), .ZN(n6043) );
  OR2_X1 U7466 ( .A1(n6037), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7467 ( .A1(n6038), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6040) );
  INV_X1 U7468 ( .A(n6040), .ZN(n6039) );
  NAND2_X1 U7469 ( .A1(n6039), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n6041) );
  INV_X1 U7470 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U7471 ( .A1(n6040), .A2(n10069), .ZN(n6056) );
  AND2_X1 U7472 ( .A1(n6041), .A2(n6056), .ZN(n7596) );
  AOI22_X1 U7473 ( .A1(n7596), .A2(n5921), .B1(n7948), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6042) );
  NAND2_X2 U7474 ( .A1(n6043), .A2(n6042), .ZN(n9459) );
  XNOR2_X1 U7475 ( .A(n9459), .B(n6231), .ZN(n6053) );
  AND2_X1 U7476 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .ZN(n6044) );
  AOI21_X1 U7477 ( .B1(n6045), .B2(P2_REG3_REG_13__SCAN_IN), .A(
        P2_REG3_REG_14__SCAN_IN), .ZN(n6046) );
  OR2_X1 U7478 ( .A1(n6060), .A2(n6046), .ZN(n7505) );
  INV_X1 U7479 ( .A(n7505), .ZN(n6047) );
  NAND2_X1 U7480 ( .A1(n6285), .A2(n6047), .ZN(n6051) );
  NAND2_X1 U7481 ( .A1(n5895), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7482 ( .A1(n5896), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7483 ( .A1(n6286), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7484 ( .A1(n7642), .A2(n6230), .ZN(n6052) );
  NAND2_X1 U7485 ( .A1(n6053), .A2(n6052), .ZN(n6054) );
  OAI21_X1 U7486 ( .B1(n6053), .B2(n6052), .A(n6054), .ZN(n7476) );
  INV_X1 U7487 ( .A(n6054), .ZN(n6055) );
  NAND2_X1 U7488 ( .A1(n6641), .A2(n7962), .ZN(n6059) );
  NAND2_X1 U7489 ( .A1(n6056), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6057) );
  XNOR2_X1 U7490 ( .A(n6057), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7909) );
  AOI22_X1 U7491 ( .A1(n7909), .A2(n5921), .B1(n7948), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6058) );
  XNOR2_X1 U7492 ( .A(n7677), .B(n6231), .ZN(n7665) );
  NAND2_X1 U7493 ( .A1(n5895), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6065) );
  NOR2_X1 U7494 ( .A1(n6060), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6061) );
  NOR2_X1 U7495 ( .A1(n6072), .A2(n6061), .ZN(n7639) );
  NAND2_X1 U7496 ( .A1(n6285), .A2(n7639), .ZN(n6064) );
  NAND2_X1 U7497 ( .A1(n5896), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7498 ( .A1(n6286), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6062) );
  OR2_X1 U7499 ( .A1(n7688), .A2(n6741), .ZN(n7666) );
  NAND2_X1 U7500 ( .A1(n6737), .A2(n7962), .ZN(n6071) );
  NAND2_X1 U7501 ( .A1(n6066), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6067) );
  MUX2_X1 U7502 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6067), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6069) );
  AND2_X1 U7503 ( .A1(n6069), .A2(n6068), .ZN(n7902) );
  AOI22_X1 U7504 ( .A1(n7948), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5921), .B2(
        n7902), .ZN(n6070) );
  XNOR2_X1 U7505 ( .A(n8899), .B(n6186), .ZN(n6078) );
  OR2_X1 U7506 ( .A1(n6072), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7507 ( .A1(n6072), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6087) );
  AND2_X1 U7508 ( .A1(n6073), .A2(n6087), .ZN(n7693) );
  NAND2_X1 U7509 ( .A1(n6285), .A2(n7693), .ZN(n6077) );
  NAND2_X1 U7510 ( .A1(n5895), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7511 ( .A1(n5896), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7512 ( .A1(n6286), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6074) );
  NOR2_X1 U7513 ( .A1(n7680), .A2(n6741), .ZN(n6079) );
  NOR2_X1 U7514 ( .A1(n6078), .A2(n6079), .ZN(n7669) );
  AOI21_X1 U7515 ( .B1(n7665), .B2(n7666), .A(n7669), .ZN(n6083) );
  NOR3_X1 U7516 ( .A1(n7669), .A2(n7665), .A3(n7666), .ZN(n6082) );
  INV_X1 U7517 ( .A(n6078), .ZN(n6081) );
  INV_X1 U7518 ( .A(n6079), .ZN(n6080) );
  NOR2_X1 U7519 ( .A1(n6081), .A2(n6080), .ZN(n7668) );
  NAND2_X1 U7520 ( .A1(n6785), .A2(n7962), .ZN(n6086) );
  NAND2_X1 U7521 ( .A1(n6068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7522 ( .A(n6084), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7915) );
  AOI22_X1 U7523 ( .A1(n7948), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5921), .B2(
        n7915), .ZN(n6085) );
  XNOR2_X1 U7524 ( .A(n8895), .B(n6186), .ZN(n6092) );
  NAND2_X1 U7525 ( .A1(n5895), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6091) );
  INV_X1 U7526 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10004) );
  NOR2_X1 U7527 ( .A1(n10004), .A2(n6087), .ZN(n6100) );
  AOI21_X1 U7528 ( .B1(n10004), .B2(n6087), .A(n6100), .ZN(n7718) );
  NAND2_X1 U7529 ( .A1(n6285), .A2(n7718), .ZN(n6090) );
  NAND2_X1 U7530 ( .A1(n5896), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7531 ( .A1(n6286), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6088) );
  AND4_X1 U7532 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n7708)
         );
  NOR2_X1 U7533 ( .A1(n7708), .A2(n6230), .ZN(n6093) );
  XNOR2_X1 U7534 ( .A(n6092), .B(n6093), .ZN(n7572) );
  INV_X1 U7535 ( .A(n6092), .ZN(n6095) );
  INV_X1 U7536 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7537 ( .A1(n6844), .A2(n7962), .ZN(n6099) );
  NAND2_X1 U7538 ( .A1(n6096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6097) );
  XNOR2_X1 U7539 ( .A(n6097), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8640) );
  AOI22_X1 U7540 ( .A1(n7948), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5921), .B2(
        n8640), .ZN(n6098) );
  XNOR2_X1 U7541 ( .A(n7847), .B(n6186), .ZN(n6105) );
  NAND2_X1 U7542 ( .A1(n5895), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7543 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n6100), .ZN(n6109) );
  OAI21_X1 U7544 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n6100), .A(n6109), .ZN(
        n7620) );
  INV_X1 U7545 ( .A(n7620), .ZN(n7811) );
  NAND2_X1 U7546 ( .A1(n6285), .A2(n7811), .ZN(n6103) );
  NAND2_X1 U7547 ( .A1(n5896), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7548 ( .A1(n6286), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6101) );
  AND4_X1 U7549 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n7846)
         );
  NOR2_X1 U7550 ( .A1(n7846), .A2(n6741), .ZN(n6107) );
  XNOR2_X1 U7551 ( .A(n6105), .B(n6107), .ZN(n7617) );
  INV_X1 U7552 ( .A(n6105), .ZN(n6106) );
  INV_X1 U7553 ( .A(n6109), .ZN(n6108) );
  NAND2_X1 U7554 ( .A1(n6108), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6124) );
  INV_X1 U7555 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U7556 ( .A1(n6109), .A2(n9948), .ZN(n6110) );
  AND2_X1 U7557 ( .A1(n6124), .A2(n6110), .ZN(n7857) );
  NAND2_X1 U7558 ( .A1(n6285), .A2(n7857), .ZN(n6114) );
  NAND2_X1 U7559 ( .A1(n5895), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7560 ( .A1(n5896), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7561 ( .A1(n5897), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6111) );
  NAND4_X1 U7562 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n8552)
         );
  AND2_X1 U7563 ( .A1(n8552), .A2(n7969), .ZN(n6118) );
  NAND2_X1 U7564 ( .A1(n6908), .A2(n7962), .ZN(n6116) );
  AOI22_X1 U7565 ( .A1(n7948), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5921), .B2(
        n7966), .ZN(n6115) );
  XNOR2_X1 U7566 ( .A(n8884), .B(n6186), .ZN(n6117) );
  NOR2_X1 U7567 ( .A1(n6117), .A2(n6118), .ZN(n6119) );
  AOI21_X1 U7568 ( .B1(n6118), .B2(n6117), .A(n6119), .ZN(n7725) );
  NAND2_X1 U7569 ( .A1(n7726), .A2(n7725), .ZN(n7724) );
  INV_X1 U7570 ( .A(n6119), .ZN(n6120) );
  NAND2_X1 U7571 ( .A1(n7724), .A2(n6120), .ZN(n7770) );
  NAND2_X1 U7572 ( .A1(n7018), .A2(n7962), .ZN(n6122) );
  NAND2_X1 U7573 ( .A1(n7948), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U7574 ( .A(n8878), .B(n6186), .ZN(n6130) );
  INV_X1 U7575 ( .A(n6124), .ZN(n6123) );
  NAND2_X1 U7576 ( .A1(n6123), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6137) );
  INV_X1 U7577 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U7578 ( .A1(n6124), .A2(n7771), .ZN(n6125) );
  AND2_X1 U7579 ( .A1(n6137), .A2(n6125), .ZN(n8792) );
  NAND2_X1 U7580 ( .A1(n6285), .A2(n8792), .ZN(n6129) );
  NAND2_X1 U7581 ( .A1(n5895), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7582 ( .A1(n5896), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7583 ( .A1(n5897), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6126) );
  AND4_X1 U7584 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), .ZN(n8456)
         );
  NOR2_X1 U7585 ( .A1(n8456), .A2(n6230), .ZN(n6131) );
  XNOR2_X1 U7586 ( .A(n6130), .B(n6131), .ZN(n7769) );
  INV_X1 U7587 ( .A(n6130), .ZN(n6133) );
  INV_X1 U7588 ( .A(n6131), .ZN(n6132) );
  NAND2_X1 U7589 ( .A1(n7147), .A2(n7962), .ZN(n6135) );
  NAND2_X1 U7590 ( .A1(n7948), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6134) );
  XNOR2_X1 U7591 ( .A(n8778), .B(n6186), .ZN(n6143) );
  INV_X1 U7592 ( .A(n6137), .ZN(n6136) );
  NAND2_X1 U7593 ( .A1(n6136), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6162) );
  INV_X1 U7594 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U7595 ( .A1(n6137), .A2(n7779), .ZN(n6138) );
  AND2_X1 U7596 ( .A1(n6162), .A2(n6138), .ZN(n8776) );
  NAND2_X1 U7597 ( .A1(n6285), .A2(n8776), .ZN(n6142) );
  NAND2_X1 U7598 ( .A1(n5895), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7599 ( .A1(n6286), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7600 ( .A1(n5896), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6139) );
  NOR2_X1 U7601 ( .A1(n8799), .A2(n6741), .ZN(n6144) );
  XNOR2_X1 U7602 ( .A(n6143), .B(n6144), .ZN(n7778) );
  INV_X1 U7603 ( .A(n6143), .ZN(n6145) );
  NAND2_X1 U7604 ( .A1(n7215), .A2(n7962), .ZN(n6147) );
  NAND2_X1 U7605 ( .A1(n7948), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6146) );
  XNOR2_X1 U7606 ( .A(n8868), .B(n6186), .ZN(n6153) );
  NAND2_X1 U7607 ( .A1(n5895), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6152) );
  XNOR2_X1 U7608 ( .A(n6162), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U7609 ( .A1(n6285), .A2(n8761), .ZN(n6151) );
  NAND2_X1 U7610 ( .A1(n5896), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7611 ( .A1(n5897), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6149) );
  AND4_X1 U7612 ( .A1(n6152), .A2(n6151), .A3(n6150), .A4(n6149), .ZN(n8493)
         );
  INV_X1 U7613 ( .A(n8493), .ZN(n8782) );
  NAND2_X1 U7614 ( .A1(n8782), .A2(n7969), .ZN(n8525) );
  NAND2_X1 U7615 ( .A1(n8526), .A2(n8525), .ZN(n8524) );
  NAND2_X1 U7616 ( .A1(n8524), .A2(n6155), .ZN(n6169) );
  NAND2_X1 U7617 ( .A1(n7235), .A2(n7962), .ZN(n6157) );
  NAND2_X1 U7618 ( .A1(n7948), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6156) );
  XNOR2_X1 U7619 ( .A(n8748), .B(n6186), .ZN(n6168) );
  NOR2_X1 U7620 ( .A1(n6169), .A2(n6168), .ZN(n8488) );
  INV_X1 U7621 ( .A(n6162), .ZN(n6159) );
  AND2_X1 U7622 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6158) );
  NAND2_X1 U7623 ( .A1(n6159), .A2(n6158), .ZN(n6173) );
  INV_X1 U7624 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6161) );
  INV_X1 U7625 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6160) );
  OAI21_X1 U7626 ( .B1(n6162), .B2(n6161), .A(n6160), .ZN(n6163) );
  AND2_X1 U7627 ( .A1(n6173), .A2(n6163), .ZN(n8754) );
  NAND2_X1 U7628 ( .A1(n6285), .A2(n8754), .ZN(n6167) );
  NAND2_X1 U7629 ( .A1(n5895), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7630 ( .A1(n5897), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7631 ( .A1(n5896), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U7632 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n8737)
         );
  INV_X1 U7633 ( .A(n8737), .ZN(n8768) );
  NAND2_X1 U7634 ( .A1(n6169), .A2(n6168), .ZN(n8489) );
  OAI21_X2 U7635 ( .B1(n8488), .B2(n8491), .A(n8489), .ZN(n6179) );
  NAND2_X1 U7636 ( .A1(n7342), .A2(n7962), .ZN(n6171) );
  NAND2_X1 U7637 ( .A1(n7948), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6170) );
  XNOR2_X1 U7638 ( .A(n8858), .B(n6231), .ZN(n6180) );
  XNOR2_X1 U7639 ( .A(n6179), .B(n6180), .ZN(n8511) );
  INV_X1 U7640 ( .A(n6173), .ZN(n6172) );
  NAND2_X1 U7641 ( .A1(n6172), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6195) );
  INV_X1 U7642 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U7643 ( .A1(n6173), .A2(n8513), .ZN(n6174) );
  AND2_X1 U7644 ( .A1(n6195), .A2(n6174), .ZN(n8732) );
  NAND2_X1 U7645 ( .A1(n6285), .A2(n8732), .ZN(n6178) );
  NAND2_X1 U7646 ( .A1(n5895), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7647 ( .A1(n5897), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7648 ( .A1(n5896), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6175) );
  OR2_X1 U7649 ( .A1(n8504), .A2(n6741), .ZN(n8512) );
  OAI21_X2 U7650 ( .B1(n8511), .B2(n8512), .A(n6183), .ZN(n8499) );
  NAND2_X1 U7651 ( .A1(n7408), .A2(n7962), .ZN(n6185) );
  NAND2_X1 U7652 ( .A1(n7948), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6184) );
  XNOR2_X1 U7653 ( .A(n8854), .B(n6186), .ZN(n8501) );
  XNOR2_X1 U7654 ( .A(n6195), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U7655 ( .A1(n6285), .A2(n8717), .ZN(n6190) );
  NAND2_X1 U7656 ( .A1(n5895), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7657 ( .A1(n6286), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7658 ( .A1(n5896), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6187) );
  AND4_X1 U7659 ( .A1(n6190), .A2(n6189), .A3(n6188), .A4(n6187), .ZN(n8538)
         );
  INV_X1 U7660 ( .A(n8538), .ZN(n8738) );
  NAND2_X1 U7661 ( .A1(n8738), .A2(n7969), .ZN(n8500) );
  INV_X1 U7662 ( .A(n8501), .ZN(n6191) );
  NAND2_X1 U7663 ( .A1(n7536), .A2(n7962), .ZN(n6193) );
  NAND2_X1 U7664 ( .A1(n7948), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6192) );
  XNOR2_X1 U7665 ( .A(n8849), .B(n6231), .ZN(n6202) );
  INV_X1 U7666 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6194) );
  INV_X1 U7667 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8539) );
  OAI21_X1 U7668 ( .B1(n6195), .B2(n6194), .A(n8539), .ZN(n6196) );
  AND2_X1 U7669 ( .A1(n6196), .A2(n6208), .ZN(n8706) );
  NAND2_X1 U7670 ( .A1(n6285), .A2(n8706), .ZN(n6200) );
  NAND2_X1 U7671 ( .A1(n5895), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7672 ( .A1(n5897), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7673 ( .A1(n5896), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6197) );
  OR2_X1 U7674 ( .A1(n8503), .A2(n6230), .ZN(n6201) );
  NOR2_X1 U7675 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  AOI21_X1 U7676 ( .B1(n6202), .B2(n6201), .A(n6203), .ZN(n8537) );
  NAND2_X1 U7677 ( .A1(n7948), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6204) );
  XNOR2_X1 U7678 ( .A(n8843), .B(n6231), .ZN(n6215) );
  INV_X1 U7679 ( .A(n6208), .ZN(n6206) );
  NAND2_X1 U7680 ( .A1(n6206), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6224) );
  INV_X1 U7681 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7682 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  AND2_X1 U7683 ( .A1(n6224), .A2(n6209), .ZN(n8682) );
  NAND2_X1 U7684 ( .A1(n6285), .A2(n8682), .ZN(n6213) );
  NAND2_X1 U7685 ( .A1(n5895), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7686 ( .A1(n6286), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7687 ( .A1(n5896), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6210) );
  NAND4_X1 U7688 ( .A1(n6213), .A2(n6212), .A3(n6211), .A4(n6210), .ZN(n8550)
         );
  NAND2_X1 U7689 ( .A1(n8550), .A2(n7969), .ZN(n6214) );
  NOR2_X1 U7690 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  AOI21_X1 U7691 ( .B1(n6215), .B2(n6214), .A(n6216), .ZN(n8481) );
  NAND2_X1 U7692 ( .A1(n8482), .A2(n8481), .ZN(n8480) );
  INV_X1 U7693 ( .A(n6216), .ZN(n6217) );
  NAND2_X1 U7694 ( .A1(n8480), .A2(n6217), .ZN(n6278) );
  MUX2_X1 U7695 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5497), .Z(n7700) );
  INV_X1 U7696 ( .A(SI_28_), .ZN(n7701) );
  XNOR2_X1 U7697 ( .A(n7700), .B(n7701), .ZN(n7698) );
  NAND2_X1 U7698 ( .A1(n7875), .A2(n7962), .ZN(n6221) );
  NAND2_X1 U7699 ( .A1(n7948), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6220) );
  INV_X1 U7700 ( .A(n6224), .ZN(n6222) );
  NAND2_X1 U7701 ( .A1(n6222), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6284) );
  INV_X1 U7702 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7703 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  AND2_X1 U7704 ( .A1(n6284), .A2(n6225), .ZN(n8664) );
  NAND2_X1 U7705 ( .A1(n6285), .A2(n8664), .ZN(n6229) );
  NAND2_X1 U7706 ( .A1(n5895), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7707 ( .A1(n5897), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7708 ( .A1(n5896), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6226) );
  OR2_X1 U7709 ( .A1(n8483), .A2(n6230), .ZN(n6232) );
  XNOR2_X1 U7710 ( .A(n6232), .B(n6231), .ZN(n6270) );
  INV_X1 U7711 ( .A(n6270), .ZN(n6271) );
  INV_X1 U7712 ( .A(n6233), .ZN(n6234) );
  OAI21_X1 U7713 ( .B1(n6234), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6262) );
  INV_X1 U7714 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7715 ( .A1(n6262), .A2(n6261), .ZN(n6264) );
  NAND2_X1 U7716 ( .A1(n6264), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6236) );
  INV_X1 U7717 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6235) );
  XNOR2_X1 U7718 ( .A(n6236), .B(n6235), .ZN(n7344) );
  XNOR2_X1 U7719 ( .A(n7344), .B(P2_B_REG_SCAN_IN), .ZN(n6242) );
  NOR2_X1 U7720 ( .A1(n4472), .A2(n6238), .ZN(n6237) );
  MUX2_X1 U7721 ( .A(n6238), .B(n6237), .S(P2_IR_REG_25__SCAN_IN), .Z(n6239)
         );
  INV_X1 U7722 ( .A(n6239), .ZN(n6241) );
  NAND2_X1 U7723 ( .A1(n6241), .A2(n6240), .ZN(n7411) );
  NAND2_X1 U7724 ( .A1(n6242), .A2(n7411), .ZN(n6247) );
  NAND2_X1 U7725 ( .A1(n6240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6243) );
  MUX2_X1 U7726 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6243), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6245) );
  NAND2_X1 U7727 ( .A1(n6245), .A2(n6244), .ZN(n7540) );
  INV_X1 U7728 ( .A(n7540), .ZN(n6246) );
  INV_X1 U7729 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U7730 ( .A1(n9779), .A2(n10082), .ZN(n6249) );
  AND2_X1 U7731 ( .A1(n7344), .A2(n7540), .ZN(n9782) );
  INV_X1 U7732 ( .A(n9782), .ZN(n6248) );
  NAND2_X1 U7733 ( .A1(n6249), .A2(n6248), .ZN(n7199) );
  NOR4_X1 U7734 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6258) );
  OR4_X1 U7735 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6255) );
  NOR4_X1 U7736 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6253) );
  NOR4_X1 U7737 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6252) );
  NOR4_X1 U7738 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6251) );
  NOR4_X1 U7739 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6250) );
  NAND4_X1 U7740 ( .A1(n6253), .A2(n6252), .A3(n6251), .A4(n6250), .ZN(n6254)
         );
  NOR4_X1 U7741 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n6255), .A4(n6254), .ZN(n6257) );
  NOR4_X1 U7742 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6256) );
  NAND3_X1 U7743 ( .A1(n6258), .A2(n6257), .A3(n6256), .ZN(n6259) );
  NAND2_X1 U7744 ( .A1(n9779), .A2(n6259), .ZN(n6545) );
  INV_X1 U7745 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9783) );
  AND2_X1 U7746 ( .A1(n7411), .A2(n7540), .ZN(n9784) );
  AOI21_X1 U7747 ( .B1(n9779), .B2(n9783), .A(n9784), .ZN(n6547) );
  AND2_X1 U7748 ( .A1(n6545), .A2(n6547), .ZN(n7195) );
  INV_X1 U7749 ( .A(n7195), .ZN(n6260) );
  OR2_X1 U7750 ( .A1(n7199), .A2(n6260), .ZN(n6293) );
  OR2_X1 U7751 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  NAND2_X1 U7752 ( .A1(n6264), .A2(n6263), .ZN(n6391) );
  NAND2_X1 U7753 ( .A1(n6571), .A2(n9785), .ZN(n9780) );
  INV_X1 U7754 ( .A(n7021), .ZN(n8151) );
  NAND2_X1 U7755 ( .A1(n6265), .A2(n8151), .ZN(n7206) );
  OR2_X1 U7756 ( .A1(n6282), .A2(n7206), .ZN(n6267) );
  NAND2_X1 U7757 ( .A1(n6266), .A2(n7966), .ZN(n6543) );
  NAND2_X1 U7758 ( .A1(n6267), .A2(n8817), .ZN(n8520) );
  NOR3_X1 U7759 ( .A1(n8666), .A2(n6271), .A3(n8520), .ZN(n6268) );
  AOI21_X1 U7760 ( .B1(n8666), .B2(n6271), .A(n6268), .ZN(n6269) );
  NOR3_X1 U7761 ( .A1(n8666), .A2(n6270), .A3(n8520), .ZN(n6273) );
  NOR2_X1 U7762 ( .A1(n8838), .A2(n6271), .ZN(n6272) );
  OR2_X1 U7763 ( .A1(n6273), .A2(n6272), .ZN(n6277) );
  AND2_X1 U7764 ( .A1(n7021), .A2(n8707), .ZN(n6294) );
  INV_X1 U7765 ( .A(n6294), .ZN(n6281) );
  NAND2_X1 U7766 ( .A1(n8159), .A2(n8152), .ZN(n6390) );
  NAND2_X1 U7767 ( .A1(n9850), .A2(n6390), .ZN(n6274) );
  OAI21_X1 U7768 ( .B1(n8666), .B2(n8546), .A(n8522), .ZN(n6275) );
  AOI21_X1 U7769 ( .B1(n6278), .B2(n6277), .A(n6276), .ZN(n6279) );
  NAND2_X1 U7770 ( .A1(n6280), .A2(n6279), .ZN(n6303) );
  INV_X1 U7771 ( .A(n6390), .ZN(n6574) );
  AND2_X1 U7772 ( .A1(n6574), .A2(n6283), .ZN(n8781) );
  INV_X1 U7773 ( .A(n8781), .ZN(n9761) );
  NOR2_X1 U7774 ( .A1(n8541), .A2(n9761), .ZN(n8528) );
  INV_X1 U7775 ( .A(n6284), .ZN(n8460) );
  NAND2_X1 U7776 ( .A1(n6285), .A2(n8460), .ZN(n6290) );
  NAND2_X1 U7777 ( .A1(n5895), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7778 ( .A1(n6286), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7779 ( .A1(n5896), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6287) );
  AND4_X1 U7780 ( .A1(n6290), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(n8670)
         );
  INV_X1 U7781 ( .A(n8670), .ZN(n8548) );
  INV_X1 U7782 ( .A(n6283), .ZN(n6291) );
  AND2_X1 U7783 ( .A1(n6574), .A2(n6291), .ZN(n8783) );
  INV_X2 U7784 ( .A(n8783), .ZN(n9763) );
  AOI22_X1 U7785 ( .A1(n8528), .A2(n8548), .B1(n8527), .B2(n8550), .ZN(n6292)
         );
  INV_X1 U7786 ( .A(n6292), .ZN(n6301) );
  NAND2_X1 U7787 ( .A1(n6293), .A2(n6543), .ZN(n6297) );
  OR2_X1 U7788 ( .A1(n6390), .A2(n6294), .ZN(n7196) );
  AND2_X1 U7789 ( .A1(n7196), .A2(n6391), .ZN(n6295) );
  NAND2_X1 U7790 ( .A1(n6571), .A2(n6295), .ZN(n8158) );
  INV_X1 U7791 ( .A(n8158), .ZN(n6296) );
  NAND2_X1 U7792 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  AOI22_X1 U7793 ( .A1(n8543), .A2(n8664), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6299) );
  NAND2_X1 U7794 ( .A1(n6303), .A2(n6302), .ZN(P2_U3222) );
  INV_X1 U7795 ( .A(n7212), .ZN(n6306) );
  OR2_X1 U7796 ( .A1(n6304), .A2(n6306), .ZN(n6342) );
  NOR2_X1 U7797 ( .A1(n6342), .A2(P1_U3084), .ZN(P1_U4006) );
  INV_X1 U7798 ( .A(n9785), .ZN(n6305) );
  NOR2_X2 U7799 ( .A1(n6571), .A2(n6305), .ZN(P2_U3966) );
  OR2_X1 U7800 ( .A1(n6887), .A2(n6306), .ZN(n6307) );
  AND2_X1 U7801 ( .A1(n6342), .A2(n6307), .ZN(n9501) );
  NAND2_X1 U7802 ( .A1(n9501), .A2(n6308), .ZN(n6309) );
  NAND2_X1 U7803 ( .A1(n6309), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7804 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6975) );
  XNOR2_X1 U7805 ( .A(n6631), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6322) );
  NOR2_X1 U7806 ( .A1(n9531), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6310) );
  AOI21_X1 U7807 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9531), .A(n6310), .ZN(
        n9527) );
  INV_X1 U7808 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7010) );
  XNOR2_X1 U7809 ( .A(n6470), .B(n7010), .ZN(n6466) );
  INV_X1 U7810 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6311) );
  MUX2_X1 U7811 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6311), .S(n6364), .Z(n6488)
         );
  AND2_X1 U7812 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6487) );
  NAND2_X1 U7813 ( .A1(n6488), .A2(n6487), .ZN(n6486) );
  NAND2_X1 U7814 ( .A1(n6364), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7815 ( .A1(n6486), .A2(n6312), .ZN(n6465) );
  NAND2_X1 U7816 ( .A1(n6466), .A2(n6465), .ZN(n6464) );
  NAND2_X1 U7817 ( .A1(n6470), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7818 ( .A1(n6464), .A2(n6313), .ZN(n6412) );
  INV_X1 U7819 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6994) );
  XNOR2_X1 U7820 ( .A(n7867), .B(n6994), .ZN(n6413) );
  NAND2_X1 U7821 ( .A1(n6412), .A2(n6413), .ZN(n6411) );
  NAND2_X1 U7822 ( .A1(n7867), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7823 ( .A1(n6411), .A2(n6314), .ZN(n6473) );
  XNOR2_X1 U7824 ( .A(n7871), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6472) );
  OR2_X1 U7825 ( .A1(n7871), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6315) );
  XNOR2_X1 U7826 ( .A(n6372), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U7827 ( .A1(n6425), .A2(n6426), .ZN(n6424) );
  NAND2_X1 U7828 ( .A1(n6372), .A2(n6316), .ZN(n6317) );
  NAND2_X1 U7829 ( .A1(n6424), .A2(n6317), .ZN(n6508) );
  MUX2_X1 U7830 ( .A(n6318), .B(P1_REG2_REG_6__SCAN_IN), .S(n6334), .Z(n6509)
         );
  XNOR2_X1 U7831 ( .A(n9516), .B(n6957), .ZN(n9511) );
  NAND2_X1 U7832 ( .A1(n6334), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9512) );
  AND2_X1 U7833 ( .A1(n9511), .A2(n9512), .ZN(n6319) );
  NAND2_X1 U7834 ( .A1(n9527), .A2(n9528), .ZN(n9526) );
  OAI21_X1 U7835 ( .B1(n9531), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9526), .ZN(
        n6321) );
  NOR2_X1 U7836 ( .A1(n6321), .A2(n6322), .ZN(n6630) );
  INV_X1 U7837 ( .A(n9501), .ZN(n6320) );
  INV_X1 U7838 ( .A(n9067), .ZN(n8447) );
  NAND2_X1 U7839 ( .A1(n8447), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7584) );
  NOR2_X1 U7840 ( .A1(n6320), .A2(n7584), .ZN(n9499) );
  AND2_X1 U7841 ( .A1(n9499), .A2(n9500), .ZN(n9619) );
  INV_X1 U7842 ( .A(n9619), .ZN(n9587) );
  AOI211_X1 U7843 ( .C1(n6322), .C2(n6321), .A(n6630), .B(n9587), .ZN(n6347)
         );
  NOR2_X1 U7844 ( .A1(n9531), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9533) );
  INV_X1 U7845 ( .A(n9531), .ZN(n6377) );
  INV_X1 U7846 ( .A(n6334), .ZN(n6510) );
  MUX2_X1 U7847 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5130), .S(n6372), .Z(n6428)
         );
  MUX2_X1 U7848 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6323), .S(n6470), .Z(n6326)
         );
  MUX2_X1 U7849 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6324), .S(n6364), .Z(n6492)
         );
  AND2_X1 U7850 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6493) );
  NAND2_X1 U7851 ( .A1(n6492), .A2(n6493), .ZN(n6491) );
  NAND2_X1 U7852 ( .A1(n6364), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U7853 ( .A1(n6491), .A2(n6459), .ZN(n6325) );
  NAND2_X1 U7854 ( .A1(n6326), .A2(n6325), .ZN(n6462) );
  NAND2_X1 U7855 ( .A1(n6470), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U7856 ( .A1(n6462), .A2(n6406), .ZN(n6329) );
  MUX2_X1 U7857 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6327), .S(n7867), .Z(n6328)
         );
  NAND2_X1 U7858 ( .A1(n6329), .A2(n6328), .ZN(n6408) );
  NAND2_X1 U7859 ( .A1(n7867), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6330) );
  MUX2_X1 U7860 ( .A(n5098), .B(P1_REG1_REG_4__SCAN_IN), .S(n7871), .Z(n6331)
         );
  OR2_X1 U7861 ( .A1(n7871), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7862 ( .A1(n6477), .A2(n6332), .ZN(n6429) );
  NAND2_X1 U7863 ( .A1(n6427), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7864 ( .A1(n6431), .A2(n6333), .ZN(n6503) );
  MUX2_X1 U7865 ( .A(n6335), .B(P1_REG1_REG_6__SCAN_IN), .S(n6334), .Z(n6502)
         );
  INV_X1 U7866 ( .A(n9516), .ZN(n6336) );
  OAI21_X1 U7867 ( .B1(n5191), .B2(n6336), .A(n4459), .ZN(n9508) );
  INV_X1 U7868 ( .A(n9532), .ZN(n9524) );
  INV_X1 U7869 ( .A(n6631), .ZN(n6344) );
  NOR2_X1 U7870 ( .A1(n6631), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6625) );
  INV_X1 U7871 ( .A(n6625), .ZN(n6337) );
  OAI21_X1 U7872 ( .B1(n5243), .B2(n6344), .A(n6337), .ZN(n6338) );
  AOI21_X1 U7873 ( .B1(n6339), .B2(n6338), .A(n6624), .ZN(n6341) );
  NOR2_X1 U7874 ( .A1(n5777), .A2(n8447), .ZN(n6458) );
  AND2_X1 U7875 ( .A1(n6458), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6340) );
  AND2_X1 U7876 ( .A1(n6340), .A2(n9501), .ZN(n9625) );
  INV_X1 U7877 ( .A(n9625), .ZN(n9575) );
  NOR2_X1 U7878 ( .A1(n6341), .A2(n9575), .ZN(n6346) );
  INV_X1 U7879 ( .A(n6342), .ZN(n6343) );
  NOR2_X1 U7880 ( .A1(P1_U3083), .A2(n6343), .ZN(n9571) );
  INV_X1 U7881 ( .A(n9571), .ZN(n9631) );
  INV_X1 U7882 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10223) );
  AND2_X1 U7883 ( .A1(n9499), .A2(n5777), .ZN(n9621) );
  INV_X1 U7884 ( .A(n9621), .ZN(n6697) );
  OAI22_X1 U7885 ( .A1(n9631), .A2(n10223), .B1(n6344), .B2(n6697), .ZN(n6345)
         );
  OR4_X1 U7886 ( .A1(n6975), .A2(n6347), .A3(n6346), .A4(n6345), .ZN(P1_U3250)
         );
  AND2_X1 U7887 ( .A1(n6348), .A2(n6761), .ZN(n6349) );
  AOI211_X1 U7888 ( .C1(n6350), .C2(n6349), .A(n8522), .B(n4475), .ZN(n6354)
         );
  INV_X1 U7889 ( .A(n8528), .ZN(n8516) );
  OAI22_X1 U7890 ( .A1(n8516), .A2(n7297), .B1(n7336), .B2(n8546), .ZN(n6353)
         );
  INV_X1 U7891 ( .A(n8527), .ZN(n8517) );
  NOR2_X1 U7892 ( .A1(n8517), .A2(n6718), .ZN(n6352) );
  OAI22_X1 U7893 ( .A1(n8515), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n5875), .ZN(n6351) );
  OR4_X1 U7894 ( .A1(n6354), .A2(n6353), .A3(n6352), .A4(n6351), .ZN(P2_U3220)
         );
  NAND2_X1 U7895 ( .A1(n5497), .A2(P2_U3152), .ZN(n8475) );
  AND2_X1 U7896 ( .A1(n7833), .A2(P2_U3152), .ZN(n7234) );
  INV_X2 U7897 ( .A(n7234), .ZN(n8478) );
  INV_X1 U7898 ( .A(n6598), .ZN(n9406) );
  OAI222_X1 U7899 ( .A1(n8475), .A2(n6355), .B1(n8478), .B2(n6366), .C1(n9406), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  NAND2_X1 U7900 ( .A1(n6356), .A2(n9633), .ZN(n6357) );
  OAI21_X1 U7901 ( .B1(n9633), .B2(n10011), .A(n6357), .ZN(P1_U3441) );
  NAND2_X1 U7902 ( .A1(n7833), .A2(P1_U3084), .ZN(n7863) );
  INV_X1 U7903 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9972) );
  AND2_X1 U7904 ( .A1(n5497), .A2(P1_U3084), .ZN(n7582) );
  INV_X2 U7905 ( .A(n7582), .ZN(n7873) );
  INV_X1 U7906 ( .A(n6358), .ZN(n6362) );
  OAI222_X1 U7907 ( .A1(n7863), .A2(n9972), .B1(n7873), .B2(n6362), .C1(
        P1_U3084), .C2(n6510), .ZN(P1_U3347) );
  INV_X1 U7908 ( .A(n7863), .ZN(n7870) );
  AOI22_X1 U7909 ( .A1(n6470), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n7870), .ZN(n6359) );
  OAI21_X1 U7910 ( .B1(n6361), .B2(n7873), .A(n6359), .ZN(P1_U3351) );
  INV_X1 U7911 ( .A(n8475), .ZN(n7578) );
  INV_X1 U7912 ( .A(n7578), .ZN(n7837) );
  INV_X1 U7913 ( .A(n9419), .ZN(n6360) );
  OAI222_X1 U7914 ( .A1(n7837), .A2(n9907), .B1(n8478), .B2(n6361), .C1(
        P2_U3152), .C2(n6360), .ZN(P2_U3356) );
  INV_X1 U7915 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6363) );
  INV_X1 U7916 ( .A(n8571), .ZN(n6586) );
  OAI222_X1 U7917 ( .A1(n7837), .A2(n6363), .B1(n8478), .B2(n6362), .C1(
        P2_U3152), .C2(n6586), .ZN(P2_U3352) );
  INV_X1 U7918 ( .A(n6364), .ZN(n6490) );
  INV_X1 U7919 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6365) );
  OAI222_X1 U7920 ( .A1(P1_U3084), .A2(n6490), .B1(n7873), .B2(n6366), .C1(
        n6365), .C2(n7863), .ZN(P1_U3352) );
  INV_X1 U7921 ( .A(n6367), .ZN(n6370) );
  AOI22_X1 U7922 ( .A1(n6735), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n7578), .ZN(n6368) );
  OAI21_X1 U7923 ( .B1(n6370), .B2(n8478), .A(n6368), .ZN(P2_U3351) );
  AOI22_X1 U7924 ( .A1(n9516), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7870), .ZN(n6369) );
  OAI21_X1 U7925 ( .B1(n6370), .B2(n7873), .A(n6369), .ZN(P1_U3346) );
  INV_X1 U7926 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6371) );
  INV_X1 U7927 ( .A(n5907), .ZN(n6373) );
  INV_X1 U7928 ( .A(n6604), .ZN(n6669) );
  OAI222_X1 U7929 ( .A1(n7837), .A2(n6371), .B1(n8478), .B2(n6373), .C1(
        P2_U3152), .C2(n6669), .ZN(P2_U3353) );
  INV_X1 U7930 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6374) );
  OAI222_X1 U7931 ( .A1(n7863), .A2(n6374), .B1(n7873), .B2(n6373), .C1(
        P1_U3084), .C2(n6372), .ZN(P1_U3348) );
  INV_X1 U7932 ( .A(n6603), .ZN(n6657) );
  OAI222_X1 U7933 ( .A1(n7837), .A2(n6375), .B1(n8478), .B2(n7874), .C1(
        P2_U3152), .C2(n6657), .ZN(P2_U3354) );
  OAI222_X1 U7934 ( .A1(n7837), .A2(n9968), .B1(n8478), .B2(n7869), .C1(
        P2_U3152), .C2(n6681), .ZN(P2_U3355) );
  INV_X1 U7935 ( .A(n6376), .ZN(n6379) );
  OAI222_X1 U7936 ( .A1(n7863), .A2(n9973), .B1(n7873), .B2(n6379), .C1(
        P1_U3084), .C2(n6377), .ZN(P1_U3345) );
  INV_X1 U7937 ( .A(n8587), .ZN(n6378) );
  OAI222_X1 U7938 ( .A1(n7837), .A2(n9951), .B1(n8478), .B2(n6379), .C1(
        P2_U3152), .C2(n6378), .ZN(P2_U3350) );
  INV_X1 U7939 ( .A(n6380), .ZN(n6385) );
  AOI22_X1 U7940 ( .A1(n6631), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7870), .ZN(n6381) );
  OAI21_X1 U7941 ( .B1(n6385), .B2(n7873), .A(n6381), .ZN(P1_U3344) );
  INV_X1 U7942 ( .A(n6382), .ZN(n6383) );
  INV_X1 U7943 ( .A(n6700), .ZN(n6694) );
  OAI222_X1 U7944 ( .A1(n7863), .A2(n9985), .B1(n7873), .B2(n6383), .C1(n6694), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U7945 ( .A(n7151), .ZN(n7159) );
  OAI222_X1 U7946 ( .A1(P2_U3152), .A2(n7159), .B1(n8478), .B2(n6383), .C1(
        n6500), .C2(n7837), .ZN(P2_U3348) );
  INV_X1 U7947 ( .A(n6770), .ZN(n6774) );
  OAI222_X1 U7948 ( .A1(P2_U3152), .A2(n6774), .B1(n8478), .B2(n6385), .C1(
        n6384), .C2(n7837), .ZN(P2_U3349) );
  INV_X1 U7949 ( .A(n6386), .ZN(n6388) );
  INV_X1 U7950 ( .A(n9042), .ZN(n9030) );
  OAI222_X1 U7951 ( .A1(n7863), .A2(n6387), .B1(n7873), .B2(n6388), .C1(n9030), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7952 ( .A(n8596), .ZN(n6389) );
  OAI222_X1 U7953 ( .A1(P2_U3152), .A2(n6389), .B1(n8478), .B2(n6388), .C1(
        n10104), .C2(n7837), .ZN(P2_U3347) );
  OAI21_X1 U7954 ( .B1(n9780), .B2(n6390), .A(n6575), .ZN(n6394) );
  INV_X1 U7955 ( .A(n6391), .ZN(n6392) );
  NAND2_X1 U7956 ( .A1(n6392), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8161) );
  NAND2_X1 U7957 ( .A1(n9780), .A2(n8161), .ZN(n6393) );
  NAND2_X1 U7958 ( .A1(n6394), .A2(n6393), .ZN(n9402) );
  INV_X1 U7959 ( .A(n9402), .ZN(n9715) );
  NOR2_X1 U7960 ( .A1(n9715), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7961 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U7962 ( .A1(n5895), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U7963 ( .A1(n5897), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U7964 ( .A1(n5896), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6395) );
  NAND3_X1 U7965 ( .A1(n6397), .A2(n6396), .A3(n6395), .ZN(n8649) );
  NAND2_X1 U7966 ( .A1(P2_U3966), .A2(n8649), .ZN(n6398) );
  OAI21_X1 U7967 ( .B1(P2_U3966), .B2(n6399), .A(n6398), .ZN(P2_U3583) );
  NAND2_X1 U7968 ( .A1(P2_U3966), .A2(n6751), .ZN(n6400) );
  OAI21_X1 U7969 ( .B1(P2_U3966), .B2(n5003), .A(n6400), .ZN(P2_U3552) );
  INV_X1 U7970 ( .A(n6401), .ZN(n6404) );
  AOI22_X1 U7971 ( .A1(n7227), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n7578), .ZN(n6402) );
  OAI21_X1 U7972 ( .B1(n6404), .B2(n8478), .A(n6402), .ZN(P2_U3346) );
  AOI22_X1 U7973 ( .A1(n9543), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7870), .ZN(n6403) );
  OAI21_X1 U7974 ( .B1(n6404), .B2(n7873), .A(n6403), .ZN(P1_U3341) );
  INV_X1 U7975 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6416) );
  MUX2_X1 U7976 ( .A(n6327), .B(P1_REG1_REG_3__SCAN_IN), .S(n7867), .Z(n6405)
         );
  NAND3_X1 U7977 ( .A1(n6462), .A2(n6406), .A3(n6405), .ZN(n6407) );
  NAND3_X1 U7978 ( .A1(n9625), .A2(n6408), .A3(n6407), .ZN(n6409) );
  OAI21_X1 U7979 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6618), .A(n6409), .ZN(n6410) );
  AOI21_X1 U7980 ( .B1(n7867), .B2(n9621), .A(n6410), .ZN(n6415) );
  OAI211_X1 U7981 ( .C1(n6413), .C2(n6412), .A(n9619), .B(n6411), .ZN(n6414)
         );
  OAI211_X1 U7982 ( .C1(n9631), .C2(n6416), .A(n6415), .B(n6414), .ZN(P1_U3244) );
  INV_X1 U7983 ( .A(P1_U4006), .ZN(n9026) );
  INV_X1 U7984 ( .A(n9026), .ZN(n9019) );
  INV_X1 U7985 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6422) );
  INV_X1 U7986 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U7987 ( .A1(n5017), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6419) );
  INV_X1 U7988 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6417) );
  OR2_X1 U7989 ( .A1(n5100), .A2(n6417), .ZN(n6418) );
  OAI211_X1 U7990 ( .C1(n8172), .C2(n6420), .A(n6419), .B(n6418), .ZN(n9069)
         );
  NAND2_X1 U7991 ( .A1(n9069), .A2(n9019), .ZN(n6421) );
  OAI21_X1 U7992 ( .B1(n9019), .B2(n6422), .A(n6421), .ZN(P1_U3586) );
  NAND2_X1 U7993 ( .A1(n6888), .A2(n9019), .ZN(n6423) );
  OAI21_X1 U7994 ( .B1(n9019), .B2(n4492), .A(n6423), .ZN(P1_U3555) );
  INV_X1 U7995 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6437) );
  OAI21_X1 U7996 ( .B1(n6426), .B2(n6425), .A(n6424), .ZN(n6435) );
  NAND2_X1 U7997 ( .A1(n9621), .A2(n6427), .ZN(n6433) );
  NAND2_X1 U7998 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U7999 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  NAND3_X1 U8000 ( .A1(n9625), .A2(n6431), .A3(n6430), .ZN(n6432) );
  NAND3_X1 U8001 ( .A1(n6433), .A2(n6864), .A3(n6432), .ZN(n6434) );
  AOI21_X1 U8002 ( .B1(n9619), .B2(n6435), .A(n6434), .ZN(n6436) );
  OAI21_X1 U8003 ( .B1(n9631), .B2(n6437), .A(n6436), .ZN(P1_U3246) );
  AND2_X1 U8004 ( .A1(n6439), .A2(n7020), .ZN(n9366) );
  NAND2_X1 U8005 ( .A1(n9366), .A2(n9275), .ZN(n6438) );
  NAND4_X1 U8006 ( .A1(n6899), .A2(n6897), .A3(n6896), .A4(n6438), .ZN(n6446)
         );
  INV_X2 U8007 ( .A(n9694), .ZN(n9696) );
  INV_X1 U8008 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6445) );
  INV_X1 U8009 ( .A(n6904), .ZN(n6891) );
  INV_X1 U8010 ( .A(n6439), .ZN(n6443) );
  AND2_X1 U8011 ( .A1(n6888), .A2(n6891), .ZN(n8190) );
  NOR2_X1 U8012 ( .A1(n6947), .A2(n8190), .ZN(n8242) );
  OR3_X1 U8013 ( .A1(n8242), .A2(n6440), .A3(n6439), .ZN(n6442) );
  OR2_X1 U8014 ( .A1(n6887), .A2(n9500), .ZN(n9269) );
  INV_X1 U8015 ( .A(n9269), .ZN(n9218) );
  NAND2_X1 U8016 ( .A1(n9027), .A2(n9218), .ZN(n6441) );
  AND2_X1 U8017 ( .A1(n6442), .A2(n6441), .ZN(n6907) );
  OAI21_X1 U8018 ( .B1(n6891), .B2(n6443), .A(n6907), .ZN(n6447) );
  NAND2_X1 U8019 ( .A1(n6447), .A2(n9696), .ZN(n6444) );
  OAI21_X1 U8020 ( .B1(n9696), .B2(n6445), .A(n6444), .ZN(P1_U3454) );
  INV_X2 U8021 ( .A(n9705), .ZN(n9707) );
  NAND2_X1 U8022 ( .A1(n6447), .A2(n9707), .ZN(n6448) );
  OAI21_X1 U8023 ( .B1(n9707), .B2(n5011), .A(n6448), .ZN(P1_U3523) );
  INV_X1 U8024 ( .A(n6449), .ZN(n6515) );
  AOI22_X1 U8025 ( .A1(n9552), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7870), .ZN(n6450) );
  OAI21_X1 U8026 ( .B1(n6515), .B2(n7873), .A(n6450), .ZN(P1_U3340) );
  INV_X1 U8027 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U8028 ( .A1(n8447), .A2(n6451), .ZN(n6452) );
  NAND2_X1 U8029 ( .A1(n9500), .A2(n6452), .ZN(n6453) );
  XNOR2_X1 U8030 ( .A(n6453), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9503) );
  INV_X1 U8031 ( .A(n6539), .ZN(n6456) );
  NAND2_X1 U8032 ( .A1(n6456), .A2(n6458), .ZN(n6457) );
  OAI211_X1 U8033 ( .C1(n6458), .C2(n9503), .A(n6457), .B(n9019), .ZN(n6485)
         );
  MUX2_X1 U8034 ( .A(n6323), .B(P1_REG1_REG_2__SCAN_IN), .S(n6470), .Z(n6460)
         );
  NAND3_X1 U8035 ( .A1(n6460), .A2(n6491), .A3(n6459), .ZN(n6461) );
  NAND3_X1 U8036 ( .A1(n9625), .A2(n6462), .A3(n6461), .ZN(n6463) );
  OAI21_X1 U8037 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7009), .A(n6463), .ZN(n6469) );
  OAI211_X1 U8038 ( .C1(n6466), .C2(n6465), .A(n9619), .B(n6464), .ZN(n6467)
         );
  INV_X1 U8039 ( .A(n6467), .ZN(n6468) );
  AOI211_X1 U8040 ( .C1(n9621), .C2(n6470), .A(n6469), .B(n6468), .ZN(n6471)
         );
  OAI211_X1 U8041 ( .C1(n7546), .C2(n9631), .A(n6485), .B(n6471), .ZN(P1_U3243) );
  INV_X1 U8042 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U8043 ( .A1(n9621), .A2(n7871), .ZN(n6483) );
  NAND2_X1 U8044 ( .A1(n6473), .A2(n6472), .ZN(n6474) );
  NAND2_X1 U8045 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  NAND2_X1 U8046 ( .A1(n9619), .A2(n6476), .ZN(n6482) );
  NAND2_X1 U8047 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n6687) );
  MUX2_X1 U8048 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n5098), .S(n7871), .Z(n6478)
         );
  OAI21_X1 U8049 ( .B1(n6479), .B2(n6478), .A(n6477), .ZN(n6480) );
  NAND2_X1 U8050 ( .A1(n9625), .A2(n6480), .ZN(n6481) );
  AND4_X1 U8051 ( .A1(n6483), .A2(n6482), .A3(n6687), .A4(n6481), .ZN(n6484)
         );
  OAI211_X1 U8052 ( .C1(n9986), .C2(n9631), .A(n6485), .B(n6484), .ZN(P1_U3245) );
  OAI211_X1 U8053 ( .C1(n6488), .C2(n6487), .A(n9619), .B(n6486), .ZN(n6489)
         );
  OAI21_X1 U8054 ( .B1(n6697), .B2(n6490), .A(n6489), .ZN(n6496) );
  OAI211_X1 U8055 ( .C1(n6493), .C2(n6492), .A(n9625), .B(n6491), .ZN(n6494)
         );
  OAI21_X1 U8056 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n5018), .A(n6494), .ZN(n6495) );
  AOI211_X1 U8057 ( .C1(n9571), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6496), .B(
        n6495), .ZN(n6497) );
  INV_X1 U8058 ( .A(n6497), .ZN(P1_U3242) );
  MUX2_X1 U8059 ( .A(n6498), .B(n7516), .S(n9019), .Z(n6499) );
  INV_X1 U8060 ( .A(n6499), .ZN(P1_U3567) );
  MUX2_X1 U8061 ( .A(n6500), .B(n7177), .S(n9019), .Z(n6501) );
  INV_X1 U8062 ( .A(n6501), .ZN(P1_U3565) );
  AND2_X1 U8063 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  NOR2_X1 U8064 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  NAND2_X1 U8065 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6919) );
  OAI21_X1 U8066 ( .B1(n6506), .B2(n9575), .A(n6919), .ZN(n6514) );
  INV_X1 U8067 ( .A(n9513), .ZN(n6507) );
  AOI211_X1 U8068 ( .C1(n6509), .C2(n6508), .A(n6507), .B(n9587), .ZN(n6513)
         );
  INV_X1 U8069 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6511) );
  OAI22_X1 U8070 ( .A1(n9631), .A2(n6511), .B1(n6510), .B2(n6697), .ZN(n6512)
         );
  OR3_X1 U8071 ( .A1(n6514), .A2(n6513), .A3(n6512), .ZN(P1_U3247) );
  INV_X1 U8072 ( .A(n7399), .ZN(n7394) );
  OAI222_X1 U8073 ( .A1(n7837), .A2(n6516), .B1(n8478), .B2(n6515), .C1(n7394), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8074 ( .A(P2_U3966), .ZN(n8549) );
  NAND2_X1 U8075 ( .A1(n8549), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6517) );
  OAI21_X1 U8076 ( .B1(n8549), .B2(n8504), .A(n6517), .ZN(P2_U3576) );
  XNOR2_X1 U8077 ( .A(n6519), .B(n6518), .ZN(n6521) );
  XNOR2_X1 U8078 ( .A(n6521), .B(n6520), .ZN(n6525) );
  INV_X1 U8079 ( .A(n9435), .ZN(n8980) );
  INV_X1 U8080 ( .A(n8983), .ZN(n9438) );
  AOI22_X1 U8081 ( .A1(n8980), .A2(n6888), .B1(n9438), .B2(n9025), .ZN(n6523)
         );
  NAND2_X1 U8082 ( .A1(n9445), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6522) );
  OAI211_X1 U8083 ( .C1(n9010), .C2(n9640), .A(n6523), .B(n6522), .ZN(n6524)
         );
  AOI21_X1 U8084 ( .B1(n6525), .B2(n9002), .A(n6524), .ZN(n6526) );
  INV_X1 U8085 ( .A(n6526), .ZN(P1_U3220) );
  INV_X1 U8086 ( .A(n6527), .ZN(n6529) );
  INV_X1 U8087 ( .A(n9568), .ZN(n9049) );
  OAI222_X1 U8088 ( .A1(n7863), .A2(n6528), .B1(n7873), .B2(n6529), .C1(n9049), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8089 ( .A(n7596), .ZN(n7599) );
  OAI222_X1 U8090 ( .A1(n8475), .A2(n6530), .B1(n8478), .B2(n6529), .C1(n7599), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8091 ( .A(n6532), .ZN(n6533) );
  AOI21_X1 U8092 ( .B1(n6534), .B2(n6531), .A(n6533), .ZN(n6538) );
  INV_X1 U8093 ( .A(n9445), .ZN(n6797) );
  AOI22_X1 U8094 ( .A1(n8980), .A2(n9027), .B1(n9438), .B2(n9024), .ZN(n6535)
         );
  OAI21_X1 U8095 ( .B1(n6797), .B2(n7009), .A(n6535), .ZN(n6536) );
  AOI21_X1 U8096 ( .B1(n5797), .B2(n7015), .A(n6536), .ZN(n6537) );
  OAI21_X1 U8097 ( .B1(n6538), .B2(n9446), .A(n6537), .ZN(P1_U3235) );
  AOI22_X1 U8098 ( .A1(n6539), .A2(n9002), .B1(n9438), .B2(n9027), .ZN(n6541)
         );
  NAND2_X1 U8099 ( .A1(n5797), .A2(n6904), .ZN(n6540) );
  OAI211_X1 U8100 ( .C1(n6797), .C2(n6542), .A(n6541), .B(n6540), .ZN(P1_U3230) );
  INV_X1 U8101 ( .A(n9780), .ZN(n6544) );
  NAND4_X1 U8102 ( .A1(n6545), .A2(n6544), .A3(n7196), .A4(n6543), .ZN(n6546)
         );
  OR2_X1 U8103 ( .A1(n6547), .A2(n6546), .ZN(n6567) );
  INV_X1 U8104 ( .A(n7199), .ZN(n6548) );
  INV_X2 U8105 ( .A(n9855), .ZN(n9856) );
  INV_X1 U8106 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6556) );
  INV_X1 U8107 ( .A(n6751), .ZN(n6549) );
  NAND2_X1 U8108 ( .A1(n6549), .A2(n7208), .ZN(n6715) );
  INV_X1 U8109 ( .A(n7208), .ZN(n6747) );
  NAND2_X1 U8110 ( .A1(n6751), .A2(n6747), .ZN(n8121) );
  NAND2_X1 U8111 ( .A1(n6715), .A2(n8121), .ZN(n7194) );
  NAND2_X1 U8112 ( .A1(n8152), .A2(n8151), .ZN(n7968) );
  NAND2_X1 U8113 ( .A1(n6550), .A2(n7968), .ZN(n9766) );
  AOI22_X1 U8114 ( .A1(n7194), .A2(n9766), .B1(n8781), .B2(n6557), .ZN(n7204)
         );
  XNOR2_X1 U8115 ( .A(n8159), .B(n7200), .ZN(n6551) );
  NAND2_X1 U8116 ( .A1(n6551), .A2(n8707), .ZN(n9769) );
  AND2_X1 U8117 ( .A1(n7021), .A2(n7966), .ZN(n6553) );
  NAND2_X1 U8118 ( .A1(n6552), .A2(n6553), .ZN(n9827) );
  AND2_X1 U8119 ( .A1(n9769), .A2(n9827), .ZN(n8897) );
  INV_X1 U8120 ( .A(n8897), .ZN(n9854) );
  AOI22_X1 U8121 ( .A1(n7194), .A2(n9854), .B1(n6265), .B2(n7208), .ZN(n6554)
         );
  NAND2_X1 U8122 ( .A1(n7204), .A2(n6554), .ZN(n6569) );
  NAND2_X1 U8123 ( .A1(n9856), .A2(n6569), .ZN(n6555) );
  OAI21_X1 U8124 ( .B1(n9856), .B2(n6556), .A(n6555), .ZN(P2_U3451) );
  OAI21_X1 U8125 ( .B1(n6558), .B2(n6559), .A(n6710), .ZN(n7242) );
  NAND2_X1 U8126 ( .A1(n7241), .A2(n7208), .ZN(n6560) );
  NAND2_X1 U8127 ( .A1(n6560), .A2(n6266), .ZN(n6561) );
  OR2_X1 U8128 ( .A1(n6561), .A2(n7279), .ZN(n7237) );
  OAI21_X1 U8129 ( .B1(n6708), .B2(n9850), .A(n7237), .ZN(n6566) );
  INV_X1 U8130 ( .A(n6715), .ZN(n6744) );
  NOR2_X1 U8131 ( .A1(n6558), .A2(n6744), .ZN(n8123) );
  NAND2_X1 U8132 ( .A1(n6558), .A2(n6744), .ZN(n6562) );
  NAND2_X1 U8133 ( .A1(n6562), .A2(n9766), .ZN(n6563) );
  OR2_X1 U8134 ( .A1(n8123), .A2(n6563), .ZN(n6565) );
  AOI22_X1 U8135 ( .A1(n8570), .A2(n8781), .B1(n8783), .B2(n6751), .ZN(n6564)
         );
  NAND2_X1 U8136 ( .A1(n6565), .A2(n6564), .ZN(n7240) );
  AOI211_X1 U8137 ( .C1(n9854), .C2(n7242), .A(n6566), .B(n7240), .ZN(n6638)
         );
  NAND2_X1 U8138 ( .A1(n9870), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6568) );
  OAI21_X1 U8139 ( .B1(n6638), .B2(n9870), .A(n6568), .ZN(P2_U3521) );
  INV_X2 U8140 ( .A(n9870), .ZN(n9873) );
  INV_X1 U8141 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U8142 ( .A1(n9873), .A2(n6569), .ZN(n6570) );
  OAI21_X1 U8143 ( .B1(n9873), .B2(n9408), .A(n6570), .ZN(P2_U3520) );
  INV_X1 U8144 ( .A(n6571), .ZN(n6572) );
  NAND2_X1 U8145 ( .A1(n6572), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6573) );
  OAI211_X1 U8146 ( .C1(n9780), .C2(n6574), .A(n8161), .B(n6573), .ZN(n6576)
         );
  NAND2_X1 U8147 ( .A1(n6576), .A2(n6575), .ZN(n6591) );
  NAND2_X1 U8148 ( .A1(n6591), .A2(n8549), .ZN(n6611) );
  NAND2_X1 U8149 ( .A1(n6611), .A2(n6283), .ZN(n9711) );
  INV_X1 U8150 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6853) );
  NOR2_X1 U8151 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6853), .ZN(n6595) );
  MUX2_X1 U8152 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9863), .S(n8587), .Z(n8591)
         );
  NAND2_X1 U8153 ( .A1(n6735), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6589) );
  INV_X1 U8154 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U8155 ( .A1(n6604), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6585) );
  INV_X1 U8156 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6577) );
  MUX2_X1 U8157 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6577), .S(n6604), .Z(n6664)
         );
  NAND2_X1 U8158 ( .A1(n6603), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6584) );
  INV_X1 U8159 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6578) );
  MUX2_X1 U8160 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6578), .S(n6603), .Z(n6652)
         );
  NAND2_X1 U8161 ( .A1(n6601), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6583) );
  INV_X1 U8162 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6579) );
  MUX2_X1 U8163 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6579), .S(n6601), .Z(n6676)
         );
  NAND2_X1 U8164 ( .A1(n9419), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6582) );
  INV_X1 U8165 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6580) );
  MUX2_X1 U8166 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6580), .S(n9419), .Z(n9422)
         );
  INV_X1 U8167 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6581) );
  MUX2_X1 U8168 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6581), .S(n6598), .Z(n9410)
         );
  NAND3_X1 U8169 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9410), .ZN(n9409) );
  OAI21_X1 U8170 ( .B1(n9406), .B2(n6581), .A(n9409), .ZN(n9423) );
  NAND2_X1 U8171 ( .A1(n9422), .A2(n9423), .ZN(n9421) );
  NAND2_X1 U8172 ( .A1(n6582), .A2(n9421), .ZN(n6677) );
  NAND2_X1 U8173 ( .A1(n6676), .A2(n6677), .ZN(n6675) );
  NAND2_X1 U8174 ( .A1(n6583), .A2(n6675), .ZN(n6653) );
  NAND2_X1 U8175 ( .A1(n6652), .A2(n6653), .ZN(n6651) );
  NAND2_X1 U8176 ( .A1(n6584), .A2(n6651), .ZN(n6665) );
  NAND2_X1 U8177 ( .A1(n6664), .A2(n6665), .ZN(n6663) );
  NAND2_X1 U8178 ( .A1(n6585), .A2(n6663), .ZN(n8578) );
  MUX2_X1 U8179 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9860), .S(n8571), .Z(n8577)
         );
  NAND2_X1 U8180 ( .A1(n8578), .A2(n8577), .ZN(n8576) );
  OAI21_X1 U8181 ( .B1(n9860), .B2(n6586), .A(n8576), .ZN(n6725) );
  INV_X1 U8182 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9967) );
  MUX2_X1 U8183 ( .A(n9967), .B(P2_REG1_REG_7__SCAN_IN), .S(n6735), .Z(n6726)
         );
  INV_X1 U8184 ( .A(n6726), .ZN(n6587) );
  NAND2_X1 U8185 ( .A1(n6725), .A2(n6587), .ZN(n6588) );
  NAND2_X1 U8186 ( .A1(n6589), .A2(n6588), .ZN(n8592) );
  NAND2_X1 U8187 ( .A1(n8591), .A2(n8592), .ZN(n8590) );
  INV_X1 U8188 ( .A(n8590), .ZN(n6590) );
  AOI21_X1 U8189 ( .B1(n8587), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6590), .ZN(
        n6593) );
  INV_X1 U8190 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9865) );
  MUX2_X1 U8191 ( .A(n9865), .B(P2_REG1_REG_9__SCAN_IN), .S(n6770), .Z(n6592)
         );
  NOR2_X1 U8192 ( .A1(n6592), .A2(n6593), .ZN(n6780) );
  INV_X1 U8193 ( .A(n8467), .ZN(n7579) );
  OR2_X1 U8194 ( .A1(n6591), .A2(n7579), .ZN(n9713) );
  AOI211_X1 U8195 ( .C1(n6593), .C2(n6592), .A(n6780), .B(n9713), .ZN(n6594)
         );
  AOI211_X1 U8196 ( .C1(n9715), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n6595), .B(
        n6594), .ZN(n6614) );
  XOR2_X1 U8197 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6770), .Z(n6612) );
  INV_X1 U8198 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6596) );
  MUX2_X1 U8199 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6596), .S(n8571), .Z(n8574)
         );
  NAND2_X1 U8200 ( .A1(n6604), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6606) );
  INV_X1 U8201 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10016) );
  INV_X1 U8202 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9709) );
  INV_X1 U8203 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6597) );
  NOR3_X1 U8204 ( .A1(n10016), .A2(n9709), .A3(n9399), .ZN(n9397) );
  AOI21_X1 U8205 ( .B1(n6598), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9397), .ZN(
        n9417) );
  NAND2_X1 U8206 ( .A1(n9419), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6599) );
  OAI21_X1 U8207 ( .B1(n9419), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6599), .ZN(
        n9416) );
  NOR2_X1 U8208 ( .A1(n9417), .A2(n9416), .ZN(n9415) );
  AOI21_X1 U8209 ( .B1(n9419), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9415), .ZN(
        n6674) );
  NAND2_X1 U8210 ( .A1(n6601), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6600) );
  OAI21_X1 U8211 ( .B1(n6601), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6600), .ZN(
        n6673) );
  NOR2_X1 U8212 ( .A1(n6674), .A2(n6673), .ZN(n6672) );
  AOI21_X1 U8213 ( .B1(n6601), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6672), .ZN(
        n6650) );
  NAND2_X1 U8214 ( .A1(n6603), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6602) );
  OAI21_X1 U8215 ( .B1(n6603), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6602), .ZN(
        n6649) );
  NOR2_X1 U8216 ( .A1(n6650), .A2(n6649), .ZN(n6648) );
  AOI21_X1 U8217 ( .B1(n6603), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6648), .ZN(
        n6662) );
  OAI21_X1 U8218 ( .B1(n6604), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6606), .ZN(
        n6661) );
  NOR2_X1 U8219 ( .A1(n6662), .A2(n6661), .ZN(n6660) );
  INV_X1 U8220 ( .A(n6660), .ZN(n6605) );
  NAND2_X1 U8221 ( .A1(n6606), .A2(n6605), .ZN(n8573) );
  NAND2_X1 U8222 ( .A1(n8571), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U8223 ( .A1(n6735), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6608) );
  OAI21_X1 U8224 ( .B1(n6735), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6608), .ZN(
        n6731) );
  NAND2_X1 U8225 ( .A1(n8587), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6609) );
  OAI21_X1 U8226 ( .B1(n8587), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6609), .ZN(
        n8584) );
  NOR2_X1 U8227 ( .A1(n8585), .A2(n8584), .ZN(n8583) );
  NOR2_X1 U8228 ( .A1(n6283), .A2(n8467), .ZN(n6610) );
  OAI211_X1 U8229 ( .C1(n6612), .C2(n4619), .A(n9710), .B(n6769), .ZN(n6613)
         );
  OAI211_X1 U8230 ( .C1(n9711), .C2(n6774), .A(n6614), .B(n6613), .ZN(P2_U3254) );
  OAI21_X1 U8231 ( .B1(n6617), .B2(n6616), .A(n6615), .ZN(n6622) );
  MUX2_X1 U8232 ( .A(P1_STATE_REG_SCAN_IN), .B(n9452), .S(n6618), .Z(n6620) );
  AOI22_X1 U8233 ( .A1(n8980), .A2(n9025), .B1(n9438), .B2(n9023), .ZN(n6619)
         );
  OAI211_X1 U8234 ( .C1(n6926), .C2(n9010), .A(n6620), .B(n6619), .ZN(n6621)
         );
  AOI21_X1 U8235 ( .B1(n6622), .B2(n9002), .A(n6621), .ZN(n6623) );
  INV_X1 U8236 ( .A(n6623), .ZN(P1_U3216) );
  NOR2_X1 U8237 ( .A1(n6625), .A2(n6624), .ZN(n6627) );
  AOI22_X1 U8238 ( .A1(n6700), .A2(n5288), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n6694), .ZN(n6626) );
  AOI21_X1 U8239 ( .B1(n6627), .B2(n6626), .A(n6693), .ZN(n6628) );
  NAND2_X1 U8240 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7096) );
  OAI21_X1 U8241 ( .B1(n6628), .B2(n9575), .A(n7096), .ZN(n6629) );
  INV_X1 U8242 ( .A(n6629), .ZN(n6637) );
  NAND2_X1 U8243 ( .A1(n6700), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6632) );
  OAI21_X1 U8244 ( .B1(n6700), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6632), .ZN(
        n6633) );
  NOR2_X1 U8245 ( .A1(n6634), .A2(n6633), .ZN(n6699) );
  AOI211_X1 U8246 ( .C1(n6634), .C2(n6633), .A(n9587), .B(n6699), .ZN(n6635)
         );
  AOI21_X1 U8247 ( .B1(n9621), .B2(n6700), .A(n6635), .ZN(n6636) );
  OAI211_X1 U8248 ( .C1(n9631), .C2(n10043), .A(n6637), .B(n6636), .ZN(
        P1_U3251) );
  INV_X1 U8249 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6640) );
  OR2_X1 U8250 ( .A1(n6638), .A2(n9855), .ZN(n6639) );
  OAI21_X1 U8251 ( .B1(n9856), .B2(n6640), .A(n6639), .ZN(P2_U3454) );
  INV_X1 U8252 ( .A(n6641), .ZN(n6643) );
  INV_X1 U8253 ( .A(n9581), .ZN(n9052) );
  OAI222_X1 U8254 ( .A1(n7863), .A2(n6642), .B1(n7873), .B2(n6643), .C1(
        P1_U3084), .C2(n9052), .ZN(P1_U3338) );
  INV_X1 U8255 ( .A(n7909), .ZN(n7899) );
  OAI222_X1 U8256 ( .A1(n8475), .A2(n6644), .B1(n8478), .B2(n6643), .C1(
        P2_U3152), .C2(n7899), .ZN(P2_U3343) );
  XNOR2_X1 U8257 ( .A(n6809), .B(n6808), .ZN(n6647) );
  INV_X1 U8258 ( .A(n8541), .ZN(n8505) );
  INV_X1 U8259 ( .A(n8565), .ZN(n7383) );
  OAI22_X1 U8260 ( .A1(n7383), .A2(n9761), .B1(n7297), .B2(n9763), .ZN(n7305)
         );
  AOI22_X1 U8261 ( .A1(n8505), .A2(n7305), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6646) );
  INV_X1 U8262 ( .A(n9799), .ZN(n7299) );
  AOI22_X1 U8263 ( .A1(n7299), .A2(n8520), .B1(n8543), .B2(n7301), .ZN(n6645)
         );
  OAI211_X1 U8264 ( .C1(n6647), .C2(n8522), .A(n6646), .B(n6645), .ZN(P2_U3229) );
  INV_X1 U8265 ( .A(n9710), .ZN(n9414) );
  AOI211_X1 U8266 ( .C1(n6650), .C2(n6649), .A(n6648), .B(n9414), .ZN(n6659)
         );
  INV_X1 U8267 ( .A(n9713), .ZN(n9708) );
  OAI211_X1 U8268 ( .C1(n6653), .C2(n6652), .A(n9708), .B(n6651), .ZN(n6656)
         );
  NAND2_X1 U8269 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6827) );
  INV_X1 U8270 ( .A(n6827), .ZN(n6654) );
  AOI21_X1 U8271 ( .B1(n9715), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6654), .ZN(
        n6655) );
  OAI211_X1 U8272 ( .C1(n9711), .C2(n6657), .A(n6656), .B(n6655), .ZN(n6658)
         );
  OR2_X1 U8273 ( .A1(n6659), .A2(n6658), .ZN(P2_U3249) );
  AOI211_X1 U8274 ( .C1(n6662), .C2(n6661), .A(n6660), .B(n9414), .ZN(n6671)
         );
  OAI211_X1 U8275 ( .C1(n6665), .C2(n6664), .A(n9708), .B(n6663), .ZN(n6668)
         );
  AND2_X1 U8276 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6666) );
  AOI21_X1 U8277 ( .B1(n9715), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6666), .ZN(
        n6667) );
  OAI211_X1 U8278 ( .C1(n9711), .C2(n6669), .A(n6668), .B(n6667), .ZN(n6670)
         );
  OR2_X1 U8279 ( .A1(n6671), .A2(n6670), .ZN(P2_U3250) );
  AOI211_X1 U8280 ( .C1(n6674), .C2(n6673), .A(n6672), .B(n9414), .ZN(n6683)
         );
  OAI211_X1 U8281 ( .C1(n6677), .C2(n6676), .A(n9708), .B(n6675), .ZN(n6680)
         );
  NOR2_X1 U8282 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5875), .ZN(n6678) );
  AOI21_X1 U8283 ( .B1(n9715), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6678), .ZN(
        n6679) );
  OAI211_X1 U8284 ( .C1(n9711), .C2(n6681), .A(n6680), .B(n6679), .ZN(n6682)
         );
  OR2_X1 U8285 ( .A1(n6683), .A2(n6682), .ZN(P2_U3248) );
  OAI211_X1 U8286 ( .C1(n6686), .C2(n6685), .A(n6684), .B(n9002), .ZN(n6692)
         );
  INV_X1 U8287 ( .A(n9022), .ZN(n6689) );
  NAND2_X1 U8288 ( .A1(n8980), .A2(n9024), .ZN(n6688) );
  OAI211_X1 U8289 ( .C1(n6689), .C2(n8983), .A(n6688), .B(n6687), .ZN(n6690)
         );
  AOI21_X1 U8290 ( .B1(n5797), .B2(n6938), .A(n6690), .ZN(n6691) );
  OAI211_X1 U8291 ( .C1(n9452), .C2(n7082), .A(n6692), .B(n6691), .ZN(P1_U3228) );
  AOI22_X1 U8292 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9030), .B1(n9042), .B2(
        n5311), .ZN(n6695) );
  AOI21_X1 U8293 ( .B1(n6696), .B2(n6695), .A(n9029), .ZN(n6707) );
  AND2_X1 U8294 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7175) );
  NOR2_X1 U8295 ( .A1(n6697), .A2(n9030), .ZN(n6698) );
  AOI211_X1 U8296 ( .C1(n9571), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7175), .B(
        n6698), .ZN(n6706) );
  MUX2_X1 U8297 ( .A(n7142), .B(P1_REG2_REG_11__SCAN_IN), .S(n9042), .Z(n6701)
         );
  INV_X1 U8298 ( .A(n6701), .ZN(n6702) );
  NAND2_X1 U8299 ( .A1(n6702), .A2(n6703), .ZN(n9043) );
  OAI21_X1 U8300 ( .B1(n6703), .B2(n6702), .A(n9043), .ZN(n6704) );
  NAND2_X1 U8301 ( .A1(n6704), .A2(n9619), .ZN(n6705) );
  OAI211_X1 U8302 ( .C1(n6707), .C2(n9575), .A(n6706), .B(n6705), .ZN(P1_U3252) );
  INV_X1 U8303 ( .A(n9827), .ZN(n9839) );
  NAND2_X1 U8304 ( .A1(n7286), .A2(n6708), .ZN(n6709) );
  NAND2_X1 U8305 ( .A1(n6718), .A2(n6765), .ZN(n7987) );
  NAND2_X1 U8306 ( .A1(n6718), .A2(n9786), .ZN(n6711) );
  NAND2_X1 U8307 ( .A1(n7277), .A2(n6711), .ZN(n6712) );
  NAND2_X1 U8308 ( .A1(n7348), .A2(n6713), .ZN(n7972) );
  INV_X1 U8309 ( .A(n7348), .ZN(n8569) );
  NAND2_X1 U8310 ( .A1(n8569), .A2(n7336), .ZN(n7993) );
  NAND2_X1 U8311 ( .A1(n7972), .A2(n7993), .ZN(n8124) );
  NAND2_X1 U8312 ( .A1(n6712), .A2(n8124), .ZN(n7296) );
  OAI21_X1 U8313 ( .B1(n6712), .B2(n8124), .A(n7296), .ZN(n6723) );
  NAND2_X1 U8314 ( .A1(n7279), .A2(n9786), .ZN(n7281) );
  INV_X1 U8315 ( .A(n6266), .ZN(n9842) );
  AOI21_X1 U8316 ( .B1(n7281), .B2(n6713), .A(n9842), .ZN(n6714) );
  OR2_X1 U8317 ( .A1(n7281), .A2(n6713), .ZN(n7354) );
  NAND2_X1 U8318 ( .A1(n6714), .A2(n7354), .ZN(n7334) );
  OAI21_X1 U8319 ( .B1(n7336), .B2(n9850), .A(n7334), .ZN(n6722) );
  INV_X1 U8320 ( .A(n6723), .ZN(n7337) );
  INV_X1 U8321 ( .A(n8124), .ZN(n7981) );
  NAND2_X1 U8322 ( .A1(n6715), .A2(n7986), .ZN(n7978) );
  NAND2_X1 U8323 ( .A1(n7978), .A2(n7984), .ZN(n7283) );
  OAI21_X1 U8324 ( .B1(n7981), .B2(n6717), .A(n7303), .ZN(n6720) );
  OAI22_X1 U8325 ( .A1(n6718), .A2(n9763), .B1(n7297), .B2(n9761), .ZN(n6719)
         );
  AOI21_X1 U8326 ( .B1(n6720), .B2(n9766), .A(n6719), .ZN(n6721) );
  OAI21_X1 U8327 ( .B1(n7337), .B2(n9769), .A(n6721), .ZN(n7333) );
  AOI211_X1 U8328 ( .C1(n9839), .C2(n6723), .A(n6722), .B(n7333), .ZN(n6748)
         );
  NAND2_X1 U8329 ( .A1(n9870), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6724) );
  OAI21_X1 U8330 ( .B1(n6748), .B2(n9870), .A(n6724), .ZN(P2_U3523) );
  INV_X1 U8331 ( .A(n9711), .ZN(n9420) );
  XOR2_X1 U8332 ( .A(n6726), .B(n6725), .Z(n6729) );
  INV_X1 U8333 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6873) );
  NOR2_X1 U8334 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6873), .ZN(n6727) );
  AOI21_X1 U8335 ( .B1(n9715), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6727), .ZN(
        n6728) );
  OAI21_X1 U8336 ( .B1(n9713), .B2(n6729), .A(n6728), .ZN(n6734) );
  AOI211_X1 U8337 ( .C1(n6732), .C2(n6731), .A(n6730), .B(n9414), .ZN(n6733)
         );
  AOI211_X1 U8338 ( .C1(n9420), .C2(n6735), .A(n6734), .B(n6733), .ZN(n6736)
         );
  INV_X1 U8339 ( .A(n6736), .ZN(P2_U3252) );
  INV_X1 U8340 ( .A(n7902), .ZN(n8617) );
  INV_X1 U8341 ( .A(n6737), .ZN(n6739) );
  OAI222_X1 U8342 ( .A1(P2_U3152), .A2(n8617), .B1(n8478), .B2(n6739), .C1(
        n6738), .C2(n7837), .ZN(P2_U3342) );
  INV_X1 U8343 ( .A(n9593), .ZN(n9036) );
  OAI222_X1 U8344 ( .A1(n7863), .A2(n6740), .B1(n7873), .B2(n6739), .C1(n9036), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  NAND2_X1 U8345 ( .A1(n8515), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6764) );
  AOI22_X1 U8346 ( .A1(n6764), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n8528), .B2(
        n6557), .ZN(n6746) );
  INV_X1 U8347 ( .A(n8121), .ZN(n6742) );
  MUX2_X1 U8348 ( .A(n6742), .B(n7208), .S(n6741), .Z(n6743) );
  INV_X1 U8349 ( .A(n8522), .ZN(n8535) );
  OAI21_X1 U8350 ( .B1(n6744), .B2(n6743), .A(n8535), .ZN(n6745) );
  OAI211_X1 U8351 ( .C1(n8546), .C2(n6747), .A(n6746), .B(n6745), .ZN(P2_U3234) );
  INV_X1 U8352 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6750) );
  OR2_X1 U8353 ( .A1(n6748), .A2(n9855), .ZN(n6749) );
  OAI21_X1 U8354 ( .B1(n9856), .B2(n6750), .A(n6749), .ZN(P2_U3460) );
  INV_X1 U8355 ( .A(n6764), .ZN(n6758) );
  INV_X1 U8356 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9401) );
  AOI22_X1 U8357 ( .A1(n8527), .A2(n6751), .B1(n8528), .B2(n8570), .ZN(n6757)
         );
  OAI21_X1 U8358 ( .B1(n6754), .B2(n6753), .A(n6752), .ZN(n6755) );
  AOI22_X1 U8359 ( .A1(n8535), .A2(n6755), .B1(n8520), .B2(n7241), .ZN(n6756)
         );
  OAI211_X1 U8360 ( .C1(n6758), .C2(n9401), .A(n6757), .B(n6756), .ZN(P2_U3224) );
  NAND2_X1 U8361 ( .A1(n6752), .A2(n6759), .ZN(n6763) );
  NAND2_X1 U8362 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  XNOR2_X1 U8363 ( .A(n6763), .B(n6762), .ZN(n6768) );
  AOI22_X1 U8364 ( .A1(n6764), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8527), .B2(
        n6557), .ZN(n6767) );
  AOI22_X1 U8365 ( .A1(n8528), .A2(n8569), .B1(n6765), .B2(n8520), .ZN(n6766)
         );
  OAI211_X1 U8366 ( .C1(n8522), .C2(n6768), .A(n6767), .B(n6766), .ZN(P2_U3239) );
  NAND2_X1 U8367 ( .A1(n7151), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6771) );
  OAI21_X1 U8368 ( .B1(n7151), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6771), .ZN(
        n6772) );
  NOR2_X1 U8369 ( .A1(n6773), .A2(n6772), .ZN(n7150) );
  AOI211_X1 U8370 ( .C1(n6773), .C2(n6772), .A(n7150), .B(n9414), .ZN(n6784)
         );
  INV_X1 U8371 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9867) );
  MUX2_X1 U8372 ( .A(n9867), .B(P2_REG1_REG_10__SCAN_IN), .S(n7151), .Z(n6776)
         );
  NOR2_X1 U8373 ( .A1(n6774), .A2(n9865), .ZN(n6778) );
  INV_X1 U8374 ( .A(n6778), .ZN(n6775) );
  NAND2_X1 U8375 ( .A1(n6776), .A2(n6775), .ZN(n6779) );
  MUX2_X1 U8376 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9867), .S(n7151), .Z(n6777)
         );
  OAI21_X1 U8377 ( .B1(n6780), .B2(n6778), .A(n6777), .ZN(n7158) );
  OAI211_X1 U8378 ( .C1(n6780), .C2(n6779), .A(n9708), .B(n7158), .ZN(n6782)
         );
  AND2_X1 U8379 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n6967) );
  AOI21_X1 U8380 ( .B1(n9715), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6967), .ZN(
        n6781) );
  OAI211_X1 U8381 ( .C1(n9711), .C2(n7159), .A(n6782), .B(n6781), .ZN(n6783)
         );
  OR2_X1 U8382 ( .A1(n6784), .A2(n6783), .ZN(P2_U3255) );
  INV_X1 U8383 ( .A(n6785), .ZN(n6786) );
  INV_X1 U8384 ( .A(n9601), .ZN(n9038) );
  OAI222_X1 U8385 ( .A1(n7863), .A2(n10053), .B1(n7873), .B2(n6786), .C1(n9038), .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U8386 ( .A(n7915), .ZN(n8627) );
  OAI222_X1 U8387 ( .A1(n8475), .A2(n6787), .B1(n8478), .B2(n6786), .C1(n8627), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  XNOR2_X1 U8388 ( .A(n6789), .B(n6788), .ZN(n6790) );
  XNOR2_X1 U8389 ( .A(n6791), .B(n6790), .ZN(n6799) );
  NAND2_X1 U8390 ( .A1(n7029), .A2(n9443), .ZN(n9673) );
  INV_X1 U8391 ( .A(n9673), .ZN(n6796) );
  INV_X1 U8392 ( .A(n9268), .ZN(n9021) );
  NAND2_X1 U8393 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9520) );
  INV_X1 U8394 ( .A(n9520), .ZN(n6792) );
  AOI21_X1 U8395 ( .B1(n8980), .B2(n9021), .A(n6792), .ZN(n6794) );
  INV_X1 U8396 ( .A(n7046), .ZN(n9018) );
  NAND2_X1 U8397 ( .A1(n9438), .A2(n9018), .ZN(n6793) );
  OAI211_X1 U8398 ( .C1(n9452), .C2(n6956), .A(n6794), .B(n6793), .ZN(n6795)
         );
  AOI21_X1 U8399 ( .B1(n6797), .B2(n6796), .A(n6795), .ZN(n6798) );
  OAI21_X1 U8400 ( .B1(n6799), .B2(n9446), .A(n6798), .ZN(P1_U3211) );
  XNOR2_X1 U8401 ( .A(n6801), .B(n6800), .ZN(n6806) );
  INV_X1 U8402 ( .A(n9764), .ZN(n8564) );
  AOI22_X1 U8403 ( .A1(n8527), .A2(n8564), .B1(n8528), .B2(n8562), .ZN(n6802)
         );
  NAND2_X1 U8404 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8588) );
  OAI211_X1 U8405 ( .C1(n6803), .C2(n8515), .A(n6802), .B(n8588), .ZN(n6804)
         );
  AOI21_X1 U8406 ( .B1(n9770), .B2(n8520), .A(n6804), .ZN(n6805) );
  OAI21_X1 U8407 ( .B1(n6806), .B2(n8522), .A(n6805), .ZN(P2_U3223) );
  NOR2_X1 U8408 ( .A1(n6809), .A2(n6808), .ZN(n6812) );
  NOR2_X1 U8409 ( .A1(n6812), .A2(n6810), .ZN(n6814) );
  OR2_X1 U8410 ( .A1(n6812), .A2(n6811), .ZN(n6813) );
  OAI21_X1 U8411 ( .B1(n6815), .B2(n6814), .A(n6813), .ZN(n6821) );
  OAI22_X1 U8412 ( .A1(n8516), .A2(n9764), .B1(n9806), .B2(n8546), .ZN(n6820)
         );
  INV_X1 U8413 ( .A(n6816), .ZN(n8566) );
  NAND2_X1 U8414 ( .A1(n8527), .A2(n8566), .ZN(n6818) );
  INV_X1 U8415 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10019) );
  NOR2_X1 U8416 ( .A1(n10019), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8575) );
  INV_X1 U8417 ( .A(n8575), .ZN(n6817) );
  OAI211_X1 U8418 ( .C1(n8515), .C2(n8816), .A(n6818), .B(n6817), .ZN(n6819)
         );
  AOI211_X1 U8419 ( .C1(n6821), .C2(n8535), .A(n6820), .B(n6819), .ZN(n6822)
         );
  INV_X1 U8420 ( .A(n6822), .ZN(P2_U3241) );
  NOR2_X1 U8421 ( .A1(n6824), .A2(n4799), .ZN(n6825) );
  XNOR2_X1 U8422 ( .A(n6826), .B(n6825), .ZN(n6832) );
  INV_X1 U8423 ( .A(n7359), .ZN(n6828) );
  OAI21_X1 U8424 ( .B1(n8515), .B2(n6828), .A(n6827), .ZN(n6830) );
  INV_X1 U8425 ( .A(n7358), .ZN(n9792) );
  OAI22_X1 U8426 ( .A1(n8516), .A2(n6816), .B1(n9792), .B2(n8546), .ZN(n6829)
         );
  AOI211_X1 U8427 ( .C1(n8527), .C2(n8569), .A(n6830), .B(n6829), .ZN(n6831)
         );
  OAI21_X1 U8428 ( .B1(n6832), .B2(n8522), .A(n6831), .ZN(P2_U3232) );
  XNOR2_X1 U8429 ( .A(n6835), .B(n6834), .ZN(n6836) );
  XNOR2_X1 U8430 ( .A(n6833), .B(n6836), .ZN(n6843) );
  INV_X1 U8431 ( .A(n7032), .ZN(n6841) );
  INV_X1 U8432 ( .A(n9017), .ZN(n7043) );
  INV_X1 U8433 ( .A(n6943), .ZN(n9020) );
  NAND2_X1 U8434 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9535) );
  INV_X1 U8435 ( .A(n9535), .ZN(n6837) );
  AOI21_X1 U8436 ( .B1(n8980), .B2(n9020), .A(n6837), .ZN(n6838) );
  OAI21_X1 U8437 ( .B1(n7043), .B2(n8983), .A(n6838), .ZN(n6840) );
  NAND2_X1 U8438 ( .A1(n7044), .A2(n9443), .ZN(n9678) );
  NOR2_X1 U8439 ( .A1(n9678), .A2(n9445), .ZN(n6839) );
  AOI211_X1 U8440 ( .C1(n6841), .C2(n9003), .A(n6840), .B(n6839), .ZN(n6842)
         );
  OAI21_X1 U8441 ( .B1(n6843), .B2(n9446), .A(n6842), .ZN(P1_U3219) );
  INV_X1 U8442 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6845) );
  INV_X1 U8443 ( .A(n6844), .ZN(n6846) );
  INV_X1 U8444 ( .A(n8640), .ZN(n7920) );
  OAI222_X1 U8445 ( .A1(n8475), .A2(n6845), .B1(n8478), .B2(n6846), .C1(
        P2_U3152), .C2(n7920), .ZN(P2_U3340) );
  INV_X1 U8446 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6847) );
  INV_X1 U8447 ( .A(n9620), .ZN(n9040) );
  OAI222_X1 U8448 ( .A1(n7863), .A2(n6847), .B1(n7873), .B2(n6846), .C1(
        P1_U3084), .C2(n9040), .ZN(P1_U3335) );
  XNOR2_X1 U8449 ( .A(n6850), .B(n6849), .ZN(n6851) );
  XNOR2_X1 U8450 ( .A(n6848), .B(n6851), .ZN(n6858) );
  OR2_X1 U8451 ( .A1(n7384), .A2(n9763), .ZN(n6852) );
  OAI21_X1 U8452 ( .B1(n7367), .B2(n9761), .A(n6852), .ZN(n7328) );
  INV_X1 U8453 ( .A(n7328), .ZN(n6854) );
  OAI22_X1 U8454 ( .A1(n8541), .A2(n6854), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6853), .ZN(n6856) );
  INV_X1 U8455 ( .A(n9823), .ZN(n7322) );
  NOR2_X1 U8456 ( .A1(n8546), .A2(n7322), .ZN(n6855) );
  AOI211_X1 U8457 ( .C1(n8543), .C2(n7320), .A(n6856), .B(n6855), .ZN(n6857)
         );
  OAI21_X1 U8458 ( .B1(n6858), .B2(n8522), .A(n6857), .ZN(P2_U3233) );
  INV_X1 U8459 ( .A(n6859), .ZN(n6861) );
  NAND2_X1 U8460 ( .A1(n6861), .A2(n6860), .ZN(n6914) );
  OAI21_X1 U8461 ( .B1(n6861), .B2(n6860), .A(n6914), .ZN(n6862) );
  NOR2_X1 U8462 ( .A1(n6862), .A2(n6863), .ZN(n6916) );
  AOI21_X1 U8463 ( .B1(n6863), .B2(n6862), .A(n6916), .ZN(n6870) );
  INV_X1 U8464 ( .A(n9663), .ZN(n9279) );
  INV_X1 U8465 ( .A(n6864), .ZN(n6865) );
  AOI21_X1 U8466 ( .B1(n8980), .B2(n9023), .A(n6865), .ZN(n6867) );
  NAND2_X1 U8467 ( .A1(n9438), .A2(n9021), .ZN(n6866) );
  OAI211_X1 U8468 ( .C1(n9452), .C2(n9273), .A(n6867), .B(n6866), .ZN(n6868)
         );
  AOI21_X1 U8469 ( .B1(n5797), .B2(n9279), .A(n6868), .ZN(n6869) );
  OAI21_X1 U8470 ( .B1(n6870), .B2(n9446), .A(n6869), .ZN(P1_U3225) );
  XNOR2_X1 U8471 ( .A(n6872), .B(n6871), .ZN(n6878) );
  INV_X1 U8472 ( .A(n7387), .ZN(n6874) );
  OAI22_X1 U8473 ( .A1(n8515), .A2(n6874), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6873), .ZN(n6876) );
  OAI22_X1 U8474 ( .A1(n7383), .A2(n8517), .B1(n8516), .B2(n7384), .ZN(n6875)
         );
  AOI211_X1 U8475 ( .C1(n9810), .C2(n8520), .A(n6876), .B(n6875), .ZN(n6877)
         );
  OAI21_X1 U8476 ( .B1(n6878), .B2(n8522), .A(n6877), .ZN(P2_U3215) );
  NAND3_X1 U8477 ( .A1(n9633), .A2(n9366), .A3(n9275), .ZN(n9274) );
  INV_X1 U8478 ( .A(n9274), .ZN(n9254) );
  AND2_X1 U8479 ( .A1(n6888), .A2(n6904), .ZN(n6879) );
  NAND2_X1 U8480 ( .A1(n6884), .A2(n6879), .ZN(n7001) );
  OAI21_X1 U8481 ( .B1(n6884), .B2(n6879), .A(n7001), .ZN(n9637) );
  OR2_X1 U8482 ( .A1(n6880), .A2(n6988), .ZN(n6883) );
  OR2_X1 U8483 ( .A1(n6881), .A2(n8267), .ZN(n6882) );
  AND2_X1 U8484 ( .A1(n6883), .A2(n6882), .ZN(n9295) );
  XNOR2_X1 U8485 ( .A(n4643), .B(n6947), .ZN(n6886) );
  NAND2_X1 U8486 ( .A1(n8445), .A2(n9275), .ZN(n6885) );
  NAND2_X1 U8487 ( .A1(n5766), .A2(n8436), .ZN(n8439) );
  AND2_X1 U8488 ( .A1(n6885), .A2(n8439), .ZN(n9265) );
  INV_X1 U8489 ( .A(n9265), .ZN(n9223) );
  NAND2_X1 U8490 ( .A1(n6886), .A2(n9223), .ZN(n6890) );
  INV_X1 U8491 ( .A(n6887), .ZN(n8431) );
  AND2_X1 U8492 ( .A1(n8431), .A2(n9500), .ZN(n9220) );
  AOI22_X1 U8493 ( .A1(n9220), .A2(n6888), .B1(n9025), .B2(n9218), .ZN(n6889)
         );
  OAI211_X1 U8494 ( .C1(n9637), .C2(n9295), .A(n6890), .B(n6889), .ZN(n9641)
         );
  OAI21_X1 U8495 ( .B1(n9640), .B2(n6891), .A(n9366), .ZN(n6892) );
  NOR2_X1 U8496 ( .A1(n6932), .A2(n6904), .ZN(n7012) );
  NOR2_X1 U8497 ( .A1(n6892), .A2(n7012), .ZN(n9638) );
  NOR2_X1 U8498 ( .A1(n9637), .A2(n6893), .ZN(n6894) );
  MUX2_X1 U8499 ( .A(n9638), .B(n6894), .S(n9275), .Z(n6895) );
  AOI211_X1 U8500 ( .C1(n9254), .C2(P1_REG3_REG_1__SCAN_IN), .A(n9641), .B(
        n6895), .ZN(n6903) );
  NAND3_X1 U8501 ( .A1(n6898), .A2(n6897), .A3(n6896), .ZN(n6900) );
  OR2_X1 U8502 ( .A1(n6900), .A2(n6899), .ZN(n6955) );
  INV_X1 U8503 ( .A(n9276), .ZN(n9253) );
  INV_X1 U8504 ( .A(n9276), .ZN(n9278) );
  AOI22_X1 U8505 ( .A1(n9280), .A2(n6932), .B1(n9278), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6902) );
  OAI21_X1 U8506 ( .B1(n6903), .B2(n9253), .A(n6902), .ZN(P1_U3290) );
  AOI22_X1 U8507 ( .A1(n9278), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9254), .ZN(n6906) );
  AND2_X1 U8508 ( .A1(n9276), .A2(n6909), .ZN(n9252) );
  AND2_X1 U8509 ( .A1(n9252), .A2(n9366), .ZN(n9226) );
  OAI21_X1 U8510 ( .B1(n9226), .B2(n9280), .A(n6904), .ZN(n6905) );
  OAI211_X1 U8511 ( .C1(n6907), .C2(n9253), .A(n6906), .B(n6905), .ZN(P1_U3291) );
  INV_X1 U8512 ( .A(n6908), .ZN(n6911) );
  OAI222_X1 U8513 ( .A1(n7863), .A2(n6910), .B1(n7873), .B2(n6911), .C1(n6909), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8514 ( .A1(n8475), .A2(n9924), .B1(n8478), .B2(n6911), .C1(
        P2_U3152), .C2(n8707), .ZN(P2_U3339) );
  NAND2_X1 U8515 ( .A1(n6913), .A2(n6912), .ZN(n6918) );
  INV_X1 U8516 ( .A(n6914), .ZN(n6915) );
  NOR2_X1 U8517 ( .A1(n6916), .A2(n6915), .ZN(n6917) );
  XOR2_X1 U8518 ( .A(n6918), .B(n6917), .Z(n6925) );
  INV_X1 U8519 ( .A(n6919), .ZN(n6920) );
  AOI21_X1 U8520 ( .B1(n8980), .B2(n9022), .A(n6920), .ZN(n6922) );
  NAND2_X1 U8521 ( .A1(n9438), .A2(n9020), .ZN(n6921) );
  OAI211_X1 U8522 ( .C1(n9452), .C2(n7062), .A(n6922), .B(n6921), .ZN(n6923)
         );
  AOI21_X1 U8523 ( .B1(n5797), .B2(n7064), .A(n6923), .ZN(n6924) );
  OAI21_X1 U8524 ( .B1(n6925), .B2(n9446), .A(n6924), .ZN(P1_U3237) );
  NAND2_X1 U8525 ( .A1(n9024), .A2(n6926), .ZN(n8199) );
  OR2_X1 U8526 ( .A1(n6927), .A2(n9024), .ZN(n6935) );
  NAND2_X1 U8527 ( .A1(n8240), .A2(n6935), .ZN(n7076) );
  INV_X1 U8528 ( .A(n9023), .ZN(n9266) );
  NAND2_X1 U8529 ( .A1(n6938), .A2(n9266), .ZN(n8313) );
  AND3_X1 U8530 ( .A1(n6930), .A2(n6929), .A3(n6928), .ZN(n6931) );
  NAND2_X1 U8531 ( .A1(n6931), .A2(n9023), .ZN(n8307) );
  NAND2_X1 U8532 ( .A1(n8313), .A2(n8307), .ZN(n7077) );
  AND2_X1 U8533 ( .A1(n7076), .A2(n7077), .ZN(n6937) );
  NAND2_X1 U8534 ( .A1(n9025), .A2(n9645), .ZN(n8195) );
  NAND2_X1 U8535 ( .A1(n8193), .A2(n8195), .ZN(n6933) );
  NAND2_X1 U8536 ( .A1(n9027), .A2(n6932), .ZN(n7000) );
  AND2_X1 U8537 ( .A1(n6933), .A2(n7000), .ZN(n6934) );
  NAND2_X1 U8538 ( .A1(n7001), .A2(n6934), .ZN(n7002) );
  OR2_X1 U8539 ( .A1(n9025), .A2(n7015), .ZN(n6986) );
  AND2_X1 U8540 ( .A1(n6935), .A2(n6986), .ZN(n6936) );
  NAND2_X1 U8541 ( .A1(n7002), .A2(n6936), .ZN(n7075) );
  NAND2_X1 U8542 ( .A1(n6937), .A2(n7075), .ZN(n6940) );
  OR2_X1 U8543 ( .A1(n9023), .A2(n6938), .ZN(n6939) );
  OR2_X1 U8544 ( .A1(n9022), .A2(n9663), .ZN(n7066) );
  NAND2_X1 U8545 ( .A1(n9663), .A2(n9022), .ZN(n8308) );
  AND2_X1 U8546 ( .A1(n7066), .A2(n8308), .ZN(n9281) );
  OR2_X1 U8547 ( .A1(n7064), .A2(n9268), .ZN(n8203) );
  NAND2_X1 U8548 ( .A1(n7064), .A2(n9268), .ZN(n8316) );
  NAND2_X1 U8549 ( .A1(n8203), .A2(n8316), .ZN(n8238) );
  OR2_X1 U8550 ( .A1(n7064), .A2(n9021), .ZN(n6942) );
  NAND2_X1 U8551 ( .A1(n7058), .A2(n6942), .ZN(n7028) );
  OR2_X1 U8552 ( .A1(n7029), .A2(n6943), .ZN(n8320) );
  NAND2_X1 U8553 ( .A1(n7029), .A2(n6943), .ZN(n8322) );
  NAND2_X1 U8554 ( .A1(n8320), .A2(n8322), .ZN(n8239) );
  XNOR2_X1 U8555 ( .A(n7028), .B(n8239), .ZN(n9677) );
  INV_X1 U8556 ( .A(n9677), .ZN(n6962) );
  AND2_X1 U8557 ( .A1(n6945), .A2(n6944), .ZN(n6946) );
  NAND2_X1 U8558 ( .A1(n9276), .A2(n6946), .ZN(n9262) );
  INV_X1 U8559 ( .A(n9220), .ZN(n9267) );
  OR2_X1 U8560 ( .A1(n9027), .A2(n9640), .ZN(n6948) );
  AND2_X1 U8561 ( .A1(n8193), .A2(n8195), .ZN(n8241) );
  NAND2_X1 U8562 ( .A1(n7005), .A2(n8193), .ZN(n8276) );
  INV_X1 U8563 ( .A(n8313), .ZN(n6949) );
  AND2_X1 U8564 ( .A1(n8316), .A2(n7066), .ZN(n8201) );
  INV_X1 U8565 ( .A(n8308), .ZN(n7067) );
  NAND2_X1 U8566 ( .A1(n8316), .A2(n7067), .ZN(n8318) );
  AND2_X1 U8567 ( .A1(n8318), .A2(n8203), .ZN(n6950) );
  INV_X1 U8568 ( .A(n7024), .ZN(n6951) );
  AOI21_X1 U8569 ( .B1(n8239), .B2(n6952), .A(n6951), .ZN(n6953) );
  OAI222_X1 U8570 ( .A1(n9267), .A2(n9268), .B1(n9269), .B2(n7046), .C1(n9265), 
        .C2(n6953), .ZN(n9675) );
  NAND2_X1 U8571 ( .A1(n7012), .A2(n9645), .ZN(n7011) );
  INV_X1 U8572 ( .A(n7064), .ZN(n9667) );
  NAND2_X1 U8573 ( .A1(n9270), .A2(n9667), .ZN(n7061) );
  INV_X1 U8574 ( .A(n9366), .ZN(n9688) );
  AOI21_X1 U8575 ( .B1(n7061), .B2(n7029), .A(n9688), .ZN(n6954) );
  NAND2_X1 U8576 ( .A1(n6954), .A2(n7034), .ZN(n9674) );
  NOR2_X1 U8577 ( .A1(n6955), .A2(n9275), .ZN(n7635) );
  INV_X1 U8578 ( .A(n7635), .ZN(n7450) );
  OAI22_X1 U8579 ( .A1(n9276), .A2(n6957), .B1(n6956), .B2(n9274), .ZN(n6958)
         );
  AOI21_X1 U8580 ( .B1(n7029), .B2(n9280), .A(n6958), .ZN(n6959) );
  OAI21_X1 U8581 ( .B1(n9674), .B2(n7450), .A(n6959), .ZN(n6960) );
  AOI21_X1 U8582 ( .B1(n9675), .B2(n9276), .A(n6960), .ZN(n6961) );
  OAI21_X1 U8583 ( .B1(n6962), .B2(n9262), .A(n6961), .ZN(P1_U3284) );
  INV_X1 U8584 ( .A(n7434), .ZN(n9834) );
  OAI211_X1 U8585 ( .C1(n6965), .C2(n6964), .A(n6963), .B(n8535), .ZN(n6969)
         );
  OAI22_X1 U8586 ( .A1(n7455), .A2(n8516), .B1(n8517), .B2(n9762), .ZN(n6966)
         );
  AOI211_X1 U8587 ( .C1(n7427), .C2(n8543), .A(n6967), .B(n6966), .ZN(n6968)
         );
  OAI211_X1 U8588 ( .C1(n9834), .C2(n8546), .A(n6969), .B(n6968), .ZN(P2_U3219) );
  INV_X1 U8589 ( .A(n6971), .ZN(n6972) );
  AOI21_X1 U8590 ( .B1(n6973), .B2(n6970), .A(n6972), .ZN(n6979) );
  NOR2_X1 U8591 ( .A1(n8983), .A2(n7177), .ZN(n6974) );
  AOI211_X1 U8592 ( .C1(n8980), .C2(n9018), .A(n6975), .B(n6974), .ZN(n6976)
         );
  OAI21_X1 U8593 ( .B1(n9452), .B2(n7050), .A(n6976), .ZN(n6977) );
  AOI21_X1 U8594 ( .B1(n5797), .B2(n7103), .A(n6977), .ZN(n6978) );
  OAI21_X1 U8595 ( .B1(n6979), .B2(n9446), .A(n6978), .ZN(P1_U3229) );
  INV_X1 U8596 ( .A(n9116), .ZN(n6984) );
  INV_X1 U8597 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U8598 ( .A1(n5017), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6981) );
  INV_X1 U8599 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10107) );
  OR2_X1 U8600 ( .A1(n5100), .A2(n10107), .ZN(n6980) );
  OAI211_X1 U8601 ( .C1(n8172), .C2(n9952), .A(n6981), .B(n6980), .ZN(n6982)
         );
  AOI21_X1 U8602 ( .B1(n6984), .B2(n6983), .A(n6982), .ZN(n9129) );
  NAND2_X1 U8603 ( .A1(n9026), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6985) );
  OAI21_X1 U8604 ( .B1(n9129), .B2(n9026), .A(n6985), .ZN(P1_U3584) );
  NAND2_X1 U8605 ( .A1(n7002), .A2(n6986), .ZN(n6987) );
  XNOR2_X1 U8606 ( .A(n6987), .B(n8240), .ZN(n9650) );
  AND2_X1 U8607 ( .A1(n6988), .A2(n9275), .ZN(n6989) );
  AND2_X1 U8608 ( .A1(n9276), .A2(n6989), .ZN(n7659) );
  INV_X1 U8609 ( .A(n7659), .ZN(n7090) );
  AOI22_X1 U8610 ( .A1(n9220), .A2(n9025), .B1(n9023), .B2(n9218), .ZN(n6993)
         );
  OAI21_X1 U8611 ( .B1(n8240), .B2(n8276), .A(n6990), .ZN(n6991) );
  NAND2_X1 U8612 ( .A1(n6991), .A2(n9223), .ZN(n6992) );
  OAI211_X1 U8613 ( .C1(n9650), .C2(n9295), .A(n6993), .B(n6992), .ZN(n9652)
         );
  NAND2_X1 U8614 ( .A1(n9652), .A2(n9276), .ZN(n6999) );
  OAI22_X1 U8615 ( .A1(n9276), .A2(n6994), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9274), .ZN(n6997) );
  INV_X1 U8616 ( .A(n9226), .ZN(n9163) );
  NAND2_X1 U8617 ( .A1(n7011), .A2(n6927), .ZN(n6995) );
  NAND2_X1 U8618 ( .A1(n7084), .A2(n6995), .ZN(n9651) );
  NOR2_X1 U8619 ( .A1(n9163), .A2(n9651), .ZN(n6996) );
  AOI211_X1 U8620 ( .C1(n9280), .C2(n6927), .A(n6997), .B(n6996), .ZN(n6998)
         );
  OAI211_X1 U8621 ( .C1(n9650), .C2(n7090), .A(n6999), .B(n6998), .ZN(P1_U3288) );
  NAND2_X1 U8622 ( .A1(n7001), .A2(n7000), .ZN(n7004) );
  INV_X1 U8623 ( .A(n7002), .ZN(n7003) );
  AOI21_X1 U8624 ( .B1(n8241), .B2(n7004), .A(n7003), .ZN(n9644) );
  AOI22_X1 U8625 ( .A1(n9220), .A2(n9027), .B1(n9024), .B2(n9218), .ZN(n7008)
         );
  OAI21_X1 U8626 ( .B1(n8241), .B2(n8197), .A(n7005), .ZN(n7006) );
  NAND2_X1 U8627 ( .A1(n7006), .A2(n9223), .ZN(n7007) );
  OAI211_X1 U8628 ( .C1(n9644), .C2(n9295), .A(n7008), .B(n7007), .ZN(n9647)
         );
  NAND2_X1 U8629 ( .A1(n9647), .A2(n9276), .ZN(n7017) );
  OAI22_X1 U8630 ( .A1(n9276), .A2(n7010), .B1(n7009), .B2(n9274), .ZN(n7014)
         );
  OAI21_X1 U8631 ( .B1(n7012), .B2(n9645), .A(n7011), .ZN(n9646) );
  NOR2_X1 U8632 ( .A1(n9163), .A2(n9646), .ZN(n7013) );
  AOI211_X1 U8633 ( .C1(n9280), .C2(n7015), .A(n7014), .B(n7013), .ZN(n7016)
         );
  OAI211_X1 U8634 ( .C1(n9644), .C2(n7090), .A(n7017), .B(n7016), .ZN(P1_U3289) );
  INV_X1 U8635 ( .A(n7018), .ZN(n7022) );
  OAI222_X1 U8636 ( .A1(P1_U3084), .A2(n7020), .B1(n7873), .B2(n7022), .C1(
        n7019), .C2(n7863), .ZN(P1_U3333) );
  OAI222_X1 U8637 ( .A1(n8475), .A2(n9936), .B1(n8478), .B2(n7022), .C1(n7021), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OR2_X1 U8638 ( .A1(n7044), .A2(n7046), .ZN(n8208) );
  NAND2_X1 U8639 ( .A1(n7044), .A2(n7046), .ZN(n8329) );
  INV_X1 U8640 ( .A(n8322), .ZN(n8310) );
  NOR2_X1 U8641 ( .A1(n4936), .A2(n8310), .ZN(n7023) );
  NAND2_X1 U8642 ( .A1(n7024), .A2(n7023), .ZN(n7045) );
  NAND2_X1 U8643 ( .A1(n7045), .A2(n9223), .ZN(n7027) );
  AOI21_X1 U8644 ( .B1(n7024), .B2(n8322), .A(n8245), .ZN(n7026) );
  AOI22_X1 U8645 ( .A1(n9020), .A2(n9220), .B1(n9218), .B2(n9017), .ZN(n7025)
         );
  OAI21_X1 U8646 ( .B1(n7027), .B2(n7026), .A(n7025), .ZN(n9681) );
  INV_X1 U8647 ( .A(n9681), .ZN(n7042) );
  OR2_X1 U8648 ( .A1(n7029), .A2(n9020), .ZN(n7030) );
  AOI21_X1 U8649 ( .B1(n8245), .B2(n7031), .A(n4470), .ZN(n9683) );
  INV_X1 U8650 ( .A(n9262), .ZN(n9283) );
  NAND2_X1 U8651 ( .A1(n9683), .A2(n9283), .ZN(n7041) );
  OAI22_X1 U8652 ( .A1(n9276), .A2(n7033), .B1(n7032), .B2(n9274), .ZN(n7039)
         );
  INV_X1 U8653 ( .A(n7044), .ZN(n7037) );
  INV_X1 U8654 ( .A(n7034), .ZN(n7036) );
  NOR2_X1 U8655 ( .A1(n7034), .A2(n7044), .ZN(n7052) );
  INV_X1 U8656 ( .A(n7052), .ZN(n7035) );
  OAI21_X1 U8657 ( .B1(n7037), .B2(n7036), .A(n7035), .ZN(n9679) );
  NOR2_X1 U8658 ( .A1(n9679), .A2(n9163), .ZN(n7038) );
  AOI211_X1 U8659 ( .C1(n9280), .C2(n7044), .A(n7039), .B(n7038), .ZN(n7040)
         );
  OAI211_X1 U8660 ( .C1(n9278), .C2(n7042), .A(n7041), .B(n7040), .ZN(P1_U3283) );
  OR2_X1 U8661 ( .A1(n7103), .A2(n7043), .ZN(n7131) );
  NAND2_X1 U8662 ( .A1(n7103), .A2(n7043), .ZN(n8330) );
  AND2_X1 U8663 ( .A1(n7131), .A2(n8330), .ZN(n8250) );
  XOR2_X1 U8664 ( .A(n8250), .B(n7106), .Z(n9685) );
  XNOR2_X1 U8665 ( .A(n7134), .B(n8250), .ZN(n7048) );
  OAI22_X1 U8666 ( .A1(n7177), .A2(n9269), .B1(n7046), .B2(n9267), .ZN(n7047)
         );
  AOI21_X1 U8667 ( .B1(n7048), .B2(n9223), .A(n7047), .ZN(n7049) );
  OAI21_X1 U8668 ( .B1(n9685), .B2(n9295), .A(n7049), .ZN(n9690) );
  NAND2_X1 U8669 ( .A1(n9690), .A2(n9276), .ZN(n7057) );
  OAI22_X1 U8670 ( .A1(n9276), .A2(n7051), .B1(n7050), .B2(n9274), .ZN(n7055)
         );
  INV_X1 U8671 ( .A(n7103), .ZN(n9687) );
  NOR2_X1 U8672 ( .A1(n7052), .A2(n9687), .ZN(n7053) );
  OR2_X1 U8673 ( .A1(n7114), .A2(n7053), .ZN(n9689) );
  NOR2_X1 U8674 ( .A1(n9689), .A2(n9163), .ZN(n7054) );
  AOI211_X1 U8675 ( .C1(n9280), .C2(n7103), .A(n7055), .B(n7054), .ZN(n7056)
         );
  OAI211_X1 U8676 ( .C1(n9685), .C2(n7090), .A(n7057), .B(n7056), .ZN(P1_U3282) );
  OAI21_X1 U8677 ( .B1(n7059), .B2(n8238), .A(n7058), .ZN(n9671) );
  OR2_X1 U8678 ( .A1(n9270), .A2(n9667), .ZN(n7060) );
  NAND2_X1 U8679 ( .A1(n7061), .A2(n7060), .ZN(n9668) );
  INV_X1 U8680 ( .A(n7062), .ZN(n7063) );
  AOI22_X1 U8681 ( .A1(n9280), .A2(n7064), .B1(n9254), .B2(n7063), .ZN(n7065)
         );
  OAI21_X1 U8682 ( .B1(n9668), .B2(n9163), .A(n7065), .ZN(n7073) );
  OAI21_X1 U8683 ( .B1(n9263), .B2(n7067), .A(n7066), .ZN(n7068) );
  XNOR2_X1 U8684 ( .A(n7068), .B(n8238), .ZN(n7071) );
  INV_X1 U8685 ( .A(n9295), .ZN(n7139) );
  NAND2_X1 U8686 ( .A1(n9671), .A2(n7139), .ZN(n7070) );
  AOI22_X1 U8687 ( .A1(n9020), .A2(n9218), .B1(n9220), .B2(n9022), .ZN(n7069)
         );
  OAI211_X1 U8688 ( .C1(n9265), .C2(n7071), .A(n7070), .B(n7069), .ZN(n9669)
         );
  MUX2_X1 U8689 ( .A(n9669), .B(P1_REG2_REG_6__SCAN_IN), .S(n9278), .Z(n7072)
         );
  AOI211_X1 U8690 ( .C1(n7659), .C2(n9671), .A(n7073), .B(n7072), .ZN(n7074)
         );
  INV_X1 U8691 ( .A(n7074), .ZN(P1_U3285) );
  AND2_X1 U8692 ( .A1(n7076), .A2(n7075), .ZN(n7078) );
  XNOR2_X1 U8693 ( .A(n7078), .B(n7077), .ZN(n9658) );
  INV_X1 U8694 ( .A(n9658), .ZN(n7091) );
  XNOR2_X1 U8695 ( .A(n8304), .B(n7077), .ZN(n7081) );
  NAND2_X1 U8696 ( .A1(n9658), .A2(n7139), .ZN(n7080) );
  AOI22_X1 U8697 ( .A1(n9220), .A2(n9024), .B1(n9022), .B2(n9218), .ZN(n7079)
         );
  OAI211_X1 U8698 ( .C1(n9265), .C2(n7081), .A(n7080), .B(n7079), .ZN(n9656)
         );
  NAND2_X1 U8699 ( .A1(n9656), .A2(n9276), .ZN(n7089) );
  OAI22_X1 U8700 ( .A1(n9276), .A2(n7083), .B1(n7082), .B2(n9274), .ZN(n7087)
         );
  AND2_X1 U8701 ( .A1(n7084), .A2(n6938), .ZN(n7085) );
  OR2_X1 U8702 ( .A1(n7085), .A2(n9272), .ZN(n9655) );
  NOR2_X1 U8703 ( .A1(n9655), .A2(n9163), .ZN(n7086) );
  AOI211_X1 U8704 ( .C1(n9280), .C2(n6938), .A(n7087), .B(n7086), .ZN(n7088)
         );
  OAI211_X1 U8705 ( .C1(n7091), .C2(n7090), .A(n7089), .B(n7088), .ZN(P1_U3287) );
  NAND2_X1 U8706 ( .A1(n7094), .A2(n7093), .ZN(n7095) );
  XNOR2_X1 U8707 ( .A(n7092), .B(n7095), .ZN(n7102) );
  INV_X1 U8708 ( .A(n7096), .ZN(n7097) );
  AOI21_X1 U8709 ( .B1(n8980), .B2(n9017), .A(n7097), .ZN(n7099) );
  NAND2_X1 U8710 ( .A1(n9438), .A2(n9016), .ZN(n7098) );
  OAI211_X1 U8711 ( .C1(n9452), .C2(n7115), .A(n7099), .B(n7098), .ZN(n7100)
         );
  AOI21_X1 U8712 ( .B1(n5797), .B2(n7128), .A(n7100), .ZN(n7101) );
  OAI21_X1 U8713 ( .B1(n7102), .B2(n9446), .A(n7101), .ZN(P1_U3215) );
  OR2_X1 U8714 ( .A1(n7103), .A2(n9017), .ZN(n7105) );
  AND2_X1 U8715 ( .A1(n7103), .A2(n9017), .ZN(n7104) );
  AOI21_X1 U8716 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n7107) );
  OR2_X1 U8717 ( .A1(n7128), .A2(n7177), .ZN(n7132) );
  NAND2_X1 U8718 ( .A1(n7128), .A2(n7177), .ZN(n8331) );
  NAND2_X1 U8719 ( .A1(n7132), .A2(n8331), .ZN(n8246) );
  NAND2_X1 U8720 ( .A1(n7107), .A2(n8246), .ZN(n7130) );
  OR2_X1 U8721 ( .A1(n7107), .A2(n8246), .ZN(n7108) );
  NAND2_X1 U8722 ( .A1(n7130), .A2(n7108), .ZN(n9430) );
  NAND2_X1 U8723 ( .A1(n7134), .A2(n7131), .ZN(n7109) );
  NAND2_X1 U8724 ( .A1(n7109), .A2(n8330), .ZN(n7110) );
  XNOR2_X1 U8725 ( .A(n7110), .B(n8246), .ZN(n7112) );
  AOI22_X1 U8726 ( .A1(n9220), .A2(n9017), .B1(n9016), .B2(n9218), .ZN(n7111)
         );
  OAI21_X1 U8727 ( .B1(n7112), .B2(n9265), .A(n7111), .ZN(n7113) );
  AOI21_X1 U8728 ( .B1(n9430), .B2(n7139), .A(n7113), .ZN(n9432) );
  INV_X1 U8729 ( .A(n7128), .ZN(n9428) );
  OAI211_X1 U8730 ( .C1(n7114), .C2(n9428), .A(n9366), .B(n7140), .ZN(n9427)
         );
  INV_X1 U8731 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7116) );
  OAI22_X1 U8732 ( .A1(n9276), .A2(n7116), .B1(n7115), .B2(n9274), .ZN(n7117)
         );
  AOI21_X1 U8733 ( .B1(n7128), .B2(n9280), .A(n7117), .ZN(n7118) );
  OAI21_X1 U8734 ( .B1(n9427), .B2(n7450), .A(n7118), .ZN(n7119) );
  AOI21_X1 U8735 ( .B1(n9430), .B2(n7659), .A(n7119), .ZN(n7120) );
  OAI21_X1 U8736 ( .B1(n9432), .B2(n9253), .A(n7120), .ZN(P1_U3281) );
  INV_X1 U8737 ( .A(n7456), .ZN(n9841) );
  OAI211_X1 U8738 ( .C1(n7123), .C2(n7122), .A(n7121), .B(n8535), .ZN(n7126)
         );
  NOR2_X1 U8739 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5996), .ZN(n8601) );
  OAI22_X1 U8740 ( .A1(n7464), .A2(n8516), .B1(n8517), .B2(n7367), .ZN(n7124)
         );
  AOI211_X1 U8741 ( .C1(n8543), .C2(n7375), .A(n8601), .B(n7124), .ZN(n7125)
         );
  OAI211_X1 U8742 ( .C1(n9841), .C2(n8546), .A(n7126), .B(n7125), .ZN(P2_U3238) );
  INV_X1 U8743 ( .A(n7177), .ZN(n7127) );
  OR2_X1 U8744 ( .A1(n7128), .A2(n7127), .ZN(n7129) );
  OR2_X1 U8745 ( .A1(n7249), .A2(n9016), .ZN(n7247) );
  NAND2_X1 U8746 ( .A1(n7249), .A2(n9016), .ZN(n7245) );
  AND2_X1 U8747 ( .A1(n7247), .A2(n7245), .ZN(n8349) );
  XNOR2_X1 U8748 ( .A(n7246), .B(n8349), .ZN(n7264) );
  AND2_X1 U8749 ( .A1(n7131), .A2(n7132), .ZN(n8334) );
  NAND2_X1 U8750 ( .A1(n8330), .A2(n8331), .ZN(n7133) );
  AND2_X1 U8751 ( .A1(n7133), .A2(n7132), .ZN(n8326) );
  INV_X1 U8752 ( .A(n8349), .ZN(n8248) );
  XNOR2_X1 U8753 ( .A(n7248), .B(n8248), .ZN(n7137) );
  OAI22_X1 U8754 ( .A1(n7177), .A2(n9267), .B1(n7516), .B2(n9269), .ZN(n7135)
         );
  INV_X1 U8755 ( .A(n7135), .ZN(n7136) );
  OAI21_X1 U8756 ( .B1(n7137), .B2(n9265), .A(n7136), .ZN(n7138) );
  AOI21_X1 U8757 ( .B1(n7264), .B2(n7139), .A(n7138), .ZN(n7266) );
  NAND2_X1 U8758 ( .A1(n7140), .A2(n7249), .ZN(n7141) );
  NAND2_X1 U8759 ( .A1(n7255), .A2(n7141), .ZN(n7262) );
  OAI22_X1 U8760 ( .A1(n9276), .A2(n7142), .B1(n7174), .B2(n9274), .ZN(n7143)
         );
  AOI21_X1 U8761 ( .B1(n7249), .B2(n9280), .A(n7143), .ZN(n7144) );
  OAI21_X1 U8762 ( .B1(n7262), .B2(n9163), .A(n7144), .ZN(n7145) );
  AOI21_X1 U8763 ( .B1(n7264), .B2(n7659), .A(n7145), .ZN(n7146) );
  OAI21_X1 U8764 ( .B1(n7266), .B2(n9253), .A(n7146), .ZN(P1_U3280) );
  INV_X1 U8765 ( .A(n7147), .ZN(n7149) );
  OAI222_X1 U8766 ( .A1(n8475), .A2(n7148), .B1(n8478), .B2(n7149), .C1(n7970), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI222_X1 U8767 ( .A1(P1_U3084), .A2(n8267), .B1(n7873), .B2(n7149), .C1(
        n10003), .C2(n7863), .ZN(P1_U3332) );
  INV_X1 U8768 ( .A(n7227), .ZN(n7169) );
  XNOR2_X1 U8769 ( .A(n7227), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7155) );
  AOI21_X1 U8770 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7151), .A(n7150), .ZN(
        n8599) );
  INV_X1 U8771 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7152) );
  MUX2_X1 U8772 ( .A(n7152), .B(P2_REG2_REG_11__SCAN_IN), .S(n8596), .Z(n7153)
         );
  INV_X1 U8773 ( .A(n7153), .ZN(n8598) );
  NAND2_X1 U8774 ( .A1(n8599), .A2(n8598), .ZN(n8597) );
  OAI21_X1 U8775 ( .B1(n8596), .B2(P2_REG2_REG_11__SCAN_IN), .A(n8597), .ZN(
        n7154) );
  NOR2_X1 U8776 ( .A1(n7154), .A2(n7155), .ZN(n7226) );
  AOI211_X1 U8777 ( .C1(n7155), .C2(n7154), .A(n7226), .B(n9414), .ZN(n7156)
         );
  INV_X1 U8778 ( .A(n7156), .ZN(n7168) );
  INV_X1 U8779 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7157) );
  MUX2_X1 U8780 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7157), .S(n8596), .Z(n8603)
         );
  OAI21_X1 U8781 ( .B1(n9867), .B2(n7159), .A(n7158), .ZN(n8604) );
  NAND2_X1 U8782 ( .A1(n8603), .A2(n8604), .ZN(n8602) );
  INV_X1 U8783 ( .A(n8602), .ZN(n7160) );
  AOI21_X1 U8784 ( .B1(n8596), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7160), .ZN(
        n7162) );
  INV_X1 U8785 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9871) );
  MUX2_X1 U8786 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9871), .S(n7227), .Z(n7161)
         );
  NAND2_X1 U8787 ( .A1(n7161), .A2(n7162), .ZN(n7220) );
  OAI21_X1 U8788 ( .B1(n7162), .B2(n7161), .A(n7220), .ZN(n7166) );
  NOR2_X1 U8789 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7188), .ZN(n7165) );
  INV_X1 U8790 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7163) );
  NOR2_X1 U8791 ( .A1(n9402), .A2(n7163), .ZN(n7164) );
  AOI211_X1 U8792 ( .C1(n9708), .C2(n7166), .A(n7165), .B(n7164), .ZN(n7167)
         );
  OAI211_X1 U8793 ( .C1(n9711), .C2(n7169), .A(n7168), .B(n7167), .ZN(P2_U3257) );
  AOI21_X1 U8794 ( .B1(n7171), .B2(n7170), .A(n9446), .ZN(n7173) );
  NAND2_X1 U8795 ( .A1(n7173), .A2(n7172), .ZN(n7181) );
  INV_X1 U8796 ( .A(n7174), .ZN(n7179) );
  INV_X1 U8797 ( .A(n7516), .ZN(n7437) );
  AOI21_X1 U8798 ( .B1(n9438), .B2(n7437), .A(n7175), .ZN(n7176) );
  OAI21_X1 U8799 ( .B1(n7177), .B2(n9435), .A(n7176), .ZN(n7178) );
  AOI21_X1 U8800 ( .B1(n9003), .B2(n7179), .A(n7178), .ZN(n7180) );
  OAI211_X1 U8801 ( .C1(n4597), .C2(n9010), .A(n7181), .B(n7180), .ZN(P1_U3234) );
  INV_X1 U8802 ( .A(n7182), .ZN(n7183) );
  NOR2_X1 U8803 ( .A1(n7184), .A2(n7183), .ZN(n7185) );
  XNOR2_X1 U8804 ( .A(n7186), .B(n7185), .ZN(n7193) );
  OR2_X1 U8805 ( .A1(n7455), .A2(n9763), .ZN(n7187) );
  OAI21_X1 U8806 ( .B1(n7499), .B2(n9761), .A(n7187), .ZN(n9727) );
  INV_X1 U8807 ( .A(n9727), .ZN(n7189) );
  OAI22_X1 U8808 ( .A1(n8541), .A2(n7189), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7188), .ZN(n7191) );
  INV_X1 U8809 ( .A(n9732), .ZN(n9851) );
  NOR2_X1 U8810 ( .A1(n9851), .A2(n8546), .ZN(n7190) );
  AOI211_X1 U8811 ( .C1(n8543), .C2(n9730), .A(n7191), .B(n7190), .ZN(n7192)
         );
  OAI21_X1 U8812 ( .B1(n7193), .B2(n8522), .A(n7192), .ZN(P2_U3226) );
  INV_X1 U8813 ( .A(n7194), .ZN(n7211) );
  NAND2_X1 U8814 ( .A1(n7196), .A2(n7195), .ZN(n7197) );
  NOR2_X1 U8815 ( .A1(n9780), .A2(n7197), .ZN(n7198) );
  NAND2_X1 U8816 ( .A1(n7199), .A2(n7198), .ZN(n7207) );
  OR2_X1 U8817 ( .A1(n7200), .A2(n8707), .ZN(n7335) );
  AND2_X1 U8818 ( .A1(n9769), .A2(n7335), .ZN(n7201) );
  INV_X1 U8819 ( .A(n9773), .ZN(n7202) );
  INV_X1 U8820 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7203) );
  OAI22_X1 U8821 ( .A1(n9773), .A2(n7204), .B1(n7203), .B2(n8817), .ZN(n7205)
         );
  AOI21_X1 U8822 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9749), .A(n7205), .ZN(
        n7210) );
  OR2_X1 U8823 ( .A1(n7207), .A2(n7966), .ZN(n8815) );
  OR2_X1 U8824 ( .A1(n8815), .A2(n9842), .ZN(n9757) );
  INV_X1 U8825 ( .A(n9757), .ZN(n8806) );
  OAI21_X1 U8826 ( .B1(n9731), .B2(n8806), .A(n7208), .ZN(n7209) );
  OAI211_X1 U8827 ( .C1(n7211), .C2(n8808), .A(n7210), .B(n7209), .ZN(P2_U3296) );
  INV_X1 U8828 ( .A(n7235), .ZN(n7214) );
  OR2_X1 U8829 ( .A1(n7212), .A2(P1_U3084), .ZN(n8444) );
  NAND2_X1 U8830 ( .A1(n7870), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7213) );
  OAI211_X1 U8831 ( .C1(n7214), .C2(n7873), .A(n8444), .B(n7213), .ZN(P1_U3330) );
  INV_X1 U8832 ( .A(n7215), .ZN(n8450) );
  OAI222_X1 U8833 ( .A1(n7863), .A2(n7216), .B1(n7873), .B2(n8450), .C1(n8441), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  INV_X1 U8834 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7218) );
  OAI22_X1 U8835 ( .A1(n9402), .A2(n7218), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7217), .ZN(n7225) );
  INV_X1 U8836 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U8837 ( .A1(n7399), .A2(n9954), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7394), .ZN(n7222) );
  OR2_X1 U8838 ( .A1(n7227), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7219) );
  AND2_X1 U8839 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  NOR2_X1 U8840 ( .A1(n7221), .A2(n7222), .ZN(n7393) );
  AOI21_X1 U8841 ( .B1(n7222), .B2(n7221), .A(n7393), .ZN(n7223) );
  NOR2_X1 U8842 ( .A1(n9713), .A2(n7223), .ZN(n7224) );
  AOI211_X1 U8843 ( .C1(n9420), .C2(n7399), .A(n7225), .B(n7224), .ZN(n7233)
         );
  NOR2_X1 U8844 ( .A1(n7399), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7228) );
  AOI21_X1 U8845 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7399), .A(n7228), .ZN(
        n7229) );
  OAI21_X1 U8846 ( .B1(n7230), .B2(n7229), .A(n7398), .ZN(n7231) );
  NAND2_X1 U8847 ( .A1(n9710), .A2(n7231), .ZN(n7232) );
  NAND2_X1 U8848 ( .A1(n7233), .A2(n7232), .ZN(P2_U3258) );
  NAND2_X1 U8849 ( .A1(n7235), .A2(n7234), .ZN(n7236) );
  OAI211_X1 U8850 ( .C1(n9940), .C2(n7837), .A(n7236), .B(n8161), .ZN(P2_U3335) );
  OAI22_X1 U8851 ( .A1(n8815), .A2(n7237), .B1(n9401), .B2(n8817), .ZN(n7239)
         );
  NOR2_X1 U8852 ( .A1(n7202), .A2(n6597), .ZN(n7238) );
  AOI211_X1 U8853 ( .C1(n7202), .C2(n7240), .A(n7239), .B(n7238), .ZN(n7244)
         );
  INV_X1 U8854 ( .A(n8808), .ZN(n9746) );
  AOI22_X1 U8855 ( .A1(n9746), .A2(n7242), .B1(n9731), .B2(n7241), .ZN(n7243)
         );
  NAND2_X1 U8856 ( .A1(n7244), .A2(n7243), .ZN(P2_U3295) );
  OR2_X1 U8857 ( .A1(n9444), .A2(n7516), .ZN(n8343) );
  NAND2_X1 U8858 ( .A1(n9444), .A2(n7516), .ZN(n8342) );
  AOI21_X1 U8859 ( .B1(n8251), .B2(n7439), .A(n4467), .ZN(n9493) );
  INV_X1 U8860 ( .A(n9016), .ZN(n9434) );
  NAND2_X1 U8861 ( .A1(n7249), .A2(n9434), .ZN(n8341) );
  OR2_X1 U8862 ( .A1(n7249), .A2(n9434), .ZN(n7441) );
  NAND2_X1 U8863 ( .A1(n7442), .A2(n7441), .ZN(n7251) );
  INV_X1 U8864 ( .A(n8251), .ZN(n7250) );
  XNOR2_X1 U8865 ( .A(n7251), .B(n7250), .ZN(n7252) );
  NAND2_X1 U8866 ( .A1(n7252), .A2(n9223), .ZN(n9491) );
  NAND2_X1 U8867 ( .A1(n9437), .A2(n9218), .ZN(n7254) );
  NAND2_X1 U8868 ( .A1(n9016), .A2(n9220), .ZN(n7253) );
  AND2_X1 U8869 ( .A1(n7254), .A2(n7253), .ZN(n9490) );
  AOI21_X1 U8870 ( .B1(n9491), .B2(n9490), .A(n9253), .ZN(n7260) );
  AOI21_X1 U8871 ( .B1(n7255), .B2(n9444), .A(n9688), .ZN(n7256) );
  NAND2_X1 U8872 ( .A1(n7256), .A2(n7488), .ZN(n9488) );
  INV_X1 U8873 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9045) );
  OAI22_X1 U8874 ( .A1(n9276), .A2(n9045), .B1(n9451), .B2(n9274), .ZN(n7257)
         );
  AOI21_X1 U8875 ( .B1(n9444), .B2(n9280), .A(n7257), .ZN(n7258) );
  OAI21_X1 U8876 ( .B1(n9488), .B2(n7450), .A(n7258), .ZN(n7259) );
  AOI211_X1 U8877 ( .C1(n9493), .C2(n9283), .A(n7260), .B(n7259), .ZN(n7261)
         );
  INV_X1 U8878 ( .A(n7261), .ZN(P1_U3279) );
  NAND2_X1 U8879 ( .A1(n8441), .A2(n9275), .ZN(n8424) );
  OR2_X1 U8880 ( .A1(n8424), .A2(n8436), .ZN(n9377) );
  INV_X1 U8881 ( .A(n9377), .ZN(n9693) );
  OAI22_X1 U8882 ( .A1(n7262), .A2(n9688), .B1(n4597), .B2(n9686), .ZN(n7263)
         );
  AOI21_X1 U8883 ( .B1(n7264), .B2(n9693), .A(n7263), .ZN(n7265) );
  AND2_X1 U8884 ( .A1(n7266), .A2(n7265), .ZN(n7268) );
  MUX2_X1 U8885 ( .A(n5311), .B(n7268), .S(n9707), .Z(n7267) );
  INV_X1 U8886 ( .A(n7267), .ZN(P1_U3534) );
  INV_X1 U8887 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10079) );
  MUX2_X1 U8888 ( .A(n10079), .B(n7268), .S(n9696), .Z(n7269) );
  INV_X1 U8889 ( .A(n7269), .ZN(P1_U3487) );
  XNOR2_X1 U8890 ( .A(n7271), .B(n7270), .ZN(n7276) );
  INV_X1 U8891 ( .A(n7469), .ZN(n7272) );
  OAI22_X1 U8892 ( .A1(n8515), .A2(n7272), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7217), .ZN(n7274) );
  OAI22_X1 U8893 ( .A1(n7464), .A2(n8517), .B1(n8516), .B2(n7642), .ZN(n7273)
         );
  AOI211_X1 U8894 ( .C1(n8037), .C2(n8520), .A(n7274), .B(n7273), .ZN(n7275)
         );
  OAI21_X1 U8895 ( .B1(n7276), .B2(n8522), .A(n7275), .ZN(P2_U3236) );
  OAI21_X1 U8896 ( .B1(n7278), .B2(n7282), .A(n7277), .ZN(n9790) );
  OR2_X1 U8897 ( .A1(n9786), .A2(n7279), .ZN(n7280) );
  NAND2_X1 U8898 ( .A1(n7281), .A2(n7280), .ZN(n9787) );
  OAI22_X1 U8899 ( .A1(n9775), .A2(n9786), .B1(n9757), .B2(n9787), .ZN(n7293)
         );
  INV_X1 U8900 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7291) );
  NAND2_X1 U8901 ( .A1(n7283), .A2(n7282), .ZN(n7284) );
  INV_X1 U8902 ( .A(n9766), .ZN(n9725) );
  AOI21_X1 U8903 ( .B1(n7285), .B2(n7284), .A(n9725), .ZN(n7288) );
  OAI22_X1 U8904 ( .A1(n7286), .A2(n9763), .B1(n7348), .B2(n9761), .ZN(n7287)
         );
  OR2_X1 U8905 ( .A1(n7288), .A2(n7287), .ZN(n9788) );
  INV_X1 U8906 ( .A(n8817), .ZN(n9771) );
  AND2_X1 U8907 ( .A1(n9771), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7289) );
  AOI21_X1 U8908 ( .B1(n9788), .B2(n7202), .A(n7289), .ZN(n7290) );
  OAI21_X1 U8909 ( .B1(n7291), .B2(n7202), .A(n7290), .ZN(n7292) );
  AOI211_X1 U8910 ( .C1(n9746), .C2(n9790), .A(n7293), .B(n7292), .ZN(n7294)
         );
  INV_X1 U8911 ( .A(n7294), .ZN(P2_U3294) );
  NAND2_X1 U8912 ( .A1(n7348), .A2(n7336), .ZN(n7295) );
  NAND2_X1 U8913 ( .A1(n7296), .A2(n7295), .ZN(n7353) );
  NAND2_X1 U8914 ( .A1(n7297), .A2(n7358), .ZN(n7973) );
  INV_X1 U8915 ( .A(n7297), .ZN(n8568) );
  NAND2_X1 U8916 ( .A1(n8568), .A2(n9792), .ZN(n7323) );
  NAND2_X1 U8917 ( .A1(n7973), .A2(n7323), .ZN(n8125) );
  NAND2_X1 U8918 ( .A1(n7297), .A2(n9792), .ZN(n7298) );
  NAND2_X1 U8919 ( .A1(n6816), .A2(n7299), .ZN(n7974) );
  NAND2_X1 U8920 ( .A1(n8566), .A2(n9799), .ZN(n7992) );
  NAND2_X1 U8921 ( .A1(n7974), .A2(n7992), .ZN(n8126) );
  XNOR2_X1 U8922 ( .A(n7312), .B(n8126), .ZN(n9801) );
  INV_X1 U8923 ( .A(n9801), .ZN(n7311) );
  OAI21_X1 U8924 ( .B1(n7355), .B2(n9799), .A(n6266), .ZN(n7300) );
  OR2_X1 U8925 ( .A1(n7300), .A2(n8814), .ZN(n9797) );
  INV_X1 U8926 ( .A(n9797), .ZN(n7309) );
  INV_X1 U8927 ( .A(n8815), .ZN(n9745) );
  AOI22_X1 U8928 ( .A1(n9773), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n7301), .B2(
        n9771), .ZN(n7302) );
  OAI21_X1 U8929 ( .B1(n9775), .B2(n9799), .A(n7302), .ZN(n7308) );
  NAND2_X1 U8930 ( .A1(n7324), .A2(n7323), .ZN(n7304) );
  XNOR2_X1 U8931 ( .A(n7304), .B(n8126), .ZN(n7306) );
  AOI21_X1 U8932 ( .B1(n7306), .B2(n9766), .A(n7305), .ZN(n9798) );
  INV_X1 U8933 ( .A(n7202), .ZN(n8740) );
  NOR2_X1 U8934 ( .A1(n9798), .A2(n8740), .ZN(n7307) );
  AOI211_X1 U8935 ( .C1(n7309), .C2(n9745), .A(n7308), .B(n7307), .ZN(n7310)
         );
  OAI21_X1 U8936 ( .B1(n7311), .B2(n8808), .A(n7310), .ZN(P2_U3291) );
  INV_X1 U8937 ( .A(n8821), .ZN(n7313) );
  NAND2_X1 U8938 ( .A1(n9806), .A2(n8565), .ZN(n7998) );
  INV_X1 U8939 ( .A(n9806), .ZN(n7314) );
  NAND2_X1 U8940 ( .A1(n7314), .A2(n8565), .ZN(n7315) );
  OR2_X1 U8941 ( .A1(n9810), .A2(n9764), .ZN(n8006) );
  NAND2_X1 U8942 ( .A1(n9810), .A2(n9764), .ZN(n8005) );
  INV_X1 U8943 ( .A(n9751), .ZN(n7318) );
  OR2_X1 U8944 ( .A1(n9770), .A2(n7384), .ZN(n8010) );
  NAND2_X1 U8945 ( .A1(n9770), .A2(n7384), .ZN(n8011) );
  INV_X1 U8946 ( .A(n7384), .ZN(n8563) );
  NAND2_X1 U8947 ( .A1(n9770), .A2(n8563), .ZN(n7319) );
  OR2_X1 U8948 ( .A1(n9823), .A2(n9762), .ZN(n8016) );
  NAND2_X1 U8949 ( .A1(n9823), .A2(n9762), .ZN(n8023) );
  INV_X1 U8950 ( .A(n7414), .ZN(n8132) );
  XNOR2_X1 U8951 ( .A(n7454), .B(n8132), .ZN(n9828) );
  AOI211_X1 U8952 ( .C1(n9823), .C2(n4631), .A(n9842), .B(n7429), .ZN(n9822)
         );
  AOI22_X1 U8953 ( .A1(n9773), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7320), .B2(
        n9771), .ZN(n7321) );
  OAI21_X1 U8954 ( .B1(n9775), .B2(n7322), .A(n7321), .ZN(n7331) );
  AND2_X1 U8955 ( .A1(n7992), .A2(n7323), .ZN(n7994) );
  NAND2_X1 U8956 ( .A1(n7324), .A2(n7994), .ZN(n7325) );
  NAND2_X1 U8957 ( .A1(n7325), .A2(n7974), .ZN(n8810) );
  INV_X1 U8958 ( .A(n8005), .ZN(n7326) );
  NAND2_X1 U8959 ( .A1(n7327), .A2(n7414), .ZN(n7365) );
  OAI21_X1 U8960 ( .B1(n7414), .B2(n7327), .A(n7365), .ZN(n7329) );
  AOI21_X1 U8961 ( .B1(n7329), .B2(n9766), .A(n7328), .ZN(n9826) );
  NOR2_X1 U8962 ( .A1(n9826), .A2(n8740), .ZN(n7330) );
  AOI211_X1 U8963 ( .C1(n9822), .C2(n9745), .A(n7331), .B(n7330), .ZN(n7332)
         );
  OAI21_X1 U8964 ( .B1(n8808), .B2(n9828), .A(n7332), .ZN(P2_U3287) );
  INV_X1 U8965 ( .A(n7333), .ZN(n7341) );
  OAI22_X1 U8966 ( .A1(n8815), .A2(n7334), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8817), .ZN(n7339) );
  OR2_X1 U8967 ( .A1(n9749), .A2(n7335), .ZN(n9758) );
  OAI22_X1 U8968 ( .A1(n7337), .A2(n9758), .B1(n7336), .B2(n9775), .ZN(n7338)
         );
  AOI211_X1 U8969 ( .C1(P2_REG2_REG_3__SCAN_IN), .C2(n9773), .A(n7339), .B(
        n7338), .ZN(n7340) );
  OAI21_X1 U8970 ( .B1(n9749), .B2(n7341), .A(n7340), .ZN(P2_U3293) );
  INV_X1 U8971 ( .A(n7342), .ZN(n7865) );
  OAI222_X1 U8972 ( .A1(P2_U3152), .A2(n7344), .B1(n8478), .B2(n7865), .C1(
        n7343), .C2(n7837), .ZN(P2_U3334) );
  INV_X1 U8973 ( .A(n8125), .ZN(n7345) );
  XNOR2_X1 U8974 ( .A(n7346), .B(n7345), .ZN(n7347) );
  NAND2_X1 U8975 ( .A1(n7347), .A2(n9766), .ZN(n7351) );
  OAI22_X1 U8976 ( .A1(n7348), .A2(n9763), .B1(n6816), .B2(n9761), .ZN(n7349)
         );
  INV_X1 U8977 ( .A(n7349), .ZN(n7350) );
  NAND2_X1 U8978 ( .A1(n7351), .A2(n7350), .ZN(n9793) );
  INV_X1 U8979 ( .A(n9793), .ZN(n7364) );
  OAI21_X1 U8980 ( .B1(n7353), .B2(n8125), .A(n7352), .ZN(n9795) );
  INV_X1 U8981 ( .A(n7354), .ZN(n7357) );
  INV_X1 U8982 ( .A(n7355), .ZN(n7356) );
  OAI211_X1 U8983 ( .C1(n9792), .C2(n7357), .A(n7356), .B(n6266), .ZN(n9791)
         );
  NAND2_X1 U8984 ( .A1(n9731), .A2(n7358), .ZN(n7361) );
  AOI22_X1 U8985 ( .A1(n9773), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n7359), .B2(
        n9771), .ZN(n7360) );
  OAI211_X1 U8986 ( .C1(n8815), .C2(n9791), .A(n7361), .B(n7360), .ZN(n7362)
         );
  AOI21_X1 U8987 ( .B1(n9795), .B2(n9746), .A(n7362), .ZN(n7363) );
  OAI21_X1 U8988 ( .B1(n7364), .B2(n8740), .A(n7363), .ZN(P2_U3292) );
  NAND2_X1 U8989 ( .A1(n7365), .A2(n8023), .ZN(n7420) );
  NAND2_X1 U8990 ( .A1(n7420), .A2(n8015), .ZN(n7423) );
  NAND2_X1 U8991 ( .A1(n7423), .A2(n8022), .ZN(n9719) );
  OR2_X1 U8992 ( .A1(n7456), .A2(n7455), .ZN(n9720) );
  NAND2_X1 U8993 ( .A1(n7456), .A2(n7455), .ZN(n8028) );
  NAND2_X1 U8994 ( .A1(n9720), .A2(n8028), .ZN(n8131) );
  XNOR2_X1 U8995 ( .A(n9719), .B(n8131), .ZN(n7366) );
  OAI222_X1 U8996 ( .A1(n9763), .A2(n7367), .B1(n9761), .B2(n7464), .C1(n7366), 
        .C2(n9725), .ZN(n9844) );
  INV_X1 U8997 ( .A(n9844), .ZN(n7380) );
  INV_X1 U8998 ( .A(n7367), .ZN(n8561) );
  AND2_X1 U8999 ( .A1(n7434), .A2(n8561), .ZN(n7368) );
  OR2_X1 U9000 ( .A1(n7414), .A2(n7368), .ZN(n7457) );
  OR2_X1 U9001 ( .A1(n7454), .A2(n7457), .ZN(n7371) );
  OR2_X1 U9002 ( .A1(n9823), .A2(n8562), .ZN(n7415) );
  AND2_X1 U9003 ( .A1(n8130), .A2(n7415), .ZN(n7416) );
  OR2_X1 U9004 ( .A1(n7368), .A2(n7416), .ZN(n7370) );
  AND2_X1 U9005 ( .A1(n7371), .A2(n7370), .ZN(n7369) );
  OR2_X1 U9006 ( .A1(n7369), .A2(n8131), .ZN(n7373) );
  NAND2_X1 U9007 ( .A1(n7371), .A2(n7458), .ZN(n7372) );
  AND2_X1 U9008 ( .A1(n7373), .A2(n7372), .ZN(n9846) );
  NAND2_X1 U9009 ( .A1(n7429), .A2(n9834), .ZN(n7431) );
  INV_X1 U9010 ( .A(n7431), .ZN(n7374) );
  OAI21_X1 U9011 ( .B1(n7374), .B2(n9841), .A(n9741), .ZN(n9843) );
  AOI22_X1 U9012 ( .A1(n9749), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7375), .B2(
        n9771), .ZN(n7377) );
  NAND2_X1 U9013 ( .A1(n9731), .A2(n7456), .ZN(n7376) );
  OAI211_X1 U9014 ( .C1(n9843), .C2(n9757), .A(n7377), .B(n7376), .ZN(n7378)
         );
  AOI21_X1 U9015 ( .B1(n9846), .B2(n9746), .A(n7378), .ZN(n7379) );
  OAI21_X1 U9016 ( .B1(n7380), .B2(n8740), .A(n7379), .ZN(P2_U3285) );
  XOR2_X1 U9017 ( .A(n8128), .B(n7381), .Z(n7382) );
  OAI222_X1 U9018 ( .A1(n9761), .A2(n7384), .B1(n9763), .B2(n7383), .C1(n7382), 
        .C2(n9725), .ZN(n9813) );
  INV_X1 U9019 ( .A(n9813), .ZN(n7392) );
  OAI21_X1 U9020 ( .B1(n4946), .B2(n7316), .A(n7385), .ZN(n9815) );
  NAND2_X1 U9021 ( .A1(n8813), .A2(n9810), .ZN(n7386) );
  NAND2_X1 U9022 ( .A1(n9754), .A2(n7386), .ZN(n9812) );
  AOI22_X1 U9023 ( .A1(n9773), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7387), .B2(
        n9771), .ZN(n7389) );
  NAND2_X1 U9024 ( .A1(n9731), .A2(n9810), .ZN(n7388) );
  OAI211_X1 U9025 ( .C1(n9812), .C2(n9757), .A(n7389), .B(n7388), .ZN(n7390)
         );
  AOI21_X1 U9026 ( .B1(n9815), .B2(n9746), .A(n7390), .ZN(n7391) );
  OAI21_X1 U9027 ( .B1(n7392), .B2(n8740), .A(n7391), .ZN(P2_U3289) );
  AOI21_X1 U9028 ( .B1(n7394), .B2(n9954), .A(n7393), .ZN(n7396) );
  INV_X1 U9029 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U9030 ( .A1(n7596), .A2(n10091), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7599), .ZN(n7395) );
  NOR2_X1 U9031 ( .A1(n7396), .A2(n7395), .ZN(n7598) );
  AOI21_X1 U9032 ( .B1(n7396), .B2(n7395), .A(n7598), .ZN(n7407) );
  INV_X1 U9033 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7397) );
  AOI22_X1 U9034 ( .A1(n7596), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7397), .B2(
        n7599), .ZN(n7401) );
  OAI21_X1 U9035 ( .B1(n7401), .B2(n7400), .A(n7595), .ZN(n7402) );
  NAND2_X1 U9036 ( .A1(n7402), .A2(n9710), .ZN(n7406) );
  INV_X1 U9037 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U9038 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7477) );
  OAI21_X1 U9039 ( .B1(n9402), .B2(n7403), .A(n7477), .ZN(n7404) );
  AOI21_X1 U9040 ( .B1(n9420), .B2(n7596), .A(n7404), .ZN(n7405) );
  OAI211_X1 U9041 ( .C1(n7407), .C2(n9713), .A(n7406), .B(n7405), .ZN(P2_U3259) );
  INV_X1 U9042 ( .A(n7408), .ZN(n7412) );
  OAI222_X1 U9043 ( .A1(n7863), .A2(n7410), .B1(n7873), .B2(n7412), .C1(n7409), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9044 ( .A1(n8475), .A2(n7413), .B1(n8478), .B2(n7412), .C1(
        P2_U3152), .C2(n7411), .ZN(P2_U3333) );
  OR2_X1 U9045 ( .A1(n7454), .A2(n7414), .ZN(n7417) );
  AND2_X1 U9046 ( .A1(n7417), .A2(n7415), .ZN(n7419) );
  NAND2_X1 U9047 ( .A1(n7417), .A2(n7416), .ZN(n7418) );
  OAI21_X1 U9048 ( .B1(n7419), .B2(n8130), .A(n7418), .ZN(n9833) );
  INV_X1 U9049 ( .A(n8022), .ZN(n7422) );
  INV_X1 U9050 ( .A(n8130), .ZN(n7421) );
  OAI22_X1 U9051 ( .A1(n7423), .A2(n7422), .B1(n7421), .B2(n7420), .ZN(n7425)
         );
  OAI22_X1 U9052 ( .A1(n7455), .A2(n9761), .B1(n9762), .B2(n9763), .ZN(n7424)
         );
  AOI21_X1 U9053 ( .B1(n7425), .B2(n9766), .A(n7424), .ZN(n7426) );
  OAI21_X1 U9054 ( .B1(n9833), .B2(n9769), .A(n7426), .ZN(n9836) );
  NAND2_X1 U9055 ( .A1(n9836), .A2(n7202), .ZN(n7436) );
  INV_X1 U9056 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10095) );
  INV_X1 U9057 ( .A(n7427), .ZN(n7428) );
  OAI22_X1 U9058 ( .A1(n7202), .A2(n10095), .B1(n7428), .B2(n8817), .ZN(n7433)
         );
  OR2_X1 U9059 ( .A1(n7429), .A2(n9834), .ZN(n7430) );
  NAND2_X1 U9060 ( .A1(n7431), .A2(n7430), .ZN(n9835) );
  NOR2_X1 U9061 ( .A1(n9835), .A2(n9757), .ZN(n7432) );
  AOI211_X1 U9062 ( .C1(n9731), .C2(n7434), .A(n7433), .B(n7432), .ZN(n7435)
         );
  OAI211_X1 U9063 ( .C1(n9833), .C2(n9758), .A(n7436), .B(n7435), .ZN(P2_U3286) );
  INV_X1 U9064 ( .A(n9015), .ZN(n7648) );
  OR2_X1 U9065 ( .A1(n7628), .A2(n7648), .ZN(n8354) );
  NAND2_X1 U9066 ( .A1(n7628), .A2(n7648), .ZN(n8352) );
  NAND2_X1 U9067 ( .A1(n8354), .A2(n8352), .ZN(n8253) );
  NAND2_X1 U9068 ( .A1(n9444), .A2(n7437), .ZN(n7438) );
  OAI21_X1 U9069 ( .B1(n9437), .B2(n7521), .A(n7484), .ZN(n7440) );
  INV_X1 U9070 ( .A(n7521), .ZN(n9371) );
  INV_X1 U9071 ( .A(n9437), .ZN(n7529) );
  XOR2_X1 U9072 ( .A(n8253), .B(n7629), .Z(n9487) );
  INV_X1 U9073 ( .A(n9487), .ZN(n7453) );
  AND2_X1 U9074 ( .A1(n8343), .A2(n7441), .ZN(n8206) );
  NAND2_X1 U9075 ( .A1(n7443), .A2(n8342), .ZN(n7482) );
  OR2_X1 U9076 ( .A1(n7521), .A2(n7529), .ZN(n8351) );
  NAND2_X1 U9077 ( .A1(n7521), .A2(n7529), .ZN(n8210) );
  INV_X1 U9078 ( .A(n8253), .ZN(n7444) );
  OAI211_X1 U9079 ( .C1(n4469), .C2(n7444), .A(n7624), .B(n9223), .ZN(n7446)
         );
  AOI22_X1 U9080 ( .A1(n9220), .A2(n9437), .B1(n9014), .B2(n9218), .ZN(n7445)
         );
  NAND2_X1 U9081 ( .A1(n7446), .A2(n7445), .ZN(n9486) );
  OAI211_X1 U9082 ( .C1(n9484), .C2(n7489), .A(n4457), .B(n9366), .ZN(n9483)
         );
  OAI22_X1 U9083 ( .A1(n9276), .A2(n7447), .B1(n7532), .B2(n9274), .ZN(n7448)
         );
  AOI21_X1 U9084 ( .B1(n7628), .B2(n9280), .A(n7448), .ZN(n7449) );
  OAI21_X1 U9085 ( .B1(n9483), .B2(n7450), .A(n7449), .ZN(n7451) );
  AOI21_X1 U9086 ( .B1(n9486), .B2(n9276), .A(n7451), .ZN(n7452) );
  OAI21_X1 U9087 ( .B1(n7453), .B2(n9262), .A(n7452), .ZN(P1_U3277) );
  INV_X1 U9088 ( .A(n7455), .ZN(n8560) );
  AND2_X1 U9089 ( .A1(n7456), .A2(n8560), .ZN(n7459) );
  OR2_X1 U9090 ( .A1(n7457), .A2(n7459), .ZN(n9733) );
  NAND2_X1 U9091 ( .A1(n9732), .A2(n7464), .ZN(n8033) );
  INV_X1 U9092 ( .A(n7464), .ZN(n8559) );
  OR2_X1 U9093 ( .A1(n9732), .A2(n8559), .ZN(n7460) );
  XNOR2_X1 U9094 ( .A(n8037), .B(n7499), .ZN(n8041) );
  OAI21_X1 U9095 ( .B1(n7462), .B2(n8041), .A(n7503), .ZN(n9465) );
  INV_X1 U9096 ( .A(n8028), .ZN(n9726) );
  OAI21_X1 U9097 ( .B1(n9719), .B2(n9726), .A(n9720), .ZN(n7463) );
  NAND2_X1 U9098 ( .A1(n7463), .A2(n9722), .ZN(n9728) );
  OAI21_X1 U9099 ( .B1(n4956), .B2(n4853), .A(n7497), .ZN(n7466) );
  OAI22_X1 U9100 ( .A1(n7464), .A2(n9763), .B1(n7642), .B2(n9761), .ZN(n7465)
         );
  AOI21_X1 U9101 ( .B1(n7466), .B2(n9766), .A(n7465), .ZN(n7467) );
  OAI21_X1 U9102 ( .B1(n9465), .B2(n9769), .A(n7467), .ZN(n9468) );
  NAND2_X1 U9103 ( .A1(n9468), .A2(n7202), .ZN(n7474) );
  AND2_X1 U9104 ( .A1(n9742), .A2(n8037), .ZN(n7468) );
  OR2_X1 U9105 ( .A1(n7468), .A2(n7507), .ZN(n9467) );
  INV_X1 U9106 ( .A(n9467), .ZN(n7472) );
  INV_X1 U9107 ( .A(n8037), .ZN(n9466) );
  AOI22_X1 U9108 ( .A1(n9749), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7469), .B2(
        n9771), .ZN(n7470) );
  OAI21_X1 U9109 ( .B1(n9466), .B2(n9775), .A(n7470), .ZN(n7471) );
  AOI21_X1 U9110 ( .B1(n7472), .B2(n8806), .A(n7471), .ZN(n7473) );
  OAI211_X1 U9111 ( .C1(n9465), .C2(n9758), .A(n7474), .B(n7473), .ZN(P2_U3283) );
  AOI21_X1 U9112 ( .B1(n7476), .B2(n7475), .A(n4461), .ZN(n7481) );
  INV_X1 U9113 ( .A(n7688), .ZN(n8556) );
  INV_X1 U9114 ( .A(n7499), .ZN(n8558) );
  AOI22_X1 U9115 ( .A1(n8528), .A2(n8556), .B1(n8527), .B2(n8558), .ZN(n7478)
         );
  OAI211_X1 U9116 ( .C1(n8515), .C2(n7505), .A(n7478), .B(n7477), .ZN(n7479)
         );
  AOI21_X1 U9117 ( .B1(n9459), .B2(n8520), .A(n7479), .ZN(n7480) );
  OAI21_X1 U9118 ( .B1(n7481), .B2(n8522), .A(n7480), .ZN(P2_U3217) );
  XNOR2_X1 U9119 ( .A(n7482), .B(n7483), .ZN(n7487) );
  OAI22_X1 U9120 ( .A1(n7648), .A2(n9269), .B1(n7516), .B2(n9267), .ZN(n7486)
         );
  XNOR2_X1 U9121 ( .A(n7484), .B(n4647), .ZN(n9376) );
  NOR2_X1 U9122 ( .A1(n9376), .A2(n9295), .ZN(n7485) );
  AOI211_X1 U9123 ( .C1(n7487), .C2(n9223), .A(n7486), .B(n7485), .ZN(n9375)
         );
  INV_X1 U9124 ( .A(n9376), .ZN(n7494) );
  AND2_X1 U9125 ( .A1(n7488), .A2(n7521), .ZN(n7490) );
  OR2_X1 U9126 ( .A1(n7490), .A2(n7489), .ZN(n9372) );
  OAI22_X1 U9127 ( .A1(n9276), .A2(n9047), .B1(n7519), .B2(n9274), .ZN(n7491)
         );
  AOI21_X1 U9128 ( .B1(n7521), .B2(n9280), .A(n7491), .ZN(n7492) );
  OAI21_X1 U9129 ( .B1(n9372), .B2(n9163), .A(n7492), .ZN(n7493) );
  AOI21_X1 U9130 ( .B1(n7494), .B2(n7659), .A(n7493), .ZN(n7495) );
  OAI21_X1 U9131 ( .B1(n9375), .B2(n9253), .A(n7495), .ZN(P1_U3278) );
  NAND2_X1 U9132 ( .A1(n8037), .A2(n7499), .ZN(n7496) );
  NAND2_X1 U9133 ( .A1(n9459), .A2(n7642), .ZN(n8044) );
  INV_X1 U9134 ( .A(n8135), .ZN(n7504) );
  AOI21_X1 U9135 ( .B1(n7498), .B2(n7504), .A(n9725), .ZN(n7501) );
  OAI22_X1 U9136 ( .A1(n7688), .A2(n9761), .B1(n7499), .B2(n9763), .ZN(n7500)
         );
  AOI21_X1 U9137 ( .B1(n7501), .B2(n7608), .A(n7500), .ZN(n9461) );
  NAND2_X1 U9138 ( .A1(n8037), .A2(n8558), .ZN(n7502) );
  OAI21_X1 U9139 ( .B1(n4468), .B2(n7504), .A(n7607), .ZN(n9464) );
  NAND2_X1 U9140 ( .A1(n9464), .A2(n9746), .ZN(n7511) );
  OAI22_X1 U9141 ( .A1(n7202), .A2(n7397), .B1(n7505), .B2(n8817), .ZN(n7509)
         );
  INV_X1 U9142 ( .A(n9459), .ZN(n7506) );
  OAI21_X1 U9143 ( .B1(n7507), .B2(n7506), .A(n7610), .ZN(n9462) );
  NOR2_X1 U9144 ( .A1(n9462), .A2(n9757), .ZN(n7508) );
  AOI211_X1 U9145 ( .C1(n9731), .C2(n9459), .A(n7509), .B(n7508), .ZN(n7510)
         );
  OAI211_X1 U9146 ( .C1(n9749), .C2(n9461), .A(n7511), .B(n7510), .ZN(P2_U3282) );
  XNOR2_X1 U9147 ( .A(n7513), .B(n7512), .ZN(n7514) );
  XNOR2_X1 U9148 ( .A(n7515), .B(n7514), .ZN(n7523) );
  NOR2_X1 U9149 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5375), .ZN(n9551) );
  NOR2_X1 U9150 ( .A1(n9435), .A2(n7516), .ZN(n7517) );
  AOI211_X1 U9151 ( .C1(n9438), .C2(n9015), .A(n9551), .B(n7517), .ZN(n7518)
         );
  OAI21_X1 U9152 ( .B1(n9452), .B2(n7519), .A(n7518), .ZN(n7520) );
  AOI21_X1 U9153 ( .B1(n7521), .B2(n5797), .A(n7520), .ZN(n7522) );
  OAI21_X1 U9154 ( .B1(n7523), .B2(n9446), .A(n7522), .ZN(P1_U3232) );
  XNOR2_X1 U9155 ( .A(n7525), .B(n7524), .ZN(n7526) );
  XNOR2_X1 U9156 ( .A(n7527), .B(n7526), .ZN(n7535) );
  NOR2_X1 U9157 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7528), .ZN(n9567) );
  NOR2_X1 U9158 ( .A1(n9435), .A2(n7529), .ZN(n7530) );
  AOI211_X1 U9159 ( .C1(n9438), .C2(n9014), .A(n9567), .B(n7530), .ZN(n7531)
         );
  OAI21_X1 U9160 ( .B1(n9452), .B2(n7532), .A(n7531), .ZN(n7533) );
  AOI21_X1 U9161 ( .B1(n7628), .B2(n5797), .A(n7533), .ZN(n7534) );
  OAI21_X1 U9162 ( .B1(n7535), .B2(n9446), .A(n7534), .ZN(P1_U3213) );
  INV_X1 U9163 ( .A(n7536), .ZN(n7539) );
  OAI222_X1 U9164 ( .A1(n7537), .A2(P1_U3084), .B1(n7873), .B2(n7539), .C1(
        n9934), .C2(n7863), .ZN(P1_U3327) );
  OAI222_X1 U9165 ( .A1(P2_U3152), .A2(n7540), .B1(n8478), .B2(n7539), .C1(
        n7538), .C2(n7837), .ZN(P2_U3332) );
  INV_X1 U9166 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U9167 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7541) );
  AOI21_X1 U9168 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7541), .ZN(n9881) );
  NOR2_X1 U9169 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7542) );
  AOI21_X1 U9170 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7542), .ZN(n9884) );
  NOR2_X1 U9171 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7543) );
  AOI21_X1 U9172 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7543), .ZN(n9887) );
  NOR2_X1 U9173 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7544) );
  AOI21_X1 U9174 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7544), .ZN(n9890) );
  NOR2_X1 U9175 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7545) );
  AOI21_X1 U9176 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7545), .ZN(n9893) );
  NOR2_X1 U9177 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7552) );
  XOR2_X1 U9178 ( .A(n9986), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10229) );
  NAND2_X1 U9179 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7550) );
  INV_X1 U9180 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10030) );
  XNOR2_X1 U9181 ( .A(n10030), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U9182 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7548) );
  XNOR2_X1 U9183 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n7546), .ZN(n10225) );
  AOI21_X1 U9184 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9874) );
  INV_X1 U9185 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9878) );
  NAND3_X1 U9186 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9876) );
  OAI21_X1 U9187 ( .B1(n9874), .B2(n9878), .A(n9876), .ZN(n10224) );
  NAND2_X1 U9188 ( .A1(n10225), .A2(n10224), .ZN(n7547) );
  NAND2_X1 U9189 ( .A1(n7548), .A2(n7547), .ZN(n10226) );
  NAND2_X1 U9190 ( .A1(n10227), .A2(n10226), .ZN(n7549) );
  NAND2_X1 U9191 ( .A1(n7550), .A2(n7549), .ZN(n10228) );
  NOR2_X1 U9192 ( .A1(n10229), .A2(n10228), .ZN(n7551) );
  NOR2_X1 U9193 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  NOR2_X1 U9194 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7553), .ZN(n10211) );
  AND2_X1 U9195 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7553), .ZN(n10212) );
  NOR2_X1 U9196 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10212), .ZN(n7554) );
  NOR2_X1 U9197 ( .A1(n10211), .A2(n7554), .ZN(n7555) );
  NAND2_X1 U9198 ( .A1(n7555), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7557) );
  XOR2_X1 U9199 ( .A(n7555), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10210) );
  NAND2_X1 U9200 ( .A1(n10210), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7556) );
  NAND2_X1 U9201 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  NAND2_X1 U9202 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7558), .ZN(n7560) );
  INV_X1 U9203 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9908) );
  XNOR2_X1 U9204 ( .A(n9908), .B(n7558), .ZN(n10214) );
  NAND2_X1 U9205 ( .A1(n10214), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U9206 ( .A1(n7560), .A2(n7559), .ZN(n7561) );
  NAND2_X1 U9207 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7561), .ZN(n7563) );
  XOR2_X1 U9208 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7561), .Z(n10220) );
  NAND2_X1 U9209 ( .A1(n10220), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7562) );
  NAND2_X1 U9210 ( .A1(n7563), .A2(n7562), .ZN(n7564) );
  AND2_X1 U9211 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7564), .ZN(n7565) );
  XNOR2_X1 U9212 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7564), .ZN(n10222) );
  NOR2_X1 U9213 ( .A1(n10223), .A2(n10222), .ZN(n10221) );
  NOR2_X1 U9214 ( .A1(n7565), .A2(n10221), .ZN(n9902) );
  NAND2_X1 U9215 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7566) );
  OAI21_X1 U9216 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7566), .ZN(n9901) );
  NOR2_X1 U9217 ( .A1(n9902), .A2(n9901), .ZN(n9900) );
  AOI21_X1 U9218 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9900), .ZN(n9899) );
  NAND2_X1 U9219 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7567) );
  OAI21_X1 U9220 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7567), .ZN(n9898) );
  NOR2_X1 U9221 ( .A1(n9899), .A2(n9898), .ZN(n9897) );
  AOI21_X1 U9222 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9897), .ZN(n9896) );
  NOR2_X1 U9223 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7568) );
  AOI21_X1 U9224 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7568), .ZN(n9895) );
  NAND2_X1 U9225 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  OAI21_X1 U9226 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9894), .ZN(n9892) );
  NAND2_X1 U9227 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  OAI21_X1 U9228 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9891), .ZN(n9889) );
  NAND2_X1 U9229 ( .A1(n9890), .A2(n9889), .ZN(n9888) );
  OAI21_X1 U9230 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9888), .ZN(n9886) );
  NAND2_X1 U9231 ( .A1(n9887), .A2(n9886), .ZN(n9885) );
  OAI21_X1 U9232 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9885), .ZN(n9883) );
  NAND2_X1 U9233 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  OAI21_X1 U9234 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9882), .ZN(n9880) );
  NAND2_X1 U9235 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  OAI21_X1 U9236 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9879), .ZN(n10216) );
  NOR2_X1 U9237 ( .A1(n10217), .A2(n10216), .ZN(n7569) );
  NAND2_X1 U9238 ( .A1(n10217), .A2(n10216), .ZN(n10215) );
  OAI21_X1 U9239 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7569), .A(n10215), .ZN(
        n7571) );
  XNOR2_X1 U9240 ( .A(n4733), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7570) );
  XNOR2_X1 U9241 ( .A(n7571), .B(n7570), .ZN(ADD_1071_U4) );
  XNOR2_X1 U9242 ( .A(n7573), .B(n7572), .ZN(n7577) );
  INV_X1 U9243 ( .A(n7680), .ZN(n8555) );
  INV_X1 U9244 ( .A(n7846), .ZN(n8553) );
  AOI22_X1 U9245 ( .A1(n8783), .A2(n8555), .B1(n8553), .B2(n8781), .ZN(n7714)
         );
  OAI22_X1 U9246 ( .A1(n8541), .A2(n7714), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10004), .ZN(n7575) );
  NOR2_X1 U9247 ( .A1(n4829), .A2(n8546), .ZN(n7574) );
  AOI211_X1 U9248 ( .C1(n8543), .C2(n7718), .A(n7575), .B(n7574), .ZN(n7576)
         );
  OAI21_X1 U9249 ( .B1(n7577), .B2(n8522), .A(n7576), .ZN(P2_U3230) );
  INV_X1 U9250 ( .A(n7583), .ZN(n7581) );
  NAND2_X1 U9251 ( .A1(n7578), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U9252 ( .A1(n7579), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8157) );
  OAI211_X1 U9253 ( .C1(n7581), .C2(n8478), .A(n7580), .B(n8157), .ZN(P2_U3331) );
  NAND2_X1 U9254 ( .A1(n7583), .A2(n7582), .ZN(n7585) );
  OAI211_X1 U9255 ( .C1(n7863), .C2(n9923), .A(n7585), .B(n7584), .ZN(P1_U3326) );
  XOR2_X1 U9256 ( .A(n7587), .B(n7586), .Z(n7588) );
  XNOR2_X1 U9257 ( .A(n7589), .B(n7588), .ZN(n7594) );
  INV_X1 U9258 ( .A(n7649), .ZN(n9013) );
  AND2_X1 U9259 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9580) );
  NOR2_X1 U9260 ( .A1(n9435), .A2(n7648), .ZN(n7590) );
  AOI211_X1 U9261 ( .C1(n9438), .C2(n9013), .A(n9580), .B(n7590), .ZN(n7591)
         );
  OAI21_X1 U9262 ( .B1(n9452), .B2(n7656), .A(n7591), .ZN(n7592) );
  AOI21_X1 U9263 ( .B1(n9365), .B2(n5797), .A(n7592), .ZN(n7593) );
  OAI21_X1 U9264 ( .B1(n7594), .B2(n9446), .A(n7593), .ZN(P1_U3239) );
  OAI21_X1 U9265 ( .B1(n7596), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7595), .ZN(
        n7898) );
  XNOR2_X1 U9266 ( .A(n7898), .B(n7909), .ZN(n7597) );
  INV_X1 U9267 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U9268 ( .A1(n7597), .A2(n10120), .ZN(n7900) );
  OAI21_X1 U9269 ( .B1(n7597), .B2(n10120), .A(n7900), .ZN(n7605) );
  AOI21_X1 U9270 ( .B1(n7599), .B2(n10091), .A(n7598), .ZN(n7908) );
  XNOR2_X1 U9271 ( .A(n7908), .B(n7899), .ZN(n7600) );
  NAND2_X1 U9272 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7600), .ZN(n7910) );
  OAI211_X1 U9273 ( .C1(n7600), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9708), .B(
        n7910), .ZN(n7603) );
  INV_X1 U9274 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7640) );
  NOR2_X1 U9275 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7640), .ZN(n7601) );
  AOI21_X1 U9276 ( .B1(n9715), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7601), .ZN(
        n7602) );
  OAI211_X1 U9277 ( .C1(n9711), .C2(n7899), .A(n7603), .B(n7602), .ZN(n7604)
         );
  AOI21_X1 U9278 ( .B1(n9710), .B2(n7605), .A(n7604), .ZN(n7606) );
  INV_X1 U9279 ( .A(n7606), .ZN(P2_U3260) );
  INV_X1 U9280 ( .A(n7642), .ZN(n8557) );
  NAND2_X1 U9281 ( .A1(n7677), .A2(n7688), .ZN(n8047) );
  NAND2_X1 U9282 ( .A1(n8048), .A2(n8047), .ZN(n8137) );
  XNOR2_X1 U9283 ( .A(n7679), .B(n8137), .ZN(n9457) );
  INV_X1 U9284 ( .A(n9457), .ZN(n7616) );
  NAND2_X1 U9285 ( .A1(n7608), .A2(n8043), .ZN(n7683) );
  INV_X1 U9286 ( .A(n8137), .ZN(n8046) );
  XNOR2_X1 U9287 ( .A(n7683), .B(n8046), .ZN(n7609) );
  OAI222_X1 U9288 ( .A1(n9763), .A2(n7642), .B1(n9761), .B2(n7680), .C1(n9725), 
        .C2(n7609), .ZN(n9455) );
  INV_X1 U9289 ( .A(n7610), .ZN(n7611) );
  INV_X1 U9290 ( .A(n7677), .ZN(n9453) );
  OAI21_X1 U9291 ( .B1(n7611), .B2(n9453), .A(n7692), .ZN(n9454) );
  AOI22_X1 U9292 ( .A1(n9749), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7639), .B2(
        n9771), .ZN(n7613) );
  NAND2_X1 U9293 ( .A1(n7677), .A2(n9731), .ZN(n7612) );
  OAI211_X1 U9294 ( .C1(n9454), .C2(n9757), .A(n7613), .B(n7612), .ZN(n7614)
         );
  AOI21_X1 U9295 ( .B1(n9455), .B2(n7202), .A(n7614), .ZN(n7615) );
  OAI21_X1 U9296 ( .B1(n7616), .B2(n8808), .A(n7615), .ZN(P2_U3281) );
  XNOR2_X1 U9297 ( .A(n7618), .B(n7617), .ZN(n7623) );
  INV_X1 U9298 ( .A(n7708), .ZN(n8554) );
  AOI22_X1 U9299 ( .A1(n8527), .A2(n8554), .B1(n8528), .B2(n8552), .ZN(n7619)
         );
  NAND2_X1 U9300 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3152), .ZN(n8638) );
  OAI211_X1 U9301 ( .C1(n7620), .C2(n8515), .A(n7619), .B(n8638), .ZN(n7621)
         );
  AOI21_X1 U9302 ( .B1(n8888), .B2(n8520), .A(n7621), .ZN(n7622) );
  OAI21_X1 U9303 ( .B1(n7623), .B2(n8522), .A(n7622), .ZN(P2_U3240) );
  INV_X1 U9304 ( .A(n9014), .ZN(n7631) );
  NAND2_X1 U9305 ( .A1(n9365), .A2(n7631), .ZN(n8214) );
  NAND2_X1 U9306 ( .A1(n7647), .A2(n8214), .ZN(n7750) );
  OR2_X1 U9307 ( .A1(n9365), .A2(n7631), .ZN(n7749) );
  NAND2_X1 U9308 ( .A1(n7750), .A2(n7749), .ZN(n7625) );
  OR2_X1 U9309 ( .A1(n7743), .A2(n7649), .ZN(n8365) );
  NAND2_X1 U9310 ( .A1(n7743), .A2(n7649), .ZN(n8217) );
  NAND2_X1 U9311 ( .A1(n8365), .A2(n8217), .ZN(n7744) );
  XNOR2_X1 U9312 ( .A(n7625), .B(n7744), .ZN(n7627) );
  OAI22_X1 U9313 ( .A1(n8992), .A2(n9269), .B1(n7631), .B2(n9267), .ZN(n7626)
         );
  AOI21_X1 U9314 ( .B1(n7627), .B2(n9223), .A(n7626), .ZN(n9478) );
  INV_X1 U9315 ( .A(n9365), .ZN(n7655) );
  INV_X1 U9316 ( .A(n7744), .ZN(n8257) );
  XNOR2_X1 U9317 ( .A(n7745), .B(n8257), .ZN(n9481) );
  NAND2_X1 U9318 ( .A1(n9481), .A2(n9283), .ZN(n7638) );
  INV_X1 U9319 ( .A(n7743), .ZN(n9479) );
  OAI211_X1 U9320 ( .C1(n7654), .C2(n9479), .A(n9366), .B(n7761), .ZN(n9477)
         );
  INV_X1 U9321 ( .A(n9477), .ZN(n7636) );
  INV_X1 U9322 ( .A(n9280), .ZN(n9258) );
  AOI22_X1 U9323 ( .A1(n9278), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7736), .B2(
        n9254), .ZN(n7633) );
  OAI21_X1 U9324 ( .B1(n9479), .B2(n9258), .A(n7633), .ZN(n7634) );
  AOI21_X1 U9325 ( .B1(n7636), .B2(n7635), .A(n7634), .ZN(n7637) );
  OAI211_X1 U9326 ( .C1(n9278), .C2(n9478), .A(n7638), .B(n7637), .ZN(P1_U3275) );
  XOR2_X1 U9327 ( .A(n7665), .B(n7663), .Z(n7667) );
  XNOR2_X1 U9328 ( .A(n7667), .B(n7666), .ZN(n7646) );
  INV_X1 U9329 ( .A(n7639), .ZN(n7641) );
  OAI22_X1 U9330 ( .A1(n8515), .A2(n7641), .B1(n7640), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n7644) );
  OAI22_X1 U9331 ( .A1(n7680), .A2(n8516), .B1(n8517), .B2(n7642), .ZN(n7643)
         );
  AOI211_X1 U9332 ( .C1(n7677), .C2(n8520), .A(n7644), .B(n7643), .ZN(n7645)
         );
  OAI21_X1 U9333 ( .B1(n7646), .B2(n8522), .A(n7645), .ZN(P2_U3243) );
  AND2_X1 U9334 ( .A1(n7749), .A2(n8214), .ZN(n8359) );
  INV_X1 U9335 ( .A(n8359), .ZN(n8255) );
  XNOR2_X1 U9336 ( .A(n7647), .B(n8255), .ZN(n7653) );
  OAI22_X1 U9337 ( .A1(n7649), .A2(n9269), .B1(n7648), .B2(n9267), .ZN(n7652)
         );
  XNOR2_X1 U9338 ( .A(n7650), .B(n8255), .ZN(n9370) );
  NOR2_X1 U9339 ( .A1(n9370), .A2(n9295), .ZN(n7651) );
  AOI211_X1 U9340 ( .C1(n9223), .C2(n7653), .A(n7652), .B(n7651), .ZN(n9369)
         );
  AOI21_X1 U9341 ( .B1(n9365), .B2(n4457), .A(n7654), .ZN(n9367) );
  NOR2_X1 U9342 ( .A1(n7655), .A2(n9258), .ZN(n7658) );
  OAI22_X1 U9343 ( .A1(n9276), .A2(n5432), .B1(n7656), .B2(n9274), .ZN(n7657)
         );
  AOI211_X1 U9344 ( .C1(n9367), .C2(n9226), .A(n7658), .B(n7657), .ZN(n7662)
         );
  INV_X1 U9345 ( .A(n9370), .ZN(n7660) );
  NAND2_X1 U9346 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  OAI211_X1 U9347 ( .C1(n9369), .C2(n9253), .A(n7662), .B(n7661), .ZN(P1_U3276) );
  INV_X1 U9348 ( .A(n7663), .ZN(n7664) );
  OAI22_X1 U9349 ( .A1(n7667), .A2(n7666), .B1(n7665), .B2(n7664), .ZN(n7671)
         );
  NOR2_X1 U9350 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  XNOR2_X1 U9351 ( .A(n7671), .B(n7670), .ZN(n7676) );
  INV_X1 U9352 ( .A(n7693), .ZN(n7673) );
  AOI22_X1 U9353 ( .A1(n8527), .A2(n8556), .B1(n8528), .B2(n8554), .ZN(n7672)
         );
  NAND2_X1 U9354 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8616) );
  OAI211_X1 U9355 ( .C1(n7673), .C2(n8515), .A(n7672), .B(n8616), .ZN(n7674)
         );
  AOI21_X1 U9356 ( .B1(n8899), .B2(n8520), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9357 ( .B1(n7676), .B2(n8522), .A(n7675), .ZN(P2_U3228) );
  NOR2_X1 U9358 ( .A1(n7677), .A2(n8556), .ZN(n7678) );
  OR2_X1 U9359 ( .A1(n8899), .A2(n7680), .ZN(n8051) );
  NAND2_X1 U9360 ( .A1(n8899), .A2(n7680), .ZN(n8050) );
  NAND2_X1 U9361 ( .A1(n8051), .A2(n8050), .ZN(n8138) );
  AND2_X2 U9362 ( .A1(n7681), .A2(n8138), .ZN(n7707) );
  NOR2_X1 U9363 ( .A1(n7681), .A2(n8138), .ZN(n7682) );
  OR2_X1 U9364 ( .A1(n7707), .A2(n7682), .ZN(n8903) );
  INV_X1 U9365 ( .A(n8903), .ZN(n7691) );
  INV_X1 U9366 ( .A(n9769), .ZN(n9831) );
  NAND2_X1 U9367 ( .A1(n7683), .A2(n8046), .ZN(n7684) );
  NAND2_X1 U9368 ( .A1(n7686), .A2(n8138), .ZN(n7687) );
  AOI21_X1 U9369 ( .B1(n7713), .B2(n7687), .A(n9725), .ZN(n7690) );
  OAI22_X1 U9370 ( .A1(n7688), .A2(n9763), .B1(n7708), .B2(n9761), .ZN(n7689)
         );
  AOI211_X1 U9371 ( .C1(n7691), .C2(n9831), .A(n7690), .B(n7689), .ZN(n8902)
         );
  AOI21_X1 U9372 ( .B1(n8899), .B2(n7692), .A(n7717), .ZN(n8900) );
  AOI22_X1 U9373 ( .A1(n9773), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7693), .B2(
        n9771), .ZN(n7694) );
  OAI21_X1 U9374 ( .B1(n4626), .B2(n9775), .A(n7694), .ZN(n7696) );
  NOR2_X1 U9375 ( .A1(n8903), .A2(n9758), .ZN(n7695) );
  AOI211_X1 U9376 ( .C1(n8900), .C2(n8806), .A(n7696), .B(n7695), .ZN(n7697)
         );
  OAI21_X1 U9377 ( .B1(n9749), .B2(n8902), .A(n7697), .ZN(P2_U3280) );
  INV_X1 U9378 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7705) );
  INV_X1 U9379 ( .A(n7700), .ZN(n7702) );
  NAND2_X1 U9380 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  INV_X1 U9381 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7931) );
  MUX2_X1 U9382 ( .A(n7931), .B(n7705), .S(n5497), .Z(n7821) );
  XNOR2_X1 U9383 ( .A(n7821), .B(SI_29_), .ZN(n7704) );
  INV_X1 U9384 ( .A(n8174), .ZN(n7932) );
  OAI222_X1 U9385 ( .A1(n7863), .A2(n7705), .B1(P1_U3084), .B2(n4997), .C1(
        n7873), .C2(n7932), .ZN(P1_U3324) );
  OR2_X1 U9386 ( .A1(n8895), .A2(n7708), .ZN(n8057) );
  NAND2_X1 U9387 ( .A1(n8895), .A2(n7708), .ZN(n8055) );
  NAND2_X1 U9388 ( .A1(n8057), .A2(n8055), .ZN(n8139) );
  OAI21_X1 U9389 ( .B1(n7709), .B2(n8139), .A(n7807), .ZN(n7710) );
  INV_X1 U9390 ( .A(n7710), .ZN(n8898) );
  INV_X1 U9391 ( .A(n8050), .ZN(n7711) );
  NOR2_X1 U9392 ( .A1(n8139), .A2(n7711), .ZN(n7712) );
  NAND2_X1 U9393 ( .A1(n7813), .A2(n9766), .ZN(n7716) );
  INV_X1 U9394 ( .A(n8139), .ZN(n8053) );
  AOI21_X1 U9395 ( .B1(n7713), .B2(n8050), .A(n8053), .ZN(n7715) );
  OAI21_X1 U9396 ( .B1(n7716), .B2(n7715), .A(n7714), .ZN(n8893) );
  AOI211_X1 U9397 ( .C1(n8895), .C2(n4628), .A(n9842), .B(n7808), .ZN(n8894)
         );
  NAND2_X1 U9398 ( .A1(n8894), .A2(n9745), .ZN(n7720) );
  AOI22_X1 U9399 ( .A1(n9749), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n7718), .B2(
        n9771), .ZN(n7719) );
  OAI211_X1 U9400 ( .C1(n4829), .C2(n9775), .A(n7720), .B(n7719), .ZN(n7721)
         );
  AOI21_X1 U9401 ( .B1(n8893), .B2(n7202), .A(n7721), .ZN(n7722) );
  OAI21_X1 U9402 ( .B1(n8898), .B2(n8808), .A(n7722), .ZN(P2_U3279) );
  INV_X1 U9403 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7723) );
  INV_X1 U9404 ( .A(n7875), .ZN(n7934) );
  OAI222_X1 U9405 ( .A1(n7863), .A2(n7723), .B1(P1_U3084), .B2(n5777), .C1(
        n7873), .C2(n7934), .ZN(P1_U3325) );
  INV_X1 U9406 ( .A(n8884), .ZN(n8455) );
  OAI21_X1 U9407 ( .B1(n7726), .B2(n7725), .A(n7724), .ZN(n7727) );
  NAND2_X1 U9408 ( .A1(n7727), .A2(n8535), .ZN(n7731) );
  OAI22_X1 U9409 ( .A1(n7846), .A2(n9763), .B1(n8456), .B2(n9761), .ZN(n7851)
         );
  INV_X1 U9410 ( .A(n7851), .ZN(n7728) );
  NAND2_X1 U9411 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7928) );
  OAI21_X1 U9412 ( .B1(n8541), .B2(n7728), .A(n7928), .ZN(n7729) );
  AOI21_X1 U9413 ( .B1(n7857), .B2(n8543), .A(n7729), .ZN(n7730) );
  OAI211_X1 U9414 ( .C1(n8455), .C2(n8546), .A(n7731), .B(n7730), .ZN(P2_U3221) );
  INV_X1 U9415 ( .A(n7732), .ZN(n7733) );
  AOI21_X1 U9416 ( .B1(n7735), .B2(n7734), .A(n7733), .ZN(n7742) );
  NAND2_X1 U9417 ( .A1(n9003), .A2(n7736), .ZN(n7739) );
  NOR2_X1 U9418 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7737), .ZN(n9592) );
  AOI21_X1 U9419 ( .B1(n8980), .B2(n9014), .A(n9592), .ZN(n7738) );
  OAI211_X1 U9420 ( .C1(n8992), .C2(n8983), .A(n7739), .B(n7738), .ZN(n7740)
         );
  AOI21_X1 U9421 ( .B1(n7743), .B2(n5797), .A(n7740), .ZN(n7741) );
  OAI21_X1 U9422 ( .B1(n7742), .B2(n9446), .A(n7741), .ZN(P1_U3224) );
  NAND2_X1 U9423 ( .A1(n9356), .A2(n7800), .ZN(n8186) );
  OAI21_X1 U9424 ( .B1(n7794), .B2(n8992), .A(n7758), .ZN(n7746) );
  OAI21_X1 U9425 ( .B1(n9012), .B2(n9359), .A(n7746), .ZN(n7747) );
  AOI21_X1 U9426 ( .B1(n8259), .B2(n7747), .A(n7795), .ZN(n7748) );
  INV_X1 U9427 ( .A(n7748), .ZN(n9358) );
  INV_X1 U9428 ( .A(n9077), .ZN(n9247) );
  AND2_X1 U9429 ( .A1(n8365), .A2(n7749), .ZN(n8362) );
  INV_X1 U9430 ( .A(n8217), .ZN(n8366) );
  NAND2_X1 U9431 ( .A1(n9359), .A2(n8992), .ZN(n8185) );
  NAND2_X1 U9432 ( .A1(n7764), .A2(n8185), .ZN(n7798) );
  OR2_X1 U9433 ( .A1(n9359), .A2(n8992), .ZN(n7796) );
  NAND2_X1 U9434 ( .A1(n7798), .A2(n7796), .ZN(n7751) );
  XNOR2_X1 U9435 ( .A(n7751), .B(n8259), .ZN(n7752) );
  OAI222_X1 U9436 ( .A1(n9267), .A2(n8992), .B1(n9269), .B2(n9247), .C1(n9265), 
        .C2(n7752), .ZN(n9354) );
  INV_X1 U9437 ( .A(n9356), .ZN(n7755) );
  AOI211_X1 U9438 ( .C1(n9356), .C2(n7759), .A(n9688), .B(n7801), .ZN(n9355)
         );
  NAND2_X1 U9439 ( .A1(n9355), .A2(n9252), .ZN(n7754) );
  AOI22_X1 U9440 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9253), .B1(n8994), .B2(
        n9254), .ZN(n7753) );
  OAI211_X1 U9441 ( .C1(n7755), .C2(n9258), .A(n7754), .B(n7753), .ZN(n7756)
         );
  AOI21_X1 U9442 ( .B1(n9354), .B2(n9276), .A(n7756), .ZN(n7757) );
  OAI21_X1 U9443 ( .B1(n9358), .B2(n9262), .A(n7757), .ZN(P1_U3273) );
  NAND2_X1 U9444 ( .A1(n7796), .A2(n8185), .ZN(n8368) );
  INV_X1 U9445 ( .A(n8368), .ZN(n8258) );
  XNOR2_X1 U9446 ( .A(n7758), .B(n8258), .ZN(n9364) );
  INV_X1 U9447 ( .A(n7759), .ZN(n7760) );
  AOI21_X1 U9448 ( .B1(n9359), .B2(n7761), .A(n7760), .ZN(n9360) );
  INV_X1 U9449 ( .A(n7762), .ZN(n7791) );
  AOI22_X1 U9450 ( .A1(n9278), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n7791), .B2(
        n9254), .ZN(n7763) );
  OAI21_X1 U9451 ( .B1(n7794), .B2(n9258), .A(n7763), .ZN(n7767) );
  XNOR2_X1 U9452 ( .A(n7764), .B(n8368), .ZN(n7765) );
  AOI222_X1 U9453 ( .A1(n9223), .A2(n7765), .B1(n9011), .B2(n9218), .C1(n9013), 
        .C2(n9220), .ZN(n9362) );
  NOR2_X1 U9454 ( .A1(n9362), .A2(n9253), .ZN(n7766) );
  AOI211_X1 U9455 ( .C1(n9360), .C2(n9226), .A(n7767), .B(n7766), .ZN(n7768)
         );
  OAI21_X1 U9456 ( .B1(n9364), .B2(n9262), .A(n7768), .ZN(P1_U3274) );
  XNOR2_X1 U9457 ( .A(n7770), .B(n7769), .ZN(n7776) );
  INV_X1 U9458 ( .A(n8792), .ZN(n7772) );
  OAI22_X1 U9459 ( .A1(n8515), .A2(n7772), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7771), .ZN(n7774) );
  INV_X1 U9460 ( .A(n8552), .ZN(n8800) );
  OAI22_X1 U9461 ( .A1(n8800), .A2(n8517), .B1(n8516), .B2(n8799), .ZN(n7773)
         );
  AOI211_X1 U9462 ( .C1(n8878), .C2(n8520), .A(n7774), .B(n7773), .ZN(n7775)
         );
  OAI21_X1 U9463 ( .B1(n7776), .B2(n8522), .A(n7775), .ZN(P2_U3235) );
  XNOR2_X1 U9464 ( .A(n7777), .B(n7778), .ZN(n7784) );
  INV_X1 U9465 ( .A(n8776), .ZN(n7780) );
  OAI22_X1 U9466 ( .A1(n8515), .A2(n7780), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7779), .ZN(n7782) );
  OAI22_X1 U9467 ( .A1(n8493), .A2(n8516), .B1(n8517), .B2(n8456), .ZN(n7781)
         );
  AOI211_X1 U9468 ( .C1(n8873), .C2(n8520), .A(n7782), .B(n7781), .ZN(n7783)
         );
  OAI21_X1 U9469 ( .B1(n7784), .B2(n8522), .A(n7783), .ZN(P2_U3225) );
  OAI21_X1 U9470 ( .B1(n7787), .B2(n7785), .A(n7786), .ZN(n7788) );
  NAND2_X1 U9471 ( .A1(n7788), .A2(n9002), .ZN(n7793) );
  AND2_X1 U9472 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9600) );
  AOI21_X1 U9473 ( .B1(n9013), .B2(n8980), .A(n9600), .ZN(n7789) );
  OAI21_X1 U9474 ( .B1(n7800), .B2(n8983), .A(n7789), .ZN(n7790) );
  AOI21_X1 U9475 ( .B1(n9003), .B2(n7791), .A(n7790), .ZN(n7792) );
  OAI211_X1 U9476 ( .C1(n7794), .C2(n9010), .A(n7793), .B(n7792), .ZN(P1_U3226) );
  OR2_X1 U9477 ( .A1(n9351), .A2(n9247), .ZN(n8376) );
  NAND2_X1 U9478 ( .A1(n9351), .A2(n9247), .ZN(n9093) );
  NAND2_X1 U9479 ( .A1(n8376), .A2(n9093), .ZN(n9094) );
  XOR2_X1 U9480 ( .A(n9094), .B(n9080), .Z(n9353) );
  AOI22_X1 U9481 ( .A1(n9351), .A2(n9280), .B1(n9278), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n7806) );
  INV_X1 U9482 ( .A(n9081), .ZN(n9234) );
  AND2_X1 U9483 ( .A1(n8377), .A2(n7796), .ZN(n8372) );
  INV_X1 U9484 ( .A(n8186), .ZN(n7797) );
  XOR2_X1 U9485 ( .A(n9094), .B(n9095), .Z(n7799) );
  OAI222_X1 U9486 ( .A1(n9267), .A2(n7800), .B1(n9269), .B2(n9234), .C1(n7799), 
        .C2(n9265), .ZN(n9349) );
  INV_X1 U9487 ( .A(n7801), .ZN(n7802) );
  AOI211_X1 U9488 ( .C1(n9351), .C2(n7802), .A(n9688), .B(n9248), .ZN(n9350)
         );
  INV_X1 U9489 ( .A(n9350), .ZN(n7803) );
  OAI22_X1 U9490 ( .A1(n7803), .A2(n9275), .B1(n9274), .B2(n8935), .ZN(n7804)
         );
  OAI21_X1 U9491 ( .B1(n9349), .B2(n7804), .A(n9276), .ZN(n7805) );
  OAI211_X1 U9492 ( .C1(n9353), .C2(n9262), .A(n7806), .B(n7805), .ZN(P1_U3272) );
  NAND2_X1 U9493 ( .A1(n8888), .A2(n7846), .ZN(n8060) );
  NAND2_X1 U9494 ( .A1(n8063), .A2(n8060), .ZN(n7848) );
  INV_X1 U9495 ( .A(n7848), .ZN(n8141) );
  XNOR2_X1 U9496 ( .A(n7849), .B(n8141), .ZN(n8892) );
  INV_X1 U9497 ( .A(n7808), .ZN(n7810) );
  NAND2_X1 U9498 ( .A1(n7808), .A2(n7847), .ZN(n7854) );
  INV_X1 U9499 ( .A(n7854), .ZN(n7809) );
  AOI21_X1 U9500 ( .B1(n8888), .B2(n7810), .A(n7809), .ZN(n8889) );
  AOI22_X1 U9501 ( .A1(n9749), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n7811), .B2(
        n9771), .ZN(n7812) );
  OAI21_X1 U9502 ( .B1(n7847), .B2(n9775), .A(n7812), .ZN(n7818) );
  NAND2_X1 U9503 ( .A1(n7813), .A2(n8057), .ZN(n7814) );
  OAI211_X1 U9504 ( .C1(n8141), .C2(n7814), .A(n7938), .B(n9766), .ZN(n7816)
         );
  AOI22_X1 U9505 ( .A1(n8554), .A2(n8783), .B1(n8781), .B2(n8552), .ZN(n7815)
         );
  NOR2_X1 U9506 ( .A1(n8891), .A2(n8740), .ZN(n7817) );
  AOI211_X1 U9507 ( .C1(n8889), .C2(n8806), .A(n7818), .B(n7817), .ZN(n7819)
         );
  OAI21_X1 U9508 ( .B1(n8892), .B2(n8808), .A(n7819), .ZN(P2_U3278) );
  INV_X1 U9509 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7828) );
  INV_X1 U9510 ( .A(SI_29_), .ZN(n7820) );
  AND2_X1 U9511 ( .A1(n7821), .A2(n7820), .ZN(n7824) );
  INV_X1 U9512 ( .A(n7821), .ZN(n7822) );
  NAND2_X1 U9513 ( .A1(n7822), .A2(SI_29_), .ZN(n7823) );
  MUX2_X1 U9514 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7826), .Z(n7830) );
  INV_X1 U9515 ( .A(n8165), .ZN(n8477) );
  OAI222_X1 U9516 ( .A1(n7863), .A2(n7828), .B1(n7873), .B2(n8477), .C1(n7827), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  NAND2_X1 U9517 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  MUX2_X1 U9518 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7833), .Z(n7834) );
  XNOR2_X1 U9519 ( .A(n7834), .B(SI_31_), .ZN(n7835) );
  INV_X1 U9520 ( .A(n8162), .ZN(n7845) );
  NAND3_X1 U9521 ( .A1(n7836), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n7838) );
  OAI22_X1 U9522 ( .A1(n5816), .A2(n7838), .B1(n6422), .B2(n7837), .ZN(n7839)
         );
  INV_X1 U9523 ( .A(n7839), .ZN(n7840) );
  OAI21_X1 U9524 ( .B1(n7845), .B2(n8478), .A(n7840), .ZN(P2_U3327) );
  NOR4_X1 U9525 ( .A1(n7841), .A2(P1_IR_REG_30__SCAN_IN), .A3(n7842), .A4(
        P1_U3084), .ZN(n7843) );
  AOI21_X1 U9526 ( .B1(n7870), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n7843), .ZN(
        n7844) );
  OAI21_X1 U9527 ( .B1(n7845), .B2(n7873), .A(n7844), .ZN(P1_U3322) );
  OR2_X1 U9528 ( .A1(n8884), .A2(n8800), .ZN(n8066) );
  NAND2_X1 U9529 ( .A1(n8884), .A2(n8800), .ZN(n8795) );
  NAND2_X1 U9530 ( .A1(n8066), .A2(n8795), .ZN(n8120) );
  XNOR2_X1 U9531 ( .A(n8453), .B(n8120), .ZN(n8887) );
  NAND2_X1 U9532 ( .A1(n7938), .A2(n8063), .ZN(n7850) );
  XNOR2_X1 U9533 ( .A(n7850), .B(n8120), .ZN(n7852) );
  AOI21_X1 U9534 ( .B1(n7852), .B2(n9766), .A(n7851), .ZN(n8886) );
  INV_X1 U9535 ( .A(n8791), .ZN(n7853) );
  AOI211_X1 U9536 ( .C1(n8884), .C2(n7854), .A(n9842), .B(n7853), .ZN(n8883)
         );
  NAND2_X1 U9537 ( .A1(n8883), .A2(n8707), .ZN(n7855) );
  OAI211_X1 U9538 ( .C1(n8887), .C2(n9769), .A(n8886), .B(n7855), .ZN(n7856)
         );
  NAND2_X1 U9539 ( .A1(n7856), .A2(n7202), .ZN(n7862) );
  INV_X1 U9540 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n7859) );
  INV_X1 U9541 ( .A(n7857), .ZN(n7858) );
  OAI22_X1 U9542 ( .A1(n7202), .A2(n7859), .B1(n7858), .B2(n8817), .ZN(n7860)
         );
  AOI21_X1 U9543 ( .B1(n8884), .B2(n9731), .A(n7860), .ZN(n7861) );
  OAI211_X1 U9544 ( .C1(n8887), .C2(n9758), .A(n7862), .B(n7861), .ZN(P2_U3277) );
  OAI222_X1 U9545 ( .A1(n7866), .A2(P1_U3084), .B1(n7873), .B2(n7865), .C1(
        n7864), .C2(n7863), .ZN(P1_U3329) );
  AOI22_X1 U9546 ( .A1(n7867), .A2(P1_STATE_REG_SCAN_IN), .B1(n7870), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n7868) );
  OAI21_X1 U9547 ( .B1(n7869), .B2(n7873), .A(n7868), .ZN(P1_U3350) );
  AOI22_X1 U9548 ( .A1(n7871), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n7870), .ZN(n7872) );
  OAI21_X1 U9549 ( .B1(n7874), .B2(n7873), .A(n7872), .ZN(P1_U3349) );
  NAND2_X1 U9550 ( .A1(n7875), .A2(n5306), .ZN(n7877) );
  NAND2_X1 U9551 ( .A1(n5732), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U9552 ( .A1(n9303), .A2(n7878), .ZN(n7880) );
  NAND2_X1 U9553 ( .A1(n9147), .A2(n5167), .ZN(n7879) );
  NAND2_X1 U9554 ( .A1(n7880), .A2(n7879), .ZN(n7882) );
  XNOR2_X1 U9555 ( .A(n7882), .B(n7881), .ZN(n7886) );
  NAND2_X1 U9556 ( .A1(n9303), .A2(n5167), .ZN(n7883) );
  OAI21_X1 U9557 ( .B1(n9092), .B2(n7884), .A(n7883), .ZN(n7885) );
  XNOR2_X1 U9558 ( .A(n7886), .B(n7885), .ZN(n7887) );
  INV_X1 U9559 ( .A(n7887), .ZN(n7892) );
  NAND3_X1 U9560 ( .A1(n7892), .A2(n9002), .A3(n7891), .ZN(n7896) );
  INV_X1 U9561 ( .A(n7888), .ZN(n9133) );
  AOI22_X1 U9562 ( .A1(n9133), .A2(n9003), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7890) );
  NAND2_X1 U9563 ( .A1(n9157), .A2(n8980), .ZN(n7889) );
  OAI211_X1 U9564 ( .C1(n9129), .C2(n8983), .A(n7890), .B(n7889), .ZN(n7894)
         );
  NOR3_X1 U9565 ( .A1(n7892), .A2(n7891), .A3(n9446), .ZN(n7893) );
  AOI211_X1 U9566 ( .C1(n5797), .C2(n9303), .A(n7894), .B(n7893), .ZN(n7895)
         );
  NAND2_X1 U9567 ( .A1(n7899), .A2(n7898), .ZN(n7901) );
  NAND2_X1 U9568 ( .A1(n7901), .A2(n7900), .ZN(n8614) );
  XNOR2_X1 U9569 ( .A(n7902), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8613) );
  NOR2_X1 U9570 ( .A1(n8614), .A2(n8613), .ZN(n8612) );
  NAND2_X1 U9571 ( .A1(n7915), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7903) );
  OAI21_X1 U9572 ( .B1(n7915), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7903), .ZN(
        n8629) );
  NOR2_X1 U9573 ( .A1(n7904), .A2(n7920), .ZN(n7906) );
  INV_X1 U9574 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9913) );
  XNOR2_X1 U9575 ( .A(n8640), .B(n7905), .ZN(n8642) );
  NOR2_X1 U9576 ( .A1(n9913), .A2(n8642), .ZN(n8641) );
  NOR2_X1 U9577 ( .A1(n7906), .A2(n8641), .ZN(n7907) );
  XNOR2_X1 U9578 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n7907), .ZN(n7925) );
  INV_X1 U9579 ( .A(n7925), .ZN(n7923) );
  INV_X1 U9580 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7919) );
  INV_X1 U9581 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U9582 ( .A1(n7909), .A2(n7908), .ZN(n7911) );
  NAND2_X1 U9583 ( .A1(n7911), .A2(n7910), .ZN(n8611) );
  INV_X1 U9584 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7912) );
  NAND2_X1 U9585 ( .A1(n8617), .A2(n7912), .ZN(n7913) );
  OAI21_X1 U9586 ( .B1(n8617), .B2(n7912), .A(n7913), .ZN(n8610) );
  NOR2_X1 U9587 ( .A1(n8611), .A2(n8610), .ZN(n8609) );
  INV_X1 U9588 ( .A(n7913), .ZN(n7914) );
  NOR2_X1 U9589 ( .A1(n8609), .A2(n7914), .ZN(n8624) );
  XNOR2_X1 U9590 ( .A(n7915), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8623) );
  INV_X1 U9591 ( .A(n8623), .ZN(n7916) );
  NAND2_X1 U9592 ( .A1(n8624), .A2(n7916), .ZN(n7917) );
  OAI21_X1 U9593 ( .B1(n7918), .B2(n8627), .A(n7917), .ZN(n8637) );
  AOI22_X1 U9594 ( .A1(n8640), .A2(n7919), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n7920), .ZN(n8636) );
  NOR2_X1 U9595 ( .A1(n8637), .A2(n8636), .ZN(n8635) );
  AOI21_X1 U9596 ( .B1(n7920), .B2(n7919), .A(n8635), .ZN(n7921) );
  XOR2_X1 U9597 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n7921), .Z(n7924) );
  OAI21_X1 U9598 ( .B1(n7924), .B2(n9713), .A(n9711), .ZN(n7922) );
  AOI21_X1 U9599 ( .B1(n7923), .B2(n9710), .A(n7922), .ZN(n7927) );
  AOI22_X1 U9600 ( .A1(n7925), .A2(n9710), .B1(n9708), .B2(n7924), .ZN(n7926)
         );
  MUX2_X1 U9601 ( .A(n7927), .B(n7926), .S(n8707), .Z(n7929) );
  OAI211_X1 U9602 ( .C1(n7930), .C2(n9402), .A(n7929), .B(n7928), .ZN(P2_U3264) );
  OAI222_X1 U9603 ( .A1(n7933), .A2(P2_U3152), .B1(n8478), .B2(n7932), .C1(
        n7931), .C2(n8475), .ZN(P2_U3329) );
  INV_X1 U9604 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7935) );
  OAI222_X1 U9605 ( .A1(n8475), .A2(n7935), .B1(n8478), .B2(n7934), .C1(n6283), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  INV_X1 U9606 ( .A(n8063), .ZN(n7936) );
  NOR2_X1 U9607 ( .A1(n8120), .A2(n7936), .ZN(n7937) );
  NAND2_X1 U9608 ( .A1(n8878), .A2(n8456), .ZN(n8069) );
  NAND2_X1 U9609 ( .A1(n8067), .A2(n8069), .ZN(n8797) );
  INV_X1 U9610 ( .A(n8797), .ZN(n8143) );
  AND2_X1 U9611 ( .A1(n8795), .A2(n8143), .ZN(n7939) );
  NAND2_X1 U9612 ( .A1(n8796), .A2(n7939), .ZN(n8802) );
  NAND2_X1 U9613 ( .A1(n8802), .A2(n8067), .ZN(n8780) );
  NAND2_X1 U9614 ( .A1(n8873), .A2(n8799), .ZN(n8764) );
  NAND2_X1 U9615 ( .A1(n8071), .A2(n8764), .ZN(n8779) );
  NAND2_X1 U9616 ( .A1(n8868), .A2(n8493), .ZN(n8073) );
  INV_X1 U9617 ( .A(n8766), .ZN(n7940) );
  AND2_X1 U9618 ( .A1(n7940), .A2(n8764), .ZN(n7941) );
  NAND2_X1 U9619 ( .A1(n8748), .A2(n8737), .ZN(n8078) );
  NAND2_X1 U9620 ( .A1(n8863), .A2(n8768), .ZN(n8076) );
  INV_X1 U9621 ( .A(n8749), .ZN(n7942) );
  NOR2_X1 U9622 ( .A1(n8750), .A2(n7942), .ZN(n7944) );
  INV_X1 U9623 ( .A(n8076), .ZN(n7943) );
  NAND2_X1 U9624 ( .A1(n8858), .A2(n8504), .ZN(n8081) );
  NAND2_X1 U9625 ( .A1(n8723), .A2(n8079), .ZN(n7945) );
  NAND2_X1 U9626 ( .A1(n8854), .A2(n8538), .ZN(n8082) );
  NAND2_X1 U9627 ( .A1(n7945), .A2(n8721), .ZN(n8696) );
  NAND2_X1 U9628 ( .A1(n8849), .A2(n8503), .ZN(n8089) );
  INV_X1 U9629 ( .A(n8085), .ZN(n8698) );
  NOR2_X1 U9630 ( .A1(n8697), .A2(n8698), .ZN(n7946) );
  INV_X1 U9631 ( .A(n8843), .ZN(n8684) );
  NAND2_X1 U9632 ( .A1(n8684), .A2(n8550), .ZN(n8092) );
  NAND2_X1 U9633 ( .A1(n7947), .A2(n8092), .ZN(n8667) );
  NAND2_X1 U9634 ( .A1(n8838), .A2(n8483), .ZN(n8097) );
  NAND2_X1 U9635 ( .A1(n8094), .A2(n8097), .ZN(n8668) );
  NAND2_X1 U9636 ( .A1(n8174), .A2(n7962), .ZN(n7950) );
  NAND2_X1 U9637 ( .A1(n7948), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U9638 ( .A1(n8833), .A2(n8670), .ZN(n8104) );
  INV_X1 U9639 ( .A(n7957), .ZN(n7959) );
  NAND2_X1 U9640 ( .A1(n8165), .A2(n7962), .ZN(n7952) );
  INV_X1 U9641 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8476) );
  OR2_X1 U9642 ( .A1(n7960), .A2(n8476), .ZN(n7951) );
  INV_X1 U9643 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U9644 ( .A1(n5895), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U9645 ( .A1(n5896), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7954) );
  OAI211_X1 U9646 ( .C1(n7956), .C2(n10001), .A(n7955), .B(n7954), .ZN(n8547)
         );
  INV_X1 U9647 ( .A(n8547), .ZN(n7964) );
  NOR2_X1 U9648 ( .A1(n8830), .A2(n7964), .ZN(n8106) );
  OAI22_X1 U9649 ( .A1(n7957), .A2(n8106), .B1(n7970), .B2(n8649), .ZN(n7958)
         );
  OAI21_X1 U9650 ( .B1(n7959), .B2(n8830), .A(n7958), .ZN(n7965) );
  NOR2_X1 U9651 ( .A1(n7960), .A2(n6422), .ZN(n7961) );
  INV_X1 U9652 ( .A(n8649), .ZN(n7963) );
  NAND2_X1 U9653 ( .A1(n8830), .A2(n7964), .ZN(n8107) );
  NOR2_X1 U9654 ( .A1(n8651), .A2(n8649), .ZN(n8114) );
  AOI21_X1 U9655 ( .B1(n7965), .B2(n8148), .A(n8114), .ZN(n7967) );
  NOR2_X1 U9656 ( .A1(n8114), .A2(n8106), .ZN(n8149) );
  MUX2_X1 U9657 ( .A(n8148), .B(n8149), .S(n8112), .Z(n8117) );
  INV_X1 U9658 ( .A(n8112), .ZN(n8098) );
  AND2_X1 U9659 ( .A1(n7974), .A2(n7973), .ZN(n7971) );
  MUX2_X1 U9660 ( .A(n7994), .B(n7971), .S(n8098), .Z(n7997) );
  NAND2_X1 U9661 ( .A1(n7973), .A2(n7972), .ZN(n7976) );
  NAND2_X1 U9662 ( .A1(n8001), .A2(n7974), .ZN(n7975) );
  AOI21_X1 U9663 ( .B1(n7997), .B2(n7976), .A(n7975), .ZN(n7983) );
  AND2_X1 U9664 ( .A1(n8121), .A2(n8152), .ZN(n7977) );
  OAI211_X1 U9665 ( .C1(n7978), .C2(n7977), .A(n7988), .B(n7984), .ZN(n7979)
         );
  NAND3_X1 U9666 ( .A1(n7979), .A2(n7987), .A3(n8112), .ZN(n7980) );
  NAND3_X1 U9667 ( .A1(n7997), .A2(n7981), .A3(n7980), .ZN(n7982) );
  OAI21_X1 U9668 ( .B1(n7983), .B2(n8098), .A(n7982), .ZN(n7991) );
  NAND2_X1 U9669 ( .A1(n7984), .A2(n8121), .ZN(n7985) );
  NAND3_X1 U9670 ( .A1(n7987), .A2(n7986), .A3(n7985), .ZN(n7989) );
  NAND3_X1 U9671 ( .A1(n7989), .A2(n8098), .A3(n7988), .ZN(n7990) );
  NAND3_X1 U9672 ( .A1(n7991), .A2(n7998), .A3(n7990), .ZN(n8004) );
  INV_X1 U9673 ( .A(n7992), .ZN(n7996) );
  NAND2_X1 U9674 ( .A1(n7994), .A2(n7993), .ZN(n7995) );
  OAI21_X1 U9675 ( .B1(n7997), .B2(n7996), .A(n7995), .ZN(n7999) );
  NAND2_X1 U9676 ( .A1(n7999), .A2(n7998), .ZN(n8000) );
  NAND2_X1 U9677 ( .A1(n8000), .A2(n8098), .ZN(n8003) );
  OAI21_X1 U9678 ( .B1(n8001), .B2(n8112), .A(n8128), .ZN(n8002) );
  AOI21_X1 U9679 ( .B1(n8004), .B2(n8003), .A(n8002), .ZN(n8009) );
  MUX2_X1 U9680 ( .A(n8006), .B(n8005), .S(n8112), .Z(n8007) );
  NAND2_X1 U9681 ( .A1(n9750), .A2(n8007), .ZN(n8008) );
  OR2_X1 U9682 ( .A1(n8009), .A2(n8008), .ZN(n8014) );
  MUX2_X1 U9683 ( .A(n8011), .B(n8010), .S(n8112), .Z(n8012) );
  AND2_X1 U9684 ( .A1(n8023), .A2(n8012), .ZN(n8013) );
  NAND2_X1 U9685 ( .A1(n8014), .A2(n8013), .ZN(n8025) );
  AND2_X1 U9686 ( .A1(n8016), .A2(n8015), .ZN(n8024) );
  NAND2_X1 U9687 ( .A1(n8028), .A2(n8022), .ZN(n8017) );
  AOI21_X1 U9688 ( .B1(n8025), .B2(n8024), .A(n8017), .ZN(n8021) );
  INV_X1 U9689 ( .A(n8024), .ZN(n8018) );
  NAND2_X1 U9690 ( .A1(n8018), .A2(n8022), .ZN(n8019) );
  AND2_X1 U9691 ( .A1(n8019), .A2(n9720), .ZN(n8020) );
  MUX2_X1 U9692 ( .A(n8021), .B(n8020), .S(n8112), .Z(n8027) );
  NAND4_X1 U9693 ( .A1(n8025), .A2(n8024), .A3(n8023), .A4(n8022), .ZN(n8026)
         );
  NAND2_X1 U9694 ( .A1(n8027), .A2(n8026), .ZN(n8030) );
  NAND3_X1 U9695 ( .A1(n8030), .A2(n8033), .A3(n8028), .ZN(n8029) );
  NAND2_X1 U9696 ( .A1(n8029), .A2(n8031), .ZN(n8036) );
  NAND2_X1 U9697 ( .A1(n8030), .A2(n9720), .ZN(n8034) );
  INV_X1 U9698 ( .A(n8031), .ZN(n8032) );
  AOI21_X1 U9699 ( .B1(n8034), .B2(n8033), .A(n8032), .ZN(n8035) );
  MUX2_X1 U9700 ( .A(n8036), .B(n8035), .S(n8098), .Z(n8042) );
  MUX2_X1 U9701 ( .A(n8558), .B(n8037), .S(n8098), .Z(n8039) );
  NOR2_X1 U9702 ( .A1(n8037), .A2(n8558), .ZN(n8038) );
  OR2_X1 U9703 ( .A1(n8039), .A2(n8038), .ZN(n8040) );
  MUX2_X1 U9704 ( .A(n8044), .B(n8043), .S(n8112), .Z(n8045) );
  MUX2_X1 U9705 ( .A(n8048), .B(n8047), .S(n8112), .Z(n8049) );
  MUX2_X1 U9706 ( .A(n8051), .B(n8050), .S(n8112), .Z(n8052) );
  NAND3_X1 U9707 ( .A1(n8054), .A2(n8053), .A3(n8052), .ZN(n8059) );
  AND2_X1 U9708 ( .A1(n8060), .A2(n8055), .ZN(n8056) );
  MUX2_X1 U9709 ( .A(n8057), .B(n8056), .S(n8098), .Z(n8058) );
  NAND2_X1 U9710 ( .A1(n8059), .A2(n8058), .ZN(n8064) );
  NAND4_X1 U9711 ( .A1(n8061), .A2(n8073), .A3(n8764), .A4(n8112), .ZN(n8062)
         );
  OAI211_X1 U9712 ( .C1(n8098), .C2(n8749), .A(n4839), .B(n8062), .ZN(n8077)
         );
  NAND2_X1 U9713 ( .A1(n8064), .A2(n8063), .ZN(n8065) );
  NAND2_X1 U9714 ( .A1(n8065), .A2(n8795), .ZN(n8068) );
  NAND3_X1 U9715 ( .A1(n8068), .A2(n8067), .A3(n8066), .ZN(n8070) );
  NAND3_X1 U9716 ( .A1(n8070), .A2(n8764), .A3(n8069), .ZN(n8072) );
  NAND3_X1 U9717 ( .A1(n8072), .A2(n8749), .A3(n8071), .ZN(n8074) );
  NAND2_X1 U9718 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  INV_X1 U9719 ( .A(n8079), .ZN(n8720) );
  AOI21_X1 U9720 ( .B1(n8079), .B2(n8078), .A(n8112), .ZN(n8080) );
  INV_X1 U9721 ( .A(n8721), .ZN(n8712) );
  INV_X1 U9722 ( .A(n8082), .ZN(n8083) );
  OAI21_X1 U9723 ( .B1(n8697), .B2(n8083), .A(n8112), .ZN(n8084) );
  AOI21_X1 U9724 ( .B1(n8087), .B2(n8085), .A(n8112), .ZN(n8086) );
  AOI21_X1 U9725 ( .B1(n8088), .B2(n8087), .A(n8086), .ZN(n8096) );
  OAI21_X1 U9726 ( .B1(n8089), .B2(n8112), .A(n8685), .ZN(n8095) );
  INV_X1 U9727 ( .A(n8550), .ZN(n8671) );
  NAND2_X1 U9728 ( .A1(n8843), .A2(n8671), .ZN(n8090) );
  AND2_X1 U9729 ( .A1(n8097), .A2(n8090), .ZN(n8091) );
  MUX2_X1 U9730 ( .A(n8092), .B(n8091), .S(n8112), .Z(n8093) );
  OAI211_X1 U9731 ( .C1(n8096), .C2(n8095), .A(n8094), .B(n8093), .ZN(n8102)
         );
  OAI21_X1 U9732 ( .B1(n8098), .B2(n8838), .A(n8097), .ZN(n8100) );
  NAND2_X1 U9733 ( .A1(n8483), .A2(n8112), .ZN(n8099) );
  NAND2_X1 U9734 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  AOI21_X1 U9735 ( .B1(n8102), .B2(n8101), .A(n8463), .ZN(n8110) );
  MUX2_X1 U9736 ( .A(n8104), .B(n8103), .S(n8112), .Z(n8105) );
  INV_X1 U9737 ( .A(n8105), .ZN(n8109) );
  INV_X1 U9738 ( .A(n8106), .ZN(n8108) );
  OAI211_X1 U9739 ( .C1(n8110), .C2(n8109), .A(n8108), .B(n8107), .ZN(n8116)
         );
  INV_X1 U9740 ( .A(n8111), .ZN(n8113) );
  MUX2_X1 U9741 ( .A(n8114), .B(n8113), .S(n8112), .Z(n8115) );
  AOI21_X1 U9742 ( .B1(n8117), .B2(n8116), .A(n8115), .ZN(n8118) );
  INV_X1 U9743 ( .A(n6550), .ZN(n8119) );
  NOR3_X1 U9744 ( .A1(n8155), .A2(n8119), .A3(n6265), .ZN(n8156) );
  INV_X1 U9745 ( .A(n8697), .ZN(n8693) );
  INV_X1 U9746 ( .A(n8120), .ZN(n8142) );
  NAND4_X1 U9747 ( .A1(n8123), .A2(n8122), .A3(n8151), .A4(n8121), .ZN(n8127)
         );
  NOR4_X1 U9748 ( .A1(n8127), .A2(n8126), .A3(n8125), .A4(n8124), .ZN(n8129)
         );
  NAND4_X1 U9749 ( .A1(n8129), .A2(n9750), .A3(n8128), .A4(n8820), .ZN(n8133)
         );
  NOR4_X1 U9750 ( .A1(n8133), .A2(n8132), .A3(n8131), .A4(n8130), .ZN(n8134)
         );
  NAND4_X1 U9751 ( .A1(n8135), .A2(n9722), .A3(n8134), .A4(n4853), .ZN(n8136)
         );
  NOR4_X1 U9752 ( .A1(n8139), .A2(n8138), .A3(n8137), .A4(n8136), .ZN(n8140)
         );
  NAND4_X1 U9753 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n8144)
         );
  NOR4_X1 U9754 ( .A1(n8750), .A2(n8766), .A3(n8779), .A4(n8144), .ZN(n8145)
         );
  NAND4_X1 U9755 ( .A1(n8693), .A2(n8721), .A3(n8736), .A4(n8145), .ZN(n8146)
         );
  NOR4_X1 U9756 ( .A1(n8463), .A2(n8668), .A3(n8678), .A4(n8146), .ZN(n8147)
         );
  NAND3_X1 U9757 ( .A1(n8149), .A2(n8148), .A3(n8147), .ZN(n8150) );
  XNOR2_X1 U9758 ( .A(n8150), .B(n8707), .ZN(n8153) );
  OAI22_X1 U9759 ( .A1(n8153), .A2(n8152), .B1(n8151), .B2(n6550), .ZN(n8154)
         );
  OAI21_X1 U9760 ( .B1(n8161), .B2(n8159), .A(P2_B_REG_SCAN_IN), .ZN(n8160) );
  NAND2_X1 U9761 ( .A1(n8162), .A2(n5306), .ZN(n8164) );
  NAND2_X1 U9762 ( .A1(n5732), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8163) );
  INV_X1 U9763 ( .A(n9069), .ZN(n8233) );
  NAND2_X1 U9764 ( .A1(n9287), .A2(n8233), .ZN(n8423) );
  NAND2_X1 U9765 ( .A1(n8165), .A2(n5306), .ZN(n8167) );
  NAND2_X1 U9766 ( .A1(n5732), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8166) );
  INV_X1 U9767 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8171) );
  NAND2_X1 U9768 ( .A1(n5017), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U9769 ( .A1(n8168), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8169) );
  OAI211_X1 U9770 ( .C1(n8172), .C2(n8171), .A(n8170), .B(n8169), .ZN(n9111)
         );
  INV_X1 U9771 ( .A(n9111), .ZN(n8226) );
  NAND2_X1 U9772 ( .A1(n8174), .A2(n5306), .ZN(n8176) );
  NAND2_X1 U9773 ( .A1(n5732), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U9774 ( .A1(n8418), .A2(n9107), .ZN(n8292) );
  NAND2_X1 U9775 ( .A1(n9334), .A2(n9233), .ZN(n9101) );
  NAND2_X1 U9776 ( .A1(n9341), .A2(n9246), .ZN(n9098) );
  AND2_X1 U9777 ( .A1(n9101), .A2(n9098), .ZN(n8386) );
  INV_X1 U9778 ( .A(n8386), .ZN(n8178) );
  AND2_X1 U9779 ( .A1(n9346), .A2(n9234), .ZN(n9097) );
  AND2_X1 U9780 ( .A1(n8398), .A2(n9097), .ZN(n8177) );
  OR2_X1 U9781 ( .A1(n8178), .A2(n8177), .ZN(n8397) );
  INV_X1 U9782 ( .A(n8397), .ZN(n8181) );
  AND2_X1 U9783 ( .A1(n9093), .A2(n8186), .ZN(n8380) );
  INV_X1 U9784 ( .A(n8380), .ZN(n8179) );
  OR2_X1 U9785 ( .A1(n9346), .A2(n9234), .ZN(n9096) );
  AND2_X1 U9786 ( .A1(n9096), .A2(n8376), .ZN(n8382) );
  OAI211_X1 U9787 ( .C1(n8372), .C2(n8179), .A(n8398), .B(n8382), .ZN(n8180)
         );
  AOI21_X1 U9788 ( .B1(n8181), .B2(n8180), .A(n9100), .ZN(n8183) );
  INV_X1 U9789 ( .A(n9219), .ZN(n9086) );
  NAND2_X1 U9790 ( .A1(n9331), .A2(n9086), .ZN(n8400) );
  INV_X1 U9791 ( .A(n8400), .ZN(n8182) );
  NAND2_X1 U9792 ( .A1(n9208), .A2(n9219), .ZN(n8402) );
  NAND2_X1 U9793 ( .A1(n8395), .A2(n8402), .ZN(n9102) );
  INV_X1 U9794 ( .A(n9102), .ZN(n8389) );
  OAI21_X1 U9795 ( .B1(n8183), .B2(n8182), .A(n8389), .ZN(n8287) );
  NAND2_X1 U9796 ( .A1(n8400), .A2(n9093), .ZN(n8184) );
  OR2_X1 U9797 ( .A1(n8184), .A2(n8397), .ZN(n8285) );
  AND2_X1 U9798 ( .A1(n8186), .A2(n8185), .ZN(n8373) );
  INV_X1 U9799 ( .A(n8373), .ZN(n8220) );
  AND2_X1 U9800 ( .A1(n8217), .A2(n8214), .ZN(n8361) );
  INV_X1 U9801 ( .A(n8361), .ZN(n8189) );
  NAND2_X1 U9802 ( .A1(n8352), .A2(n8210), .ZN(n8355) );
  INV_X1 U9803 ( .A(n8342), .ZN(n8205) );
  OR3_X1 U9804 ( .A1(n8205), .A2(n4667), .A3(n8326), .ZN(n8209) );
  INV_X1 U9805 ( .A(n8329), .ZN(n8187) );
  OR4_X1 U9806 ( .A1(n8355), .A2(n8209), .A3(n8187), .A4(n8310), .ZN(n8188) );
  OR3_X1 U9807 ( .A1(n8220), .A2(n8189), .A3(n8188), .ZN(n8282) );
  INV_X1 U9808 ( .A(n8190), .ZN(n8192) );
  NAND2_X1 U9809 ( .A1(n9027), .A2(n9640), .ZN(n8191) );
  NAND3_X1 U9810 ( .A1(n8192), .A2(n5766), .A3(n8191), .ZN(n8194) );
  NAND2_X1 U9811 ( .A1(n8194), .A2(n8193), .ZN(n8196) );
  OAI21_X1 U9812 ( .B1(n8197), .B2(n8196), .A(n8195), .ZN(n8198) );
  NAND2_X1 U9813 ( .A1(n8198), .A2(n8270), .ZN(n8200) );
  AND2_X1 U9814 ( .A1(n8307), .A2(n8199), .ZN(n8275) );
  NAND2_X1 U9815 ( .A1(n8200), .A2(n8275), .ZN(n8202) );
  NAND3_X1 U9816 ( .A1(n8202), .A2(n8201), .A3(n8313), .ZN(n8204) );
  AND2_X1 U9817 ( .A1(n8320), .A2(n8203), .ZN(n8311) );
  AND3_X1 U9818 ( .A1(n8204), .A2(n8311), .A3(n8318), .ZN(n8221) );
  OR2_X1 U9819 ( .A1(n8206), .A2(n8205), .ZN(n8207) );
  AND2_X1 U9820 ( .A1(n8207), .A2(n8351), .ZN(n8340) );
  INV_X1 U9821 ( .A(n8340), .ZN(n8212) );
  NAND2_X1 U9822 ( .A1(n8334), .A2(n8208), .ZN(n8336) );
  NOR2_X1 U9823 ( .A1(n8209), .A2(n4669), .ZN(n8211) );
  OAI21_X1 U9824 ( .B1(n8212), .B2(n8211), .A(n8210), .ZN(n8213) );
  NAND2_X1 U9825 ( .A1(n8213), .A2(n8354), .ZN(n8215) );
  NAND3_X1 U9826 ( .A1(n8215), .A2(n8214), .A3(n8352), .ZN(n8216) );
  NAND2_X1 U9827 ( .A1(n8362), .A2(n8216), .ZN(n8218) );
  NAND2_X1 U9828 ( .A1(n8218), .A2(n8217), .ZN(n8219) );
  OR2_X1 U9829 ( .A1(n8220), .A2(n8219), .ZN(n8280) );
  OAI21_X1 U9830 ( .B1(n8282), .B2(n8221), .A(n8280), .ZN(n8222) );
  INV_X1 U9831 ( .A(n8222), .ZN(n8223) );
  NOR2_X1 U9832 ( .A1(n8285), .A2(n8223), .ZN(n8224) );
  NAND2_X1 U9833 ( .A1(n9317), .A2(n9006), .ZN(n8299) );
  NAND2_X1 U9834 ( .A1(n8299), .A2(n9168), .ZN(n9103) );
  INV_X1 U9835 ( .A(n9103), .ZN(n8391) );
  OAI21_X1 U9836 ( .B1(n8287), .B2(n8224), .A(n8391), .ZN(n8225) );
  NAND3_X1 U9837 ( .A1(n9145), .A2(n4408), .A3(n8225), .ZN(n8231) );
  NAND2_X1 U9838 ( .A1(n9073), .A2(n8226), .ZN(n8265) );
  NAND2_X1 U9839 ( .A1(n9303), .A2(n9092), .ZN(n9108) );
  NAND2_X1 U9840 ( .A1(n9312), .A2(n9089), .ZN(n9104) );
  NAND2_X1 U9841 ( .A1(n8411), .A2(n9104), .ZN(n8227) );
  NAND2_X1 U9842 ( .A1(n8227), .A2(n9105), .ZN(n8228) );
  AND2_X1 U9843 ( .A1(n9108), .A2(n8228), .ZN(n8229) );
  OR2_X1 U9844 ( .A1(n8292), .A2(n8229), .ZN(n8230) );
  NAND2_X1 U9845 ( .A1(n9299), .A2(n9129), .ZN(n8415) );
  AND2_X1 U9846 ( .A1(n8230), .A2(n8415), .ZN(n8290) );
  OAI211_X1 U9847 ( .C1(n8292), .C2(n8231), .A(n8265), .B(n8290), .ZN(n8232)
         );
  NAND2_X1 U9848 ( .A1(n4392), .A2(n8232), .ZN(n8234) );
  NAND2_X1 U9849 ( .A1(n8234), .A2(n8440), .ZN(n8235) );
  XNOR2_X1 U9850 ( .A(n8235), .B(n9275), .ZN(n8437) );
  INV_X1 U9851 ( .A(n9101), .ZN(n8237) );
  NOR2_X1 U9852 ( .A1(n9100), .A2(n8237), .ZN(n9217) );
  INV_X1 U9853 ( .A(n9097), .ZN(n8378) );
  NAND4_X1 U9854 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n4643), .ZN(n8243)
         );
  NOR3_X1 U9855 ( .A1(n8243), .A2(n6941), .A3(n7077), .ZN(n8244) );
  NAND4_X1 U9856 ( .A1(n8245), .A2(n4908), .A3(n4933), .A4(n8244), .ZN(n8247)
         );
  NOR2_X1 U9857 ( .A1(n8247), .A2(n8246), .ZN(n8249) );
  NAND4_X1 U9858 ( .A1(n8251), .A2(n8250), .A3(n8249), .A4(n8248), .ZN(n8252)
         );
  OR3_X1 U9859 ( .A1(n4647), .A2(n8253), .A3(n8252), .ZN(n8254) );
  NOR2_X1 U9860 ( .A1(n8255), .A2(n8254), .ZN(n8256) );
  NAND4_X1 U9861 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n8260)
         );
  NOR2_X1 U9862 ( .A1(n9094), .A2(n8260), .ZN(n8261) );
  NAND4_X1 U9863 ( .A1(n9217), .A2(n4691), .A3(n9244), .A4(n8261), .ZN(n8262)
         );
  XNOR2_X1 U9864 ( .A(n9331), .B(n9086), .ZN(n9199) );
  NOR3_X1 U9865 ( .A1(n9187), .A2(n8262), .A3(n9199), .ZN(n8263) );
  NAND4_X1 U9866 ( .A1(n9145), .A2(n9155), .A3(n9172), .A4(n8263), .ZN(n8264)
         );
  NOR2_X1 U9867 ( .A1(n9123), .A2(n8264), .ZN(n8266) );
  INV_X1 U9868 ( .A(n8432), .ZN(n8296) );
  NAND2_X1 U9869 ( .A1(n8268), .A2(n9069), .ZN(n8269) );
  NAND2_X1 U9870 ( .A1(n8313), .A2(n8270), .ZN(n8271) );
  NAND2_X1 U9871 ( .A1(n8271), .A2(n8307), .ZN(n8272) );
  NAND2_X1 U9872 ( .A1(n8272), .A2(n8316), .ZN(n8274) );
  INV_X1 U9873 ( .A(n7066), .ZN(n8273) );
  AOI21_X1 U9874 ( .B1(n8318), .B2(n8274), .A(n8273), .ZN(n8279) );
  INV_X1 U9875 ( .A(n8311), .ZN(n8278) );
  NAND4_X1 U9876 ( .A1(n8276), .A2(n8311), .A3(n8275), .A4(n8318), .ZN(n8277)
         );
  OAI21_X1 U9877 ( .B1(n8279), .B2(n8278), .A(n8277), .ZN(n8281) );
  OAI21_X1 U9878 ( .B1(n8282), .B2(n8281), .A(n8280), .ZN(n8283) );
  INV_X1 U9879 ( .A(n8283), .ZN(n8284) );
  NOR2_X1 U9880 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  OAI21_X1 U9881 ( .B1(n8287), .B2(n8286), .A(n8391), .ZN(n8288) );
  NAND3_X1 U9882 ( .A1(n4408), .A2(n9105), .A3(n8288), .ZN(n8291) );
  NAND2_X1 U9883 ( .A1(n9111), .A2(n9069), .ZN(n8289) );
  NAND2_X1 U9884 ( .A1(n9073), .A2(n8289), .ZN(n8429) );
  OAI211_X1 U9885 ( .C1(n8292), .C2(n8291), .A(n8429), .B(n8290), .ZN(n8293)
         );
  NAND2_X1 U9886 ( .A1(n8422), .A2(n8293), .ZN(n8294) );
  NAND3_X1 U9887 ( .A1(n8294), .A2(n5766), .A3(n8440), .ZN(n8295) );
  NAND2_X1 U9888 ( .A1(n8296), .A2(n8295), .ZN(n8435) );
  INV_X1 U9889 ( .A(n9108), .ZN(n8298) );
  NAND2_X1 U9890 ( .A1(n8422), .A2(n9107), .ZN(n8297) );
  MUX2_X1 U9891 ( .A(n8298), .B(n8297), .S(n8424), .Z(n8421) );
  MUX2_X1 U9892 ( .A(n9089), .B(n9160), .S(n8424), .Z(n8302) );
  OAI21_X1 U9893 ( .B1(n8302), .B2(n9312), .A(n9153), .ZN(n8301) );
  OAI21_X1 U9894 ( .B1(n8302), .B2(n9174), .A(n8299), .ZN(n8300) );
  MUX2_X1 U9895 ( .A(n8301), .B(n8300), .S(n8424), .Z(n8303) );
  NAND2_X1 U9896 ( .A1(n8302), .A2(n9090), .ZN(n8407) );
  NAND2_X1 U9897 ( .A1(n8303), .A2(n8407), .ZN(n8410) );
  INV_X1 U9898 ( .A(n8395), .ZN(n8392) );
  NAND2_X1 U9899 ( .A1(n8304), .A2(n8307), .ZN(n8305) );
  NAND3_X1 U9900 ( .A1(n8314), .A2(n8308), .A3(n8307), .ZN(n8309) );
  NAND3_X1 U9901 ( .A1(n8309), .A2(n4908), .A3(n7066), .ZN(n8312) );
  AOI21_X1 U9902 ( .B1(n8312), .B2(n8311), .A(n8310), .ZN(n8325) );
  NAND3_X1 U9903 ( .A1(n8314), .A2(n8313), .A3(n7066), .ZN(n8315) );
  NAND2_X1 U9904 ( .A1(n8315), .A2(n4908), .ZN(n8317) );
  NAND2_X1 U9905 ( .A1(n8317), .A2(n8316), .ZN(n8319) );
  NAND2_X1 U9906 ( .A1(n8319), .A2(n8318), .ZN(n8323) );
  INV_X1 U9907 ( .A(n8320), .ZN(n8321) );
  AOI21_X1 U9908 ( .B1(n8323), .B2(n8322), .A(n8321), .ZN(n8324) );
  AOI21_X1 U9909 ( .B1(n8328), .B2(n8329), .A(n8336), .ZN(n8327) );
  OAI21_X1 U9910 ( .B1(n8327), .B2(n8326), .A(n8343), .ZN(n8339) );
  INV_X1 U9911 ( .A(n8328), .ZN(n8337) );
  NAND2_X1 U9912 ( .A1(n8330), .A2(n8329), .ZN(n8333) );
  INV_X1 U9913 ( .A(n8331), .ZN(n8332) );
  AOI21_X1 U9914 ( .B1(n8334), .B2(n8333), .A(n8332), .ZN(n8335) );
  OAI211_X1 U9915 ( .C1(n8337), .C2(n8336), .A(n8335), .B(n8342), .ZN(n8338)
         );
  AND2_X1 U9916 ( .A1(n8340), .A2(n8354), .ZN(n8347) );
  NAND2_X1 U9917 ( .A1(n8342), .A2(n8341), .ZN(n8344) );
  AND2_X1 U9918 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  NOR2_X1 U9919 ( .A1(n8355), .A2(n8345), .ZN(n8346) );
  INV_X1 U9920 ( .A(n8424), .ZN(n8393) );
  MUX2_X1 U9921 ( .A(n8347), .B(n8346), .S(n8393), .Z(n8348) );
  NAND2_X1 U9922 ( .A1(n8354), .A2(n8351), .ZN(n8353) );
  NAND2_X1 U9923 ( .A1(n8353), .A2(n8352), .ZN(n8357) );
  NAND2_X1 U9924 ( .A1(n8355), .A2(n8354), .ZN(n8356) );
  MUX2_X1 U9925 ( .A(n8357), .B(n8356), .S(n8424), .Z(n8358) );
  NAND3_X1 U9926 ( .A1(n8360), .A2(n8359), .A3(n8358), .ZN(n8364) );
  MUX2_X1 U9927 ( .A(n8362), .B(n8361), .S(n8393), .Z(n8363) );
  NAND2_X1 U9928 ( .A1(n8364), .A2(n8363), .ZN(n8371) );
  INV_X1 U9929 ( .A(n8365), .ZN(n8367) );
  MUX2_X1 U9930 ( .A(n8367), .B(n8366), .S(n8424), .Z(n8369) );
  NOR2_X1 U9931 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  NAND2_X1 U9932 ( .A1(n8371), .A2(n8370), .ZN(n8375) );
  MUX2_X1 U9933 ( .A(n8373), .B(n8372), .S(n8424), .Z(n8374) );
  NAND2_X1 U9934 ( .A1(n8375), .A2(n8374), .ZN(n8381) );
  NAND3_X1 U9935 ( .A1(n8381), .A2(n8377), .A3(n8376), .ZN(n8379) );
  NAND3_X1 U9936 ( .A1(n8379), .A2(n9093), .A3(n8378), .ZN(n8385) );
  NAND2_X1 U9937 ( .A1(n8381), .A2(n8380), .ZN(n8383) );
  NAND2_X1 U9938 ( .A1(n8383), .A2(n8382), .ZN(n8384) );
  MUX2_X1 U9939 ( .A(n8385), .B(n8384), .S(n8424), .Z(n8396) );
  INV_X1 U9940 ( .A(n9100), .ZN(n8387) );
  NAND3_X1 U9941 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(n8390) );
  MUX2_X1 U9942 ( .A(n8395), .B(n8394), .S(n8393), .Z(n8408) );
  INV_X1 U9943 ( .A(n8396), .ZN(n8399) );
  AOI21_X1 U9944 ( .B1(n8399), .B2(n8398), .A(n8397), .ZN(n8401) );
  OAI211_X1 U9945 ( .C1(n8401), .C2(n9100), .A(n8400), .B(n9168), .ZN(n8404)
         );
  INV_X1 U9946 ( .A(n8402), .ZN(n9182) );
  NAND2_X1 U9947 ( .A1(n9168), .A2(n9182), .ZN(n8403) );
  NAND3_X1 U9948 ( .A1(n8404), .A2(n9153), .A3(n8403), .ZN(n8405) );
  NAND2_X1 U9949 ( .A1(n8405), .A2(n8424), .ZN(n8406) );
  NAND3_X1 U9950 ( .A1(n8408), .A2(n8407), .A3(n8406), .ZN(n8409) );
  MUX2_X1 U9951 ( .A(n8411), .B(n9105), .S(n8424), .Z(n8412) );
  INV_X1 U9952 ( .A(n9123), .ZN(n9125) );
  NAND2_X1 U9953 ( .A1(n8413), .A2(n9125), .ZN(n8414) );
  NAND2_X1 U9954 ( .A1(n8414), .A2(n9109), .ZN(n8420) );
  INV_X1 U9955 ( .A(n8415), .ZN(n8416) );
  NAND2_X1 U9956 ( .A1(n8422), .A2(n8416), .ZN(n8417) );
  OAI21_X1 U9957 ( .B1(n8421), .B2(n8420), .A(n8419), .ZN(n8430) );
  AND2_X1 U9958 ( .A1(n8424), .A2(n8423), .ZN(n8426) );
  AOI21_X2 U9959 ( .B1(n8430), .B2(n8429), .A(n8428), .ZN(n8438) );
  AND2_X1 U9960 ( .A1(n8440), .A2(n8431), .ZN(n8433) );
  AOI21_X1 U9961 ( .B1(n8438), .B2(n8433), .A(n8432), .ZN(n8434) );
  INV_X1 U9962 ( .A(n8438), .ZN(n8443) );
  INV_X1 U9963 ( .A(n8439), .ZN(n8442) );
  OAI21_X1 U9964 ( .B1(n8445), .B2(n8444), .A(P1_B_REG_SCAN_IN), .ZN(n8446) );
  AOI21_X1 U9965 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(n8449) );
  OAI222_X1 U9966 ( .A1(n8475), .A2(n8451), .B1(n8478), .B2(n8450), .C1(
        P2_U3152), .C2(n6552), .ZN(P2_U3336) );
  INV_X1 U9967 ( .A(n8858), .ZN(n8734) );
  INV_X1 U9968 ( .A(n8799), .ZN(n8551) );
  OR2_X1 U9969 ( .A1(n8884), .A2(n8552), .ZN(n8452) );
  INV_X1 U9970 ( .A(n8456), .ZN(n8784) );
  AOI22_X2 U9971 ( .A1(n8789), .A2(n8797), .B1(n8878), .B2(n8784), .ZN(n8775)
         );
  NAND2_X1 U9972 ( .A1(n8863), .A2(n8737), .ZN(n8457) );
  OAI22_X1 U9973 ( .A1(n8713), .A2(n8721), .B1(n8738), .B2(n8854), .ZN(n8694)
         );
  AOI22_X1 U9974 ( .A1(n8694), .A2(n8697), .B1(n8695), .B2(n8503), .ZN(n8679)
         );
  AOI22_X1 U9975 ( .A1(n8662), .A2(n8668), .B1(n8666), .B2(n8483), .ZN(n8458)
         );
  XNOR2_X1 U9976 ( .A(n8458), .B(n8463), .ZN(n8837) );
  INV_X1 U9977 ( .A(n8854), .ZN(n8719) );
  NOR2_X2 U9978 ( .A1(n8838), .A2(n8680), .ZN(n8663) );
  INV_X1 U9979 ( .A(n8663), .ZN(n8459) );
  INV_X1 U9980 ( .A(n8833), .ZN(n8462) );
  AOI21_X1 U9981 ( .B1(n8833), .B2(n8459), .A(n8647), .ZN(n8834) );
  AOI22_X1 U9982 ( .A1(n9749), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8460), .B2(
        n9771), .ZN(n8461) );
  OAI21_X1 U9983 ( .B1(n8462), .B2(n9775), .A(n8461), .ZN(n8473) );
  XNOR2_X1 U9984 ( .A(n8464), .B(n8463), .ZN(n8465) );
  INV_X1 U9985 ( .A(n8465), .ZN(n8470) );
  INV_X1 U9986 ( .A(P2_B_REG_SCAN_IN), .ZN(n8466) );
  NOR2_X1 U9987 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  NOR2_X1 U9988 ( .A1(n9761), .A2(n8468), .ZN(n8648) );
  INV_X1 U9989 ( .A(n8648), .ZN(n8469) );
  INV_X1 U9990 ( .A(n8471), .ZN(n8836) );
  NOR2_X1 U9991 ( .A1(n8836), .A2(n8740), .ZN(n8472) );
  OAI21_X1 U9992 ( .B1(n8837), .B2(n8808), .A(n8474), .ZN(P2_U3267) );
  OAI222_X1 U9993 ( .A1(P2_U3152), .A2(n8479), .B1(n8478), .B2(n8477), .C1(
        n8476), .C2(n8475), .ZN(P2_U3328) );
  OAI211_X1 U9994 ( .C1(n8482), .C2(n8481), .A(n8480), .B(n8535), .ZN(n8487)
         );
  AOI22_X1 U9995 ( .A1(n8543), .A2(n8682), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8486) );
  INV_X1 U9996 ( .A(n8483), .ZN(n8687) );
  INV_X1 U9997 ( .A(n8503), .ZN(n8688) );
  AOI22_X1 U9998 ( .A1(n8528), .A2(n8687), .B1(n8527), .B2(n8688), .ZN(n8485)
         );
  NAND2_X1 U9999 ( .A1(n8843), .A2(n8520), .ZN(n8484) );
  NAND4_X1 U10000 ( .A1(n8487), .A2(n8486), .A3(n8485), .A4(n8484), .ZN(
        P2_U3216) );
  INV_X1 U10001 ( .A(n8489), .ZN(n8490) );
  NOR2_X1 U10002 ( .A1(n8488), .A2(n8490), .ZN(n8492) );
  XNOR2_X1 U10003 ( .A(n8492), .B(n8491), .ZN(n8498) );
  INV_X1 U10004 ( .A(n8754), .ZN(n8495) );
  OAI22_X1 U10005 ( .A1(n8504), .A2(n9761), .B1(n8493), .B2(n9763), .ZN(n8752)
         );
  AOI22_X1 U10006 ( .A1(n8505), .A2(n8752), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8494) );
  OAI21_X1 U10007 ( .B1(n8495), .B2(n8515), .A(n8494), .ZN(n8496) );
  AOI21_X1 U10008 ( .B1(n8863), .B2(n8520), .A(n8496), .ZN(n8497) );
  OAI21_X1 U10009 ( .B1(n8498), .B2(n8522), .A(n8497), .ZN(P2_U3218) );
  XNOR2_X1 U10010 ( .A(n8501), .B(n8500), .ZN(n8502) );
  XNOR2_X1 U10011 ( .A(n8499), .B(n8502), .ZN(n8510) );
  INV_X1 U10012 ( .A(n8717), .ZN(n8507) );
  OAI22_X1 U10013 ( .A1(n8504), .A2(n9763), .B1(n8503), .B2(n9761), .ZN(n8725)
         );
  AOI22_X1 U10014 ( .A1(n8505), .A2(n8725), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8506) );
  OAI21_X1 U10015 ( .B1(n8507), .B2(n8515), .A(n8506), .ZN(n8508) );
  AOI21_X1 U10016 ( .B1(n8854), .B2(n8520), .A(n8508), .ZN(n8509) );
  OAI21_X1 U10017 ( .B1(n8510), .B2(n8522), .A(n8509), .ZN(P2_U3227) );
  XNOR2_X1 U10018 ( .A(n8511), .B(n8512), .ZN(n8523) );
  INV_X1 U10019 ( .A(n8732), .ZN(n8514) );
  OAI22_X1 U10020 ( .A1(n8515), .A2(n8514), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8513), .ZN(n8519) );
  OAI22_X1 U10021 ( .A1(n8768), .A2(n8517), .B1(n8516), .B2(n8538), .ZN(n8518)
         );
  AOI211_X1 U10022 ( .C1(n8858), .C2(n8520), .A(n8519), .B(n8518), .ZN(n8521)
         );
  OAI21_X1 U10023 ( .B1(n8523), .B2(n8522), .A(n8521), .ZN(P2_U3231) );
  OAI21_X1 U10024 ( .B1(n8526), .B2(n8525), .A(n8524), .ZN(n8532) );
  AOI22_X1 U10025 ( .A1(n8543), .A2(n8761), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8530) );
  AOI22_X1 U10026 ( .A1(n8528), .A2(n8737), .B1(n8527), .B2(n8551), .ZN(n8529)
         );
  OAI211_X1 U10027 ( .C1(n8763), .C2(n8546), .A(n8530), .B(n8529), .ZN(n8531)
         );
  AOI21_X1 U10028 ( .B1(n8532), .B2(n8535), .A(n8531), .ZN(n8533) );
  INV_X1 U10029 ( .A(n8533), .ZN(P2_U3237) );
  OAI211_X1 U10030 ( .C1(n8534), .C2(n8537), .A(n8536), .B(n8535), .ZN(n8545)
         );
  OAI22_X1 U10031 ( .A1(n8671), .A2(n9761), .B1(n8538), .B2(n9763), .ZN(n8701)
         );
  INV_X1 U10032 ( .A(n8701), .ZN(n8540) );
  OAI22_X1 U10033 ( .A1(n8541), .A2(n8540), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8539), .ZN(n8542) );
  AOI21_X1 U10034 ( .B1(n8706), .B2(n8543), .A(n8542), .ZN(n8544) );
  OAI211_X1 U10035 ( .C1(n8695), .C2(n8546), .A(n8545), .B(n8544), .ZN(
        P2_U3242) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8547), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8548), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10038 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8687), .S(n8567), .Z(
        P2_U3580) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8550), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8688), .S(n8567), .Z(
        P2_U3578) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8738), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8737), .S(n8567), .Z(
        P2_U3575) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8782), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10044 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8551), .S(n8567), .Z(
        P2_U3573) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8784), .S(n8567), .Z(
        P2_U3572) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8552), .S(n8567), .Z(
        P2_U3571) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8553), .S(n8567), .Z(
        P2_U3570) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8554), .S(n8567), .Z(
        P2_U3569) );
  MUX2_X1 U10049 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8555), .S(n8567), .Z(
        P2_U3568) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8556), .S(n8567), .Z(
        P2_U3567) );
  MUX2_X1 U10051 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8557), .S(n8567), .Z(
        P2_U3566) );
  MUX2_X1 U10052 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8558), .S(n8567), .Z(
        P2_U3565) );
  MUX2_X1 U10053 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8559), .S(n8567), .Z(
        P2_U3564) );
  MUX2_X1 U10054 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8560), .S(n8567), .Z(
        P2_U3563) );
  MUX2_X1 U10055 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8561), .S(n8567), .Z(
        P2_U3562) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8562), .S(n8567), .Z(
        P2_U3561) );
  MUX2_X1 U10057 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8563), .S(n8567), .Z(
        P2_U3560) );
  MUX2_X1 U10058 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8564), .S(n8567), .Z(
        P2_U3559) );
  MUX2_X1 U10059 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8565), .S(n8567), .Z(
        P2_U3558) );
  MUX2_X1 U10060 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8566), .S(n8567), .Z(
        P2_U3557) );
  MUX2_X1 U10061 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8568), .S(n8567), .Z(
        P2_U3556) );
  MUX2_X1 U10062 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8569), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10063 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8570), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10064 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6557), .S(P2_U3966), .Z(
        P2_U3553) );
  NAND2_X1 U10065 ( .A1(n9420), .A2(n8571), .ZN(n8582) );
  OAI211_X1 U10066 ( .C1(n8574), .C2(n8573), .A(n9710), .B(n8572), .ZN(n8581)
         );
  AOI21_X1 U10067 ( .B1(n9715), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8575), .ZN(
        n8580) );
  OAI211_X1 U10068 ( .C1(n8578), .C2(n8577), .A(n9708), .B(n8576), .ZN(n8579)
         );
  NAND4_X1 U10069 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(
        P2_U3251) );
  AOI211_X1 U10070 ( .C1(n8585), .C2(n8584), .A(n8583), .B(n9414), .ZN(n8586)
         );
  AOI21_X1 U10071 ( .B1(n9420), .B2(n8587), .A(n8586), .ZN(n8595) );
  INV_X1 U10072 ( .A(n8588), .ZN(n8589) );
  AOI21_X1 U10073 ( .B1(n9715), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8589), .ZN(
        n8594) );
  OAI211_X1 U10074 ( .C1(n8592), .C2(n8591), .A(n9708), .B(n8590), .ZN(n8593)
         );
  NAND3_X1 U10075 ( .A1(n8595), .A2(n8594), .A3(n8593), .ZN(P2_U3253) );
  NAND2_X1 U10076 ( .A1(n9420), .A2(n8596), .ZN(n8608) );
  OAI21_X1 U10077 ( .B1(n8599), .B2(n8598), .A(n8597), .ZN(n8600) );
  NAND2_X1 U10078 ( .A1(n8600), .A2(n9710), .ZN(n8607) );
  AOI21_X1 U10079 ( .B1(n9715), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8601), .ZN(
        n8606) );
  OAI211_X1 U10080 ( .C1(n8604), .C2(n8603), .A(n9708), .B(n8602), .ZN(n8605)
         );
  NAND4_X1 U10081 ( .A1(n8608), .A2(n8607), .A3(n8606), .A4(n8605), .ZN(
        P2_U3256) );
  AOI21_X1 U10082 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8622) );
  AOI211_X1 U10083 ( .C1(n8614), .C2(n8613), .A(n9414), .B(n8612), .ZN(n8615)
         );
  INV_X1 U10084 ( .A(n8615), .ZN(n8621) );
  INV_X1 U10085 ( .A(n8616), .ZN(n8619) );
  NOR2_X1 U10086 ( .A1(n9711), .A2(n8617), .ZN(n8618) );
  AOI211_X1 U10087 ( .C1(n9715), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8619), .B(
        n8618), .ZN(n8620) );
  OAI211_X1 U10088 ( .C1(n8622), .C2(n9713), .A(n8621), .B(n8620), .ZN(
        P2_U3261) );
  XNOR2_X1 U10089 ( .A(n8624), .B(n8623), .ZN(n8633) );
  NOR2_X1 U10090 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10004), .ZN(n8625) );
  AOI21_X1 U10091 ( .B1(n9715), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8625), .ZN(
        n8626) );
  OAI21_X1 U10092 ( .B1(n9711), .B2(n8627), .A(n8626), .ZN(n8632) );
  AOI211_X1 U10093 ( .C1(n8630), .C2(n8629), .A(n9414), .B(n8628), .ZN(n8631)
         );
  AOI211_X1 U10094 ( .C1(n8633), .C2(n9708), .A(n8632), .B(n8631), .ZN(n8634)
         );
  INV_X1 U10095 ( .A(n8634), .ZN(P2_U3262) );
  AOI21_X1 U10096 ( .B1(n8637), .B2(n8636), .A(n8635), .ZN(n8646) );
  OAI21_X1 U10097 ( .B1(n9402), .B2(n10217), .A(n8638), .ZN(n8639) );
  AOI21_X1 U10098 ( .B1(n9420), .B2(n8640), .A(n8639), .ZN(n8645) );
  AOI21_X1 U10099 ( .B1(n8642), .B2(n9913), .A(n8641), .ZN(n8643) );
  NAND2_X1 U10100 ( .A1(n9710), .A2(n8643), .ZN(n8644) );
  OAI211_X1 U10101 ( .C1(n8646), .C2(n9713), .A(n8645), .B(n8644), .ZN(
        P2_U3263) );
  AND2_X1 U10102 ( .A1(n8649), .A2(n8648), .ZN(n8829) );
  INV_X1 U10103 ( .A(n8829), .ZN(n8650) );
  NOR2_X1 U10104 ( .A1(n9749), .A2(n8650), .ZN(n8658) );
  NOR2_X1 U10105 ( .A1(n8651), .A2(n9775), .ZN(n8652) );
  AOI211_X1 U10106 ( .C1(n9773), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8658), .B(
        n8652), .ZN(n8653) );
  OAI21_X1 U10107 ( .B1(n8827), .B2(n9757), .A(n8653), .ZN(P2_U3265) );
  NAND2_X1 U10108 ( .A1(n8830), .A2(n8654), .ZN(n8655) );
  NAND2_X1 U10109 ( .A1(n8656), .A2(n8655), .ZN(n8828) );
  AND2_X1 U10110 ( .A1(n9773), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8657) );
  NOR2_X1 U10111 ( .A1(n8658), .A2(n8657), .ZN(n8660) );
  NAND2_X1 U10112 ( .A1(n8830), .A2(n9731), .ZN(n8659) );
  OAI211_X1 U10113 ( .C1(n8828), .C2(n9757), .A(n8660), .B(n8659), .ZN(
        P2_U3266) );
  XNOR2_X1 U10114 ( .A(n8662), .B(n8661), .ZN(n8842) );
  AOI21_X1 U10115 ( .B1(n8838), .B2(n8680), .A(n8663), .ZN(n8839) );
  AOI22_X1 U10116 ( .A1(n9773), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8664), .B2(
        n9771), .ZN(n8665) );
  OAI21_X1 U10117 ( .B1(n8666), .B2(n9775), .A(n8665), .ZN(n8676) );
  INV_X1 U10118 ( .A(n8667), .ZN(n8669) );
  AOI21_X1 U10119 ( .B1(n8669), .B2(n8668), .A(n9725), .ZN(n8674) );
  OAI22_X1 U10120 ( .A1(n8671), .A2(n9763), .B1(n8670), .B2(n9761), .ZN(n8672)
         );
  AOI21_X1 U10121 ( .B1(n8674), .B2(n8673), .A(n8672), .ZN(n8841) );
  NOR2_X1 U10122 ( .A1(n8841), .A2(n9749), .ZN(n8675) );
  AOI211_X1 U10123 ( .C1(n8806), .C2(n8839), .A(n8676), .B(n8675), .ZN(n8677)
         );
  OAI21_X1 U10124 ( .B1(n8842), .B2(n8808), .A(n8677), .ZN(P2_U3268) );
  XNOR2_X1 U10125 ( .A(n8679), .B(n8678), .ZN(n8847) );
  INV_X1 U10126 ( .A(n8680), .ZN(n8681) );
  AOI21_X1 U10127 ( .B1(n8843), .B2(n8703), .A(n8681), .ZN(n8844) );
  AOI22_X1 U10128 ( .A1(n9773), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8682), .B2(
        n9771), .ZN(n8683) );
  OAI21_X1 U10129 ( .B1(n8684), .B2(n9775), .A(n8683), .ZN(n8691) );
  XNOR2_X1 U10130 ( .A(n8686), .B(n8685), .ZN(n8689) );
  AOI222_X1 U10131 ( .A1(n9766), .A2(n8689), .B1(n8688), .B2(n8783), .C1(n8687), .C2(n8781), .ZN(n8846) );
  NOR2_X1 U10132 ( .A1(n8846), .A2(n9749), .ZN(n8690) );
  AOI211_X1 U10133 ( .C1(n8806), .C2(n8844), .A(n8691), .B(n8690), .ZN(n8692)
         );
  OAI21_X1 U10134 ( .B1(n8847), .B2(n8808), .A(n8692), .ZN(P2_U3269) );
  XNOR2_X1 U10135 ( .A(n8694), .B(n8693), .ZN(n8852) );
  NOR2_X1 U10136 ( .A1(n8695), .A2(n9775), .ZN(n8710) );
  INV_X1 U10137 ( .A(n8696), .ZN(n8722) );
  OAI21_X1 U10138 ( .B1(n8722), .B2(n8698), .A(n8697), .ZN(n8700) );
  AOI21_X1 U10139 ( .B1(n8700), .B2(n8699), .A(n9725), .ZN(n8702) );
  NOR2_X1 U10140 ( .A1(n8702), .A2(n8701), .ZN(n8851) );
  INV_X1 U10141 ( .A(n8715), .ZN(n8705) );
  INV_X1 U10142 ( .A(n8703), .ZN(n8704) );
  AOI211_X1 U10143 ( .C1(n8849), .C2(n8705), .A(n9842), .B(n8704), .ZN(n8848)
         );
  AOI22_X1 U10144 ( .A1(n8848), .A2(n8707), .B1(n9771), .B2(n8706), .ZN(n8708)
         );
  AOI21_X1 U10145 ( .B1(n8851), .B2(n8708), .A(n9773), .ZN(n8709) );
  AOI211_X1 U10146 ( .C1(n9749), .C2(P2_REG2_REG_26__SCAN_IN), .A(n8710), .B(
        n8709), .ZN(n8711) );
  OAI21_X1 U10147 ( .B1(n8852), .B2(n8808), .A(n8711), .ZN(P2_U3270) );
  XNOR2_X1 U10148 ( .A(n8713), .B(n8712), .ZN(n8857) );
  INV_X1 U10149 ( .A(n8714), .ZN(n8716) );
  AOI211_X1 U10150 ( .C1(n8854), .C2(n8716), .A(n9842), .B(n8715), .ZN(n8853)
         );
  AOI22_X1 U10151 ( .A1(n9749), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8717), .B2(
        n9771), .ZN(n8718) );
  OAI21_X1 U10152 ( .B1(n8719), .B2(n9775), .A(n8718), .ZN(n8728) );
  NOR2_X1 U10153 ( .A1(n8721), .A2(n8720), .ZN(n8724) );
  AOI211_X1 U10154 ( .C1(n8724), .C2(n8723), .A(n9725), .B(n8722), .ZN(n8726)
         );
  NOR2_X1 U10155 ( .A1(n8726), .A2(n8725), .ZN(n8856) );
  NOR2_X1 U10156 ( .A1(n8856), .A2(n8740), .ZN(n8727) );
  AOI211_X1 U10157 ( .C1(n8853), .C2(n9745), .A(n8728), .B(n8727), .ZN(n8729)
         );
  OAI21_X1 U10158 ( .B1(n8857), .B2(n8808), .A(n8729), .ZN(P2_U3271) );
  AOI21_X1 U10159 ( .B1(n8736), .B2(n8731), .A(n8730), .ZN(n8862) );
  XNOR2_X1 U10160 ( .A(n8734), .B(n8746), .ZN(n8859) );
  AOI22_X1 U10161 ( .A1(n9773), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8732), .B2(
        n9771), .ZN(n8733) );
  OAI21_X1 U10162 ( .B1(n8734), .B2(n9775), .A(n8733), .ZN(n8742) );
  XOR2_X1 U10163 ( .A(n8736), .B(n8735), .Z(n8739) );
  AOI222_X1 U10164 ( .A1(n9766), .A2(n8739), .B1(n8738), .B2(n8781), .C1(n8737), .C2(n8783), .ZN(n8861) );
  NOR2_X1 U10165 ( .A1(n8861), .A2(n8740), .ZN(n8741) );
  AOI211_X1 U10166 ( .C1(n8859), .C2(n8806), .A(n8742), .B(n8741), .ZN(n8743)
         );
  OAI21_X1 U10167 ( .B1(n8862), .B2(n8808), .A(n8743), .ZN(P2_U3272) );
  OAI21_X1 U10168 ( .B1(n8745), .B2(n8750), .A(n8744), .ZN(n8867) );
  AOI21_X1 U10169 ( .B1(n8863), .B2(n8760), .A(n4636), .ZN(n8864) );
  INV_X1 U10170 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8747) );
  OAI22_X1 U10171 ( .A1(n8748), .A2(n9775), .B1(n7202), .B2(n8747), .ZN(n8757)
         );
  NAND2_X1 U10172 ( .A1(n8770), .A2(n8749), .ZN(n8751) );
  XNOR2_X1 U10173 ( .A(n8751), .B(n8750), .ZN(n8753) );
  AOI21_X1 U10174 ( .B1(n8753), .B2(n9766), .A(n8752), .ZN(n8866) );
  NAND2_X1 U10175 ( .A1(n9771), .A2(n8754), .ZN(n8755) );
  AOI21_X1 U10176 ( .B1(n8866), .B2(n8755), .A(n9749), .ZN(n8756) );
  AOI211_X1 U10177 ( .C1(n8864), .C2(n8806), .A(n8757), .B(n8756), .ZN(n8758)
         );
  OAI21_X1 U10178 ( .B1(n8867), .B2(n8808), .A(n8758), .ZN(P2_U3273) );
  XOR2_X1 U10179 ( .A(n8759), .B(n8766), .Z(n8872) );
  AOI21_X1 U10180 ( .B1(n8868), .B2(n4405), .A(n4632), .ZN(n8869) );
  AOI22_X1 U10181 ( .A1(n9749), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8761), .B2(
        n9771), .ZN(n8762) );
  OAI21_X1 U10182 ( .B1(n8763), .B2(n9775), .A(n8762), .ZN(n8773) );
  NAND2_X1 U10183 ( .A1(n8765), .A2(n8764), .ZN(n8767) );
  AOI21_X1 U10184 ( .B1(n8767), .B2(n8766), .A(n9725), .ZN(n8771) );
  OAI22_X1 U10185 ( .A1(n8768), .A2(n9761), .B1(n8799), .B2(n9763), .ZN(n8769)
         );
  AOI21_X1 U10186 ( .B1(n8771), .B2(n8770), .A(n8769), .ZN(n8871) );
  NOR2_X1 U10187 ( .A1(n8871), .A2(n9773), .ZN(n8772) );
  AOI211_X1 U10188 ( .C1(n8869), .C2(n8806), .A(n8773), .B(n8772), .ZN(n8774)
         );
  OAI21_X1 U10189 ( .B1(n8872), .B2(n8808), .A(n8774), .ZN(P2_U3274) );
  XOR2_X1 U10190 ( .A(n8775), .B(n8779), .Z(n8877) );
  XNOR2_X1 U10191 ( .A(n8790), .B(n8873), .ZN(n8874) );
  AOI22_X1 U10192 ( .A1(n9773), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8776), .B2(
        n9771), .ZN(n8777) );
  OAI21_X1 U10193 ( .B1(n8778), .B2(n9775), .A(n8777), .ZN(n8787) );
  XNOR2_X1 U10194 ( .A(n8780), .B(n8779), .ZN(n8785) );
  AOI222_X1 U10195 ( .A1(n9766), .A2(n8785), .B1(n8784), .B2(n8783), .C1(n8782), .C2(n8781), .ZN(n8876) );
  NOR2_X1 U10196 ( .A1(n8876), .A2(n9773), .ZN(n8786) );
  AOI211_X1 U10197 ( .C1(n8874), .C2(n8806), .A(n8787), .B(n8786), .ZN(n8788)
         );
  OAI21_X1 U10198 ( .B1(n8877), .B2(n8808), .A(n8788), .ZN(P2_U3275) );
  XNOR2_X1 U10199 ( .A(n8789), .B(n8797), .ZN(n8882) );
  AOI21_X1 U10200 ( .B1(n8878), .B2(n8791), .A(n8790), .ZN(n8879) );
  INV_X1 U10201 ( .A(n8878), .ZN(n8794) );
  AOI22_X1 U10202 ( .A1(n9773), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8792), .B2(
        n9771), .ZN(n8793) );
  OAI21_X1 U10203 ( .B1(n8794), .B2(n9775), .A(n8793), .ZN(n8805) );
  NAND2_X1 U10204 ( .A1(n8796), .A2(n8795), .ZN(n8798) );
  AOI21_X1 U10205 ( .B1(n8798), .B2(n8797), .A(n9725), .ZN(n8803) );
  OAI22_X1 U10206 ( .A1(n8800), .A2(n9763), .B1(n8799), .B2(n9761), .ZN(n8801)
         );
  AOI21_X1 U10207 ( .B1(n8803), .B2(n8802), .A(n8801), .ZN(n8881) );
  NOR2_X1 U10208 ( .A1(n8881), .A2(n9773), .ZN(n8804) );
  AOI211_X1 U10209 ( .C1(n8879), .C2(n8806), .A(n8805), .B(n8804), .ZN(n8807)
         );
  OAI21_X1 U10210 ( .B1(n8882), .B2(n8808), .A(n8807), .ZN(P2_U3276) );
  OAI21_X1 U10211 ( .B1(n8820), .B2(n8810), .A(n8809), .ZN(n8812) );
  OAI22_X1 U10212 ( .A1(n6816), .A2(n9763), .B1(n9764), .B2(n9761), .ZN(n8811)
         );
  AOI21_X1 U10213 ( .B1(n8812), .B2(n9766), .A(n8811), .ZN(n9805) );
  MUX2_X1 U10214 ( .A(n6596), .B(n9805), .S(n7202), .Z(n8824) );
  OAI211_X1 U10215 ( .C1(n8814), .C2(n9806), .A(n6266), .B(n8813), .ZN(n9804)
         );
  NOR2_X1 U10216 ( .A1(n9804), .A2(n8815), .ZN(n8819) );
  OAI22_X1 U10217 ( .A1(n9775), .A2(n9806), .B1(n8817), .B2(n8816), .ZN(n8818)
         );
  NOR2_X1 U10218 ( .A1(n8819), .A2(n8818), .ZN(n8823) );
  NAND2_X1 U10219 ( .A1(n8821), .A2(n8820), .ZN(n9802) );
  NAND3_X1 U10220 ( .A1(n9803), .A2(n9802), .A3(n9746), .ZN(n8822) );
  NAND3_X1 U10221 ( .A1(n8824), .A2(n8823), .A3(n8822), .ZN(P2_U3290) );
  AOI21_X1 U10222 ( .B1(n8825), .B2(n9824), .A(n8829), .ZN(n8826) );
  OAI21_X1 U10223 ( .B1(n8827), .B2(n9842), .A(n8826), .ZN(n8904) );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8904), .S(n9873), .Z(
        P2_U3551) );
  AOI21_X1 U10225 ( .B1(n8830), .B2(n9824), .A(n8829), .ZN(n8831) );
  NAND2_X1 U10226 ( .A1(n8832), .A2(n8831), .ZN(n8905) );
  MUX2_X1 U10227 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8905), .S(n9873), .Z(
        P2_U3550) );
  AOI22_X1 U10228 ( .A1(n8834), .A2(n6266), .B1(n9824), .B2(n8833), .ZN(n8835)
         );
  OAI211_X1 U10229 ( .C1(n8837), .C2(n8897), .A(n8836), .B(n8835), .ZN(n8906)
         );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8906), .S(n9873), .Z(
        P2_U3549) );
  AOI22_X1 U10231 ( .A1(n8839), .A2(n6266), .B1(n9824), .B2(n8838), .ZN(n8840)
         );
  OAI211_X1 U10232 ( .C1(n8842), .C2(n8897), .A(n8841), .B(n8840), .ZN(n8907)
         );
  MUX2_X1 U10233 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8907), .S(n9873), .Z(
        P2_U3548) );
  AOI22_X1 U10234 ( .A1(n8844), .A2(n6266), .B1(n9824), .B2(n8843), .ZN(n8845)
         );
  OAI211_X1 U10235 ( .C1(n8847), .C2(n8897), .A(n8846), .B(n8845), .ZN(n8908)
         );
  MUX2_X1 U10236 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8908), .S(n9873), .Z(
        P2_U3547) );
  AOI21_X1 U10237 ( .B1(n9824), .B2(n8849), .A(n8848), .ZN(n8850) );
  OAI211_X1 U10238 ( .C1(n8852), .C2(n8897), .A(n8851), .B(n8850), .ZN(n8909)
         );
  MUX2_X1 U10239 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8909), .S(n9873), .Z(
        P2_U3546) );
  AOI21_X1 U10240 ( .B1(n9824), .B2(n8854), .A(n8853), .ZN(n8855) );
  OAI211_X1 U10241 ( .C1(n8857), .C2(n8897), .A(n8856), .B(n8855), .ZN(n8910)
         );
  MUX2_X1 U10242 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8910), .S(n9873), .Z(
        P2_U3545) );
  AOI22_X1 U10243 ( .A1(n8859), .A2(n6266), .B1(n9824), .B2(n8858), .ZN(n8860)
         );
  OAI211_X1 U10244 ( .C1(n8862), .C2(n8897), .A(n8861), .B(n8860), .ZN(n8911)
         );
  MUX2_X1 U10245 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8911), .S(n9873), .Z(
        P2_U3544) );
  AOI22_X1 U10246 ( .A1(n8864), .A2(n6266), .B1(n9824), .B2(n8863), .ZN(n8865)
         );
  OAI211_X1 U10247 ( .C1(n8867), .C2(n8897), .A(n8866), .B(n8865), .ZN(n8912)
         );
  MUX2_X1 U10248 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8912), .S(n9873), .Z(
        P2_U3543) );
  AOI22_X1 U10249 ( .A1(n8869), .A2(n6266), .B1(n9824), .B2(n8868), .ZN(n8870)
         );
  OAI211_X1 U10250 ( .C1(n8872), .C2(n8897), .A(n8871), .B(n8870), .ZN(n8913)
         );
  MUX2_X1 U10251 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8913), .S(n9873), .Z(
        P2_U3542) );
  AOI22_X1 U10252 ( .A1(n8874), .A2(n6266), .B1(n9824), .B2(n8873), .ZN(n8875)
         );
  OAI211_X1 U10253 ( .C1(n8877), .C2(n8897), .A(n8876), .B(n8875), .ZN(n8914)
         );
  MUX2_X1 U10254 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8914), .S(n9873), .Z(
        P2_U3541) );
  AOI22_X1 U10255 ( .A1(n8879), .A2(n6266), .B1(n9824), .B2(n8878), .ZN(n8880)
         );
  OAI211_X1 U10256 ( .C1(n8882), .C2(n8897), .A(n8881), .B(n8880), .ZN(n8915)
         );
  MUX2_X1 U10257 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8915), .S(n9873), .Z(
        P2_U3540) );
  AOI21_X1 U10258 ( .B1(n9824), .B2(n8884), .A(n8883), .ZN(n8885) );
  OAI211_X1 U10259 ( .C1(n8887), .C2(n8897), .A(n8886), .B(n8885), .ZN(n8916)
         );
  MUX2_X1 U10260 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8916), .S(n9873), .Z(
        P2_U3539) );
  AOI22_X1 U10261 ( .A1(n8889), .A2(n6266), .B1(n9824), .B2(n8888), .ZN(n8890)
         );
  OAI211_X1 U10262 ( .C1(n8892), .C2(n8897), .A(n8891), .B(n8890), .ZN(n8917)
         );
  MUX2_X1 U10263 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8917), .S(n9873), .Z(
        P2_U3538) );
  AOI211_X1 U10264 ( .C1(n9824), .C2(n8895), .A(n8894), .B(n8893), .ZN(n8896)
         );
  OAI21_X1 U10265 ( .B1(n8898), .B2(n8897), .A(n8896), .ZN(n8918) );
  MUX2_X1 U10266 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8918), .S(n9873), .Z(
        P2_U3537) );
  AOI22_X1 U10267 ( .A1(n8900), .A2(n6266), .B1(n9824), .B2(n8899), .ZN(n8901)
         );
  OAI211_X1 U10268 ( .C1(n9827), .C2(n8903), .A(n8902), .B(n8901), .ZN(n8919)
         );
  MUX2_X1 U10269 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8919), .S(n9873), .Z(
        P2_U3536) );
  MUX2_X1 U10270 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8904), .S(n9856), .Z(
        P2_U3519) );
  MUX2_X1 U10271 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8905), .S(n9856), .Z(
        P2_U3518) );
  MUX2_X1 U10272 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8906), .S(n9856), .Z(
        P2_U3517) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8907), .S(n9856), .Z(
        P2_U3516) );
  MUX2_X1 U10274 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8908), .S(n9856), .Z(
        P2_U3515) );
  MUX2_X1 U10275 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8909), .S(n9856), .Z(
        P2_U3514) );
  MUX2_X1 U10276 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8910), .S(n9856), .Z(
        P2_U3513) );
  MUX2_X1 U10277 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8911), .S(n9856), .Z(
        P2_U3512) );
  MUX2_X1 U10278 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8912), .S(n9856), .Z(
        P2_U3511) );
  MUX2_X1 U10279 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8913), .S(n9856), .Z(
        P2_U3510) );
  MUX2_X1 U10280 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8914), .S(n9856), .Z(
        P2_U3509) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8915), .S(n9856), .Z(
        P2_U3508) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8916), .S(n9856), .Z(
        P2_U3507) );
  MUX2_X1 U10283 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8917), .S(n9856), .Z(
        P2_U3505) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8918), .S(n9856), .Z(
        P2_U3502) );
  MUX2_X1 U10285 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8919), .S(n9856), .Z(
        P2_U3499) );
  MUX2_X1 U10286 ( .A(n8920), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10287 ( .A(n8921), .ZN(n8925) );
  AOI21_X1 U10288 ( .B1(n8923), .B2(n8958), .A(n8922), .ZN(n8924) );
  AOI21_X1 U10289 ( .B1(n8925), .B2(n8958), .A(n8924), .ZN(n8930) );
  NAND2_X1 U10290 ( .A1(n9173), .A2(n9438), .ZN(n8927) );
  AOI22_X1 U10291 ( .A1(n9083), .A2(n8980), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8926) );
  OAI211_X1 U10292 ( .C1(n9452), .C2(n9204), .A(n8927), .B(n8926), .ZN(n8928)
         );
  AOI21_X1 U10293 ( .B1(n9331), .B2(n5797), .A(n8928), .ZN(n8929) );
  OAI21_X1 U10294 ( .B1(n8930), .B2(n9446), .A(n8929), .ZN(P1_U3214) );
  INV_X1 U10295 ( .A(n8990), .ZN(n8932) );
  NOR3_X1 U10296 ( .A1(n4456), .A2(n8932), .A3(n8931), .ZN(n8934) );
  INV_X1 U10297 ( .A(n8933), .ZN(n8968) );
  OAI21_X1 U10298 ( .B1(n8934), .B2(n8968), .A(n9002), .ZN(n8939) );
  NOR2_X1 U10299 ( .A1(n9452), .A2(n8935), .ZN(n8937) );
  NAND2_X1 U10300 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9065) );
  OAI21_X1 U10301 ( .B1(n9234), .B2(n8983), .A(n9065), .ZN(n8936) );
  AOI211_X1 U10302 ( .C1(n8980), .C2(n9011), .A(n8937), .B(n8936), .ZN(n8938)
         );
  OAI211_X1 U10303 ( .C1(n9078), .C2(n9010), .A(n8939), .B(n8938), .ZN(
        P1_U3217) );
  INV_X1 U10304 ( .A(n9341), .ZN(n9082) );
  OAI21_X1 U10305 ( .B1(n8942), .B2(n8941), .A(n8940), .ZN(n8943) );
  NAND2_X1 U10306 ( .A1(n8943), .A2(n9002), .ZN(n8948) );
  INV_X1 U10307 ( .A(n9237), .ZN(n8946) );
  AOI22_X1 U10308 ( .A1(n9081), .A2(n8980), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8944) );
  OAI21_X1 U10309 ( .B1(n9233), .B2(n8983), .A(n8944), .ZN(n8945) );
  AOI21_X1 U10310 ( .B1(n8946), .B2(n9003), .A(n8945), .ZN(n8947) );
  OAI211_X1 U10311 ( .C1(n9082), .C2(n9010), .A(n8948), .B(n8947), .ZN(
        P1_U3221) );
  AOI21_X1 U10312 ( .B1(n8950), .B2(n8949), .A(n9000), .ZN(n8956) );
  OAI22_X1 U10313 ( .A1(n9202), .A2(n9435), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8951), .ZN(n8952) );
  AOI21_X1 U10314 ( .B1(n9176), .B2(n9003), .A(n8952), .ZN(n8953) );
  OAI21_X1 U10315 ( .B1(n9089), .B2(n8983), .A(n8953), .ZN(n8954) );
  AOI21_X1 U10316 ( .B1(n9317), .B2(n5797), .A(n8954), .ZN(n8955) );
  OAI21_X1 U10317 ( .B1(n8956), .B2(n9446), .A(n8955), .ZN(P1_U3223) );
  AND3_X1 U10318 ( .A1(n8921), .A2(n8958), .A3(n8957), .ZN(n8959) );
  OAI21_X1 U10319 ( .B1(n8960), .B2(n8959), .A(n9002), .ZN(n8964) );
  AOI22_X1 U10320 ( .A1(n9219), .A2(n8980), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8961) );
  OAI21_X1 U10321 ( .B1(n9452), .B2(n9190), .A(n8961), .ZN(n8962) );
  AOI21_X1 U10322 ( .B1(n9185), .B2(n9438), .A(n8962), .ZN(n8963) );
  OAI211_X1 U10323 ( .C1(n9192), .C2(n9010), .A(n8964), .B(n8963), .ZN(
        P1_U3227) );
  INV_X1 U10324 ( .A(n8965), .ZN(n8967) );
  NOR3_X1 U10325 ( .A1(n8968), .A2(n8967), .A3(n8966), .ZN(n8971) );
  INV_X1 U10326 ( .A(n8969), .ZN(n8970) );
  OAI21_X1 U10327 ( .B1(n8971), .B2(n8970), .A(n9002), .ZN(n8975) );
  AOI22_X1 U10328 ( .A1(n9221), .A2(n9438), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8972) );
  OAI21_X1 U10329 ( .B1(n9247), .B2(n9435), .A(n8972), .ZN(n8973) );
  AOI21_X1 U10330 ( .B1(n9255), .B2(n9003), .A(n8973), .ZN(n8974) );
  OAI211_X1 U10331 ( .C1(n9259), .C2(n9010), .A(n8975), .B(n8974), .ZN(
        P1_U3231) );
  NAND2_X1 U10332 ( .A1(n8977), .A2(n8976), .ZN(n8979) );
  XNOR2_X1 U10333 ( .A(n8979), .B(n8978), .ZN(n8986) );
  AOI22_X1 U10334 ( .A1(n9221), .A2(n8980), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8982) );
  NAND2_X1 U10335 ( .A1(n9213), .A2(n9003), .ZN(n8981) );
  OAI211_X1 U10336 ( .C1(n9086), .C2(n8983), .A(n8982), .B(n8981), .ZN(n8984)
         );
  AOI21_X1 U10337 ( .B1(n9334), .B2(n5797), .A(n8984), .ZN(n8985) );
  OAI21_X1 U10338 ( .B1(n8986), .B2(n9446), .A(n8985), .ZN(P1_U3233) );
  AOI21_X1 U10339 ( .B1(n8988), .B2(n8990), .A(n8987), .ZN(n8989) );
  AOI21_X1 U10340 ( .B1(n4456), .B2(n8990), .A(n8989), .ZN(n8997) );
  NAND2_X1 U10341 ( .A1(n9077), .A2(n9438), .ZN(n8991) );
  NAND2_X1 U10342 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9622) );
  OAI211_X1 U10343 ( .C1(n8992), .C2(n9435), .A(n8991), .B(n9622), .ZN(n8993)
         );
  AOI21_X1 U10344 ( .B1(n8994), .B2(n9003), .A(n8993), .ZN(n8996) );
  NAND2_X1 U10345 ( .A1(n9356), .A2(n5797), .ZN(n8995) );
  OAI211_X1 U10346 ( .C1(n8997), .C2(n9446), .A(n8996), .B(n8995), .ZN(
        P1_U3236) );
  OAI21_X1 U10347 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(n9001) );
  NAND3_X1 U10348 ( .A1(n4895), .A2(n9002), .A3(n9001), .ZN(n9009) );
  INV_X1 U10349 ( .A(n9159), .ZN(n9004) );
  AOI22_X1 U10350 ( .A1(n9004), .A2(n9003), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9005) );
  OAI21_X1 U10351 ( .B1(n9006), .B2(n9435), .A(n9005), .ZN(n9007) );
  AOI21_X1 U10352 ( .B1(n9438), .B2(n9157), .A(n9007), .ZN(n9008) );
  OAI211_X1 U10353 ( .C1(n9160), .C2(n9010), .A(n9009), .B(n9008), .ZN(
        P1_U3238) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9111), .S(n9019), .Z(
        P1_U3585) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9147), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10356 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9157), .S(n9019), .Z(
        P1_U3582) );
  MUX2_X1 U10357 ( .A(n9174), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9026), .Z(
        P1_U3581) );
  MUX2_X1 U10358 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9185), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10359 ( .A(n9173), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9026), .Z(
        P1_U3579) );
  MUX2_X1 U10360 ( .A(n9219), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9026), .Z(
        P1_U3578) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9083), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10362 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9221), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9081), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10364 ( .A(n9077), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9026), .Z(
        P1_U3574) );
  MUX2_X1 U10365 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9011), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9012), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9013), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9014), .S(n9019), .Z(
        P1_U3570) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9015), .S(n9019), .Z(
        P1_U3569) );
  MUX2_X1 U10370 ( .A(n9437), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9026), .Z(
        P1_U3568) );
  MUX2_X1 U10371 ( .A(n9016), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9026), .Z(
        P1_U3566) );
  MUX2_X1 U10372 ( .A(n9017), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9026), .Z(
        P1_U3564) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9018), .S(n9019), .Z(
        P1_U3563) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9020), .S(n9019), .Z(
        P1_U3562) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9021), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10376 ( .A(n9022), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9026), .Z(
        P1_U3560) );
  MUX2_X1 U10377 ( .A(n9023), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9026), .Z(
        P1_U3559) );
  MUX2_X1 U10378 ( .A(n9024), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9026), .Z(
        P1_U3558) );
  MUX2_X1 U10379 ( .A(n9025), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9026), .Z(
        P1_U3557) );
  MUX2_X1 U10380 ( .A(n9027), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9026), .Z(
        P1_U3556) );
  INV_X1 U10381 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9039) );
  AOI22_X1 U10382 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9040), .B1(n9620), .B2(
        n9039), .ZN(n9626) );
  INV_X1 U10383 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9037) );
  AOI22_X1 U10384 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(n9601), .B1(n9038), .B2(
        n9037), .ZN(n9610) );
  INV_X1 U10385 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9482) );
  AOI22_X1 U10386 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(n9593), .B1(n9036), .B2(
        n9482), .ZN(n9596) );
  INV_X1 U10387 ( .A(n9552), .ZN(n9033) );
  MUX2_X1 U10388 ( .A(n9028), .B(P1_REG1_REG_12__SCAN_IN), .S(n9543), .Z(n9539) );
  NOR2_X1 U10389 ( .A1(n9539), .A2(n9540), .ZN(n9538) );
  NOR2_X1 U10390 ( .A1(n9543), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9031) );
  NOR2_X1 U10391 ( .A1(n9538), .A2(n9031), .ZN(n9559) );
  MUX2_X1 U10392 ( .A(n9032), .B(P1_REG1_REG_13__SCAN_IN), .S(n9552), .Z(n9558) );
  AOI22_X1 U10393 ( .A1(n9568), .A2(n5398), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9049), .ZN(n9565) );
  NAND2_X1 U10394 ( .A1(n9581), .A2(n9034), .ZN(n9035) );
  NAND2_X1 U10395 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9583), .ZN(n9582) );
  NAND2_X1 U10396 ( .A1(n9035), .A2(n9582), .ZN(n9595) );
  NAND2_X1 U10397 ( .A1(n9596), .A2(n9595), .ZN(n9594) );
  OAI21_X1 U10398 ( .B1(n9036), .B2(n9482), .A(n9594), .ZN(n9609) );
  NAND2_X1 U10399 ( .A1(n9610), .A2(n9609), .ZN(n9608) );
  OAI21_X1 U10400 ( .B1(n9038), .B2(n9037), .A(n9608), .ZN(n9627) );
  NOR2_X1 U10401 ( .A1(n9626), .A2(n9627), .ZN(n9628) );
  AOI21_X1 U10402 ( .B1(n9040), .B2(n9039), .A(n9628), .ZN(n9041) );
  OR2_X1 U10403 ( .A1(n9042), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9044) );
  XNOR2_X1 U10404 ( .A(n9543), .B(n9045), .ZN(n9545) );
  NAND2_X1 U10405 ( .A1(n9543), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U10406 ( .A1(n9544), .A2(n9046), .ZN(n9554) );
  XNOR2_X1 U10407 ( .A(n9552), .B(n9047), .ZN(n9555) );
  NAND2_X1 U10408 ( .A1(n9554), .A2(n9555), .ZN(n9553) );
  INV_X1 U10409 ( .A(n9553), .ZN(n9048) );
  NAND2_X1 U10410 ( .A1(n9050), .A2(n9049), .ZN(n9051) );
  XNOR2_X1 U10411 ( .A(n9050), .B(n9568), .ZN(n9570) );
  NAND2_X1 U10412 ( .A1(n9570), .A2(n7447), .ZN(n9569) );
  NAND2_X1 U10413 ( .A1(n9051), .A2(n9569), .ZN(n9053) );
  NOR2_X1 U10414 ( .A1(n9052), .A2(n9053), .ZN(n9054) );
  XNOR2_X1 U10415 ( .A(n9053), .B(n9052), .ZN(n9578) );
  NOR2_X1 U10416 ( .A1(n5432), .A2(n9578), .ZN(n9577) );
  NAND2_X1 U10417 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9593), .ZN(n9055) );
  OAI21_X1 U10418 ( .B1(n9593), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9055), .ZN(
        n9589) );
  NOR2_X1 U10419 ( .A1(n9590), .A2(n9589), .ZN(n9588) );
  AOI21_X1 U10420 ( .B1(n9593), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9588), .ZN(
        n9603) );
  NAND2_X1 U10421 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9601), .ZN(n9056) );
  OAI21_X1 U10422 ( .B1(n9601), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9056), .ZN(
        n9604) );
  NOR2_X1 U10423 ( .A1(n9603), .A2(n9604), .ZN(n9602) );
  OR2_X1 U10424 ( .A1(n9620), .A2(n9057), .ZN(n9059) );
  NAND2_X1 U10425 ( .A1(n9620), .A2(n9057), .ZN(n9058) );
  AND2_X1 U10426 ( .A1(n9059), .A2(n9058), .ZN(n9615) );
  NOR2_X1 U10427 ( .A1(n9614), .A2(n9615), .ZN(n9616) );
  AOI21_X1 U10428 ( .B1(n9620), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9616), .ZN(
        n9060) );
  AOI22_X1 U10429 ( .A1(n9063), .A2(n9625), .B1(n9619), .B2(n9062), .ZN(n9064)
         );
  OAI211_X1 U10430 ( .C1(n4733), .C2(n9631), .A(n9066), .B(n9065), .ZN(
        P1_U3260) );
  INV_X1 U10431 ( .A(P1_B_REG_SCAN_IN), .ZN(n10017) );
  NOR2_X1 U10432 ( .A1(n9067), .A2(n10017), .ZN(n9068) );
  NOR2_X1 U10433 ( .A1(n9269), .A2(n9068), .ZN(n9112) );
  NAND2_X1 U10434 ( .A1(n9069), .A2(n9112), .ZN(n9292) );
  NOR2_X1 U10435 ( .A1(n9278), .A2(n9292), .ZN(n9074) );
  AOI21_X1 U10436 ( .B1(n9278), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9074), .ZN(
        n9071) );
  NAND2_X1 U10437 ( .A1(n9287), .A2(n9280), .ZN(n9070) );
  OAI211_X1 U10438 ( .C1(n9289), .C2(n9163), .A(n9071), .B(n9070), .ZN(
        P1_U3261) );
  INV_X1 U10439 ( .A(n9115), .ZN(n9072) );
  NAND2_X1 U10440 ( .A1(n9073), .A2(n9072), .ZN(n9290) );
  NAND3_X1 U10441 ( .A1(n9291), .A2(n9226), .A3(n9290), .ZN(n9076) );
  AOI21_X1 U10442 ( .B1(n9278), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9074), .ZN(
        n9075) );
  OAI211_X1 U10443 ( .C1(n9294), .C2(n9258), .A(n9076), .B(n9075), .ZN(
        P1_U3262) );
  NOR2_X1 U10444 ( .A1(n9351), .A2(n9077), .ZN(n9079) );
  NAND2_X1 U10445 ( .A1(n9229), .A2(n9231), .ZN(n9228) );
  NAND2_X1 U10446 ( .A1(n9215), .A2(n9233), .ZN(n9085) );
  NAND2_X1 U10447 ( .A1(n9331), .A2(n9219), .ZN(n9087) );
  AOI22_X1 U10448 ( .A1(n9198), .A2(n9087), .B1(n9208), .B2(n9086), .ZN(n9188)
         );
  NAND2_X1 U10449 ( .A1(n9091), .A2(n9090), .ZN(n9139) );
  INV_X1 U10450 ( .A(n9296), .ZN(n9121) );
  AOI22_X1 U10451 ( .A1(n9299), .A2(n9280), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9253), .ZN(n9120) );
  INV_X1 U10452 ( .A(n9098), .ZN(n9099) );
  XNOR2_X1 U10453 ( .A(n9110), .B(n4900), .ZN(n9114) );
  AOI22_X1 U10454 ( .A1(n9147), .A2(n9220), .B1(n9112), .B2(n9111), .ZN(n9113)
         );
  AOI211_X1 U10455 ( .C1(n9299), .C2(n9130), .A(n9688), .B(n9115), .ZN(n9298)
         );
  INV_X1 U10456 ( .A(n9298), .ZN(n9117) );
  OAI22_X1 U10457 ( .A1(n9117), .A2(n9275), .B1(n9274), .B2(n9116), .ZN(n9118)
         );
  OAI21_X1 U10458 ( .B1(n9297), .B2(n9118), .A(n9276), .ZN(n9119) );
  OAI211_X1 U10459 ( .C1(n9121), .C2(n9262), .A(n9120), .B(n9119), .ZN(
        P1_U3355) );
  OAI21_X1 U10460 ( .B1(n9124), .B2(n9123), .A(n9122), .ZN(n9305) );
  XNOR2_X1 U10461 ( .A(n9126), .B(n9125), .ZN(n9127) );
  OAI222_X1 U10462 ( .A1(n9269), .A2(n9129), .B1(n9267), .B2(n9128), .C1(n9265), .C2(n9127), .ZN(n9301) );
  INV_X1 U10463 ( .A(n9140), .ZN(n9132) );
  INV_X1 U10464 ( .A(n9130), .ZN(n9131) );
  AOI211_X1 U10465 ( .C1(n9303), .C2(n9132), .A(n9688), .B(n9131), .ZN(n9302)
         );
  NAND2_X1 U10466 ( .A1(n9302), .A2(n9252), .ZN(n9135) );
  AOI22_X1 U10467 ( .A1(n9133), .A2(n9254), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9253), .ZN(n9134) );
  OAI211_X1 U10468 ( .C1(n9136), .C2(n9258), .A(n9135), .B(n9134), .ZN(n9137)
         );
  AOI21_X1 U10469 ( .B1(n9301), .B2(n9276), .A(n9137), .ZN(n9138) );
  OAI21_X1 U10470 ( .B1(n9305), .B2(n9262), .A(n9138), .ZN(P1_U3263) );
  XNOR2_X1 U10471 ( .A(n9139), .B(n9145), .ZN(n9310) );
  INV_X1 U10472 ( .A(n4441), .ZN(n9141) );
  AOI21_X1 U10473 ( .B1(n9306), .B2(n9141), .A(n9140), .ZN(n9307) );
  AOI22_X1 U10474 ( .A1(n9142), .A2(n9254), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9253), .ZN(n9143) );
  OAI21_X1 U10475 ( .B1(n9144), .B2(n9258), .A(n9143), .ZN(n9150) );
  XNOR2_X1 U10476 ( .A(n9146), .B(n9145), .ZN(n9148) );
  AOI222_X1 U10477 ( .A1(n9223), .A2(n9148), .B1(n9147), .B2(n9218), .C1(n9174), .C2(n9220), .ZN(n9309) );
  NOR2_X1 U10478 ( .A1(n9309), .A2(n9253), .ZN(n9149) );
  AOI211_X1 U10479 ( .C1(n9226), .C2(n9307), .A(n9150), .B(n9149), .ZN(n9151)
         );
  OAI21_X1 U10480 ( .B1(n9310), .B2(n9262), .A(n9151), .ZN(P1_U3264) );
  XNOR2_X1 U10481 ( .A(n9152), .B(n9155), .ZN(n9316) );
  INV_X1 U10482 ( .A(n9153), .ZN(n9154) );
  NOR2_X1 U10483 ( .A1(n4418), .A2(n9154), .ZN(n9156) );
  XNOR2_X1 U10484 ( .A(n9156), .B(n9155), .ZN(n9158) );
  AOI222_X1 U10485 ( .A1(n9223), .A2(n9158), .B1(n9185), .B2(n9220), .C1(n9157), .C2(n9218), .ZN(n9315) );
  OAI21_X1 U10486 ( .B1(n9159), .B2(n9274), .A(n9315), .ZN(n9165) );
  NOR2_X1 U10487 ( .A1(n9160), .A2(n4414), .ZN(n9161) );
  OR2_X1 U10488 ( .A1(n4441), .A2(n9161), .ZN(n9311) );
  AOI22_X1 U10489 ( .A1(n9312), .A2(n9280), .B1(n9278), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n9162) );
  OAI21_X1 U10490 ( .B1(n9311), .B2(n9163), .A(n9162), .ZN(n9164) );
  AOI21_X1 U10491 ( .B1(n9165), .B2(n9276), .A(n9164), .ZN(n9166) );
  OAI21_X1 U10492 ( .B1(n9316), .B2(n9262), .A(n9166), .ZN(P1_U3265) );
  AOI21_X1 U10493 ( .B1(n9172), .B2(n9167), .A(n4424), .ZN(n9321) );
  INV_X1 U10494 ( .A(n9168), .ZN(n9169) );
  NOR2_X1 U10495 ( .A1(n9170), .A2(n9169), .ZN(n9171) );
  XOR2_X1 U10496 ( .A(n9172), .B(n9171), .Z(n9175) );
  AOI222_X1 U10497 ( .A1(n9223), .A2(n9175), .B1(n9174), .B2(n9218), .C1(n9173), .C2(n9220), .ZN(n9320) );
  INV_X1 U10498 ( .A(n9320), .ZN(n9180) );
  AOI21_X1 U10499 ( .B1(n9317), .B2(n9191), .A(n4414), .ZN(n9318) );
  NAND2_X1 U10500 ( .A1(n9318), .A2(n9226), .ZN(n9178) );
  AOI22_X1 U10501 ( .A1(n9176), .A2(n9254), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9253), .ZN(n9177) );
  OAI211_X1 U10502 ( .C1(n9088), .C2(n9258), .A(n9178), .B(n9177), .ZN(n9179)
         );
  AOI21_X1 U10503 ( .B1(n9180), .B2(n9276), .A(n9179), .ZN(n9181) );
  OAI21_X1 U10504 ( .B1(n9321), .B2(n9262), .A(n9181), .ZN(P1_U3266) );
  NOR2_X1 U10505 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  XOR2_X1 U10506 ( .A(n9187), .B(n9184), .Z(n9186) );
  AOI222_X1 U10507 ( .A1(n9223), .A2(n9186), .B1(n9185), .B2(n9218), .C1(n9219), .C2(n9220), .ZN(n9327) );
  OR2_X1 U10508 ( .A1(n9188), .A2(n9187), .ZN(n9323) );
  NAND3_X1 U10509 ( .A1(n9323), .A2(n9322), .A3(n9283), .ZN(n9197) );
  INV_X1 U10510 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9189) );
  OAI22_X1 U10511 ( .A1(n9190), .A2(n9274), .B1(n9189), .B2(n9276), .ZN(n9195)
         );
  OAI211_X1 U10512 ( .C1(n9192), .C2(n9203), .A(n9366), .B(n9191), .ZN(n9326)
         );
  INV_X1 U10513 ( .A(n9252), .ZN(n9193) );
  NOR2_X1 U10514 ( .A1(n9326), .A2(n9193), .ZN(n9194) );
  AOI211_X1 U10515 ( .C1(n9280), .C2(n9324), .A(n9195), .B(n9194), .ZN(n9196)
         );
  OAI211_X1 U10516 ( .C1(n9278), .C2(n9327), .A(n9197), .B(n9196), .ZN(
        P1_U3267) );
  XOR2_X1 U10517 ( .A(n9199), .B(n9198), .Z(n9333) );
  XNOR2_X1 U10518 ( .A(n9200), .B(n9199), .ZN(n9201) );
  OAI222_X1 U10519 ( .A1(n9269), .A2(n9202), .B1(n9267), .B2(n9233), .C1(n9201), .C2(n9265), .ZN(n9329) );
  AOI211_X1 U10520 ( .C1(n9331), .C2(n4608), .A(n9688), .B(n9203), .ZN(n9330)
         );
  NAND2_X1 U10521 ( .A1(n9330), .A2(n9252), .ZN(n9207) );
  INV_X1 U10522 ( .A(n9204), .ZN(n9205) );
  AOI22_X1 U10523 ( .A1(n9205), .A2(n9254), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9253), .ZN(n9206) );
  OAI211_X1 U10524 ( .C1(n9208), .C2(n9258), .A(n9207), .B(n9206), .ZN(n9209)
         );
  AOI21_X1 U10525 ( .B1(n9329), .B2(n9276), .A(n9209), .ZN(n9210) );
  OAI21_X1 U10526 ( .B1(n9333), .B2(n9262), .A(n9210), .ZN(P1_U3268) );
  XOR2_X1 U10527 ( .A(n9217), .B(n9211), .Z(n9338) );
  AOI21_X1 U10528 ( .B1(n9334), .B2(n9235), .A(n9212), .ZN(n9335) );
  AOI22_X1 U10529 ( .A1(n9213), .A2(n9254), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9253), .ZN(n9214) );
  OAI21_X1 U10530 ( .B1(n9215), .B2(n9258), .A(n9214), .ZN(n9225) );
  XOR2_X1 U10531 ( .A(n9217), .B(n9216), .Z(n9222) );
  AOI222_X1 U10532 ( .A1(n9223), .A2(n9222), .B1(n9221), .B2(n9220), .C1(n9219), .C2(n9218), .ZN(n9337) );
  NOR2_X1 U10533 ( .A1(n9337), .A2(n9253), .ZN(n9224) );
  AOI211_X1 U10534 ( .C1(n9335), .C2(n9226), .A(n9225), .B(n9224), .ZN(n9227)
         );
  OAI21_X1 U10535 ( .B1(n9338), .B2(n9262), .A(n9227), .ZN(P1_U3269) );
  OAI21_X1 U10536 ( .B1(n9229), .B2(n9231), .A(n9228), .ZN(n9343) );
  AOI22_X1 U10537 ( .A1(n9341), .A2(n9280), .B1(n9278), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9241) );
  AOI21_X1 U10538 ( .B1(n9231), .B2(n9230), .A(n4427), .ZN(n9232) );
  OAI222_X1 U10539 ( .A1(n9267), .A2(n9234), .B1(n9269), .B2(n9233), .C1(n9265), .C2(n9232), .ZN(n9339) );
  INV_X1 U10540 ( .A(n9235), .ZN(n9236) );
  AOI211_X1 U10541 ( .C1(n9341), .C2(n9249), .A(n9688), .B(n9236), .ZN(n9340)
         );
  INV_X1 U10542 ( .A(n9340), .ZN(n9238) );
  OAI22_X1 U10543 ( .A1(n9238), .A2(n9275), .B1(n9274), .B2(n9237), .ZN(n9239)
         );
  OAI21_X1 U10544 ( .B1(n9339), .B2(n9239), .A(n9276), .ZN(n9240) );
  OAI211_X1 U10545 ( .C1(n9343), .C2(n9262), .A(n9241), .B(n9240), .ZN(
        P1_U3270) );
  XOR2_X1 U10546 ( .A(n9244), .B(n9242), .Z(n9348) );
  XOR2_X1 U10547 ( .A(n9244), .B(n9243), .Z(n9245) );
  OAI222_X1 U10548 ( .A1(n9267), .A2(n9247), .B1(n9269), .B2(n9246), .C1(n9245), .C2(n9265), .ZN(n9344) );
  INV_X1 U10549 ( .A(n9248), .ZN(n9251) );
  INV_X1 U10550 ( .A(n9249), .ZN(n9250) );
  AOI211_X1 U10551 ( .C1(n9346), .C2(n9251), .A(n9688), .B(n9250), .ZN(n9345)
         );
  NAND2_X1 U10552 ( .A1(n9345), .A2(n9252), .ZN(n9257) );
  AOI22_X1 U10553 ( .A1(n9255), .A2(n9254), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9253), .ZN(n9256) );
  OAI211_X1 U10554 ( .C1(n9259), .C2(n9258), .A(n9257), .B(n9256), .ZN(n9260)
         );
  AOI21_X1 U10555 ( .B1(n9344), .B2(n9276), .A(n9260), .ZN(n9261) );
  OAI21_X1 U10556 ( .B1(n9348), .B2(n9262), .A(n9261), .ZN(P1_U3271) );
  XNOR2_X1 U10557 ( .A(n9263), .B(n9281), .ZN(n9264) );
  OAI222_X1 U10558 ( .A1(n9269), .A2(n9268), .B1(n9267), .B2(n9266), .C1(n9265), .C2(n9264), .ZN(n9665) );
  INV_X1 U10559 ( .A(n9270), .ZN(n9271) );
  OAI211_X1 U10560 ( .C1(n9663), .C2(n9272), .A(n9271), .B(n9366), .ZN(n9661)
         );
  OAI22_X1 U10561 ( .A1(n9661), .A2(n9275), .B1(n9274), .B2(n9273), .ZN(n9277)
         );
  OAI21_X1 U10562 ( .B1(n9665), .B2(n9277), .A(n9276), .ZN(n9286) );
  AOI22_X1 U10563 ( .A1(n9280), .A2(n9279), .B1(n9278), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n9285) );
  OR2_X1 U10564 ( .A1(n9282), .A2(n9281), .ZN(n9660) );
  NAND2_X1 U10565 ( .A1(n9282), .A2(n9281), .ZN(n9659) );
  NAND3_X1 U10566 ( .A1(n9660), .A2(n9659), .A3(n9283), .ZN(n9284) );
  NAND3_X1 U10567 ( .A1(n9286), .A2(n9285), .A3(n9284), .ZN(P1_U3286) );
  NAND2_X1 U10568 ( .A1(n9287), .A2(n9443), .ZN(n9288) );
  MUX2_X1 U10569 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9378), .S(n9707), .Z(
        P1_U3554) );
  NAND3_X1 U10570 ( .A1(n9291), .A2(n9366), .A3(n9290), .ZN(n9293) );
  OAI211_X1 U10571 ( .C1(n9294), .C2(n9686), .A(n9293), .B(n9292), .ZN(n9379)
         );
  MUX2_X1 U10572 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9379), .S(n9707), .Z(
        P1_U3553) );
  NAND2_X1 U10573 ( .A1(n9295), .A2(n9377), .ZN(n9682) );
  NAND2_X1 U10574 ( .A1(n9296), .A2(n9682), .ZN(n9300) );
  MUX2_X1 U10575 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9380), .S(n9707), .Z(
        P1_U3552) );
  INV_X1 U10576 ( .A(n9682), .ZN(n9363) );
  OAI21_X1 U10577 ( .B1(n9305), .B2(n9363), .A(n9304), .ZN(n9381) );
  MUX2_X1 U10578 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9381), .S(n9707), .Z(
        P1_U3551) );
  AOI22_X1 U10579 ( .A1(n9307), .A2(n9366), .B1(n9443), .B2(n9306), .ZN(n9308)
         );
  OAI211_X1 U10580 ( .C1(n9310), .C2(n9363), .A(n9309), .B(n9308), .ZN(n9382)
         );
  MUX2_X1 U10581 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9382), .S(n9707), .Z(
        P1_U3550) );
  INV_X1 U10582 ( .A(n9311), .ZN(n9313) );
  AOI22_X1 U10583 ( .A1(n9313), .A2(n9366), .B1(n9443), .B2(n9312), .ZN(n9314)
         );
  OAI211_X1 U10584 ( .C1(n9316), .C2(n9363), .A(n9315), .B(n9314), .ZN(n9383)
         );
  MUX2_X1 U10585 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9383), .S(n9707), .Z(
        P1_U3549) );
  AOI22_X1 U10586 ( .A1(n9318), .A2(n9366), .B1(n9443), .B2(n9317), .ZN(n9319)
         );
  OAI211_X1 U10587 ( .C1(n9321), .C2(n9363), .A(n9320), .B(n9319), .ZN(n9384)
         );
  MUX2_X1 U10588 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9384), .S(n9707), .Z(
        P1_U3548) );
  NAND3_X1 U10589 ( .A1(n9323), .A2(n9322), .A3(n9682), .ZN(n9328) );
  NAND2_X1 U10590 ( .A1(n9324), .A2(n9443), .ZN(n9325) );
  NAND4_X1 U10591 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), .ZN(n9385)
         );
  MUX2_X1 U10592 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9385), .S(n9707), .Z(
        P1_U3547) );
  AOI211_X1 U10593 ( .C1(n9443), .C2(n9331), .A(n9330), .B(n9329), .ZN(n9332)
         );
  OAI21_X1 U10594 ( .B1(n9333), .B2(n9363), .A(n9332), .ZN(n9386) );
  MUX2_X1 U10595 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9386), .S(n9707), .Z(
        P1_U3546) );
  AOI22_X1 U10596 ( .A1(n9335), .A2(n9366), .B1(n9443), .B2(n9334), .ZN(n9336)
         );
  OAI211_X1 U10597 ( .C1(n9338), .C2(n9363), .A(n9337), .B(n9336), .ZN(n9387)
         );
  MUX2_X1 U10598 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9387), .S(n9707), .Z(
        P1_U3545) );
  AOI211_X1 U10599 ( .C1(n9443), .C2(n9341), .A(n9340), .B(n9339), .ZN(n9342)
         );
  OAI21_X1 U10600 ( .B1(n9343), .B2(n9363), .A(n9342), .ZN(n9388) );
  MUX2_X1 U10601 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9388), .S(n9707), .Z(
        P1_U3544) );
  AOI211_X1 U10602 ( .C1(n9443), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9347)
         );
  OAI21_X1 U10603 ( .B1(n9348), .B2(n9363), .A(n9347), .ZN(n9389) );
  MUX2_X1 U10604 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9389), .S(n9707), .Z(
        P1_U3543) );
  AOI211_X1 U10605 ( .C1(n9443), .C2(n9351), .A(n9350), .B(n9349), .ZN(n9352)
         );
  OAI21_X1 U10606 ( .B1(n9353), .B2(n9363), .A(n9352), .ZN(n9390) );
  MUX2_X1 U10607 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9390), .S(n9707), .Z(
        P1_U3542) );
  AOI211_X1 U10608 ( .C1(n9443), .C2(n9356), .A(n9355), .B(n9354), .ZN(n9357)
         );
  OAI21_X1 U10609 ( .B1(n9358), .B2(n9363), .A(n9357), .ZN(n9391) );
  MUX2_X1 U10610 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9391), .S(n9707), .Z(
        P1_U3541) );
  AOI22_X1 U10611 ( .A1(n9360), .A2(n9366), .B1(n9443), .B2(n9359), .ZN(n9361)
         );
  OAI211_X1 U10612 ( .C1(n9364), .C2(n9363), .A(n9362), .B(n9361), .ZN(n9392)
         );
  MUX2_X1 U10613 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9392), .S(n9707), .Z(
        P1_U3540) );
  AOI22_X1 U10614 ( .A1(n9367), .A2(n9366), .B1(n9443), .B2(n9365), .ZN(n9368)
         );
  OAI211_X1 U10615 ( .C1(n9370), .C2(n9377), .A(n9369), .B(n9368), .ZN(n9393)
         );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9393), .S(n9707), .Z(
        P1_U3538) );
  OAI22_X1 U10617 ( .A1(n9372), .A2(n9688), .B1(n9371), .B2(n9686), .ZN(n9373)
         );
  INV_X1 U10618 ( .A(n9373), .ZN(n9374) );
  OAI211_X1 U10619 ( .C1(n9377), .C2(n9376), .A(n9375), .B(n9374), .ZN(n9394)
         );
  MUX2_X1 U10620 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9394), .S(n9707), .Z(
        P1_U3536) );
  MUX2_X1 U10621 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9379), .S(n9696), .Z(
        P1_U3521) );
  MUX2_X1 U10622 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9381), .S(n9696), .Z(
        P1_U3519) );
  MUX2_X1 U10623 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9382), .S(n9696), .Z(
        P1_U3518) );
  MUX2_X1 U10624 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9383), .S(n9696), .Z(
        P1_U3517) );
  MUX2_X1 U10625 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9384), .S(n9696), .Z(
        P1_U3516) );
  MUX2_X1 U10626 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9385), .S(n9696), .Z(
        P1_U3515) );
  MUX2_X1 U10627 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9386), .S(n9696), .Z(
        P1_U3514) );
  MUX2_X1 U10628 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9387), .S(n9696), .Z(
        P1_U3513) );
  MUX2_X1 U10629 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9388), .S(n9696), .Z(
        P1_U3512) );
  MUX2_X1 U10630 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9389), .S(n9696), .Z(
        P1_U3511) );
  MUX2_X1 U10631 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9390), .S(n9696), .Z(
        P1_U3510) );
  MUX2_X1 U10632 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9391), .S(n9696), .Z(
        P1_U3508) );
  MUX2_X1 U10633 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9392), .S(n9696), .Z(
        P1_U3505) );
  MUX2_X1 U10634 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9393), .S(n9696), .Z(
        P1_U3499) );
  MUX2_X1 U10635 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9394), .S(n9696), .Z(
        P1_U3493) );
  MUX2_X1 U10636 ( .A(P1_D_REG_0__SCAN_IN), .B(n9395), .S(n9633), .Z(P1_U3440)
         );
  MUX2_X1 U10637 ( .A(n9396), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NAND2_X1 U10638 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9398) );
  AOI21_X1 U10639 ( .B1(n9399), .B2(n9398), .A(n9397), .ZN(n9400) );
  NAND2_X1 U10640 ( .A1(n9710), .A2(n9400), .ZN(n9405) );
  OAI22_X1 U10641 ( .A1(n9402), .A2(n9878), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9401), .ZN(n9403) );
  INV_X1 U10642 ( .A(n9403), .ZN(n9404) );
  OAI211_X1 U10643 ( .C1(n9711), .C2(n9406), .A(n9405), .B(n9404), .ZN(n9407)
         );
  INV_X1 U10644 ( .A(n9407), .ZN(n9413) );
  NOR2_X1 U10645 ( .A1(n10016), .A2(n9408), .ZN(n9411) );
  OAI211_X1 U10646 ( .C1(n9411), .C2(n9410), .A(n9708), .B(n9409), .ZN(n9412)
         );
  NAND2_X1 U10647 ( .A1(n9413), .A2(n9412), .ZN(P2_U3246) );
  AOI22_X1 U10648 ( .A1(n9715), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9426) );
  AOI211_X1 U10649 ( .C1(n9417), .C2(n9416), .A(n9415), .B(n9414), .ZN(n9418)
         );
  AOI21_X1 U10650 ( .B1(n9420), .B2(n9419), .A(n9418), .ZN(n9425) );
  OAI211_X1 U10651 ( .C1(n9423), .C2(n9422), .A(n9708), .B(n9421), .ZN(n9424)
         );
  NAND3_X1 U10652 ( .A1(n9426), .A2(n9425), .A3(n9424), .ZN(P2_U3247) );
  OAI21_X1 U10653 ( .B1(n9428), .B2(n9686), .A(n9427), .ZN(n9429) );
  AOI21_X1 U10654 ( .B1(n9430), .B2(n9693), .A(n9429), .ZN(n9431) );
  AND2_X1 U10655 ( .A1(n9432), .A2(n9431), .ZN(n9433) );
  AOI22_X1 U10656 ( .A1(n9696), .A2(n9433), .B1(n5289), .B2(n9694), .ZN(
        P1_U3484) );
  AOI22_X1 U10657 ( .A1(n9707), .A2(n9433), .B1(n5288), .B2(n9705), .ZN(
        P1_U3533) );
  NAND2_X1 U10658 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9541) );
  OAI21_X1 U10659 ( .B1(n9435), .B2(n9434), .A(n9541), .ZN(n9436) );
  AOI21_X1 U10660 ( .B1(n9438), .B2(n9437), .A(n9436), .ZN(n9450) );
  INV_X1 U10661 ( .A(n9439), .ZN(n9440) );
  AOI21_X1 U10662 ( .B1(n9442), .B2(n9441), .A(n9440), .ZN(n9447) );
  NAND2_X1 U10663 ( .A1(n9444), .A2(n9443), .ZN(n9489) );
  OAI22_X1 U10664 ( .A1(n9447), .A2(n9446), .B1(n9445), .B2(n9489), .ZN(n9448)
         );
  INV_X1 U10665 ( .A(n9448), .ZN(n9449) );
  OAI211_X1 U10666 ( .C1(n9452), .C2(n9451), .A(n9450), .B(n9449), .ZN(
        P1_U3222) );
  OAI22_X1 U10667 ( .A1(n9454), .A2(n9842), .B1(n9453), .B2(n9850), .ZN(n9456)
         );
  AOI211_X1 U10668 ( .C1(n9854), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9472)
         );
  INV_X1 U10669 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9458) );
  AOI22_X1 U10670 ( .A1(n9873), .A2(n9472), .B1(n9458), .B2(n9870), .ZN(
        P2_U3535) );
  NAND2_X1 U10671 ( .A1(n9459), .A2(n9824), .ZN(n9460) );
  OAI211_X1 U10672 ( .C1(n9842), .C2(n9462), .A(n9461), .B(n9460), .ZN(n9463)
         );
  AOI21_X1 U10673 ( .B1(n9464), .B2(n9854), .A(n9463), .ZN(n9474) );
  AOI22_X1 U10674 ( .A1(n9873), .A2(n9474), .B1(n10091), .B2(n9870), .ZN(
        P2_U3534) );
  INV_X1 U10675 ( .A(n9465), .ZN(n9470) );
  OAI22_X1 U10676 ( .A1(n9467), .A2(n9842), .B1(n9466), .B2(n9850), .ZN(n9469)
         );
  AOI211_X1 U10677 ( .C1(n9839), .C2(n9470), .A(n9469), .B(n9468), .ZN(n9476)
         );
  AOI22_X1 U10678 ( .A1(n9873), .A2(n9476), .B1(n9954), .B2(n9870), .ZN(
        P2_U3533) );
  INV_X1 U10679 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9471) );
  AOI22_X1 U10680 ( .A1(n9856), .A2(n9472), .B1(n9471), .B2(n9855), .ZN(
        P2_U3496) );
  INV_X1 U10681 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9473) );
  AOI22_X1 U10682 ( .A1(n9856), .A2(n9474), .B1(n9473), .B2(n9855), .ZN(
        P2_U3493) );
  INV_X1 U10683 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9475) );
  AOI22_X1 U10684 ( .A1(n9856), .A2(n9476), .B1(n9475), .B2(n9855), .ZN(
        P2_U3490) );
  OAI211_X1 U10685 ( .C1(n9479), .C2(n9686), .A(n9478), .B(n9477), .ZN(n9480)
         );
  AOI21_X1 U10686 ( .B1(n9481), .B2(n9682), .A(n9480), .ZN(n9495) );
  AOI22_X1 U10687 ( .A1(n9707), .A2(n9495), .B1(n9482), .B2(n9705), .ZN(
        P1_U3539) );
  OAI21_X1 U10688 ( .B1(n9484), .B2(n9686), .A(n9483), .ZN(n9485) );
  AOI211_X1 U10689 ( .C1(n9487), .C2(n9682), .A(n9486), .B(n9485), .ZN(n9497)
         );
  AOI22_X1 U10690 ( .A1(n9707), .A2(n9497), .B1(n5398), .B2(n9705), .ZN(
        P1_U3537) );
  NAND4_X1 U10691 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n9492)
         );
  AOI21_X1 U10692 ( .B1(n9493), .B2(n9682), .A(n9492), .ZN(n9498) );
  AOI22_X1 U10693 ( .A1(n9707), .A2(n9498), .B1(n9028), .B2(n9705), .ZN(
        P1_U3535) );
  INV_X1 U10694 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9494) );
  AOI22_X1 U10695 ( .A1(n9696), .A2(n9495), .B1(n9494), .B2(n9694), .ZN(
        P1_U3502) );
  INV_X1 U10696 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9496) );
  AOI22_X1 U10697 ( .A1(n9696), .A2(n9497), .B1(n9496), .B2(n9694), .ZN(
        P1_U3496) );
  AOI22_X1 U10698 ( .A1(n9696), .A2(n9498), .B1(n5350), .B2(n9694), .ZN(
        P1_U3490) );
  XNOR2_X1 U10699 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10700 ( .A(P1_RD_REG_SCAN_IN), .B(n4736), .Z(U126) );
  NAND4_X1 U10701 ( .A1(n9501), .A2(n9500), .A3(P1_REG1_REG_0__SCAN_IN), .A4(
        P1_STATE_REG_SCAN_IN), .ZN(n9502) );
  NAND2_X1 U10702 ( .A1(n4487), .A2(n9502), .ZN(n9504) );
  AOI22_X1 U10703 ( .A1(n9571), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9504), .B2(
        n9503), .ZN(n9506) );
  NAND3_X1 U10704 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(n9625), .A3(n5011), .ZN(
        n9505) );
  OAI211_X1 U10705 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6542), .A(n9506), .B(
        n9505), .ZN(P1_U3241) );
  AOI21_X1 U10706 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9522) );
  NAND2_X1 U10707 ( .A1(n9571), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n9519) );
  INV_X1 U10708 ( .A(n9510), .ZN(n9515) );
  AOI21_X1 U10709 ( .B1(n9513), .B2(n9512), .A(n9511), .ZN(n9514) );
  OAI21_X1 U10710 ( .B1(n9515), .B2(n9514), .A(n9619), .ZN(n9518) );
  NAND2_X1 U10711 ( .A1(n9621), .A2(n9516), .ZN(n9517) );
  AND3_X1 U10712 ( .A1(n9519), .A2(n9518), .A3(n9517), .ZN(n9521) );
  OAI211_X1 U10713 ( .C1(n9522), .C2(n9575), .A(n9521), .B(n9520), .ZN(
        P1_U3248) );
  NAND2_X1 U10714 ( .A1(n9531), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9523) );
  OAI22_X1 U10715 ( .A1(n9533), .A2(n9525), .B1(n9524), .B2(n9523), .ZN(n9530)
         );
  OAI21_X1 U10716 ( .B1(n9528), .B2(n9527), .A(n9526), .ZN(n9529) );
  AOI22_X1 U10717 ( .A1(n9530), .A2(n9625), .B1(n9619), .B2(n9529), .ZN(n9537)
         );
  AOI22_X1 U10718 ( .A1(n9571), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9531), .B2(
        n9621), .ZN(n9536) );
  NAND3_X1 U10719 ( .A1(n9625), .A2(n9533), .A3(n9532), .ZN(n9534) );
  NAND4_X1 U10720 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), .ZN(
        P1_U3249) );
  AOI21_X1 U10721 ( .B1(n9540), .B2(n9539), .A(n9538), .ZN(n9550) );
  INV_X1 U10722 ( .A(n9541), .ZN(n9542) );
  AOI21_X1 U10723 ( .B1(n9621), .B2(n9543), .A(n9542), .ZN(n9549) );
  OAI211_X1 U10724 ( .C1(n9545), .C2(n4410), .A(n9619), .B(n9544), .ZN(n9546)
         );
  INV_X1 U10725 ( .A(n9546), .ZN(n9547) );
  AOI21_X1 U10726 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n9571), .A(n9547), .ZN(
        n9548) );
  OAI211_X1 U10727 ( .C1(n9550), .C2(n9575), .A(n9549), .B(n9548), .ZN(
        P1_U3253) );
  INV_X1 U10728 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9563) );
  AOI21_X1 U10729 ( .B1(n9621), .B2(n9552), .A(n9551), .ZN(n9557) );
  OAI211_X1 U10730 ( .C1(n9555), .C2(n9554), .A(n9619), .B(n9553), .ZN(n9556)
         );
  AND2_X1 U10731 ( .A1(n9557), .A2(n9556), .ZN(n9562) );
  OAI221_X1 U10732 ( .B1(n9560), .B2(n9559), .C1(n9560), .C2(n9558), .A(n9625), 
        .ZN(n9561) );
  OAI211_X1 U10733 ( .C1(n9563), .C2(n9631), .A(n9562), .B(n9561), .ZN(
        P1_U3254) );
  AOI21_X1 U10734 ( .B1(n9566), .B2(n9565), .A(n9564), .ZN(n9576) );
  AOI21_X1 U10735 ( .B1(n9621), .B2(n9568), .A(n9567), .ZN(n9574) );
  OAI21_X1 U10736 ( .B1(n9570), .B2(n7447), .A(n9569), .ZN(n9572) );
  AOI22_X1 U10737 ( .A1(n9572), .A2(n9619), .B1(n9571), .B2(
        P1_ADDR_REG_14__SCAN_IN), .ZN(n9573) );
  OAI211_X1 U10738 ( .C1(n9576), .C2(n9575), .A(n9574), .B(n9573), .ZN(
        P1_U3255) );
  INV_X1 U10739 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9586) );
  AOI211_X1 U10740 ( .C1(n9578), .C2(n5432), .A(n9577), .B(n9587), .ZN(n9579)
         );
  AOI211_X1 U10741 ( .C1(n9621), .C2(n9581), .A(n9580), .B(n9579), .ZN(n9585)
         );
  OAI211_X1 U10742 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9583), .A(n9625), .B(
        n9582), .ZN(n9584) );
  OAI211_X1 U10743 ( .C1(n9586), .C2(n9631), .A(n9585), .B(n9584), .ZN(
        P1_U3256) );
  INV_X1 U10744 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9599) );
  AOI211_X1 U10745 ( .C1(n9590), .C2(n9589), .A(n9588), .B(n9587), .ZN(n9591)
         );
  AOI211_X1 U10746 ( .C1(n9621), .C2(n9593), .A(n9592), .B(n9591), .ZN(n9598)
         );
  OAI211_X1 U10747 ( .C1(n9596), .C2(n9595), .A(n9625), .B(n9594), .ZN(n9597)
         );
  OAI211_X1 U10748 ( .C1(n9599), .C2(n9631), .A(n9598), .B(n9597), .ZN(
        P1_U3257) );
  INV_X1 U10749 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9613) );
  AOI21_X1 U10750 ( .B1(n9621), .B2(n9601), .A(n9600), .ZN(n9607) );
  AOI21_X1 U10751 ( .B1(n9604), .B2(n9603), .A(n9602), .ZN(n9605) );
  NAND2_X1 U10752 ( .A1(n9619), .A2(n9605), .ZN(n9606) );
  AND2_X1 U10753 ( .A1(n9607), .A2(n9606), .ZN(n9612) );
  OAI211_X1 U10754 ( .C1(n9610), .C2(n9609), .A(n9625), .B(n9608), .ZN(n9611)
         );
  OAI211_X1 U10755 ( .C1(n9613), .C2(n9631), .A(n9612), .B(n9611), .ZN(
        P1_U3258) );
  INV_X1 U10756 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U10757 ( .A1(n9615), .A2(n9614), .ZN(n9618) );
  INV_X1 U10758 ( .A(n9616), .ZN(n9617) );
  NAND3_X1 U10759 ( .A1(n9619), .A2(n9618), .A3(n9617), .ZN(n9624) );
  NAND2_X1 U10760 ( .A1(n9621), .A2(n9620), .ZN(n9623) );
  AND3_X1 U10761 ( .A1(n9624), .A2(n9623), .A3(n9622), .ZN(n9630) );
  OAI221_X1 U10762 ( .B1(n9628), .B2(n9627), .C1(n9628), .C2(n9626), .A(n9625), 
        .ZN(n9629) );
  OAI211_X1 U10763 ( .C1(n10218), .C2(n9631), .A(n9630), .B(n9629), .ZN(
        P1_U3259) );
  INV_X1 U10764 ( .A(n9632), .ZN(n9634) );
  AND2_X1 U10765 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  INV_X1 U10766 ( .A(n9635), .ZN(n9636) );
  AND2_X1 U10767 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9636), .ZN(P1_U3292) );
  AND2_X1 U10768 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9636), .ZN(P1_U3293) );
  AND2_X1 U10769 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9636), .ZN(P1_U3294) );
  AND2_X1 U10770 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9636), .ZN(P1_U3295) );
  NOR2_X1 U10771 ( .A1(n9635), .A2(n10105), .ZN(P1_U3296) );
  AND2_X1 U10772 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9636), .ZN(P1_U3297) );
  INV_X1 U10773 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9970) );
  NOR2_X1 U10774 ( .A1(n9635), .A2(n9970), .ZN(P1_U3298) );
  AND2_X1 U10775 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9636), .ZN(P1_U3299) );
  AND2_X1 U10776 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9636), .ZN(P1_U3300) );
  AND2_X1 U10777 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9636), .ZN(P1_U3301) );
  AND2_X1 U10778 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9636), .ZN(P1_U3302) );
  NOR2_X1 U10779 ( .A1(n9635), .A2(n9916), .ZN(P1_U3303) );
  AND2_X1 U10780 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9636), .ZN(P1_U3304) );
  AND2_X1 U10781 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9636), .ZN(P1_U3305) );
  AND2_X1 U10782 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9636), .ZN(P1_U3306) );
  NOR2_X1 U10783 ( .A1(n9635), .A2(n9914), .ZN(P1_U3307) );
  AND2_X1 U10784 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9636), .ZN(P1_U3308) );
  AND2_X1 U10785 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9636), .ZN(P1_U3309) );
  AND2_X1 U10786 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9636), .ZN(P1_U3310) );
  AND2_X1 U10787 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9636), .ZN(P1_U3311) );
  AND2_X1 U10788 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9636), .ZN(P1_U3312) );
  AND2_X1 U10789 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9636), .ZN(P1_U3313) );
  AND2_X1 U10790 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9636), .ZN(P1_U3314) );
  AND2_X1 U10791 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9636), .ZN(P1_U3315) );
  AND2_X1 U10792 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9636), .ZN(P1_U3316) );
  AND2_X1 U10793 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9636), .ZN(P1_U3317) );
  NOR2_X1 U10794 ( .A1(n9635), .A2(n9921), .ZN(P1_U3318) );
  AND2_X1 U10795 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9636), .ZN(P1_U3319) );
  AND2_X1 U10796 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9636), .ZN(P1_U3320) );
  AND2_X1 U10797 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9636), .ZN(P1_U3321) );
  INV_X1 U10798 ( .A(n9637), .ZN(n9643) );
  INV_X1 U10799 ( .A(n9638), .ZN(n9639) );
  OAI21_X1 U10800 ( .B1(n9640), .B2(n9686), .A(n9639), .ZN(n9642) );
  AOI211_X1 U10801 ( .C1(n9693), .C2(n9643), .A(n9642), .B(n9641), .ZN(n9697)
         );
  AOI22_X1 U10802 ( .A1(n9696), .A2(n9697), .B1(n5019), .B2(n9694), .ZN(
        P1_U3457) );
  INV_X1 U10803 ( .A(n9644), .ZN(n9649) );
  OAI22_X1 U10804 ( .A1(n9646), .A2(n9688), .B1(n9645), .B2(n9686), .ZN(n9648)
         );
  AOI211_X1 U10805 ( .C1(n9693), .C2(n9649), .A(n9648), .B(n9647), .ZN(n9698)
         );
  AOI22_X1 U10806 ( .A1(n9696), .A2(n9698), .B1(n5037), .B2(n9694), .ZN(
        P1_U3460) );
  INV_X1 U10807 ( .A(n9650), .ZN(n9654) );
  OAI22_X1 U10808 ( .A1(n9651), .A2(n9688), .B1(n6926), .B2(n9686), .ZN(n9653)
         );
  AOI211_X1 U10809 ( .C1(n9693), .C2(n9654), .A(n9653), .B(n9652), .ZN(n9699)
         );
  AOI22_X1 U10810 ( .A1(n9696), .A2(n9699), .B1(n5068), .B2(n9694), .ZN(
        P1_U3463) );
  OAI22_X1 U10811 ( .A1(n9655), .A2(n9688), .B1(n6931), .B2(n9686), .ZN(n9657)
         );
  AOI211_X1 U10812 ( .C1(n9693), .C2(n9658), .A(n9657), .B(n9656), .ZN(n9700)
         );
  AOI22_X1 U10813 ( .A1(n9696), .A2(n9700), .B1(n5099), .B2(n9694), .ZN(
        P1_U3466) );
  NAND3_X1 U10814 ( .A1(n9660), .A2(n9659), .A3(n9682), .ZN(n9662) );
  OAI211_X1 U10815 ( .C1(n9663), .C2(n9686), .A(n9662), .B(n9661), .ZN(n9664)
         );
  NOR2_X1 U10816 ( .A1(n9665), .A2(n9664), .ZN(n9701) );
  INV_X1 U10817 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9666) );
  AOI22_X1 U10818 ( .A1(n9696), .A2(n9701), .B1(n9666), .B2(n9694), .ZN(
        P1_U3469) );
  OAI22_X1 U10819 ( .A1(n9668), .A2(n9688), .B1(n9667), .B2(n9686), .ZN(n9670)
         );
  AOI211_X1 U10820 ( .C1(n9693), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9702)
         );
  INV_X1 U10821 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U10822 ( .A1(n9696), .A2(n9702), .B1(n9672), .B2(n9694), .ZN(
        P1_U3472) );
  NAND2_X1 U10823 ( .A1(n9674), .A2(n9673), .ZN(n9676) );
  AOI211_X1 U10824 ( .C1(n9682), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9703)
         );
  INV_X1 U10825 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U10826 ( .A1(n9696), .A2(n9703), .B1(n9983), .B2(n9694), .ZN(
        P1_U3475) );
  OAI21_X1 U10827 ( .B1(n9679), .B2(n9688), .A(n9678), .ZN(n9680) );
  AOI211_X1 U10828 ( .C1(n9683), .C2(n9682), .A(n9681), .B(n9680), .ZN(n9704)
         );
  INV_X1 U10829 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9684) );
  AOI22_X1 U10830 ( .A1(n9696), .A2(n9704), .B1(n9684), .B2(n9694), .ZN(
        P1_U3478) );
  INV_X1 U10831 ( .A(n9685), .ZN(n9692) );
  OAI22_X1 U10832 ( .A1(n9689), .A2(n9688), .B1(n9687), .B2(n9686), .ZN(n9691)
         );
  AOI211_X1 U10833 ( .C1(n9693), .C2(n9692), .A(n9691), .B(n9690), .ZN(n9706)
         );
  INV_X1 U10834 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U10835 ( .A1(n9696), .A2(n9706), .B1(n9695), .B2(n9694), .ZN(
        P1_U3481) );
  AOI22_X1 U10836 ( .A1(n9707), .A2(n9697), .B1(n6324), .B2(n9705), .ZN(
        P1_U3524) );
  AOI22_X1 U10837 ( .A1(n9707), .A2(n9698), .B1(n6323), .B2(n9705), .ZN(
        P1_U3525) );
  AOI22_X1 U10838 ( .A1(n9707), .A2(n9699), .B1(n6327), .B2(n9705), .ZN(
        P1_U3526) );
  AOI22_X1 U10839 ( .A1(n9707), .A2(n9700), .B1(n5098), .B2(n9705), .ZN(
        P1_U3527) );
  AOI22_X1 U10840 ( .A1(n9707), .A2(n9701), .B1(n5130), .B2(n9705), .ZN(
        P1_U3528) );
  AOI22_X1 U10841 ( .A1(n9707), .A2(n9702), .B1(n6335), .B2(n9705), .ZN(
        P1_U3529) );
  AOI22_X1 U10842 ( .A1(n9707), .A2(n9703), .B1(n5191), .B2(n9705), .ZN(
        P1_U3530) );
  AOI22_X1 U10843 ( .A1(n9707), .A2(n9704), .B1(n5217), .B2(n9705), .ZN(
        P1_U3531) );
  AOI22_X1 U10844 ( .A1(n9707), .A2(n9706), .B1(n5243), .B2(n9705), .ZN(
        P1_U3532) );
  AOI22_X1 U10845 ( .A1(n9710), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9708), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U10846 ( .A1(n9710), .A2(n9709), .ZN(n9712) );
  OAI211_X1 U10847 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9713), .A(n9712), .B(
        n9711), .ZN(n9714) );
  INV_X1 U10848 ( .A(n9714), .ZN(n9717) );
  AOI22_X1 U10849 ( .A1(n9715), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9716) );
  OAI221_X1 U10850 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9718), .C1(n10016), .C2(
        n9717), .A(n9716), .ZN(P2_U3245) );
  INV_X1 U10851 ( .A(n9722), .ZN(n9739) );
  INV_X1 U10852 ( .A(n9719), .ZN(n9723) );
  INV_X1 U10853 ( .A(n9720), .ZN(n9721) );
  NOR3_X1 U10854 ( .A1(n9723), .A2(n9722), .A3(n9721), .ZN(n9724) );
  AOI211_X1 U10855 ( .C1(n9726), .C2(n9739), .A(n9725), .B(n9724), .ZN(n9729)
         );
  AOI21_X1 U10856 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9849) );
  AOI222_X1 U10857 ( .A1(n9732), .A2(n9731), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n9773), .C1(n9771), .C2(n9730), .ZN(n9748) );
  OR2_X1 U10858 ( .A1(n7454), .A2(n9733), .ZN(n9735) );
  NAND2_X1 U10859 ( .A1(n9735), .A2(n9734), .ZN(n9740) );
  AND2_X1 U10860 ( .A1(n9737), .A2(n9736), .ZN(n9738) );
  OAI21_X1 U10861 ( .B1(n9740), .B2(n9739), .A(n9738), .ZN(n9853) );
  INV_X1 U10862 ( .A(n9741), .ZN(n9743) );
  OAI211_X1 U10863 ( .C1(n9743), .C2(n9851), .A(n6266), .B(n9742), .ZN(n9848)
         );
  INV_X1 U10864 ( .A(n9848), .ZN(n9744) );
  AOI22_X1 U10865 ( .A1(n9853), .A2(n9746), .B1(n9745), .B2(n9744), .ZN(n9747)
         );
  OAI211_X1 U10866 ( .C1(n9749), .C2(n9849), .A(n9748), .B(n9747), .ZN(
        P2_U3284) );
  NAND2_X1 U10867 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  NAND2_X1 U10868 ( .A1(n9753), .A2(n9752), .ZN(n9817) );
  AND2_X1 U10869 ( .A1(n9754), .A2(n9770), .ZN(n9756) );
  OR2_X1 U10870 ( .A1(n9756), .A2(n9755), .ZN(n9818) );
  OAI22_X1 U10871 ( .A1(n9817), .A2(n9758), .B1(n9757), .B2(n9818), .ZN(n9759)
         );
  INV_X1 U10872 ( .A(n9759), .ZN(n9778) );
  XNOR2_X1 U10873 ( .A(n9760), .B(n7317), .ZN(n9767) );
  OAI22_X1 U10874 ( .A1(n9764), .A2(n9763), .B1(n9762), .B2(n9761), .ZN(n9765)
         );
  AOI21_X1 U10875 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9768) );
  OAI21_X1 U10876 ( .B1(n9817), .B2(n9769), .A(n9768), .ZN(n9819) );
  AOI22_X1 U10877 ( .A1(n9773), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n9772), .B2(
        n9771), .ZN(n9774) );
  OAI21_X1 U10878 ( .B1(n9775), .B2(n4629), .A(n9774), .ZN(n9776) );
  AOI21_X1 U10879 ( .B1(n9819), .B2(n7202), .A(n9776), .ZN(n9777) );
  NAND2_X1 U10880 ( .A1(n9778), .A2(n9777), .ZN(P2_U3288) );
  NOR2_X1 U10881 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  AND2_X1 U10882 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9903), .ZN(P2_U3297) );
  AND2_X1 U10883 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9903), .ZN(P2_U3299) );
  INV_X1 U10884 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U10885 ( .A1(n9781), .A2(n9955), .ZN(P2_U3300) );
  INV_X1 U10886 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U10887 ( .A1(n9781), .A2(n9996), .ZN(P2_U3301) );
  AND2_X1 U10888 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9903), .ZN(P2_U3302) );
  INV_X1 U10889 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10010) );
  NOR2_X1 U10890 ( .A1(n9781), .A2(n10010), .ZN(P2_U3303) );
  AND2_X1 U10891 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9903), .ZN(P2_U3304) );
  AND2_X1 U10892 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9903), .ZN(P2_U3305) );
  AND2_X1 U10893 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9903), .ZN(P2_U3306) );
  INV_X1 U10894 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U10895 ( .A1(n9781), .A2(n10055), .ZN(P2_U3307) );
  AND2_X1 U10896 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9903), .ZN(P2_U3308) );
  AND2_X1 U10897 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9903), .ZN(P2_U3309) );
  INV_X1 U10898 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9957) );
  NOR2_X1 U10899 ( .A1(n9781), .A2(n9957), .ZN(P2_U3310) );
  INV_X1 U10900 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U10901 ( .A1(n9781), .A2(n10014), .ZN(P2_U3311) );
  AND2_X1 U10902 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9903), .ZN(P2_U3312) );
  AND2_X1 U10903 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9903), .ZN(P2_U3313) );
  AND2_X1 U10904 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9903), .ZN(P2_U3314) );
  AND2_X1 U10905 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9903), .ZN(P2_U3315) );
  INV_X1 U10906 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10065) );
  NOR2_X1 U10907 ( .A1(n9781), .A2(n10065), .ZN(P2_U3316) );
  AND2_X1 U10908 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9903), .ZN(P2_U3317) );
  AND2_X1 U10909 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9903), .ZN(P2_U3318) );
  INV_X1 U10910 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U10911 ( .A1(n9781), .A2(n9925), .ZN(P2_U3319) );
  AND2_X1 U10912 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9903), .ZN(P2_U3320) );
  AND2_X1 U10913 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9903), .ZN(P2_U3321) );
  INV_X1 U10914 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U10915 ( .A1(n9781), .A2(n9949), .ZN(P2_U3322) );
  AND2_X1 U10916 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9903), .ZN(P2_U3323) );
  AND2_X1 U10917 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9903), .ZN(P2_U3324) );
  INV_X1 U10918 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U10919 ( .A1(n9781), .A2(n10044), .ZN(P2_U3325) );
  AND2_X1 U10920 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9903), .ZN(P2_U3326) );
  AOI22_X1 U10921 ( .A1(n9785), .A2(n9782), .B1(n10082), .B2(n9903), .ZN(
        P2_U3437) );
  AOI22_X1 U10922 ( .A1(n9785), .A2(n9784), .B1(n9783), .B2(n9903), .ZN(
        P2_U3438) );
  OAI22_X1 U10923 ( .A1(n9787), .A2(n9842), .B1(n9786), .B2(n9850), .ZN(n9789)
         );
  AOI211_X1 U10924 ( .C1(n9854), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9857)
         );
  INV_X1 U10925 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U10926 ( .A1(n9856), .A2(n9857), .B1(n10052), .B2(n9855), .ZN(
        P2_U3457) );
  OAI21_X1 U10927 ( .B1(n9792), .B2(n9850), .A(n9791), .ZN(n9794) );
  AOI211_X1 U10928 ( .C1(n9854), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9858)
         );
  INV_X1 U10929 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9796) );
  AOI22_X1 U10930 ( .A1(n9856), .A2(n9858), .B1(n9796), .B2(n9855), .ZN(
        P2_U3463) );
  OAI211_X1 U10931 ( .C1(n9799), .C2(n9850), .A(n9798), .B(n9797), .ZN(n9800)
         );
  AOI21_X1 U10932 ( .B1(n9854), .B2(n9801), .A(n9800), .ZN(n9859) );
  INV_X1 U10933 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10066) );
  AOI22_X1 U10934 ( .A1(n9856), .A2(n9859), .B1(n10066), .B2(n9855), .ZN(
        P2_U3466) );
  AND3_X1 U10935 ( .A1(n9803), .A2(n9854), .A3(n9802), .ZN(n9808) );
  OAI211_X1 U10936 ( .C1(n9806), .C2(n9850), .A(n9805), .B(n9804), .ZN(n9807)
         );
  NOR2_X1 U10937 ( .A1(n9808), .A2(n9807), .ZN(n9861) );
  INV_X1 U10938 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9809) );
  AOI22_X1 U10939 ( .A1(n9856), .A2(n9861), .B1(n9809), .B2(n9855), .ZN(
        P2_U3469) );
  INV_X1 U10940 ( .A(n9810), .ZN(n9811) );
  OAI22_X1 U10941 ( .A1(n9812), .A2(n9842), .B1(n9811), .B2(n9850), .ZN(n9814)
         );
  AOI211_X1 U10942 ( .C1(n9854), .C2(n9815), .A(n9814), .B(n9813), .ZN(n9862)
         );
  INV_X1 U10943 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9816) );
  AOI22_X1 U10944 ( .A1(n9856), .A2(n9862), .B1(n9816), .B2(n9855), .ZN(
        P2_U3472) );
  INV_X1 U10945 ( .A(n9817), .ZN(n9821) );
  OAI22_X1 U10946 ( .A1(n9818), .A2(n9842), .B1(n4629), .B2(n9850), .ZN(n9820)
         );
  AOI211_X1 U10947 ( .C1(n9839), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9864)
         );
  INV_X1 U10948 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U10949 ( .A1(n9856), .A2(n9864), .B1(n10056), .B2(n9855), .ZN(
        P2_U3475) );
  INV_X1 U10950 ( .A(n9828), .ZN(n9830) );
  AOI21_X1 U10951 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9825) );
  OAI211_X1 U10952 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9829)
         );
  AOI21_X1 U10953 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9866) );
  INV_X1 U10954 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U10955 ( .A1(n9856), .A2(n9866), .B1(n9832), .B2(n9855), .ZN(
        P2_U3478) );
  INV_X1 U10956 ( .A(n9833), .ZN(n9838) );
  OAI22_X1 U10957 ( .A1(n9835), .A2(n9842), .B1(n9834), .B2(n9850), .ZN(n9837)
         );
  AOI211_X1 U10958 ( .C1(n9839), .C2(n9838), .A(n9837), .B(n9836), .ZN(n9868)
         );
  INV_X1 U10959 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U10960 ( .A1(n9856), .A2(n9868), .B1(n9840), .B2(n9855), .ZN(
        P2_U3481) );
  OAI22_X1 U10961 ( .A1(n9843), .A2(n9842), .B1(n9841), .B2(n9850), .ZN(n9845)
         );
  AOI211_X1 U10962 ( .C1(n9846), .C2(n9854), .A(n9845), .B(n9844), .ZN(n9869)
         );
  INV_X1 U10963 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9847) );
  AOI22_X1 U10964 ( .A1(n9856), .A2(n9869), .B1(n9847), .B2(n9855), .ZN(
        P2_U3484) );
  OAI211_X1 U10965 ( .C1(n9851), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9852)
         );
  AOI21_X1 U10966 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9872) );
  INV_X1 U10967 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U10968 ( .A1(n9856), .A2(n9872), .B1(n10118), .B2(n9855), .ZN(
        P2_U3487) );
  AOI22_X1 U10969 ( .A1(n9873), .A2(n9857), .B1(n6580), .B2(n9870), .ZN(
        P2_U3522) );
  AOI22_X1 U10970 ( .A1(n9873), .A2(n9858), .B1(n6578), .B2(n9870), .ZN(
        P2_U3524) );
  AOI22_X1 U10971 ( .A1(n9873), .A2(n9859), .B1(n6577), .B2(n9870), .ZN(
        P2_U3525) );
  AOI22_X1 U10972 ( .A1(n9873), .A2(n9861), .B1(n9860), .B2(n9870), .ZN(
        P2_U3526) );
  AOI22_X1 U10973 ( .A1(n9873), .A2(n9862), .B1(n9967), .B2(n9870), .ZN(
        P2_U3527) );
  INV_X1 U10974 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9863) );
  AOI22_X1 U10975 ( .A1(n9873), .A2(n9864), .B1(n9863), .B2(n9870), .ZN(
        P2_U3528) );
  AOI22_X1 U10976 ( .A1(n9873), .A2(n9866), .B1(n9865), .B2(n9870), .ZN(
        P2_U3529) );
  AOI22_X1 U10977 ( .A1(n9873), .A2(n9868), .B1(n9867), .B2(n9870), .ZN(
        P2_U3530) );
  AOI22_X1 U10978 ( .A1(n9873), .A2(n9869), .B1(n7157), .B2(n9870), .ZN(
        P2_U3531) );
  AOI22_X1 U10979 ( .A1(n9873), .A2(n9872), .B1(n9871), .B2(n9870), .ZN(
        P2_U3532) );
  INV_X1 U10980 ( .A(n9874), .ZN(n9875) );
  NAND2_X1 U10981 ( .A1(n9876), .A2(n9875), .ZN(n9877) );
  XOR2_X1 U10982 ( .A(n9878), .B(n9877), .Z(ADD_1071_U5) );
  XOR2_X1 U10983 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10984 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(ADD_1071_U56) );
  OAI21_X1 U10985 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(ADD_1071_U57) );
  OAI21_X1 U10986 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(ADD_1071_U58) );
  OAI21_X1 U10987 ( .B1(n9890), .B2(n9889), .A(n9888), .ZN(ADD_1071_U59) );
  OAI21_X1 U10988 ( .B1(n9893), .B2(n9892), .A(n9891), .ZN(ADD_1071_U60) );
  OAI21_X1 U10989 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(ADD_1071_U61) );
  AOI21_X1 U10990 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(ADD_1071_U62) );
  AOI21_X1 U10991 ( .B1(n9902), .B2(n9901), .A(n9900), .ZN(ADD_1071_U63) );
  NAND2_X1 U10992 ( .A1(n9903), .A2(P2_D_REG_30__SCAN_IN), .ZN(n10209) );
  INV_X1 U10993 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U10994 ( .A1(n9906), .A2(keyinput70), .B1(keyinput40), .B2(n9905), 
        .ZN(n9904) );
  OAI221_X1 U10995 ( .B1(n9906), .B2(keyinput70), .C1(n9905), .C2(keyinput40), 
        .A(n9904), .ZN(n9911) );
  XNOR2_X1 U10996 ( .A(n9907), .B(keyinput32), .ZN(n9910) );
  XNOR2_X1 U10997 ( .A(n9908), .B(keyinput93), .ZN(n9909) );
  OR3_X1 U10998 ( .A1(n9911), .A2(n9910), .A3(n9909), .ZN(n9919) );
  AOI22_X1 U10999 ( .A1(n9914), .A2(keyinput78), .B1(keyinput48), .B2(n9913), 
        .ZN(n9912) );
  OAI221_X1 U11000 ( .B1(n9914), .B2(keyinput78), .C1(n9913), .C2(keyinput48), 
        .A(n9912), .ZN(n9918) );
  AOI22_X1 U11001 ( .A1(n9916), .A2(keyinput0), .B1(keyinput64), .B2(n7051), 
        .ZN(n9915) );
  OAI221_X1 U11002 ( .B1(n9916), .B2(keyinput0), .C1(n7051), .C2(keyinput64), 
        .A(n9915), .ZN(n9917) );
  NOR3_X1 U11003 ( .A1(n9919), .A2(n9918), .A3(n9917), .ZN(n9965) );
  AOI22_X1 U11004 ( .A1(n9921), .A2(keyinput2), .B1(keyinput42), .B2(n6579), 
        .ZN(n9920) );
  OAI221_X1 U11005 ( .B1(n9921), .B2(keyinput2), .C1(n6579), .C2(keyinput42), 
        .A(n9920), .ZN(n9932) );
  AOI22_X1 U11006 ( .A1(n9924), .A2(keyinput55), .B1(n9923), .B2(keyinput49), 
        .ZN(n9922) );
  OAI221_X1 U11007 ( .B1(n9924), .B2(keyinput55), .C1(n9923), .C2(keyinput49), 
        .A(n9922), .ZN(n9931) );
  XNOR2_X1 U11008 ( .A(n9925), .B(keyinput18), .ZN(n9930) );
  XNOR2_X1 U11009 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput106), .ZN(n9928)
         );
  XNOR2_X1 U11010 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput115), .ZN(n9927)
         );
  XNOR2_X1 U11011 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(keyinput26), .ZN(n9926)
         );
  NAND3_X1 U11012 ( .A1(n9928), .A2(n9927), .A3(n9926), .ZN(n9929) );
  NOR4_X1 U11013 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), .ZN(n9964)
         );
  AOI22_X1 U11014 ( .A1(n9934), .A2(keyinput22), .B1(keyinput1), .B2(n6957), 
        .ZN(n9933) );
  OAI221_X1 U11015 ( .B1(n9934), .B2(keyinput22), .C1(n6957), .C2(keyinput1), 
        .A(n9933), .ZN(n9946) );
  INV_X1 U11016 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U11017 ( .A1(n9937), .A2(keyinput67), .B1(n9936), .B2(keyinput66), 
        .ZN(n9935) );
  OAI221_X1 U11018 ( .B1(n9937), .B2(keyinput67), .C1(n9936), .C2(keyinput66), 
        .A(n9935), .ZN(n9945) );
  AOI22_X1 U11019 ( .A1(n9940), .A2(keyinput86), .B1(n9938), .B2(keyinput30), 
        .ZN(n9939) );
  OAI221_X1 U11020 ( .B1(n9940), .B2(keyinput86), .C1(n9938), .C2(keyinput30), 
        .A(n9939), .ZN(n9944) );
  XNOR2_X1 U11021 ( .A(P2_REG0_REG_31__SCAN_IN), .B(keyinput21), .ZN(n9942) );
  XNOR2_X1 U11022 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput27), .ZN(n9941) );
  NAND2_X1 U11023 ( .A1(n9942), .A2(n9941), .ZN(n9943) );
  NOR4_X1 U11024 ( .A1(n9946), .A2(n9945), .A3(n9944), .A4(n9943), .ZN(n9963)
         );
  AOI22_X1 U11025 ( .A1(n9949), .A2(keyinput51), .B1(keyinput14), .B2(n9948), 
        .ZN(n9947) );
  OAI221_X1 U11026 ( .B1(n9949), .B2(keyinput51), .C1(n9948), .C2(keyinput14), 
        .A(n9947), .ZN(n9961) );
  AOI22_X1 U11027 ( .A1(n9952), .A2(keyinput17), .B1(n9951), .B2(keyinput124), 
        .ZN(n9950) );
  OAI221_X1 U11028 ( .B1(n9952), .B2(keyinput17), .C1(n9951), .C2(keyinput124), 
        .A(n9950), .ZN(n9960) );
  AOI22_X1 U11029 ( .A1(n9955), .A2(keyinput83), .B1(keyinput71), .B2(n9954), 
        .ZN(n9953) );
  OAI221_X1 U11030 ( .B1(n9955), .B2(keyinput83), .C1(n9954), .C2(keyinput71), 
        .A(n9953), .ZN(n9959) );
  AOI22_X1 U11031 ( .A1(n9047), .A2(keyinput35), .B1(keyinput99), .B2(n9957), 
        .ZN(n9956) );
  OAI221_X1 U11032 ( .B1(n9047), .B2(keyinput35), .C1(n9957), .C2(keyinput99), 
        .A(n9956), .ZN(n9958) );
  NOR4_X1 U11033 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9962)
         );
  NAND4_X1 U11034 ( .A1(n9965), .A2(n9964), .A3(n9963), .A4(n9962), .ZN(n10207) );
  AOI22_X1 U11035 ( .A1(n9968), .A2(keyinput88), .B1(keyinput8), .B2(n9967), 
        .ZN(n9966) );
  OAI221_X1 U11036 ( .B1(n9968), .B2(keyinput88), .C1(n9967), .C2(keyinput8), 
        .A(n9966), .ZN(n9980) );
  AOI22_X1 U11037 ( .A1(n6223), .A2(keyinput100), .B1(n9970), .B2(keyinput9), 
        .ZN(n9969) );
  OAI221_X1 U11038 ( .B1(n6223), .B2(keyinput100), .C1(n9970), .C2(keyinput9), 
        .A(n9969), .ZN(n9979) );
  AOI22_X1 U11039 ( .A1(n9973), .A2(keyinput109), .B1(keyinput77), .B2(n9972), 
        .ZN(n9971) );
  OAI221_X1 U11040 ( .B1(n9973), .B2(keyinput109), .C1(n9972), .C2(keyinput77), 
        .A(n9971), .ZN(n9978) );
  INV_X1 U11041 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9974) );
  XOR2_X1 U11042 ( .A(n9974), .B(keyinput7), .Z(n9976) );
  XNOR2_X1 U11043 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput94), .ZN(n9975) );
  NAND2_X1 U11044 ( .A1(n9976), .A2(n9975), .ZN(n9977) );
  NOR4_X1 U11045 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(n10028)
         );
  AOI22_X1 U11046 ( .A1(n9983), .A2(keyinput37), .B1(n9982), .B2(keyinput90), 
        .ZN(n9981) );
  OAI221_X1 U11047 ( .B1(n9983), .B2(keyinput37), .C1(n9982), .C2(keyinput90), 
        .A(n9981), .ZN(n9994) );
  AOI22_X1 U11048 ( .A1(n9986), .A2(keyinput95), .B1(n9985), .B2(keyinput50), 
        .ZN(n9984) );
  OAI221_X1 U11049 ( .B1(n9986), .B2(keyinput95), .C1(n9985), .C2(keyinput50), 
        .A(n9984), .ZN(n9993) );
  INV_X1 U11050 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U11051 ( .A1(P2_U3152), .A2(keyinput36), .B1(keyinput81), .B2(n9988), .ZN(n9987) );
  OAI221_X1 U11052 ( .B1(P2_U3152), .B2(keyinput36), .C1(n9988), .C2(
        keyinput81), .A(n9987), .ZN(n9992) );
  INV_X1 U11053 ( .A(SI_15_), .ZN(n9990) );
  AOI22_X1 U11054 ( .A1(n9990), .A2(keyinput45), .B1(keyinput52), .B2(n5350), 
        .ZN(n9989) );
  OAI221_X1 U11055 ( .B1(n9990), .B2(keyinput45), .C1(n5350), .C2(keyinput52), 
        .A(n9989), .ZN(n9991) );
  NOR4_X1 U11056 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n10027)
         );
  AOI22_X1 U11057 ( .A1(n9996), .A2(keyinput60), .B1(n7701), .B2(keyinput63), 
        .ZN(n9995) );
  OAI221_X1 U11058 ( .B1(n9996), .B2(keyinput60), .C1(n7701), .C2(keyinput63), 
        .A(n9995), .ZN(n10008) );
  INV_X1 U11059 ( .A(SI_31_), .ZN(n9999) );
  INV_X1 U11060 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9998) );
  AOI22_X1 U11061 ( .A1(n9999), .A2(keyinput92), .B1(keyinput97), .B2(n9998), 
        .ZN(n9997) );
  OAI221_X1 U11062 ( .B1(n9999), .B2(keyinput92), .C1(n9998), .C2(keyinput97), 
        .A(n9997), .ZN(n10007) );
  AOI22_X1 U11063 ( .A1(n6578), .A2(keyinput127), .B1(keyinput72), .B2(n10001), 
        .ZN(n10000) );
  OAI221_X1 U11064 ( .B1(n6578), .B2(keyinput127), .C1(n10001), .C2(keyinput72), .A(n10000), .ZN(n10006) );
  AOI22_X1 U11065 ( .A1(n10004), .A2(keyinput59), .B1(n10003), .B2(keyinput111), .ZN(n10002) );
  OAI221_X1 U11066 ( .B1(n10004), .B2(keyinput59), .C1(n10003), .C2(
        keyinput111), .A(n10002), .ZN(n10005) );
  NOR4_X1 U11067 ( .A1(n10008), .A2(n10007), .A3(n10006), .A4(n10005), .ZN(
        n10026) );
  AOI22_X1 U11068 ( .A1(n10011), .A2(keyinput89), .B1(keyinput87), .B2(n10010), 
        .ZN(n10009) );
  OAI221_X1 U11069 ( .B1(n10011), .B2(keyinput89), .C1(n10010), .C2(keyinput87), .A(n10009), .ZN(n10024) );
  INV_X1 U11070 ( .A(keyinput34), .ZN(n10013) );
  AOI22_X1 U11071 ( .A1(n10014), .A2(keyinput33), .B1(P2_WR_REG_SCAN_IN), .B2(
        n10013), .ZN(n10012) );
  OAI221_X1 U11072 ( .B1(n10014), .B2(keyinput33), .C1(n10013), .C2(
        P2_WR_REG_SCAN_IN), .A(n10012), .ZN(n10023) );
  AOI22_X1 U11073 ( .A1(n10017), .A2(keyinput15), .B1(keyinput53), .B2(n10016), 
        .ZN(n10015) );
  OAI221_X1 U11074 ( .B1(n10017), .B2(keyinput15), .C1(n10016), .C2(keyinput53), .A(n10015), .ZN(n10022) );
  INV_X1 U11075 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10020) );
  AOI22_X1 U11076 ( .A1(n10020), .A2(keyinput39), .B1(n10019), .B2(keyinput126), .ZN(n10018) );
  OAI221_X1 U11077 ( .B1(n10020), .B2(keyinput39), .C1(n10019), .C2(
        keyinput126), .A(n10018), .ZN(n10021) );
  NOR4_X1 U11078 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10025) );
  NAND4_X1 U11079 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(
        n10206) );
  AOI22_X1 U11080 ( .A1(n6316), .A2(keyinput47), .B1(keyinput80), .B2(n10030), 
        .ZN(n10029) );
  OAI221_X1 U11081 ( .B1(n6316), .B2(keyinput47), .C1(n10030), .C2(keyinput80), 
        .A(n10029), .ZN(n10038) );
  AOI22_X1 U11082 ( .A1(n5375), .A2(keyinput44), .B1(keyinput41), .B2(n6416), 
        .ZN(n10031) );
  OAI221_X1 U11083 ( .B1(n5375), .B2(keyinput44), .C1(n6416), .C2(keyinput41), 
        .A(n10031), .ZN(n10037) );
  XNOR2_X1 U11084 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput25), .ZN(n10035) );
  XNOR2_X1 U11085 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput19), .ZN(n10034)
         );
  XNOR2_X1 U11086 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput96), .ZN(n10033) );
  XNOR2_X1 U11087 ( .A(keyinput4), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n10032) );
  NAND4_X1 U11088 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n10036) );
  NOR3_X1 U11089 ( .A1(n10038), .A2(n10037), .A3(n10036), .ZN(n10204) );
  INV_X1 U11090 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11091 ( .A1(n10040), .A2(keyinput102), .B1(n9028), .B2(keyinput38), 
        .ZN(n10039) );
  OAI221_X1 U11092 ( .B1(n10040), .B2(keyinput102), .C1(n9028), .C2(keyinput38), .A(n10039), .ZN(n10050) );
  AOI22_X1 U11093 ( .A1(n5311), .A2(keyinput104), .B1(keyinput5), .B2(n6542), 
        .ZN(n10041) );
  OAI221_X1 U11094 ( .B1(n5311), .B2(keyinput104), .C1(n6542), .C2(keyinput5), 
        .A(n10041), .ZN(n10049) );
  INV_X1 U11095 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10043) );
  AOI22_X1 U11096 ( .A1(n10044), .A2(keyinput13), .B1(keyinput23), .B2(n10043), 
        .ZN(n10042) );
  OAI221_X1 U11097 ( .B1(n10044), .B2(keyinput13), .C1(n10043), .C2(keyinput23), .A(n10042), .ZN(n10048) );
  XNOR2_X1 U11098 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(keyinput3), .ZN(n10046)
         );
  XNOR2_X1 U11099 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput24), .ZN(n10045) );
  NAND2_X1 U11100 ( .A1(n10046), .A2(n10045), .ZN(n10047) );
  NOR4_X1 U11101 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10203) );
  AOI22_X1 U11102 ( .A1(n10053), .A2(keyinput73), .B1(keyinput69), .B2(n10052), 
        .ZN(n10051) );
  OAI221_X1 U11103 ( .B1(n10053), .B2(keyinput73), .C1(n10052), .C2(keyinput69), .A(n10051), .ZN(n10136) );
  AOI22_X1 U11104 ( .A1(n10056), .A2(keyinput120), .B1(n10055), .B2(
        keyinput113), .ZN(n10054) );
  OAI221_X1 U11105 ( .B1(n10056), .B2(keyinput120), .C1(n10055), .C2(
        keyinput113), .A(n10054), .ZN(n10135) );
  XOR2_X1 U11106 ( .A(P2_REG1_REG_26__SCAN_IN), .B(keyinput91), .Z(n10061) );
  INV_X1 U11107 ( .A(keyinput16), .ZN(n10057) );
  MUX2_X1 U11108 ( .A(keyinput16), .B(n10057), .S(P1_IR_REG_14__SCAN_IN), .Z(
        n10060) );
  XNOR2_X1 U11109 ( .A(n10058), .B(keyinput121), .ZN(n10059) );
  NOR3_X1 U11110 ( .A1(n10061), .A2(n10060), .A3(n10059), .ZN(n10077) );
  AOI22_X1 U11111 ( .A1(n10063), .A2(keyinput117), .B1(keyinput61), .B2(n7033), 
        .ZN(n10062) );
  OAI221_X1 U11112 ( .B1(n10063), .B2(keyinput117), .C1(n7033), .C2(keyinput61), .A(n10062), .ZN(n10075) );
  AOI22_X1 U11113 ( .A1(n10066), .A2(keyinput76), .B1(n10065), .B2(keyinput118), .ZN(n10064) );
  OAI221_X1 U11114 ( .B1(n10066), .B2(keyinput76), .C1(n10065), .C2(
        keyinput118), .A(n10064), .ZN(n10074) );
  AOI22_X1 U11115 ( .A1(n10069), .A2(keyinput12), .B1(n10068), .B2(keyinput74), 
        .ZN(n10067) );
  OAI221_X1 U11116 ( .B1(n10069), .B2(keyinput12), .C1(n10068), .C2(keyinput74), .A(n10067), .ZN(n10073) );
  XNOR2_X1 U11117 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput116), .ZN(n10071) );
  XNOR2_X1 U11118 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput46), .ZN(n10070)
         );
  NAND2_X1 U11119 ( .A1(n10071), .A2(n10070), .ZN(n10072) );
  NOR4_X1 U11120 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n10076) );
  OAI211_X1 U11121 ( .C1(keyinput6), .C2(n6437), .A(n10077), .B(n10076), .ZN(
        n10134) );
  AOI22_X1 U11122 ( .A1(n10079), .A2(keyinput110), .B1(n4492), .B2(keyinput114), .ZN(n10078) );
  OAI221_X1 U11123 ( .B1(n10079), .B2(keyinput110), .C1(n4492), .C2(
        keyinput114), .A(n10078), .ZN(n10089) );
  AOI22_X1 U11124 ( .A1(n10082), .A2(keyinput103), .B1(n10081), .B2(
        keyinput125), .ZN(n10080) );
  OAI221_X1 U11125 ( .B1(n10082), .B2(keyinput103), .C1(n10081), .C2(
        keyinput125), .A(n10080), .ZN(n10088) );
  XNOR2_X1 U11126 ( .A(SI_3_), .B(keyinput85), .ZN(n10086) );
  XNOR2_X1 U11127 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput98), .ZN(n10085) );
  XNOR2_X1 U11128 ( .A(P2_REG0_REG_27__SCAN_IN), .B(keyinput62), .ZN(n10084)
         );
  XNOR2_X1 U11129 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput58), .ZN(n10083) );
  NAND4_X1 U11130 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10087) );
  NOR3_X1 U11131 ( .A1(n10089), .A2(n10088), .A3(n10087), .ZN(n10132) );
  AOI22_X1 U11132 ( .A1(n10092), .A2(keyinput29), .B1(keyinput123), .B2(n10091), .ZN(n10090) );
  OAI221_X1 U11133 ( .B1(n10092), .B2(keyinput29), .C1(n10091), .C2(
        keyinput123), .A(n10090), .ZN(n10102) );
  AOI22_X1 U11134 ( .A1(n4736), .A2(keyinput75), .B1(keyinput82), .B2(n10094), 
        .ZN(n10093) );
  OAI221_X1 U11135 ( .B1(n4736), .B2(keyinput75), .C1(n10094), .C2(keyinput82), 
        .A(n10093), .ZN(n10101) );
  XOR2_X1 U11136 ( .A(n10095), .B(keyinput31), .Z(n10099) );
  XNOR2_X1 U11137 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput101), .ZN(n10098) );
  XNOR2_X1 U11138 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput105), .ZN(n10097) );
  XNOR2_X1 U11139 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput108), .ZN(n10096) );
  NAND4_X1 U11140 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n10100) );
  NOR3_X1 U11141 ( .A1(n10102), .A2(n10101), .A3(n10100), .ZN(n10131) );
  AOI22_X1 U11142 ( .A1(n10105), .A2(keyinput119), .B1(keyinput57), .B2(n10104), .ZN(n10103) );
  OAI221_X1 U11143 ( .B1(n10105), .B2(keyinput119), .C1(n10104), .C2(
        keyinput57), .A(n10103), .ZN(n10115) );
  INV_X1 U11144 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10108) );
  AOI22_X1 U11145 ( .A1(n10108), .A2(keyinput10), .B1(n10107), .B2(keyinput56), 
        .ZN(n10106) );
  OAI221_X1 U11146 ( .B1(n10108), .B2(keyinput10), .C1(n10107), .C2(keyinput56), .A(n10106), .ZN(n10114) );
  XNOR2_X1 U11147 ( .A(P1_REG3_REG_12__SCAN_IN), .B(keyinput79), .ZN(n10112)
         );
  XNOR2_X1 U11148 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput11), .ZN(n10111) );
  XNOR2_X1 U11149 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput107), .ZN(n10110) );
  XNOR2_X1 U11150 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput68), .ZN(n10109) );
  NAND4_X1 U11151 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n10113) );
  NOR3_X1 U11152 ( .A1(n10115), .A2(n10114), .A3(n10113), .ZN(n10130) );
  INV_X1 U11153 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U11154 ( .A1(n10118), .A2(keyinput65), .B1(keyinput20), .B2(n10117), 
        .ZN(n10116) );
  OAI221_X1 U11155 ( .B1(n10118), .B2(keyinput65), .C1(n10117), .C2(keyinput20), .A(n10116), .ZN(n10128) );
  AOI22_X1 U11156 ( .A1(n10120), .A2(keyinput43), .B1(n7083), .B2(keyinput84), 
        .ZN(n10119) );
  OAI221_X1 U11157 ( .B1(n10120), .B2(keyinput43), .C1(n7083), .C2(keyinput84), 
        .A(n10119), .ZN(n10127) );
  INV_X1 U11158 ( .A(keyinput54), .ZN(n10121) );
  XOR2_X1 U11159 ( .A(P1_WR_REG_SCAN_IN), .B(n10121), .Z(n10125) );
  XNOR2_X1 U11160 ( .A(keyinput122), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n10124)
         );
  XNOR2_X1 U11161 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput28), .ZN(n10123)
         );
  XNOR2_X1 U11162 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput112), .ZN(n10122) );
  NAND4_X1 U11163 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10126) );
  NOR3_X1 U11164 ( .A1(n10128), .A2(n10127), .A3(n10126), .ZN(n10129) );
  NAND4_X1 U11165 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n10133) );
  NOR4_X1 U11166 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10202) );
  NOR2_X1 U11167 ( .A1(keyinput32), .A2(keyinput40), .ZN(n10137) );
  NAND3_X1 U11168 ( .A1(keyinput70), .A2(keyinput78), .A3(n10137), .ZN(n10199)
         );
  INV_X1 U11169 ( .A(keyinput64), .ZN(n10138) );
  NAND4_X1 U11170 ( .A1(keyinput0), .A2(keyinput68), .A3(keyinput93), .A4(
        n10138), .ZN(n10198) );
  NAND4_X1 U11171 ( .A1(keyinput30), .A2(keyinput22), .A3(keyinput1), .A4(
        keyinput21), .ZN(n10139) );
  NOR3_X1 U11172 ( .A1(keyinput18), .A2(keyinput67), .A3(n10139), .ZN(n10148)
         );
  NOR4_X1 U11173 ( .A1(keyinput42), .A2(keyinput115), .A3(keyinput26), .A4(
        keyinput106), .ZN(n10145) );
  NAND2_X1 U11174 ( .A1(keyinput49), .A2(keyinput48), .ZN(n10140) );
  NOR3_X1 U11175 ( .A1(keyinput55), .A2(keyinput2), .A3(n10140), .ZN(n10144)
         );
  NAND2_X1 U11176 ( .A1(keyinput83), .A2(keyinput17), .ZN(n10141) );
  NOR3_X1 U11177 ( .A1(keyinput14), .A2(keyinput124), .A3(n10141), .ZN(n10143)
         );
  NOR4_X1 U11178 ( .A1(keyinput27), .A2(keyinput51), .A3(keyinput71), .A4(
        keyinput35), .ZN(n10142) );
  NAND4_X1 U11179 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10146) );
  NOR2_X1 U11180 ( .A1(n10146), .A2(keyinput86), .ZN(n10147) );
  NAND3_X1 U11181 ( .A1(keyinput66), .A2(n10148), .A3(n10147), .ZN(n10197) );
  INV_X1 U11182 ( .A(keyinput123), .ZN(n10149) );
  NOR4_X1 U11183 ( .A1(keyinput108), .A2(keyinput31), .A3(keyinput75), .A4(
        n10149), .ZN(n10195) );
  NOR4_X1 U11184 ( .A1(keyinput41), .A2(keyinput105), .A3(keyinput101), .A4(
        keyinput29), .ZN(n10194) );
  NOR2_X1 U11185 ( .A1(keyinput112), .A2(keyinput43), .ZN(n10150) );
  NAND3_X1 U11186 ( .A1(keyinput20), .A2(keyinput54), .A3(n10150), .ZN(n10161)
         );
  INV_X1 U11187 ( .A(keyinput65), .ZN(n10151) );
  NAND4_X1 U11188 ( .A1(keyinput122), .A2(keyinput85), .A3(keyinput28), .A4(
        n10151), .ZN(n10160) );
  INV_X1 U11189 ( .A(keyinput62), .ZN(n10152) );
  NOR4_X1 U11190 ( .A1(keyinput125), .A2(keyinput58), .A3(keyinput98), .A4(
        n10152), .ZN(n10158) );
  NAND2_X1 U11191 ( .A1(keyinput114), .A2(keyinput110), .ZN(n10153) );
  NOR3_X1 U11192 ( .A1(keyinput82), .A2(keyinput103), .A3(n10153), .ZN(n10157)
         );
  NOR4_X1 U11193 ( .A1(keyinput79), .A2(keyinput119), .A3(keyinput57), .A4(
        keyinput107), .ZN(n10156) );
  NAND2_X1 U11194 ( .A1(keyinput11), .A2(keyinput10), .ZN(n10154) );
  NOR3_X1 U11195 ( .A1(keyinput84), .A2(keyinput56), .A3(n10154), .ZN(n10155)
         );
  NAND4_X1 U11196 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n10159) );
  NOR3_X1 U11197 ( .A1(n10161), .A2(n10160), .A3(n10159), .ZN(n10193) );
  NAND2_X1 U11198 ( .A1(keyinput74), .A2(keyinput12), .ZN(n10162) );
  NOR3_X1 U11199 ( .A1(keyinput118), .A2(keyinput116), .A3(n10162), .ZN(n10167) );
  NOR4_X1 U11200 ( .A1(keyinput69), .A2(keyinput117), .A3(keyinput61), .A4(
        keyinput76), .ZN(n10166) );
  NAND2_X1 U11201 ( .A1(keyinput44), .A2(keyinput80), .ZN(n10163) );
  NOR3_X1 U11202 ( .A1(keyinput4), .A2(keyinput96), .A3(n10163), .ZN(n10165)
         );
  NOR4_X1 U11203 ( .A1(keyinput38), .A2(keyinput19), .A3(keyinput25), .A4(
        keyinput47), .ZN(n10164) );
  NAND4_X1 U11204 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10191) );
  INV_X1 U11205 ( .A(keyinput120), .ZN(n10168) );
  NAND4_X1 U11206 ( .A1(keyinput91), .A2(keyinput113), .A3(keyinput73), .A4(
        n10168), .ZN(n10169) );
  NOR4_X1 U11207 ( .A1(keyinput39), .A2(keyinput16), .A3(keyinput121), .A4(
        n10169), .ZN(n10173) );
  INV_X1 U11208 ( .A(keyinput13), .ZN(n10170) );
  NAND4_X1 U11209 ( .A1(keyinput5), .A2(keyinput23), .A3(keyinput24), .A4(
        n10170), .ZN(n10171) );
  NOR3_X1 U11210 ( .A1(keyinput3), .A2(keyinput102), .A3(n10171), .ZN(n10172)
         );
  NAND4_X1 U11211 ( .A1(n10173), .A2(keyinput46), .A3(keyinput104), .A4(n10172), .ZN(n10190) );
  NAND2_X1 U11212 ( .A1(keyinput59), .A2(keyinput127), .ZN(n10174) );
  NOR3_X1 U11213 ( .A1(keyinput97), .A2(keyinput72), .A3(n10174), .ZN(n10180)
         );
  INV_X1 U11214 ( .A(keyinput52), .ZN(n10175) );
  NOR4_X1 U11215 ( .A1(keyinput63), .A2(keyinput60), .A3(keyinput92), .A4(
        n10175), .ZN(n10179) );
  AND4_X1 U11216 ( .A1(keyinput87), .A2(keyinput34), .A3(keyinput33), .A4(
        keyinput15), .ZN(n10178) );
  INV_X1 U11217 ( .A(keyinput53), .ZN(n10176) );
  NOR4_X1 U11218 ( .A1(keyinput111), .A2(keyinput89), .A3(keyinput126), .A4(
        n10176), .ZN(n10177) );
  NAND4_X1 U11219 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10189) );
  NAND2_X1 U11220 ( .A1(keyinput9), .A2(keyinput7), .ZN(n10181) );
  NOR3_X1 U11221 ( .A1(keyinput77), .A2(keyinput88), .A3(n10181), .ZN(n10187)
         );
  NOR4_X1 U11222 ( .A1(keyinput99), .A2(keyinput109), .A3(keyinput94), .A4(
        keyinput100), .ZN(n10186) );
  NAND2_X1 U11223 ( .A1(keyinput45), .A2(keyinput50), .ZN(n10182) );
  NOR3_X1 U11224 ( .A1(keyinput81), .A2(keyinput36), .A3(n10182), .ZN(n10185)
         );
  INV_X1 U11225 ( .A(keyinput37), .ZN(n10183) );
  NOR4_X1 U11226 ( .A1(keyinput8), .A2(keyinput90), .A3(keyinput95), .A4(
        n10183), .ZN(n10184) );
  NAND4_X1 U11227 ( .A1(n10187), .A2(n10186), .A3(n10185), .A4(n10184), .ZN(
        n10188) );
  NOR4_X1 U11228 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10192) );
  NAND4_X1 U11229 ( .A1(n10195), .A2(n10194), .A3(n10193), .A4(n10192), .ZN(
        n10196) );
  NOR4_X1 U11230 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n10200) );
  OAI21_X1 U11231 ( .B1(keyinput6), .B2(n10200), .A(n6437), .ZN(n10201) );
  NAND4_X1 U11232 ( .A1(n10204), .A2(n10203), .A3(n10202), .A4(n10201), .ZN(
        n10205) );
  NOR3_X1 U11233 ( .A1(n10207), .A2(n10206), .A3(n10205), .ZN(n10208) );
  XNOR2_X1 U11234 ( .A(n10209), .B(n10208), .ZN(P2_U3298) );
  XOR2_X1 U11235 ( .A(n10210), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11236 ( .A1(n10212), .A2(n10211), .ZN(n10213) );
  XOR2_X1 U11237 ( .A(n10213), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11238 ( .A(n10214), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11239 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(n10219) );
  XOR2_X1 U11240 ( .A(n10219), .B(n10218), .Z(ADD_1071_U55) );
  XOR2_X1 U11241 ( .A(n10220), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  AOI21_X1 U11242 ( .B1(n10223), .B2(n10222), .A(n10221), .ZN(ADD_1071_U47) );
  XOR2_X1 U11243 ( .A(n10225), .B(n10224), .Z(ADD_1071_U54) );
  XOR2_X1 U11244 ( .A(n10227), .B(n10226), .Z(ADD_1071_U53) );
  XNOR2_X1 U11245 ( .A(n10229), .B(n10228), .ZN(ADD_1071_U52) );
  NAND4_X1 U4922 ( .A1(n4561), .A2(n4560), .A3(n4771), .A4(n4770), .ZN(n6068)
         );
  CLKBUF_X2 U4962 ( .A(n6741), .Z(n6230) );
  AND2_X1 U5194 ( .A1(n5652), .A2(n5649), .ZN(n5633) );
endmodule

