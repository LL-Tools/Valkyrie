

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2260, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4914;

  CLKBUF_X1 U2294 ( .A(n2560), .Z(n3640) );
  INV_X1 U2295 ( .A(n3054), .ZN(n3031) );
  NAND4_X1 U2296 ( .A1(n2564), .A2(n2563), .A3(n2562), .A4(n2561), .ZN(n3034)
         );
  NAND2_X1 U2298 ( .A1(n2931), .A2(IR_REG_31__SCAN_IN), .ZN(n2514) );
  CLKBUF_X1 U2299 ( .A(n4815), .Z(n2260) );
  NOR2_X1 U2300 ( .A1(n4907), .A2(n2871), .ZN(n4815) );
  INV_X1 U2302 ( .A(n4914), .ZN(n2262) );
  BUF_X1 U2303 ( .A(n3054), .Z(n3948) );
  NAND2_X1 U2304 ( .A1(n2912), .A2(n3726), .ZN(n2979) );
  INV_X2 U2305 ( .A(n3891), .ZN(n3433) );
  CLKBUF_X2 U2307 ( .A(n2552), .Z(n3642) );
  NOR2_X1 U2308 ( .A1(n4665), .A2(n4664), .ZN(n4663) );
  XOR2_X1 U2309 ( .A(n4152), .B(n4161), .Z(n4722) );
  INV_X1 U2310 ( .A(n3726), .ZN(n3012) );
  NAND4_X1 U2311 ( .A1(n2582), .A2(n2581), .A3(n2580), .A4(n2579), .ZN(n4116)
         );
  INV_X2 U2312 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2313 ( .A(n2925), .ZN(n2517) );
  OAI21_X1 U2314 ( .B1(n2882), .B2(n2522), .A(IR_REG_31__SCAN_IN), .ZN(n2834)
         );
  NOR2_X2 U2315 ( .A1(n3152), .A2(n3153), .ZN(n3183) );
  NOR3_X2 U2316 ( .A1(n3854), .A2(n3853), .A3(n3857), .ZN(n3855) );
  AND2_X2 U2317 ( .A1(n2974), .A2(REG2_REG_4__SCAN_IN), .ZN(n3245) );
  NAND2_X2 U2318 ( .A1(n4153), .A2(n4721), .ZN(n4732) );
  XNOR2_X2 U2319 ( .A(n2514), .B(IR_REG_30__SCAN_IN), .ZN(n4447) );
  XNOR2_X1 U2320 ( .A(n2413), .B(n4905), .ZN(n4741) );
  AND2_X1 U2321 ( .A1(n2351), .A2(n2356), .ZN(n3271) );
  AND2_X2 U2322 ( .A1(n3104), .A2(n4875), .ZN(n4858) );
  INV_X4 U2323 ( .A(n3433), .ZN(n3899) );
  NAND2_X1 U2324 ( .A1(n2304), .A2(n2877), .ZN(n2882) );
  INV_X2 U2325 ( .A(IR_REG_31__SCAN_IN), .ZN(n2930) );
  NAND2_X2 U2326 ( .A1(n3968), .A2(n3915), .ZN(n3971) );
  NAND2_X1 U2327 ( .A1(n4741), .A2(n3478), .ZN(n4740) );
  NAND2_X1 U2328 ( .A1(n4196), .A2(n4195), .ZN(n2413) );
  NAND2_X1 U2329 ( .A1(n4147), .A2(n4148), .ZN(n4149) );
  OAI21_X1 U2330 ( .B1(n2356), .B2(n2355), .A(n2354), .ZN(n2349) );
  CLKBUF_X3 U2332 ( .A(n3431), .Z(n3947) );
  AND2_X1 U2333 ( .A1(n4823), .A2(n3051), .ZN(n3431) );
  NAND2_X1 U2334 ( .A1(n2764), .A2(n2814), .ZN(n4828) );
  INV_X2 U2335 ( .A(n3778), .ZN(n2263) );
  NOR2_X4 U2336 ( .A1(n4447), .A2(n2517), .ZN(n2560) );
  XNOR2_X1 U2337 ( .A(n2816), .B(n2815), .ZN(n2912) );
  NAND2_X1 U2338 ( .A1(n2814), .A2(IR_REG_31__SCAN_IN), .ZN(n2816) );
  XNOR2_X1 U2339 ( .A(n2820), .B(IR_REG_21__SCAN_IN), .ZN(n3726) );
  XNOR2_X1 U2340 ( .A(n2883), .B(n2885), .ZN(n2890) );
  NAND2_X1 U2341 ( .A1(n2882), .A2(IR_REG_31__SCAN_IN), .ZN(n2883) );
  INV_X1 U2342 ( .A(n2882), .ZN(n2829) );
  NAND2_X1 U2343 ( .A1(n2549), .A2(n2277), .ZN(n4125) );
  AND2_X1 U2344 ( .A1(n2876), .A2(n2508), .ZN(n2304) );
  AND2_X1 U2345 ( .A1(n2548), .A2(n2565), .ZN(n2574) );
  NOR2_X1 U2346 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2692)
         );
  NOR2_X1 U2347 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2691)
         );
  NOR2_X1 U2348 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2694)
         );
  NOR2_X1 U2349 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2693)
         );
  INV_X1 U2350 ( .A(IR_REG_2__SCAN_IN), .ZN(n2565) );
  NOR2_X2 U2351 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2548)
         );
  NAND2_X2 U2352 ( .A1(n3992), .A2(n3887), .ZN(n4004) );
  INV_X1 U2353 ( .A(n3639), .ZN(n3646) );
  NAND2_X1 U2354 ( .A1(n2718), .A2(n2455), .ZN(n2453) );
  NOR2_X1 U2355 ( .A1(n2440), .A2(n2437), .ZN(n2436) );
  INV_X1 U2356 ( .A(n2622), .ZN(n2437) );
  INV_X1 U2357 ( .A(n2441), .ZN(n2440) );
  INV_X1 U2358 ( .A(IR_REG_19__SCAN_IN), .ZN(n2503) );
  INV_X1 U2359 ( .A(IR_REG_5__SCAN_IN), .ZN(n2607) );
  NOR2_X1 U2360 ( .A1(n2360), .A2(n2283), .ZN(n2358) );
  INV_X1 U2361 ( .A(n2270), .ZN(n2353) );
  AND2_X1 U2362 ( .A1(n4447), .A2(n2517), .ZN(n2559) );
  AOI22_X1 U2363 ( .A1(n2959), .A2(n4138), .B1(n4454), .B2(REG1_REG_2__SCAN_IN), .ZN(n2975) );
  INV_X1 U2364 ( .A(n4654), .ZN(n2418) );
  OAI21_X1 U2365 ( .B1(n4707), .B2(n2346), .A(n2345), .ZN(n4162) );
  OR2_X1 U2366 ( .A1(n4705), .A2(REG1_REG_11__SCAN_IN), .ZN(n2345) );
  AND2_X1 U2367 ( .A1(n4705), .A2(REG1_REG_11__SCAN_IN), .ZN(n2346) );
  OAI21_X1 U2368 ( .B1(n4246), .B2(n4265), .A(n2800), .ZN(n4234) );
  NAND2_X1 U2369 ( .A1(n3535), .A2(n2738), .ZN(n2428) );
  NAND2_X1 U2370 ( .A1(n2877), .A2(n2876), .ZN(n2878) );
  OR2_X1 U2371 ( .A1(n4234), .A2(n2474), .ZN(n2467) );
  AOI21_X1 U2372 ( .B1(n4234), .B2(n2472), .A(n2469), .ZN(n2468) );
  AND2_X1 U2373 ( .A1(n4241), .A2(n2478), .ZN(n2472) );
  NAND2_X1 U2374 ( .A1(n2470), .A2(n2475), .ZN(n2469) );
  NAND2_X1 U2375 ( .A1(n2476), .A2(n2478), .ZN(n2475) );
  AND2_X1 U2376 ( .A1(n2497), .A2(n2486), .ZN(n2485) );
  NOR2_X1 U2377 ( .A1(n2789), .A2(n3814), .ZN(n2497) );
  NAND2_X1 U2378 ( .A1(n2488), .A2(n2492), .ZN(n2486) );
  AND2_X1 U2379 ( .A1(n2767), .A2(REG3_REG_21__SCAN_IN), .ZN(n2774) );
  NAND2_X1 U2380 ( .A1(n4104), .A2(n4053), .ZN(n2498) );
  AND2_X1 U2381 ( .A1(n2747), .A2(REG3_REG_20__SCAN_IN), .ZN(n2767) );
  INV_X1 U2382 ( .A(n3588), .ZN(n2324) );
  INV_X1 U2383 ( .A(n3621), .ZN(n2321) );
  INV_X1 U2384 ( .A(n3592), .ZN(n2320) );
  NOR2_X1 U2385 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2523)
         );
  NAND2_X1 U2386 ( .A1(n4256), .A2(n4243), .ZN(n2479) );
  NAND2_X1 U2387 ( .A1(n4292), .A2(n2307), .ZN(n2306) );
  AND2_X1 U2388 ( .A1(n4261), .A2(n2309), .ZN(n2307) );
  AND2_X1 U2389 ( .A1(n2310), .A2(n3698), .ZN(n2309) );
  OR2_X1 U2390 ( .A1(n3701), .A2(n3716), .ZN(n2310) );
  AOI21_X1 U2391 ( .B1(n2485), .B2(n2483), .A(n4331), .ZN(n2482) );
  INV_X1 U2392 ( .A(n2488), .ZN(n2483) );
  INV_X1 U2393 ( .A(n2485), .ZN(n2484) );
  OAI21_X1 U2394 ( .B1(n3821), .B2(n2860), .A(n2863), .ZN(n4311) );
  INV_X1 U2395 ( .A(n3377), .ZN(n2456) );
  NAND2_X1 U2396 ( .A1(n3326), .A2(n2682), .ZN(n2457) );
  NOR2_X1 U2397 ( .A1(n2650), .A2(n2442), .ZN(n2441) );
  INV_X1 U2398 ( .A(n2633), .ZN(n2442) );
  OR2_X1 U2399 ( .A1(n3148), .A2(n3145), .ZN(n2840) );
  NAND2_X1 U2400 ( .A1(n2432), .A2(n2587), .ZN(n2431) );
  OR2_X1 U2401 ( .A1(n3400), .A2(n3404), .ZN(n3402) );
  NOR2_X1 U2402 ( .A1(n2512), .A2(n2511), .ZN(n2704) );
  INV_X1 U2403 ( .A(IR_REG_13__SCAN_IN), .ZN(n2510) );
  NOR2_X1 U2404 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2509)
         );
  NOR2_X1 U2405 ( .A1(n2387), .A2(n4042), .ZN(n2385) );
  INV_X1 U2406 ( .A(n2386), .ZN(n2383) );
  INV_X1 U2407 ( .A(n3760), .ZN(n2364) );
  INV_X1 U2408 ( .A(n3994), .ZN(n3885) );
  INV_X1 U2409 ( .A(n4063), .ZN(n3910) );
  NAND2_X1 U2410 ( .A1(n2266), .A2(n2365), .ZN(n2360) );
  INV_X1 U2411 ( .A(n3866), .ZN(n2365) );
  XNOR2_X1 U2412 ( .A(n3115), .B(n3948), .ZN(n3268) );
  XNOR2_X1 U2413 ( .A(n4142), .B(n2956), .ZN(n4137) );
  NOR2_X1 U2414 ( .A1(n2972), .A2(n2971), .ZN(n3244) );
  NAND2_X1 U2415 ( .A1(n2332), .A2(n2269), .ZN(n3232) );
  NAND2_X1 U2416 ( .A1(n2265), .A2(n2339), .ZN(n2332) );
  NAND2_X1 U2417 ( .A1(n2421), .A2(n3248), .ZN(n2417) );
  NAND2_X1 U2418 ( .A1(n4658), .A2(n3233), .ZN(n3234) );
  XNOR2_X1 U2419 ( .A(n4149), .B(n2422), .ZN(n4696) );
  NAND2_X1 U2420 ( .A1(n4696), .A2(REG2_REG_10__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U2421 ( .A1(n2426), .A2(REG2_REG_14__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U2422 ( .A1(n4154), .A2(n4172), .ZN(n2426) );
  NOR2_X1 U2423 ( .A1(n4212), .A2(n4213), .ZN(n4753) );
  AND2_X1 U2424 ( .A1(n3779), .A2(n2739), .ZN(n2427) );
  NAND2_X1 U2425 ( .A1(n2500), .A2(n2763), .ZN(n2814) );
  AND2_X1 U2426 ( .A1(n2762), .A2(n2761), .ZN(n2763) );
  NAND2_X1 U2427 ( .A1(n2588), .A2(REG3_REG_6__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U2428 ( .A1(n2433), .A2(n3686), .ZN(n3136) );
  OAI21_X1 U2429 ( .B1(n2467), .B2(n2466), .A(n2464), .ZN(n2461) );
  AND2_X1 U2430 ( .A1(n2477), .A2(n4849), .ZN(n2464) );
  NAND2_X1 U2431 ( .A1(n2298), .A2(n4265), .ZN(n2297) );
  NOR2_X1 U2432 ( .A1(n2300), .A2(n4243), .ZN(n2298) );
  INV_X1 U2433 ( .A(n3658), .ZN(n2300) );
  AND2_X1 U2434 ( .A1(n2912), .A2(n3127), .ZN(n4406) );
  NAND2_X1 U2435 ( .A1(n2318), .A2(IR_REG_31__SCAN_IN), .ZN(n2317) );
  AND2_X1 U2436 ( .A1(n2513), .A2(IR_REG_29__SCAN_IN), .ZN(n2313) );
  OR2_X1 U2437 ( .A1(n2513), .A2(n2317), .ZN(n2316) );
  INV_X1 U2438 ( .A(IR_REG_28__SCAN_IN), .ZN(n2832) );
  INV_X1 U2439 ( .A(IR_REG_21__SCAN_IN), .ZN(n2821) );
  NOR2_X1 U2440 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2505)
         );
  NOR2_X1 U2441 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2504)
         );
  INV_X1 U2442 ( .A(IR_REG_9__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U2443 ( .A1(n2405), .A2(n2930), .ZN(n2404) );
  INV_X1 U2444 ( .A(n2347), .ZN(n3270) );
  NAND2_X1 U2445 ( .A1(n3114), .A2(n2276), .ZN(n2350) );
  NAND2_X1 U2446 ( .A1(n2375), .A2(n4084), .ZN(n3960) );
  AOI21_X1 U2447 ( .B1(n2264), .B2(n2397), .A(n2391), .ZN(n2390) );
  INV_X1 U2448 ( .A(n3524), .ZN(n2391) );
  NAND2_X1 U2449 ( .A1(n2392), .A2(n2394), .ZN(n3525) );
  NAND2_X1 U2450 ( .A1(n3426), .A2(n2393), .ZN(n2392) );
  NAND2_X1 U2451 ( .A1(n2552), .A2(REG0_REG_3__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U2452 ( .A1(n2552), .A2(REG0_REG_2__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U2453 ( .A(n4125), .B(REG2_REG_1__SCAN_IN), .ZN(n4124) );
  XNOR2_X1 U2454 ( .A(n2975), .B(n4453), .ZN(n2976) );
  XNOR2_X1 U2455 ( .A(n3234), .B(n4801), .ZN(n4669) );
  NAND2_X1 U2456 ( .A1(n4669), .A2(REG1_REG_6__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U2457 ( .A1(n4697), .A2(n4160), .ZN(n4707) );
  XNOR2_X1 U2458 ( .A(n4162), .B(n4882), .ZN(n4717) );
  NOR2_X1 U2459 ( .A1(n4717), .A2(n4718), .ZN(n4716) );
  NAND2_X1 U2460 ( .A1(n2344), .A2(n2343), .ZN(n2342) );
  NAND2_X1 U2461 ( .A1(n4192), .A2(n2344), .ZN(n2341) );
  INV_X1 U2462 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2343) );
  NAND2_X1 U2463 ( .A1(n2463), .A2(n2462), .ZN(n2916) );
  NAND2_X1 U2464 ( .A1(n2477), .A2(n2466), .ZN(n2462) );
  AOI21_X1 U2465 ( .B1(n2491), .B2(n2490), .A(n2489), .ZN(n2488) );
  INV_X1 U2466 ( .A(n2494), .ZN(n2490) );
  INV_X1 U2467 ( .A(n3813), .ZN(n2489) );
  NOR2_X1 U2468 ( .A1(n2790), .A2(n4608), .ZN(n2537) );
  INV_X1 U2469 ( .A(n2498), .ZN(n2493) );
  NOR2_X1 U2470 ( .A1(n2765), .A2(n2273), .ZN(n2495) );
  AND2_X1 U2471 ( .A1(n3427), .A2(n2403), .ZN(n2402) );
  INV_X1 U2472 ( .A(n3501), .ZN(n2403) );
  AND2_X1 U2473 ( .A1(n3501), .A2(n2399), .ZN(n2398) );
  AOI21_X1 U2474 ( .B1(n2402), .B2(n3428), .A(n2401), .ZN(n2400) );
  INV_X1 U2475 ( .A(n3500), .ZN(n2401) );
  INV_X1 U2476 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2961) );
  OR2_X1 U2477 ( .A1(n2337), .A2(n3243), .ZN(n2331) );
  NOR2_X1 U2478 ( .A1(n3243), .A2(n2334), .ZN(n2333) );
  INV_X1 U2479 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U2480 ( .A1(n3246), .A2(n2973), .ZN(n2421) );
  OR2_X1 U2481 ( .A1(n4292), .A2(n3701), .ZN(n2308) );
  NAND2_X1 U2482 ( .A1(n2537), .A2(REG3_REG_24__SCAN_IN), .ZN(n2539) );
  AND2_X1 U2483 ( .A1(n2498), .A2(n2766), .ZN(n2494) );
  INV_X1 U2484 ( .A(n2323), .ZN(n2322) );
  AOI21_X1 U2485 ( .B1(n2323), .B2(n2321), .A(n2320), .ZN(n2319) );
  AOI21_X1 U2486 ( .B1(n3619), .B2(n3621), .A(n2324), .ZN(n2323) );
  OR2_X1 U2487 ( .A1(n3034), .A2(n3165), .ZN(n3604) );
  OR2_X1 U2488 ( .A1(n2834), .A2(n2501), .ZN(n2524) );
  NAND2_X1 U2489 ( .A1(n2834), .A2(n2523), .ZN(n2294) );
  NAND2_X1 U2490 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2501) );
  OR2_X1 U2491 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2522)
         );
  INV_X1 U2492 ( .A(IR_REG_7__SCAN_IN), .ZN(n2643) );
  INV_X1 U2493 ( .A(n2349), .ZN(n2348) );
  XOR2_X1 U2494 ( .A(n3951), .B(n3950), .Z(n3952) );
  AOI21_X1 U2495 ( .B1(n2373), .B2(n4085), .A(n2372), .ZN(n2371) );
  INV_X1 U2496 ( .A(n3945), .ZN(n2372) );
  AOI22_X1 U2497 ( .A1(n4120), .A2(n3891), .B1(n3051), .B2(n3126), .ZN(n2993)
         );
  AOI22_X1 U2498 ( .A1(n2400), .A2(n2396), .B1(n2398), .B2(n2395), .ZN(n2394)
         );
  INV_X1 U2499 ( .A(n3427), .ZN(n2395) );
  INV_X1 U2500 ( .A(n2402), .ZN(n2396) );
  AND2_X1 U2501 ( .A1(n2672), .A2(REG3_REG_12__SCAN_IN), .ZN(n2685) );
  AND2_X1 U2502 ( .A1(n2685), .A2(REG3_REG_13__SCAN_IN), .ZN(n2698) );
  AOI21_X1 U2503 ( .B1(n2383), .B2(n2382), .A(n2282), .ZN(n2381) );
  NOR2_X1 U2504 ( .A1(n2385), .A2(n2384), .ZN(n2382) );
  OAI22_X1 U2505 ( .A1(n3927), .A2(n3926), .B1(n3433), .B2(n4301), .ZN(n4018)
         );
  NAND2_X1 U2506 ( .A1(n2698), .A2(REG3_REG_14__SCAN_IN), .ZN(n2708) );
  NOR2_X1 U2507 ( .A1(n2964), .A2(n2965), .ZN(n2972) );
  INV_X1 U2508 ( .A(IR_REG_3__SCAN_IN), .ZN(n4641) );
  INV_X1 U2509 ( .A(IR_REG_4__SCAN_IN), .ZN(n4537) );
  OR2_X1 U2510 ( .A1(n3245), .A2(n2420), .ZN(n2419) );
  INV_X1 U2511 ( .A(n2421), .ZN(n2420) );
  NOR2_X1 U2512 ( .A1(n4663), .A2(n3252), .ZN(n4676) );
  NAND2_X1 U2513 ( .A1(n2415), .A2(n2414), .ZN(n3255) );
  NAND2_X1 U2514 ( .A1(n2416), .A2(REG2_REG_7__SCAN_IN), .ZN(n2415) );
  OR2_X1 U2515 ( .A1(n4676), .A2(n4810), .ZN(n2414) );
  NAND2_X1 U2516 ( .A1(n4676), .A2(n4810), .ZN(n2416) );
  NOR2_X1 U2517 ( .A1(n3237), .A2(n4685), .ZN(n4158) );
  AND2_X1 U2518 ( .A1(n2424), .A2(n2423), .ZN(n4180) );
  NAND2_X1 U2519 ( .A1(n4740), .A2(n4198), .ZN(n4199) );
  INV_X1 U2520 ( .A(n2413), .ZN(n4197) );
  INV_X1 U2521 ( .A(n4194), .ZN(n2344) );
  NAND2_X1 U2522 ( .A1(n4754), .A2(REG2_REG_18__SCAN_IN), .ZN(n2411) );
  INV_X1 U2523 ( .A(n2479), .ZN(n2476) );
  NAND2_X1 U2524 ( .A1(n2471), .A2(n2473), .ZN(n2470) );
  INV_X1 U2525 ( .A(n4241), .ZN(n2471) );
  NAND2_X1 U2526 ( .A1(n2306), .A2(n2305), .ZN(n2311) );
  AOI21_X1 U2527 ( .B1(n2307), .B2(n3701), .A(n3702), .ZN(n2305) );
  INV_X1 U2528 ( .A(n2444), .ZN(n4262) );
  OAI21_X1 U2529 ( .B1(n4272), .B2(n2446), .A(n2445), .ZN(n2444) );
  NAND2_X1 U2530 ( .A1(n2447), .A2(n4283), .ZN(n2445) );
  NOR2_X1 U2531 ( .A1(n2447), .A2(n4283), .ZN(n2446) );
  AND2_X1 U2532 ( .A1(n2308), .A2(n2307), .ZN(n4252) );
  NAND2_X1 U2533 ( .A1(n2308), .A2(n2309), .ZN(n4254) );
  AND2_X1 U2534 ( .A1(n4292), .A2(n3716), .ZN(n4275) );
  NAND2_X1 U2535 ( .A1(n2449), .A2(n2448), .ZN(n4272) );
  NAND2_X1 U2536 ( .A1(n4316), .A2(n4296), .ZN(n2448) );
  NAND2_X1 U2537 ( .A1(n4290), .A2(n2450), .ZN(n2449) );
  OR2_X1 U2538 ( .A1(n4316), .A2(n4296), .ZN(n2450) );
  OR2_X1 U2539 ( .A1(n4319), .A2(n4347), .ZN(n2797) );
  AOI21_X1 U2540 ( .B1(n2482), .B2(n2484), .A(n2279), .ZN(n2481) );
  INV_X1 U2541 ( .A(n4101), .ZN(n4319) );
  AND2_X1 U2542 ( .A1(n2783), .A2(n2777), .ZN(n3805) );
  NAND2_X1 U2543 ( .A1(n2487), .A2(n2491), .ZN(n3815) );
  NAND2_X1 U2544 ( .A1(n3556), .A2(n2494), .ZN(n2487) );
  OAI21_X1 U2545 ( .B1(n3836), .B2(n3707), .A(n3710), .ZN(n3821) );
  AND2_X1 U2546 ( .A1(n2776), .A2(n2769), .ZN(n3847) );
  INV_X1 U2547 ( .A(n3892), .ZN(n4053) );
  NOR2_X1 U2548 ( .A1(n2740), .A2(n4076), .ZN(n2748) );
  NOR2_X1 U2549 ( .A1(n2719), .A2(n4624), .ZN(n2727) );
  NAND2_X1 U2550 ( .A1(n2453), .A2(n2452), .ZN(n2451) );
  INV_X1 U2551 ( .A(n2717), .ZN(n2452) );
  NAND2_X1 U2552 ( .A1(n2457), .A2(n2454), .ZN(n3444) );
  NAND2_X1 U2553 ( .A1(n2457), .A2(n2683), .ZN(n3378) );
  OR2_X1 U2554 ( .A1(n2634), .A2(n4550), .ZN(n2651) );
  INV_X1 U2555 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3984) );
  AOI21_X1 U2556 ( .B1(n2441), .B2(n2439), .A(n2278), .ZN(n2438) );
  INV_X1 U2557 ( .A(n2632), .ZN(n2439) );
  NAND2_X1 U2558 ( .A1(n2623), .A2(REG3_REG_8__SCAN_IN), .ZN(n2634) );
  AND2_X1 U2559 ( .A1(n2431), .A2(n2598), .ZN(n2429) );
  OAI21_X1 U2560 ( .B1(n3131), .B2(n2838), .A(n3614), .ZN(n3148) );
  NAND2_X1 U2561 ( .A1(n3195), .A2(n3609), .ZN(n3131) );
  AND2_X1 U2562 ( .A1(n3091), .A2(n2557), .ZN(n3162) );
  NAND2_X1 U2563 ( .A1(n3604), .A2(n3607), .ZN(n3685) );
  NAND2_X1 U2564 ( .A1(n3600), .A2(n3603), .ZN(n3684) );
  NAND2_X1 U2565 ( .A1(n3684), .A2(n3092), .ZN(n3091) );
  AND2_X1 U2566 ( .A1(n2872), .A2(n3012), .ZN(n3127) );
  NOR2_X1 U2567 ( .A1(n2268), .A2(n4360), .ZN(n4357) );
  INV_X1 U2568 ( .A(n4819), .ZN(n4359) );
  NAND2_X1 U2569 ( .A1(n4303), .A2(n4283), .ZN(n4370) );
  AND2_X1 U2570 ( .A1(n4322), .A2(n4301), .ZN(n4303) );
  NOR2_X1 U2571 ( .A1(n4346), .A2(n4315), .ZN(n4322) );
  OR2_X1 U2572 ( .A1(n4387), .A2(n3973), .ZN(n4346) );
  NAND2_X1 U2573 ( .A1(n3827), .A2(n4064), .ZN(n4387) );
  NOR2_X1 U2574 ( .A1(n3776), .A2(n2301), .ZN(n3827) );
  NAND2_X1 U2575 ( .A1(n3881), .A2(n2302), .ZN(n2301) );
  NOR2_X1 U2576 ( .A1(n4053), .A2(n4010), .ZN(n2302) );
  NOR3_X1 U2577 ( .A1(n3776), .A2(n3998), .A3(n4053), .ZN(n3846) );
  AND2_X1 U2578 ( .A1(n2496), .A2(n2499), .ZN(n3841) );
  NAND2_X1 U2579 ( .A1(n3556), .A2(n2766), .ZN(n2496) );
  NAND2_X1 U2580 ( .A1(n3777), .A2(n3872), .ZN(n3776) );
  NOR2_X1 U2581 ( .A1(n4407), .A2(n3769), .ZN(n3777) );
  NAND2_X1 U2582 ( .A1(n3453), .A2(n2303), .ZN(n3492) );
  NOR2_X1 U2583 ( .A1(n3528), .A2(n4894), .ZN(n2303) );
  NAND2_X1 U2584 ( .A1(n3453), .A2(n3452), .ZN(n3491) );
  INV_X1 U2585 ( .A(n3509), .ZN(n3389) );
  AND2_X1 U2586 ( .A1(n3390), .A2(n3389), .ZN(n3453) );
  NOR2_X1 U2587 ( .A1(n3398), .A2(n3436), .ZN(n3390) );
  OR2_X1 U2588 ( .A1(n3397), .A2(n3370), .ZN(n3398) );
  INV_X1 U2589 ( .A(n3985), .ZN(n3339) );
  NAND2_X1 U2590 ( .A1(n3340), .A2(n3339), .ZN(n3397) );
  AND2_X1 U2591 ( .A1(n3301), .A2(n2911), .ZN(n3340) );
  NAND2_X1 U2592 ( .A1(n2293), .A2(n2292), .ZN(n4826) );
  INV_X1 U2593 ( .A(n4825), .ZN(n2293) );
  NOR2_X1 U2594 ( .A1(n4826), .A2(n3302), .ZN(n3301) );
  INV_X1 U2595 ( .A(n3176), .ZN(n3182) );
  OR2_X1 U2596 ( .A1(n3208), .A2(n3860), .ZN(n3152) );
  INV_X1 U2597 ( .A(n3199), .ZN(n3205) );
  NOR2_X1 U2598 ( .A1(n3171), .A2(n3172), .ZN(n3206) );
  INV_X1 U2599 ( .A(n4406), .ZN(n4823) );
  INV_X1 U2600 ( .A(IR_REG_20__SCAN_IN), .ZN(n2815) );
  NAND2_X1 U2601 ( .A1(n2359), .A2(n2358), .ZN(n3877) );
  NAND2_X1 U2602 ( .A1(n2371), .A2(n2370), .ZN(n2369) );
  INV_X1 U2603 ( .A(n3952), .ZN(n2370) );
  NAND2_X1 U2604 ( .A1(n3971), .A2(n2379), .ZN(n2378) );
  NAND2_X1 U2605 ( .A1(n2383), .A2(n2380), .ZN(n2379) );
  INV_X1 U2606 ( .A(n2385), .ZN(n2380) );
  INV_X1 U2607 ( .A(n2502), .ZN(n2361) );
  AOI21_X1 U2608 ( .B1(n3971), .B2(n3922), .A(n3923), .ZN(n4041) );
  INV_X1 U2609 ( .A(n3124), .ZN(n3126) );
  OR2_X1 U2610 ( .A1(n3359), .A2(n3358), .ZN(n3360) );
  INV_X1 U2611 ( .A(n3165), .ZN(n3172) );
  INV_X1 U2612 ( .A(n2360), .ZN(n2357) );
  NAND2_X1 U2613 ( .A1(n3114), .A2(n2353), .ZN(n2352) );
  CLKBUF_X1 U2614 ( .A(n4092), .Z(n4893) );
  NAND4_X1 U2615 ( .A1(n2606), .A2(n2605), .A3(n2604), .A4(n2603), .ZN(n4816)
         );
  CLKBUF_X1 U2616 ( .A(n2996), .Z(n4118) );
  AND2_X1 U2617 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4123)
         );
  OR2_X1 U2618 ( .A1(n2548), .A2(n2930), .ZN(n2340) );
  OAI21_X1 U2619 ( .B1(n3232), .B2(n3231), .A(n2335), .ZN(n4659) );
  INV_X1 U2620 ( .A(n2419), .ZN(n4655) );
  NAND2_X1 U2621 ( .A1(n4668), .A2(n3235), .ZN(n4681) );
  XNOR2_X1 U2622 ( .A(n3255), .B(n3254), .ZN(n4691) );
  NAND2_X1 U2623 ( .A1(n4691), .A2(REG2_REG_8__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U2624 ( .A1(n4695), .A2(n4150), .ZN(n4712) );
  NOR2_X1 U2625 ( .A1(n4163), .A2(n4716), .ZN(n4728) );
  NOR2_X1 U2626 ( .A1(n4177), .A2(n2424), .ZN(n4176) );
  OR2_X1 U2627 ( .A1(n2425), .A2(n4177), .ZN(n4155) );
  INV_X1 U2628 ( .A(n2426), .ZN(n2425) );
  XNOR2_X1 U2629 ( .A(n4191), .B(n4190), .ZN(n4745) );
  NOR2_X1 U2630 ( .A1(n4745), .A2(REG1_REG_16__SCAN_IN), .ZN(n4746) );
  AOI21_X1 U2631 ( .B1(n4750), .B2(n4751), .A(n2291), .ZN(n2329) );
  INV_X1 U2632 ( .A(n4752), .ZN(n2328) );
  NAND2_X1 U2633 ( .A1(n2412), .A2(n2411), .ZN(n2410) );
  INV_X1 U2634 ( .A(n4760), .ZN(n2407) );
  NAND2_X1 U2635 ( .A1(n2428), .A2(n2739), .ZN(n3787) );
  OR2_X1 U2636 ( .A1(n3492), .A2(n4034), .ZN(n4407) );
  NAND2_X1 U2637 ( .A1(n3294), .A2(n2632), .ZN(n2443) );
  NAND2_X1 U2638 ( .A1(n3136), .A2(n2587), .ZN(n3146) );
  NOR2_X1 U2639 ( .A1(n2915), .A2(n3101), .ZN(n4846) );
  INV_X1 U2640 ( .A(n4411), .ZN(n4844) );
  INV_X1 U2641 ( .A(n2468), .ZN(n2465) );
  AND2_X1 U2642 ( .A1(n2513), .A2(n2318), .ZN(n2434) );
  AND2_X1 U2643 ( .A1(n2316), .A2(n2315), .ZN(n2314) );
  NAND2_X1 U2644 ( .A1(n2829), .A2(n2313), .ZN(n2312) );
  NAND2_X1 U2645 ( .A1(IR_REG_29__SCAN_IN), .A2(n2930), .ZN(n2315) );
  NAND2_X1 U2646 ( .A1(n2829), .A2(n2885), .ZN(n2886) );
  NAND2_X1 U2647 ( .A1(n2879), .A2(IR_REG_31__SCAN_IN), .ZN(n2881) );
  XNOR2_X1 U2648 ( .A(n2824), .B(IR_REG_22__SCAN_IN), .ZN(n4448) );
  INV_X1 U2649 ( .A(n4190), .ZN(n4905) );
  AND2_X1 U2650 ( .A1(n2649), .A2(n2668), .ZN(n4452) );
  NAND2_X1 U2651 ( .A1(n2280), .A2(IR_REG_0__SCAN_IN), .ZN(n2406) );
  NAND2_X1 U2652 ( .A1(n2375), .A2(n2373), .ZN(n3965) );
  NAND2_X1 U2653 ( .A1(n2326), .A2(n2325), .ZN(U3259) );
  NAND2_X1 U2654 ( .A1(n2327), .A2(n4744), .ZN(n2326) );
  AND2_X1 U2655 ( .A1(n2408), .A2(n2407), .ZN(n2325) );
  XNOR2_X1 U2656 ( .A(n2329), .B(n2328), .ZN(n2327) );
  OR2_X1 U2657 ( .A1(n4229), .A2(n4396), .ZN(n2918) );
  AND2_X1 U2658 ( .A1(n2394), .A2(n2288), .ZN(n2264) );
  AND2_X1 U2659 ( .A1(n2337), .A2(n3243), .ZN(n2265) );
  OR2_X1 U2660 ( .A1(n2363), .A2(n3759), .ZN(n2266) );
  NAND4_X1 U2661 ( .A1(n2532), .A2(n2531), .A3(n2530), .A4(n2529), .ZN(n4297)
         );
  INV_X1 U2662 ( .A(n4297), .ZN(n2447) );
  NOR2_X1 U2663 ( .A1(n3959), .A2(n2374), .ZN(n2373) );
  INV_X1 U2664 ( .A(n3686), .ZN(n2432) );
  OR2_X1 U2665 ( .A1(n4849), .A2(REG0_REG_29__SCAN_IN), .ZN(n2267) );
  INV_X1 U2666 ( .A(n3924), .ZN(n3051) );
  NAND4_X1 U2667 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .ZN(n3050)
         );
  OR2_X1 U2668 ( .A1(n4370), .A2(n2297), .ZN(n2268) );
  AND2_X1 U2669 ( .A1(n2818), .A2(n2507), .ZN(n2876) );
  AND2_X1 U2670 ( .A1(n2331), .A2(n2330), .ZN(n2269) );
  AND4_X1 U2671 ( .A1(n2733), .A2(n2505), .A3(n2504), .A4(n2503), .ZN(n2818)
         );
  OAI211_X1 U2672 ( .C1(n2829), .C2(n2317), .A(n2314), .B(n2312), .ZN(n2925)
         );
  AND2_X1 U2673 ( .A1(n3077), .A2(n3078), .ZN(n2270) );
  NAND3_X1 U2674 ( .A1(n2923), .A2(n2893), .A3(n2892), .ZN(n2980) );
  AND2_X1 U2675 ( .A1(n2574), .A2(n2509), .ZN(n2705) );
  AND2_X1 U2676 ( .A1(n3971), .A2(n2386), .ZN(n2271) );
  INV_X1 U2677 ( .A(n3269), .ZN(n2355) );
  AOI22_X1 U2678 ( .A1(n4816), .A2(n3947), .B1(n3899), .B2(n3176), .ZN(n3269)
         );
  NAND2_X1 U2679 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2761) );
  NOR2_X1 U2680 ( .A1(n4746), .A2(n4192), .ZN(n2272) );
  INV_X1 U2681 ( .A(n2397), .ZN(n2393) );
  NOR2_X1 U2682 ( .A1(n2400), .A2(n2398), .ZN(n2397) );
  AND2_X1 U2683 ( .A1(n3995), .A2(n3892), .ZN(n2273) );
  INV_X1 U2684 ( .A(n2492), .ZN(n2491) );
  NOR2_X1 U2685 ( .A1(n2495), .A2(n2493), .ZN(n2492) );
  NAND2_X1 U2686 ( .A1(n3891), .A2(n2998), .ZN(n2274) );
  AND2_X1 U2687 ( .A1(n2467), .A2(n2468), .ZN(n2275) );
  AND2_X1 U2688 ( .A1(n2353), .A2(n3269), .ZN(n2276) );
  AND2_X1 U2689 ( .A1(n2406), .A2(n2404), .ZN(n2277) );
  NOR2_X1 U2690 ( .A1(n4113), .A2(n3319), .ZN(n2278) );
  INV_X1 U2691 ( .A(n2455), .ZN(n2454) );
  NAND2_X1 U2692 ( .A1(n2683), .A2(n2456), .ZN(n2455) );
  INV_X1 U2693 ( .A(n2299), .ZN(n4264) );
  NOR2_X1 U2694 ( .A1(n4370), .A2(n4255), .ZN(n2299) );
  NAND2_X1 U2695 ( .A1(n2378), .A2(n2377), .ZN(n4017) );
  INV_X1 U2696 ( .A(n3248), .ZN(n3249) );
  NOR2_X1 U2697 ( .A1(n4101), .A2(n3973), .ZN(n2279) );
  INV_X1 U2698 ( .A(n3922), .ZN(n2387) );
  AND2_X1 U2699 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2280)
         );
  AND2_X1 U2700 ( .A1(n2718), .A2(n2682), .ZN(n2281) );
  NOR2_X1 U2701 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2733)
         );
  INV_X1 U2702 ( .A(IR_REG_29__SCAN_IN), .ZN(n2318) );
  XNOR2_X1 U2703 ( .A(n2881), .B(n2880), .ZN(n2891) );
  INV_X1 U2704 ( .A(n4824), .ZN(n2292) );
  XNOR2_X1 U2705 ( .A(n3948), .B(n3925), .ZN(n2282) );
  AND2_X1 U2706 ( .A1(n2359), .A2(n2357), .ZN(n4072) );
  NOR2_X1 U2707 ( .A1(n2388), .A2(n4042), .ZN(n2384) );
  INV_X1 U2708 ( .A(n2384), .ZN(n2377) );
  INV_X1 U2709 ( .A(n4084), .ZN(n2374) );
  AND2_X1 U2710 ( .A1(n4074), .A2(n4073), .ZN(n2283) );
  OR2_X1 U2711 ( .A1(n3776), .A2(n3998), .ZN(n2284) );
  AND2_X1 U2712 ( .A1(n3915), .A2(n2377), .ZN(n2285) );
  AND2_X1 U2713 ( .A1(n2373), .A2(n3952), .ZN(n2286) );
  AND2_X1 U2714 ( .A1(n2364), .A2(n3867), .ZN(n2287) );
  INV_X1 U2715 ( .A(n3695), .ZN(n2478) );
  INV_X1 U2716 ( .A(n2474), .ZN(n2473) );
  NAND2_X1 U2717 ( .A1(n3695), .A2(n2479), .ZN(n2474) );
  INV_X1 U2718 ( .A(n2765), .ZN(n2499) );
  NAND2_X1 U2719 ( .A1(n4832), .A2(n2622), .ZN(n3294) );
  NAND2_X1 U2720 ( .A1(n2878), .A2(IR_REG_31__SCAN_IN), .ZN(n2894) );
  NAND2_X1 U2721 ( .A1(n2443), .A2(n2633), .ZN(n3217) );
  OR2_X1 U2722 ( .A1(n3507), .A2(n3506), .ZN(n2288) );
  NOR2_X1 U2723 ( .A1(n3855), .A2(n2270), .ZN(n2289) );
  INV_X1 U2724 ( .A(n4840), .ZN(n2466) );
  AND2_X1 U2725 ( .A1(n2419), .A2(n2418), .ZN(n2290) );
  INV_X1 U2726 ( .A(IR_REG_0__SCAN_IN), .ZN(n2295) );
  INV_X1 U2727 ( .A(IR_REG_1__SCAN_IN), .ZN(n2405) );
  INV_X1 U2728 ( .A(n4694), .ZN(n2422) );
  AND2_X1 U2729 ( .A1(n4754), .A2(REG1_REG_18__SCAN_IN), .ZN(n2291) );
  INV_X1 U2730 ( .A(DATAI_0_), .ZN(n2296) );
  AND2_X1 U2731 ( .A1(n2980), .A2(n2939), .ZN(n3013) );
  MUX2_X1 U2732 ( .A(n2296), .B(n2295), .S(n2566), .Z(n3124) );
  NAND2_X2 U2733 ( .A1(n2524), .A2(n2294), .ZN(n2566) );
  NOR3_X2 U2734 ( .A1(n4370), .A2(n4255), .A3(n4243), .ZN(n4236) );
  AND2_X2 U2735 ( .A1(n2705), .A2(n2704), .ZN(n2877) );
  NAND2_X1 U2736 ( .A1(n2311), .A2(n3636), .ZN(n2867) );
  OAI21_X1 U2737 ( .B1(n3222), .B2(n2322), .A(n2319), .ZN(n3405) );
  OAI21_X1 U2738 ( .B1(n3222), .B2(n3619), .A(n3621), .ZN(n3342) );
  NAND2_X1 U2739 ( .A1(n2976), .A2(n2333), .ZN(n2330) );
  NAND2_X1 U2740 ( .A1(n2976), .A2(REG1_REG_3__SCAN_IN), .ZN(n2339) );
  NAND2_X1 U2741 ( .A1(n2339), .A2(n2337), .ZN(n2336) );
  NAND2_X1 U2742 ( .A1(n2336), .A2(n2973), .ZN(n2335) );
  OR2_X1 U2743 ( .A1(n2975), .A2(n2338), .ZN(n2337) );
  INV_X1 U2744 ( .A(n4453), .ZN(n2338) );
  XNOR2_X2 U2745 ( .A(n2340), .B(n2565), .ZN(n4142) );
  OAI21_X1 U2746 ( .B1(n4745), .B2(n2342), .A(n2341), .ZN(n4216) );
  NOR2_X1 U2747 ( .A1(n4687), .A2(n4686), .ZN(n4685) );
  INV_X1 U2748 ( .A(n3113), .ZN(n2356) );
  OR2_X1 U2749 ( .A1(n3855), .A2(n2352), .ZN(n2351) );
  OAI21_X1 U2750 ( .B1(n3855), .B2(n2350), .A(n2348), .ZN(n2347) );
  INV_X1 U2751 ( .A(n3268), .ZN(n2354) );
  NAND3_X1 U2752 ( .A1(n2502), .A2(n3743), .A3(n2287), .ZN(n2359) );
  NAND2_X1 U2753 ( .A1(n2502), .A2(n3743), .ZN(n4026) );
  OAI21_X1 U2754 ( .B1(n2362), .B2(n2361), .A(n3759), .ZN(n3868) );
  NAND2_X1 U2755 ( .A1(n3743), .A2(n2364), .ZN(n2362) );
  INV_X1 U2756 ( .A(n3867), .ZN(n2363) );
  OAI211_X1 U2757 ( .C1(n4087), .C2(n2369), .A(n2367), .B(n2366), .ZN(n3958)
         );
  NAND2_X1 U2758 ( .A1(n4087), .A2(n2286), .ZN(n2366) );
  OAI21_X1 U2759 ( .B1(n3952), .B2(n2371), .A(n2368), .ZN(n2367) );
  OAI21_X1 U2760 ( .B1(n2373), .B2(n3952), .A(n2371), .ZN(n2368) );
  OR2_X2 U2761 ( .A1(n4087), .A2(n4085), .ZN(n2375) );
  NAND2_X1 U2762 ( .A1(n2376), .A2(n2381), .ZN(n3928) );
  NAND2_X1 U2763 ( .A1(n3968), .A2(n2285), .ZN(n2376) );
  NOR2_X1 U2764 ( .A1(n2387), .A2(n2388), .ZN(n2386) );
  INV_X1 U2765 ( .A(n3923), .ZN(n2388) );
  NAND2_X1 U2766 ( .A1(n3429), .A2(n2264), .ZN(n2389) );
  NAND2_X2 U2767 ( .A1(n2389), .A2(n2390), .ZN(n3742) );
  OAI21_X1 U2768 ( .B1(n3429), .B2(n3428), .A(n3427), .ZN(n3502) );
  NAND2_X1 U2769 ( .A1(n3428), .A2(n3427), .ZN(n2399) );
  NAND2_X1 U2770 ( .A1(n2409), .A2(n4761), .ZN(n2408) );
  XNOR2_X1 U2771 ( .A(n2410), .B(n4755), .ZN(n2409) );
  INV_X1 U2772 ( .A(n4753), .ZN(n2412) );
  INV_X1 U2775 ( .A(n4177), .ZN(n2423) );
  NAND2_X1 U2776 ( .A1(n2428), .A2(n2427), .ZN(n3785) );
  INV_X1 U2777 ( .A(n3134), .ZN(n2433) );
  NAND2_X1 U2778 ( .A1(n2430), .A2(n2429), .ZN(n2600) );
  NAND2_X1 U2779 ( .A1(n3134), .A2(n2587), .ZN(n2430) );
  NAND2_X1 U2780 ( .A1(n2829), .A2(n2434), .ZN(n2931) );
  NAND2_X1 U2781 ( .A1(n4832), .A2(n2436), .ZN(n2435) );
  NAND2_X1 U2782 ( .A1(n2435), .A2(n2438), .ZN(n3341) );
  AOI21_X1 U2783 ( .B1(n3326), .B2(n2281), .A(n2451), .ZN(n3476) );
  NAND2_X1 U2784 ( .A1(n2458), .A2(n2267), .ZN(n2914) );
  NAND2_X1 U2785 ( .A1(n2460), .A2(n2459), .ZN(n2458) );
  NAND2_X1 U2786 ( .A1(n2465), .A2(n4840), .ZN(n2459) );
  INV_X1 U2787 ( .A(n2461), .ZN(n2460) );
  NAND3_X1 U2788 ( .A1(n2468), .A2(n2467), .A3(n2477), .ZN(n2463) );
  INV_X1 U2789 ( .A(n4231), .ZN(n2477) );
  NAND2_X1 U2790 ( .A1(n2480), .A2(n2481), .ZN(n2798) );
  NAND2_X1 U2791 ( .A1(n3556), .A2(n2482), .ZN(n2480) );
  XNOR2_X1 U2792 ( .A(n3244), .B(n2973), .ZN(n2974) );
  OAI22_X2 U2793 ( .A1(n3280), .A2(n3279), .B1(n3278), .B2(n3277), .ZN(n3315)
         );
  AOI21_X2 U2794 ( .B1(n3271), .B2(n2355), .A(n3270), .ZN(n3280) );
  NAND2_X1 U2795 ( .A1(n2560), .A2(REG1_REG_1__SCAN_IN), .ZN(n2544) );
  OAI21_X1 U2796 ( .B1(n2961), .B2(n4142), .A(n4134), .ZN(n2970) );
  NAND2_X1 U2797 ( .A1(n2552), .A2(REG0_REG_0__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U2798 ( .A1(n2552), .A2(REG0_REG_1__SCAN_IN), .ZN(n2545) );
  NOR2_X2 U2799 ( .A1(n3057), .A2(n3056), .ZN(n3854) );
  NOR2_X1 U2800 ( .A1(n2760), .A2(n2759), .ZN(n2500) );
  OAI22_X1 U2801 ( .A1(n3174), .A2(n2609), .B1(n3176), .B2(n4816), .ZN(n4829)
         );
  INV_X1 U2802 ( .A(n2980), .ZN(n2982) );
  AND2_X2 U2803 ( .A1(n4447), .A2(n2925), .ZN(n2558) );
  OR2_X1 U2804 ( .A1(n3742), .A2(n3741), .ZN(n2502) );
  INV_X1 U2805 ( .A(IR_REG_22__SCAN_IN), .ZN(n2506) );
  AND2_X1 U2806 ( .A1(n2821), .A2(n2506), .ZN(n2507) );
  AND2_X1 U2807 ( .A1(n2970), .A2(n4453), .ZN(n2971) );
  AND2_X1 U2808 ( .A1(n4273), .A2(n3691), .ZN(n3652) );
  INV_X1 U2809 ( .A(n3243), .ZN(n2973) );
  AND2_X1 U2810 ( .A1(REG3_REG_19__SCAN_IN), .A2(n2748), .ZN(n2747) );
  AND2_X1 U2811 ( .A1(n2832), .A2(n2830), .ZN(n2513) );
  AND2_X1 U2812 ( .A1(n3758), .A2(n4030), .ZN(n3759) );
  NAND2_X1 U2813 ( .A1(n2982), .A2(REG1_REG_0__SCAN_IN), .ZN(n2983) );
  NAND2_X1 U2814 ( .A1(n2774), .A2(REG3_REG_22__SCAN_IN), .ZN(n2790) );
  OR2_X1 U2815 ( .A1(n4278), .A2(n4265), .ZN(n4239) );
  OR3_X1 U2816 ( .A1(n2539), .A2(n2526), .A3(n2525), .ZN(n2527) );
  NAND2_X1 U2817 ( .A1(n2855), .A2(n3704), .ZN(n3836) );
  NAND2_X1 U2818 ( .A1(n2727), .A2(REG3_REG_17__SCAN_IN), .ZN(n2740) );
  NOR2_X1 U2819 ( .A1(n2661), .A2(n2660), .ZN(n2672) );
  INV_X1 U2820 ( .A(n3678), .ZN(n3404) );
  AND3_X1 U2821 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2588) );
  INV_X1 U2822 ( .A(n3540), .ZN(n3769) );
  NAND2_X1 U2823 ( .A1(n3183), .A2(n3182), .ZN(n4825) );
  OR2_X1 U2824 ( .A1(n2668), .A2(IR_REG_10__SCAN_IN), .ZN(n2669) );
  AND2_X1 U2825 ( .A1(n3982), .A2(n3979), .ZN(n3357) );
  INV_X1 U2826 ( .A(n3133), .ZN(n3860) );
  INV_X1 U2827 ( .A(n3023), .ZN(n3026) );
  AND2_X1 U2828 ( .A1(n2792), .A2(n2791), .ZN(n4349) );
  INV_X1 U2829 ( .A(n3253), .ZN(n3254) );
  NAND2_X1 U2830 ( .A1(n4151), .A2(n4711), .ZN(n4152) );
  NOR2_X1 U2831 ( .A1(n2735), .A2(n2759), .ZN(n2745) );
  AND2_X1 U2832 ( .A1(n4239), .A2(n3649), .ZN(n4261) );
  OR2_X1 U2833 ( .A1(n4102), .A2(n4064), .ZN(n4334) );
  INV_X1 U2834 ( .A(n3471), .ZN(n4034) );
  NAND2_X1 U2835 ( .A1(n3402), .A2(n2671), .ZN(n3326) );
  OR2_X1 U2836 ( .A1(n2651), .A2(n3984), .ZN(n2661) );
  INV_X1 U2837 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2610) );
  INV_X1 U2838 ( .A(n3408), .ZN(n3370) );
  AND2_X1 U2839 ( .A1(n2888), .A2(n2892), .ZN(n2936) );
  INV_X1 U2840 ( .A(IR_REG_23__SCAN_IN), .ZN(n2895) );
  INV_X1 U2841 ( .A(n3881), .ZN(n3998) );
  INV_X1 U2842 ( .A(n4060), .ZN(n4062) );
  INV_X1 U2843 ( .A(n4097), .ZN(n4898) );
  OR2_X1 U2844 ( .A1(n2708), .A2(n2707), .ZN(n2719) );
  INV_X1 U2845 ( .A(n4125), .ZN(n4121) );
  AND2_X1 U2846 ( .A1(n4228), .A2(n2804), .ZN(n4235) );
  AND2_X1 U2847 ( .A1(n2803), .A2(n2516), .ZN(n4260) );
  NOR2_X1 U2848 ( .A1(n2611), .A2(n2610), .ZN(n2623) );
  INV_X1 U2849 ( .A(n4871), .ZN(n4908) );
  AND2_X1 U2850 ( .A1(n4765), .A2(n2872), .ZN(n4794) );
  AND2_X1 U2851 ( .A1(n2946), .A2(n2949), .ZN(n4757) );
  NAND4_X1 U2852 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n4278)
         );
  NAND4_X1 U2853 ( .A1(n2796), .A2(n2795), .A3(n2794), .A4(n2793), .ZN(n4101)
         );
  OR2_X1 U2854 ( .A1(n4229), .A2(n4442), .ZN(n2913) );
  OR2_X1 U2855 ( .A1(n2915), .A2(n3005), .ZN(n4414) );
  INV_X1 U2856 ( .A(n4828), .ZN(n4450) );
  INV_X1 U2857 ( .A(n4705), .ZN(n4867) );
  XNOR2_X1 U2858 ( .A(n2583), .B(IR_REG_3__SCAN_IN), .ZN(n4453) );
  NOR2_X1 U2859 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2508)
         );
  NAND3_X1 U2860 ( .A1(n2694), .A2(n2691), .A3(n2510), .ZN(n2512) );
  NAND2_X1 U2861 ( .A1(n2692), .A2(n2693), .ZN(n2511) );
  NOR2_X1 U2862 ( .A1(n2522), .A2(IR_REG_27__SCAN_IN), .ZN(n2830) );
  CLKBUF_X3 U2863 ( .A(n2559), .Z(n3641) );
  NAND2_X1 U2864 ( .A1(n3641), .A2(REG2_REG_27__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U2865 ( .A1(n3640), .A2(REG1_REG_27__SCAN_IN), .ZN(n2520) );
  INV_X1 U2866 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2660) );
  INV_X1 U2867 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2707) );
  INV_X1 U2868 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4624) );
  INV_X1 U2869 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4076) );
  INV_X1 U2870 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4608) );
  INV_X1 U2871 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2526) );
  INV_X1 U2872 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2525) );
  INV_X1 U2873 ( .A(n2527), .ZN(n2515) );
  NAND2_X1 U2874 ( .A1(n2515), .A2(REG3_REG_27__SCAN_IN), .ZN(n2803) );
  INV_X1 U2875 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U2876 ( .A1(n2527), .A2(n4503), .ZN(n2516) );
  NAND2_X1 U2877 ( .A1(n2684), .A2(n4260), .ZN(n2519) );
  NOR2_X2 U2878 ( .A1(n4447), .A2(n2925), .ZN(n2552) );
  NAND2_X1 U2879 ( .A1(n3642), .A2(REG0_REG_27__SCAN_IN), .ZN(n2518) );
  INV_X1 U2880 ( .A(n4278), .ZN(n4246) );
  NAND2_X1 U2882 ( .A1(n3646), .A2(DATAI_27_), .ZN(n4265) );
  INV_X1 U2883 ( .A(n4265), .ZN(n4255) );
  NAND2_X1 U2884 ( .A1(n3641), .A2(REG2_REG_26__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U2885 ( .A1(n3640), .A2(REG1_REG_26__SCAN_IN), .ZN(n2531) );
  OAI21_X1 U2886 ( .B1(n2539), .B2(n2526), .A(n2525), .ZN(n2528) );
  AND2_X1 U2887 ( .A1(n2528), .A2(n2527), .ZN(n4088) );
  NAND2_X1 U2888 ( .A1(n2684), .A2(n4088), .ZN(n2530) );
  NAND2_X1 U2889 ( .A1(n3642), .A2(REG0_REG_26__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U2890 ( .A1(n3646), .A2(DATAI_26_), .ZN(n4283) );
  INV_X1 U2891 ( .A(n4283), .ZN(n4091) );
  NAND2_X1 U2892 ( .A1(n3641), .A2(REG2_REG_25__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U2893 ( .A1(n3640), .A2(REG1_REG_25__SCAN_IN), .ZN(n2535) );
  XNOR2_X1 U2894 ( .A(n2539), .B(REG3_REG_25__SCAN_IN), .ZN(n4304) );
  NAND2_X1 U2895 ( .A1(n2684), .A2(n4304), .ZN(n2534) );
  NAND2_X1 U2896 ( .A1(n3642), .A2(REG0_REG_25__SCAN_IN), .ZN(n2533) );
  NAND4_X1 U2897 ( .A1(n2536), .A2(n2535), .A3(n2534), .A4(n2533), .ZN(n4316)
         );
  INV_X1 U2898 ( .A(n4316), .ZN(n3927) );
  NAND2_X1 U2899 ( .A1(n3646), .A2(DATAI_25_), .ZN(n4301) );
  INV_X1 U2900 ( .A(n4301), .ZN(n4296) );
  NAND2_X1 U2901 ( .A1(n3641), .A2(REG2_REG_24__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U2902 ( .A1(n3640), .A2(REG1_REG_24__SCAN_IN), .ZN(n2542) );
  INV_X1 U2903 ( .A(n2537), .ZN(n2792) );
  INV_X1 U2904 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U2905 ( .A1(n2792), .A2(n4523), .ZN(n2538) );
  AND2_X1 U2906 ( .A1(n2539), .A2(n2538), .ZN(n4044) );
  NAND2_X1 U2907 ( .A1(n2684), .A2(n4044), .ZN(n2541) );
  NAND2_X1 U2908 ( .A1(n3642), .A2(REG0_REG_24__SCAN_IN), .ZN(n2540) );
  NAND4_X1 U2909 ( .A1(n2543), .A2(n2542), .A3(n2541), .A4(n2540), .ZN(n4342)
         );
  INV_X1 U2910 ( .A(n4342), .ZN(n4300) );
  NAND2_X1 U2911 ( .A1(n3646), .A2(DATAI_24_), .ZN(n4324) );
  INV_X1 U2912 ( .A(n4324), .ZN(n4315) );
  NAND2_X1 U2913 ( .A1(n2559), .A2(REG2_REG_1__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U2914 ( .A1(n2558), .A2(REG3_REG_1__SCAN_IN), .ZN(n2546) );
  NAND4_X2 U2915 ( .A1(n2547), .A2(n2546), .A3(n2545), .A4(n2544), .ZN(n2996)
         );
  INV_X1 U2916 ( .A(DATAI_1_), .ZN(n2550) );
  INV_X1 U2917 ( .A(n2548), .ZN(n2549) );
  MUX2_X1 U2918 ( .A(n2550), .B(n4125), .S(n2566), .Z(n2997) );
  NAND2_X1 U2919 ( .A1(n2996), .A2(n2997), .ZN(n3600) );
  INV_X1 U2920 ( .A(n2996), .ZN(n2551) );
  NAND2_X1 U2921 ( .A1(n2998), .A2(n2551), .ZN(n3603) );
  NAND2_X1 U2922 ( .A1(n2560), .A2(REG1_REG_0__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U2923 ( .A1(n2558), .A2(REG3_REG_0__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U2924 ( .A1(n2559), .A2(REG2_REG_0__SCAN_IN), .ZN(n2553) );
  NAND4_X2 U2925 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n4120)
         );
  AND2_X1 U2926 ( .A1(n4120), .A2(n3126), .ZN(n3092) );
  NAND2_X1 U2927 ( .A1(n4118), .A2(n2998), .ZN(n2557) );
  NAND2_X1 U2928 ( .A1(n2558), .A2(REG3_REG_2__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U2929 ( .A1(n2559), .A2(REG2_REG_2__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U2930 ( .A1(n2560), .A2(REG1_REG_2__SCAN_IN), .ZN(n2561) );
  INV_X1 U2931 ( .A(DATAI_2_), .ZN(n2567) );
  MUX2_X1 U2932 ( .A(n2567), .B(n4142), .S(n2566), .Z(n3165) );
  NAND2_X1 U2933 ( .A1(n3034), .A2(n3165), .ZN(n3607) );
  NAND2_X1 U2934 ( .A1(n3162), .A2(n3685), .ZN(n3161) );
  OR2_X1 U2935 ( .A1(n3034), .A2(n3172), .ZN(n2568) );
  NAND2_X1 U2936 ( .A1(n3161), .A2(n2568), .ZN(n3194) );
  NAND2_X1 U2937 ( .A1(n2560), .A2(REG1_REG_3__SCAN_IN), .ZN(n2573) );
  INV_X1 U2938 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U2939 ( .A1(n2558), .A2(n2569), .ZN(n2572) );
  NAND2_X1 U2940 ( .A1(n2559), .A2(REG2_REG_3__SCAN_IN), .ZN(n2570) );
  OR2_X1 U2941 ( .A1(n2574), .A2(n2930), .ZN(n2583) );
  MUX2_X1 U2942 ( .A(DATAI_3_), .B(n4453), .S(n3639), .Z(n3199) );
  NAND2_X1 U2943 ( .A1(n3050), .A2(n3199), .ZN(n2575) );
  NAND2_X1 U2944 ( .A1(n3194), .A2(n2575), .ZN(n2577) );
  OR2_X1 U2945 ( .A1(n3050), .A2(n3199), .ZN(n2576) );
  NAND2_X1 U2946 ( .A1(n2577), .A2(n2576), .ZN(n3134) );
  NAND2_X1 U2947 ( .A1(n3641), .A2(REG2_REG_4__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U2948 ( .A1(n2560), .A2(REG1_REG_4__SCAN_IN), .ZN(n2581) );
  INV_X1 U2949 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2578) );
  XNOR2_X1 U2950 ( .A(n2578), .B(REG3_REG_3__SCAN_IN), .ZN(n3858) );
  NAND2_X1 U2951 ( .A1(n2558), .A2(n3858), .ZN(n2580) );
  NAND2_X1 U2952 ( .A1(n2552), .A2(REG0_REG_4__SCAN_IN), .ZN(n2579) );
  INV_X1 U2953 ( .A(DATAI_4_), .ZN(n2586) );
  NAND2_X1 U2954 ( .A1(n2583), .A2(n4641), .ZN(n2584) );
  NAND2_X1 U2955 ( .A1(n2584), .A2(IR_REG_31__SCAN_IN), .ZN(n2585) );
  XNOR2_X1 U2956 ( .A(n2585), .B(n4537), .ZN(n3243) );
  MUX2_X1 U2957 ( .A(n2586), .B(n3243), .S(n3639), .Z(n3133) );
  OR2_X1 U2958 ( .A1(n4116), .A2(n3133), .ZN(n3610) );
  NAND2_X1 U2959 ( .A1(n4116), .A2(n3133), .ZN(n3614) );
  NAND2_X1 U2960 ( .A1(n3610), .A2(n3614), .ZN(n3686) );
  NAND2_X1 U2961 ( .A1(n4116), .A2(n3860), .ZN(n2587) );
  INV_X1 U2962 ( .A(n2588), .ZN(n2601) );
  INV_X1 U2963 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U2964 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2589) );
  NAND2_X1 U2965 ( .A1(n2590), .A2(n2589), .ZN(n2591) );
  NAND2_X1 U2966 ( .A1(n2601), .A2(n2591), .ZN(n3154) );
  INV_X1 U2967 ( .A(n3154), .ZN(n2592) );
  NAND2_X1 U2968 ( .A1(n2558), .A2(n2592), .ZN(n2596) );
  NAND2_X1 U2969 ( .A1(n3641), .A2(REG2_REG_5__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U2970 ( .A1(n3642), .A2(REG0_REG_5__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U2971 ( .A1(n2560), .A2(REG1_REG_5__SCAN_IN), .ZN(n2593) );
  NAND4_X1 U2972 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n4115)
         );
  OR2_X1 U2973 ( .A1(n2705), .A2(n2930), .ZN(n2597) );
  XNOR2_X1 U2974 ( .A(n2597), .B(IR_REG_5__SCAN_IN), .ZN(n3247) );
  MUX2_X1 U2975 ( .A(DATAI_5_), .B(n3247), .S(n3639), .Z(n3153) );
  OR2_X1 U2976 ( .A1(n4115), .A2(n3153), .ZN(n2598) );
  NAND2_X1 U2977 ( .A1(n4115), .A2(n3153), .ZN(n2599) );
  NAND2_X1 U2978 ( .A1(n2600), .A2(n2599), .ZN(n3174) );
  NAND2_X1 U2979 ( .A1(n2560), .A2(REG1_REG_6__SCAN_IN), .ZN(n2606) );
  INV_X1 U2980 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U2981 ( .A1(n2601), .A2(n3117), .ZN(n2602) );
  AND2_X1 U2982 ( .A1(n2602), .A2(n2611), .ZN(n4802) );
  NAND2_X1 U2983 ( .A1(n2558), .A2(n4802), .ZN(n2605) );
  NAND2_X1 U2984 ( .A1(n3642), .A2(REG0_REG_6__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U2985 ( .A1(n3641), .A2(REG2_REG_6__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U2986 ( .A1(n2705), .A2(n2607), .ZN(n2645) );
  NAND2_X1 U2987 ( .A1(n2645), .A2(IR_REG_31__SCAN_IN), .ZN(n2608) );
  XNOR2_X1 U2988 ( .A(n2608), .B(IR_REG_6__SCAN_IN), .ZN(n3250) );
  MUX2_X1 U2989 ( .A(DATAI_6_), .B(n3250), .S(n3639), .Z(n3176) );
  AND2_X1 U2990 ( .A1(n4816), .A2(n3176), .ZN(n2609) );
  INV_X1 U2991 ( .A(n4829), .ZN(n2621) );
  NAND2_X1 U2992 ( .A1(n2560), .A2(REG1_REG_7__SCAN_IN), .ZN(n2617) );
  AND2_X1 U2993 ( .A1(n2611), .A2(n2610), .ZN(n2612) );
  OR2_X1 U2994 ( .A1(n2612), .A2(n2623), .ZN(n4838) );
  INV_X1 U2995 ( .A(n4838), .ZN(n2613) );
  NAND2_X1 U2996 ( .A1(n2558), .A2(n2613), .ZN(n2616) );
  NAND2_X1 U2997 ( .A1(n3642), .A2(REG0_REG_7__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U2998 ( .A1(n3641), .A2(REG2_REG_7__SCAN_IN), .ZN(n2614) );
  NAND4_X1 U2999 ( .A1(n2617), .A2(n2616), .A3(n2615), .A4(n2614), .ZN(n4114)
         );
  OR2_X1 U3000 ( .A1(n2645), .A2(IR_REG_6__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U3001 ( .A1(n2618), .A2(IR_REG_31__SCAN_IN), .ZN(n2629) );
  XNOR2_X1 U3002 ( .A(n2629), .B(IR_REG_7__SCAN_IN), .ZN(n4673) );
  MUX2_X1 U3003 ( .A(DATAI_7_), .B(n4673), .S(n3639), .Z(n4824) );
  NAND2_X1 U3004 ( .A1(n4114), .A2(n4824), .ZN(n2622) );
  OR2_X1 U3005 ( .A1(n4114), .A2(n4824), .ZN(n2619) );
  NAND2_X1 U3006 ( .A1(n2622), .A2(n2619), .ZN(n4830) );
  INV_X1 U3007 ( .A(n4830), .ZN(n2620) );
  NAND2_X1 U3008 ( .A1(n2621), .A2(n2620), .ZN(n4832) );
  OR2_X1 U3009 ( .A1(n2623), .A2(REG3_REG_8__SCAN_IN), .ZN(n2624) );
  AND2_X1 U3010 ( .A1(n2634), .A2(n2624), .ZN(n4851) );
  NAND2_X1 U3011 ( .A1(n2558), .A2(n4851), .ZN(n2628) );
  NAND2_X1 U3012 ( .A1(n3641), .A2(REG2_REG_8__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U3013 ( .A1(n3642), .A2(REG0_REG_8__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U3014 ( .A1(n3640), .A2(REG1_REG_8__SCAN_IN), .ZN(n2625) );
  NAND4_X1 U3015 ( .A1(n2628), .A2(n2627), .A3(n2626), .A4(n2625), .ZN(n4814)
         );
  NAND2_X1 U3016 ( .A1(n2629), .A2(n2643), .ZN(n2630) );
  NAND2_X1 U3017 ( .A1(n2630), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  XNOR2_X1 U3018 ( .A(n2631), .B(IR_REG_8__SCAN_IN), .ZN(n3253) );
  MUX2_X1 U3019 ( .A(DATAI_8_), .B(n3253), .S(n3639), .Z(n3302) );
  OR2_X1 U3020 ( .A1(n4814), .A2(n3302), .ZN(n2632) );
  NAND2_X1 U3021 ( .A1(n4814), .A2(n3302), .ZN(n2633) );
  NAND2_X1 U3022 ( .A1(n3640), .A2(REG1_REG_9__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3023 ( .A1(n2634), .A2(n4550), .ZN(n2635) );
  NAND2_X1 U3024 ( .A1(n2651), .A2(n2635), .ZN(n3322) );
  INV_X1 U3025 ( .A(n3322), .ZN(n2636) );
  NAND2_X1 U3026 ( .A1(n2684), .A2(n2636), .ZN(n2639) );
  NAND2_X1 U3027 ( .A1(n3642), .A2(REG0_REG_9__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U3028 ( .A1(n3641), .A2(REG2_REG_9__SCAN_IN), .ZN(n2637) );
  NAND4_X1 U3029 ( .A1(n2640), .A2(n2639), .A3(n2638), .A4(n2637), .ZN(n4113)
         );
  INV_X1 U3030 ( .A(IR_REG_6__SCAN_IN), .ZN(n2642) );
  INV_X1 U3031 ( .A(IR_REG_8__SCAN_IN), .ZN(n2641) );
  NAND3_X1 U3032 ( .A1(n2643), .A2(n2642), .A3(n2641), .ZN(n2644) );
  NOR2_X1 U3033 ( .A1(n2645), .A2(n2644), .ZN(n2648) );
  OR2_X1 U3034 ( .A1(n2648), .A2(n2930), .ZN(n2646) );
  MUX2_X1 U3035 ( .A(n2646), .B(IR_REG_31__SCAN_IN), .S(n2647), .Z(n2649) );
  NAND2_X1 U3036 ( .A1(n2648), .A2(n2647), .ZN(n2668) );
  MUX2_X1 U3037 ( .A(DATAI_9_), .B(n4452), .S(n3639), .Z(n3319) );
  AND2_X1 U3038 ( .A1(n4113), .A2(n3319), .ZN(n2650) );
  NAND2_X1 U3039 ( .A1(n2651), .A2(n3984), .ZN(n2652) );
  AND2_X1 U3040 ( .A1(n2661), .A2(n2652), .ZN(n4860) );
  NAND2_X1 U3041 ( .A1(n2684), .A2(n4860), .ZN(n2656) );
  NAND2_X1 U3042 ( .A1(n3641), .A2(REG2_REG_10__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3043 ( .A1(n3642), .A2(REG0_REG_10__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3044 ( .A1(n3640), .A2(REG1_REG_10__SCAN_IN), .ZN(n2653) );
  NAND4_X1 U3045 ( .A1(n2656), .A2(n2655), .A3(n2654), .A4(n2653), .ZN(n4112)
         );
  NAND2_X1 U3046 ( .A1(n2668), .A2(IR_REG_31__SCAN_IN), .ZN(n2657) );
  XNOR2_X1 U3047 ( .A(n2657), .B(IR_REG_10__SCAN_IN), .ZN(n4694) );
  MUX2_X1 U3048 ( .A(DATAI_10_), .B(n4694), .S(n3639), .Z(n3985) );
  NOR2_X1 U3049 ( .A1(n4112), .A2(n3985), .ZN(n2659) );
  NAND2_X1 U3050 ( .A1(n4112), .A2(n3985), .ZN(n2658) );
  OAI21_X1 U3051 ( .B1(n3341), .B2(n2659), .A(n2658), .ZN(n3400) );
  AND2_X1 U3052 ( .A1(n2661), .A2(n2660), .ZN(n2662) );
  OR2_X1 U3053 ( .A1(n2662), .A2(n2672), .ZN(n4876) );
  INV_X1 U3054 ( .A(n4876), .ZN(n2663) );
  NAND2_X1 U3055 ( .A1(n2684), .A2(n2663), .ZN(n2667) );
  NAND2_X1 U3056 ( .A1(n3641), .A2(REG2_REG_11__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3057 ( .A1(n3642), .A2(REG0_REG_11__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3058 ( .A1(n3640), .A2(REG1_REG_11__SCAN_IN), .ZN(n2664) );
  NAND4_X1 U3059 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(n4111)
         );
  INV_X1 U3060 ( .A(DATAI_11_), .ZN(n2670) );
  NAND2_X1 U3061 ( .A1(n2669), .A2(IR_REG_31__SCAN_IN), .ZN(n2679) );
  XNOR2_X1 U3062 ( .A(n2679), .B(IR_REG_11__SCAN_IN), .ZN(n4705) );
  MUX2_X1 U3063 ( .A(n2670), .B(n4867), .S(n3639), .Z(n3408) );
  OR2_X1 U3064 ( .A1(n4111), .A2(n3408), .ZN(n3327) );
  NAND2_X1 U3065 ( .A1(n4111), .A2(n3408), .ZN(n3329) );
  NAND2_X1 U3066 ( .A1(n3327), .A2(n3329), .ZN(n3678) );
  OR2_X1 U3067 ( .A1(n4111), .A2(n3370), .ZN(n2671) );
  NAND2_X1 U3068 ( .A1(n3641), .A2(REG2_REG_12__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U3069 ( .A1(n3640), .A2(REG1_REG_12__SCAN_IN), .ZN(n2676) );
  NOR2_X1 U3070 ( .A1(n2672), .A2(REG3_REG_12__SCAN_IN), .ZN(n2673) );
  OR2_X1 U3071 ( .A1(n2685), .A2(n2673), .ZN(n3439) );
  INV_X1 U3072 ( .A(n3439), .ZN(n3334) );
  NAND2_X1 U3073 ( .A1(n2684), .A2(n3334), .ZN(n2675) );
  NAND2_X1 U3074 ( .A1(n3642), .A2(REG0_REG_12__SCAN_IN), .ZN(n2674) );
  NAND4_X1 U3075 ( .A1(n2677), .A2(n2676), .A3(n2675), .A4(n2674), .ZN(n4110)
         );
  INV_X1 U3076 ( .A(IR_REG_11__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U3077 ( .A1(n2679), .A2(n2678), .ZN(n2680) );
  NAND2_X1 U3078 ( .A1(n2680), .A2(IR_REG_31__SCAN_IN), .ZN(n2681) );
  XNOR2_X1 U3079 ( .A(n2681), .B(IR_REG_12__SCAN_IN), .ZN(n4161) );
  MUX2_X1 U3080 ( .A(DATAI_12_), .B(n4161), .S(n3639), .Z(n3436) );
  NAND2_X1 U3081 ( .A1(n4110), .A2(n3436), .ZN(n2682) );
  OR2_X1 U3082 ( .A1(n4110), .A2(n3436), .ZN(n2683) );
  NAND2_X1 U3083 ( .A1(n3641), .A2(REG2_REG_13__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3084 ( .A1(n3640), .A2(REG1_REG_13__SCAN_IN), .ZN(n2689) );
  NOR2_X1 U3085 ( .A1(n2685), .A2(REG3_REG_13__SCAN_IN), .ZN(n2686) );
  OR2_X1 U3086 ( .A1(n2698), .A2(n2686), .ZN(n3512) );
  INV_X1 U3087 ( .A(n3512), .ZN(n3392) );
  NAND2_X1 U3088 ( .A1(n2684), .A2(n3392), .ZN(n2688) );
  NAND2_X1 U3089 ( .A1(n3642), .A2(REG0_REG_13__SCAN_IN), .ZN(n2687) );
  NAND4_X1 U3090 ( .A1(n2690), .A2(n2689), .A3(n2688), .A4(n2687), .ZN(n4109)
         );
  AND4_X1 U3091 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), .ZN(n2695)
         );
  NAND2_X1 U3092 ( .A1(n2705), .A2(n2695), .ZN(n2696) );
  NAND2_X1 U3093 ( .A1(n2696), .A2(IR_REG_31__SCAN_IN), .ZN(n2697) );
  XNOR2_X1 U3094 ( .A(n2697), .B(IR_REG_13__SCAN_IN), .ZN(n4164) );
  MUX2_X1 U3095 ( .A(DATAI_13_), .B(n4164), .S(n3639), .Z(n3509) );
  NOR2_X1 U3096 ( .A1(n4109), .A2(n3509), .ZN(n3377) );
  NAND2_X1 U3097 ( .A1(n3640), .A2(REG1_REG_14__SCAN_IN), .ZN(n2703) );
  NAND2_X1 U3098 ( .A1(n3641), .A2(REG2_REG_14__SCAN_IN), .ZN(n2702) );
  OR2_X1 U3099 ( .A1(n2698), .A2(REG3_REG_14__SCAN_IN), .ZN(n2699) );
  AND2_X1 U3100 ( .A1(n2699), .A2(n2708), .ZN(n3454) );
  NAND2_X1 U3101 ( .A1(n2684), .A2(n3454), .ZN(n2701) );
  NAND2_X1 U3102 ( .A1(n3642), .A2(REG0_REG_14__SCAN_IN), .ZN(n2700) );
  NAND4_X1 U3103 ( .A1(n2703), .A2(n2702), .A3(n2701), .A4(n2700), .ZN(n4886)
         );
  INV_X1 U3104 ( .A(DATAI_14_), .ZN(n4480) );
  NAND2_X1 U3105 ( .A1(n2705), .A2(n2704), .ZN(n2817) );
  NAND2_X1 U3106 ( .A1(n2817), .A2(IR_REG_31__SCAN_IN), .ZN(n2762) );
  INV_X1 U3107 ( .A(IR_REG_14__SCAN_IN), .ZN(n2706) );
  XNOR2_X1 U3108 ( .A(n2762), .B(n2706), .ZN(n4172) );
  MUX2_X1 U3109 ( .A(n4480), .B(n4172), .S(n3639), .Z(n3452) );
  OR2_X1 U3110 ( .A1(n4886), .A2(n3452), .ZN(n3593) );
  NAND2_X1 U3111 ( .A1(n4886), .A2(n3452), .ZN(n3597) );
  NAND2_X1 U3112 ( .A1(n3593), .A2(n3597), .ZN(n3688) );
  NAND2_X1 U3113 ( .A1(n3640), .A2(REG1_REG_15__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U3114 ( .A1(n2708), .A2(n2707), .ZN(n2709) );
  NAND2_X1 U3115 ( .A1(n2719), .A2(n2709), .ZN(n4902) );
  INV_X1 U3116 ( .A(n4902), .ZN(n3495) );
  NAND2_X1 U3117 ( .A1(n2684), .A2(n3495), .ZN(n2712) );
  NAND2_X1 U3118 ( .A1(n3642), .A2(REG0_REG_15__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3119 ( .A1(n3641), .A2(REG2_REG_15__SCAN_IN), .ZN(n2710) );
  NAND4_X1 U3120 ( .A1(n2713), .A2(n2712), .A3(n2711), .A4(n2710), .ZN(n4108)
         );
  NAND2_X1 U3121 ( .A1(n2762), .A2(n2761), .ZN(n2735) );
  OR2_X1 U3122 ( .A1(n2735), .A2(IR_REG_15__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3123 ( .A1(n2735), .A2(IR_REG_15__SCAN_IN), .ZN(n2714) );
  AND2_X1 U3124 ( .A1(n2724), .A2(n2714), .ZN(n4186) );
  MUX2_X1 U3125 ( .A(DATAI_15_), .B(n4186), .S(n3639), .Z(n4894) );
  NAND2_X1 U3126 ( .A1(n4108), .A2(n4894), .ZN(n2715) );
  NAND2_X1 U3127 ( .A1(n4109), .A2(n3509), .ZN(n3443) );
  AND3_X1 U3128 ( .A1(n3688), .A2(n2715), .A3(n3443), .ZN(n2718) );
  INV_X1 U3129 ( .A(n2715), .ZN(n2716) );
  INV_X1 U3130 ( .A(n3452), .ZN(n3528) );
  OR2_X1 U3131 ( .A1(n4886), .A2(n3528), .ZN(n3483) );
  OAI22_X1 U3132 ( .A1(n2716), .A2(n3483), .B1(n4894), .B2(n4108), .ZN(n2717)
         );
  NAND2_X1 U3133 ( .A1(n3641), .A2(REG2_REG_16__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3134 ( .A1(n3640), .A2(REG1_REG_16__SCAN_IN), .ZN(n2722) );
  AOI21_X1 U3135 ( .B1(n2719), .B2(n4624), .A(n2727), .ZN(n3477) );
  NAND2_X1 U3136 ( .A1(n2684), .A2(n3477), .ZN(n2721) );
  NAND2_X1 U3137 ( .A1(n3642), .A2(REG0_REG_16__SCAN_IN), .ZN(n2720) );
  NAND4_X1 U3138 ( .A1(n2723), .A2(n2722), .A3(n2721), .A4(n2720), .ZN(n4885)
         );
  INV_X1 U3139 ( .A(DATAI_16_), .ZN(n4904) );
  NAND2_X1 U3140 ( .A1(n2724), .A2(IR_REG_31__SCAN_IN), .ZN(n2725) );
  XNOR2_X1 U3141 ( .A(n2725), .B(IR_REG_16__SCAN_IN), .ZN(n4190) );
  MUX2_X1 U3142 ( .A(n4904), .B(n4905), .S(n3639), .Z(n3471) );
  OR2_X1 U3143 ( .A1(n4885), .A2(n3471), .ZN(n3708) );
  NAND2_X1 U3144 ( .A1(n4885), .A2(n3471), .ZN(n3704) );
  NAND2_X1 U3145 ( .A1(n3708), .A2(n3704), .ZN(n3475) );
  NAND2_X1 U3146 ( .A1(n3476), .A2(n3475), .ZN(n3474) );
  NAND2_X1 U3147 ( .A1(n4885), .A2(n4034), .ZN(n2726) );
  NAND2_X1 U31480 ( .A1(n3474), .A2(n2726), .ZN(n3535) );
  NAND2_X1 U31490 ( .A1(n3640), .A2(REG1_REG_17__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U3150 ( .A1(n3641), .A2(REG2_REG_17__SCAN_IN), .ZN(n2731) );
  OAI21_X1 U3151 ( .B1(REG3_REG_17__SCAN_IN), .B2(n2727), .A(n2740), .ZN(n3772) );
  INV_X1 U3152 ( .A(n3772), .ZN(n2728) );
  NAND2_X1 U3153 ( .A1(n2684), .A2(n2728), .ZN(n2730) );
  NAND2_X1 U3154 ( .A1(n3642), .A2(REG0_REG_17__SCAN_IN), .ZN(n2729) );
  NAND4_X1 U3155 ( .A1(n2732), .A2(n2731), .A3(n2730), .A4(n2729), .ZN(n4107)
         );
  INV_X1 U3156 ( .A(DATAI_17_), .ZN(n2737) );
  INV_X1 U3157 ( .A(n2733), .ZN(n2734) );
  AND2_X1 U3158 ( .A1(n2734), .A2(IR_REG_31__SCAN_IN), .ZN(n2759) );
  INV_X1 U3159 ( .A(n2745), .ZN(n2736) );
  XNOR2_X1 U3160 ( .A(n2736), .B(IR_REG_17__SCAN_IN), .ZN(n4204) );
  MUX2_X1 U3161 ( .A(n2737), .B(n4204), .S(n3639), .Z(n3540) );
  OR2_X1 U3162 ( .A1(n4107), .A2(n3769), .ZN(n2738) );
  NAND2_X1 U3163 ( .A1(n4107), .A2(n3769), .ZN(n2739) );
  NAND2_X1 U3164 ( .A1(n3640), .A2(REG1_REG_18__SCAN_IN), .ZN(n2744) );
  NAND2_X1 U3165 ( .A1(n3641), .A2(REG2_REG_18__SCAN_IN), .ZN(n2743) );
  AOI21_X1 U3166 ( .B1(n4076), .B2(n2740), .A(n2748), .ZN(n3784) );
  NAND2_X1 U3167 ( .A1(n2684), .A2(n3784), .ZN(n2742) );
  NAND2_X1 U3168 ( .A1(n3642), .A2(REG0_REG_18__SCAN_IN), .ZN(n2741) );
  NAND4_X1 U3169 ( .A1(n2744), .A2(n2743), .A3(n2742), .A4(n2741), .ZN(n4106)
         );
  INV_X1 U3170 ( .A(DATAI_18_), .ZN(n4462) );
  NAND2_X1 U3171 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U3172 ( .A1(n2745), .A2(n2757), .ZN(n2753) );
  XNOR2_X1 U3173 ( .A(n2753), .B(IR_REG_18__SCAN_IN), .ZN(n4221) );
  MUX2_X1 U3174 ( .A(n4462), .B(n4221), .S(n3639), .Z(n3872) );
  OR2_X1 U3175 ( .A1(n4106), .A2(n3872), .ZN(n3560) );
  NAND2_X1 U3176 ( .A1(n4106), .A2(n3872), .ZN(n3561) );
  NAND2_X1 U3177 ( .A1(n3560), .A2(n3561), .ZN(n3779) );
  INV_X1 U3178 ( .A(n3779), .ZN(n3788) );
  INV_X1 U3179 ( .A(n3872), .ZN(n4077) );
  OR2_X1 U3180 ( .A1(n4106), .A2(n4077), .ZN(n2746) );
  NAND2_X1 U3181 ( .A1(n3785), .A2(n2746), .ZN(n3556) );
  NAND2_X1 U3182 ( .A1(n3641), .A2(REG2_REG_19__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U3183 ( .A1(n3640), .A2(REG1_REG_19__SCAN_IN), .ZN(n2751) );
  INV_X1 U3184 ( .A(n2747), .ZN(n2768) );
  OAI21_X1 U3185 ( .B1(REG3_REG_19__SCAN_IN), .B2(n2748), .A(n2768), .ZN(n3568) );
  INV_X1 U3186 ( .A(n3568), .ZN(n3999) );
  NAND2_X1 U3187 ( .A1(n2684), .A2(n3999), .ZN(n2750) );
  NAND2_X1 U3188 ( .A1(n3642), .A2(REG0_REG_19__SCAN_IN), .ZN(n2749) );
  NAND4_X1 U3189 ( .A1(n2752), .A2(n2751), .A3(n2750), .A4(n2749), .ZN(n4105)
         );
  INV_X1 U3190 ( .A(n2753), .ZN(n2754) );
  NAND2_X1 U3191 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2756) );
  NAND2_X1 U3192 ( .A1(n2754), .A2(n2756), .ZN(n2755) );
  NAND2_X1 U3193 ( .A1(n2755), .A2(IR_REG_19__SCAN_IN), .ZN(n2764) );
  AND2_X1 U3194 ( .A1(n2503), .A2(n2756), .ZN(n2758) );
  NAND2_X1 U3195 ( .A1(n2758), .A2(n2757), .ZN(n2760) );
  MUX2_X1 U3196 ( .A(n4554), .B(n4828), .S(n3639), .Z(n3881) );
  NAND2_X1 U3197 ( .A1(n4105), .A2(n3998), .ZN(n2766) );
  NOR2_X1 U3198 ( .A1(n4105), .A2(n3998), .ZN(n2765) );
  NAND2_X1 U3199 ( .A1(n3640), .A2(REG1_REG_20__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U3200 ( .A1(n3641), .A2(REG2_REG_20__SCAN_IN), .ZN(n2772) );
  INV_X1 U3201 ( .A(n2767), .ZN(n2776) );
  INV_X1 U3202 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U3203 ( .A1(n2768), .A2(n4635), .ZN(n2769) );
  NAND2_X1 U3204 ( .A1(n2684), .A2(n3847), .ZN(n2771) );
  NAND2_X1 U3205 ( .A1(n3642), .A2(REG0_REG_20__SCAN_IN), .ZN(n2770) );
  NAND4_X1 U3206 ( .A1(n2773), .A2(n2772), .A3(n2771), .A4(n2770), .ZN(n4104)
         );
  INV_X1 U3207 ( .A(n4104), .ZN(n3995) );
  NAND2_X1 U3208 ( .A1(n3646), .A2(DATAI_20_), .ZN(n3892) );
  NAND2_X1 U3209 ( .A1(n3640), .A2(REG1_REG_21__SCAN_IN), .ZN(n2781) );
  NAND2_X1 U32100 ( .A1(n3641), .A2(REG2_REG_21__SCAN_IN), .ZN(n2780) );
  INV_X1 U32110 ( .A(n2774), .ZN(n2783) );
  INV_X1 U32120 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U32130 ( .A1(n2776), .A2(n2775), .ZN(n2777) );
  NAND2_X1 U32140 ( .A1(n2684), .A2(n3805), .ZN(n2779) );
  NAND2_X1 U32150 ( .A1(n3642), .A2(REG0_REG_21__SCAN_IN), .ZN(n2778) );
  NAND4_X1 U32160 ( .A1(n2781), .A2(n2780), .A3(n2779), .A4(n2778), .ZN(n4103)
         );
  NAND2_X1 U32170 ( .A1(n3646), .A2(DATAI_21_), .ZN(n3808) );
  INV_X1 U32180 ( .A(n3808), .ZN(n4010) );
  NAND2_X1 U32190 ( .A1(n4103), .A2(n4010), .ZN(n3813) );
  NAND2_X1 U32200 ( .A1(n3641), .A2(REG2_REG_22__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U32210 ( .A1(n3640), .A2(REG1_REG_22__SCAN_IN), .ZN(n2787) );
  INV_X1 U32220 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U32230 ( .A1(n2783), .A2(n2782), .ZN(n2784) );
  AND2_X1 U32240 ( .A1(n2790), .A2(n2784), .ZN(n3826) );
  NAND2_X1 U32250 ( .A1(n2684), .A2(n3826), .ZN(n2786) );
  NAND2_X1 U32260 ( .A1(n3642), .A2(REG0_REG_22__SCAN_IN), .ZN(n2785) );
  NAND4_X1 U32270 ( .A1(n2788), .A2(n2787), .A3(n2786), .A4(n2785), .ZN(n4102)
         );
  NAND2_X1 U32280 ( .A1(n3646), .A2(DATAI_22_), .ZN(n4064) );
  NAND2_X1 U32290 ( .A1(n4102), .A2(n4064), .ZN(n2861) );
  NAND2_X1 U32300 ( .A1(n4334), .A2(n2861), .ZN(n4335) );
  INV_X1 U32310 ( .A(n4335), .ZN(n2789) );
  NOR2_X1 U32320 ( .A1(n4103), .A2(n4010), .ZN(n3814) );
  INV_X1 U32330 ( .A(n4102), .ZN(n4340) );
  NOR2_X1 U32340 ( .A1(n4340), .A2(n4064), .ZN(n4331) );
  NAND2_X1 U32350 ( .A1(n3646), .A2(DATAI_23_), .ZN(n4347) );
  INV_X1 U32360 ( .A(n4347), .ZN(n3973) );
  NAND2_X1 U32370 ( .A1(n3641), .A2(REG2_REG_23__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U32380 ( .A1(n3640), .A2(REG1_REG_23__SCAN_IN), .ZN(n2795) );
  NAND2_X1 U32390 ( .A1(n2790), .A2(n4608), .ZN(n2791) );
  NAND2_X1 U32400 ( .A1(n2684), .A2(n4349), .ZN(n2794) );
  NAND2_X1 U32410 ( .A1(n3642), .A2(REG0_REG_23__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U32420 ( .A1(n2798), .A2(n2797), .ZN(n4309) );
  AOI21_X1 U32430 ( .B1(n4315), .B2(n4342), .A(n4309), .ZN(n2799) );
  AOI21_X1 U32440 ( .B1(n4300), .B2(n4324), .A(n2799), .ZN(n4290) );
  OAI21_X1 U32450 ( .B1(n4255), .B2(n4278), .A(n4262), .ZN(n2800) );
  NAND2_X1 U32460 ( .A1(n3641), .A2(REG2_REG_28__SCAN_IN), .ZN(n2808) );
  NAND2_X1 U32470 ( .A1(n3640), .A2(REG1_REG_28__SCAN_IN), .ZN(n2807) );
  INV_X1 U32480 ( .A(n2803), .ZN(n2801) );
  NAND2_X1 U32490 ( .A1(n2801), .A2(REG3_REG_28__SCAN_IN), .ZN(n4228) );
  INV_X1 U32500 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U32510 ( .A1(n2803), .A2(n2802), .ZN(n2804) );
  NAND2_X1 U32520 ( .A1(n2684), .A2(n4235), .ZN(n2806) );
  NAND2_X1 U32530 ( .A1(n3642), .A2(REG0_REG_28__SCAN_IN), .ZN(n2805) );
  NAND4_X1 U32540 ( .A1(n2808), .A2(n2807), .A3(n2806), .A4(n2805), .ZN(n4256)
         );
  NAND2_X1 U32550 ( .A1(n3646), .A2(DATAI_28_), .ZN(n4238) );
  OR2_X1 U32560 ( .A1(n4256), .A2(n4238), .ZN(n2866) );
  NAND2_X1 U32570 ( .A1(n4256), .A2(n4238), .ZN(n3636) );
  NAND2_X1 U32580 ( .A1(n2866), .A2(n3636), .ZN(n4241) );
  INV_X1 U32590 ( .A(n4238), .ZN(n4243) );
  NAND2_X1 U32600 ( .A1(n3641), .A2(REG2_REG_29__SCAN_IN), .ZN(n2813) );
  NAND2_X1 U32610 ( .A1(n3640), .A2(REG1_REG_29__SCAN_IN), .ZN(n2812) );
  INV_X1 U32620 ( .A(n4228), .ZN(n2809) );
  NAND2_X1 U32630 ( .A1(n2684), .A2(n2809), .ZN(n2811) );
  NAND2_X1 U32640 ( .A1(n3642), .A2(REG0_REG_29__SCAN_IN), .ZN(n2810) );
  NAND4_X1 U32650 ( .A1(n2813), .A2(n2812), .A3(n2811), .A4(n2810), .ZN(n4244)
         );
  NAND2_X1 U32660 ( .A1(n3646), .A2(DATAI_29_), .ZN(n3658) );
  XNOR2_X1 U32670 ( .A(n4244), .B(n3658), .ZN(n3695) );
  NAND2_X1 U32680 ( .A1(n2877), .A2(n2818), .ZN(n2819) );
  NAND2_X1 U32690 ( .A1(n2819), .A2(IR_REG_31__SCAN_IN), .ZN(n2820) );
  AND2_X1 U32700 ( .A1(n2818), .A2(n2821), .ZN(n2822) );
  NAND2_X1 U32710 ( .A1(n2877), .A2(n2822), .ZN(n2823) );
  NAND2_X1 U32720 ( .A1(n2823), .A2(IR_REG_31__SCAN_IN), .ZN(n2824) );
  XNOR2_X1 U32730 ( .A(n2979), .B(n4448), .ZN(n2825) );
  NAND2_X1 U32740 ( .A1(n2825), .A2(n4828), .ZN(n3842) );
  AND2_X1 U32750 ( .A1(n2912), .A2(n4450), .ZN(n4765) );
  INV_X1 U32760 ( .A(n4448), .ZN(n2872) );
  INV_X1 U32770 ( .A(n4794), .ZN(n4774) );
  NAND2_X1 U32780 ( .A1(n3842), .A2(n4774), .ZN(n4840) );
  NAND2_X1 U32790 ( .A1(n3640), .A2(REG1_REG_30__SCAN_IN), .ZN(n2828) );
  NAND2_X1 U32800 ( .A1(n3641), .A2(REG2_REG_30__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U32810 ( .A1(n3642), .A2(REG0_REG_30__SCAN_IN), .ZN(n2826) );
  AND3_X1 U32820 ( .A1(n2828), .A2(n2827), .A3(n2826), .ZN(n3655) );
  AND2_X1 U32830 ( .A1(n2829), .A2(n2830), .ZN(n2831) );
  OR2_X1 U32840 ( .A1(n2831), .A2(n2930), .ZN(n2833) );
  XNOR2_X1 U32850 ( .A(n2833), .B(n2832), .ZN(n4907) );
  AND2_X1 U32860 ( .A1(n4448), .A2(n3726), .ZN(n3006) );
  NAND2_X1 U32870 ( .A1(n4907), .A2(n3006), .ZN(n3778) );
  XNOR2_X1 U32880 ( .A(n2834), .B(IR_REG_27__SCAN_IN), .ZN(n2951) );
  NAND2_X1 U32890 ( .A1(n2951), .A2(B_REG_SCAN_IN), .ZN(n2835) );
  NAND2_X1 U32900 ( .A1(n2263), .A2(n2835), .ZN(n4223) );
  INV_X1 U32910 ( .A(n3684), .ZN(n3094) );
  OR2_X1 U32920 ( .A1(n4120), .A2(n3124), .ZN(n3125) );
  INV_X1 U32930 ( .A(n3125), .ZN(n3602) );
  NAND2_X1 U32940 ( .A1(n3094), .A2(n3602), .ZN(n3093) );
  NAND2_X1 U32950 ( .A1(n3093), .A2(n3603), .ZN(n3166) );
  INV_X1 U32960 ( .A(n3685), .ZN(n2836) );
  NAND2_X1 U32970 ( .A1(n3166), .A2(n2836), .ZN(n2837) );
  NAND2_X1 U32980 ( .A1(n2837), .A2(n3604), .ZN(n3196) );
  OR2_X1 U32990 ( .A1(n3050), .A2(n3205), .ZN(n3609) );
  NAND2_X1 U33000 ( .A1(n3050), .A2(n3205), .ZN(n3606) );
  NAND2_X1 U33010 ( .A1(n3609), .A2(n3606), .ZN(n3683) );
  INV_X1 U33020 ( .A(n3683), .ZN(n3197) );
  NAND2_X1 U33030 ( .A1(n3196), .A2(n3197), .ZN(n3195) );
  INV_X1 U33040 ( .A(n3610), .ZN(n2838) );
  INV_X1 U33050 ( .A(n3153), .ZN(n2839) );
  AND2_X1 U33060 ( .A1(n4115), .A2(n2839), .ZN(n3145) );
  OR2_X1 U33070 ( .A1(n4115), .A2(n2839), .ZN(n3585) );
  NAND2_X1 U33080 ( .A1(n2840), .A2(n3585), .ZN(n3175) );
  NAND2_X1 U33090 ( .A1(n4816), .A2(n3182), .ZN(n3613) );
  NAND2_X1 U33100 ( .A1(n3175), .A2(n3613), .ZN(n4812) );
  OR2_X1 U33110 ( .A1(n4816), .A2(n3182), .ZN(n4811) );
  OR2_X1 U33120 ( .A1(n4114), .A2(n2292), .ZN(n2841) );
  AND2_X1 U33130 ( .A1(n4811), .A2(n2841), .ZN(n3617) );
  NAND2_X1 U33140 ( .A1(n4812), .A2(n3617), .ZN(n2842) );
  NAND2_X1 U33150 ( .A1(n4114), .A2(n2292), .ZN(n3582) );
  NAND2_X1 U33160 ( .A1(n2842), .A2(n3582), .ZN(n3295) );
  INV_X1 U33170 ( .A(n3302), .ZN(n2843) );
  OR2_X1 U33180 ( .A1(n4814), .A2(n2843), .ZN(n3620) );
  NAND2_X1 U33190 ( .A1(n3295), .A2(n3620), .ZN(n2844) );
  NAND2_X1 U33200 ( .A1(n4814), .A2(n2843), .ZN(n3583) );
  NAND2_X1 U33210 ( .A1(n2844), .A2(n3583), .ZN(n3222) );
  INV_X1 U33220 ( .A(n3319), .ZN(n2911) );
  AND2_X1 U33230 ( .A1(n4113), .A2(n2911), .ZN(n3619) );
  OR2_X1 U33240 ( .A1(n4113), .A2(n2911), .ZN(n3621) );
  NAND2_X1 U33250 ( .A1(n4112), .A2(n3339), .ZN(n3588) );
  OR2_X1 U33260 ( .A1(n4112), .A2(n3339), .ZN(n3592) );
  INV_X1 U33270 ( .A(n3436), .ZN(n3432) );
  NAND2_X1 U33280 ( .A1(n4110), .A2(n3432), .ZN(n3379) );
  NAND2_X1 U33290 ( .A1(n4109), .A2(n3389), .ZN(n2845) );
  NAND2_X1 U33300 ( .A1(n3379), .A2(n2845), .ZN(n2847) );
  INV_X1 U33310 ( .A(n3329), .ZN(n2846) );
  NOR2_X1 U33320 ( .A1(n2847), .A2(n2846), .ZN(n3589) );
  NAND2_X1 U33330 ( .A1(n3405), .A2(n3589), .ZN(n2851) );
  INV_X1 U33340 ( .A(n2847), .ZN(n2850) );
  OR2_X1 U33350 ( .A1(n4110), .A2(n3432), .ZN(n3381) );
  NAND2_X1 U33360 ( .A1(n3327), .A2(n3381), .ZN(n2849) );
  NOR2_X1 U33370 ( .A1(n4109), .A2(n3389), .ZN(n2848) );
  AOI21_X1 U33380 ( .B1(n2850), .B2(n2849), .A(n2848), .ZN(n3594) );
  NAND2_X1 U33390 ( .A1(n2851), .A2(n3594), .ZN(n3706) );
  INV_X1 U33400 ( .A(n3688), .ZN(n3446) );
  NAND2_X1 U33410 ( .A1(n3706), .A2(n3446), .ZN(n3486) );
  INV_X1 U33420 ( .A(n4894), .ZN(n3493) );
  OR2_X1 U33430 ( .A1(n4108), .A2(n3493), .ZN(n3599) );
  NAND2_X1 U33440 ( .A1(n4108), .A2(n3493), .ZN(n3598) );
  NAND2_X1 U33450 ( .A1(n3599), .A2(n3598), .ZN(n3687) );
  INV_X1 U33460 ( .A(n3593), .ZN(n2852) );
  NOR2_X1 U33470 ( .A1(n3687), .A2(n2852), .ZN(n2853) );
  NAND2_X1 U33480 ( .A1(n3486), .A2(n2853), .ZN(n2854) );
  NAND2_X1 U33490 ( .A1(n2854), .A2(n3598), .ZN(n3468) );
  INV_X1 U33500 ( .A(n3475), .ZN(n3693) );
  NAND2_X1 U33510 ( .A1(n3468), .A2(n3693), .ZN(n2855) );
  NAND2_X1 U33520 ( .A1(n4105), .A2(n3881), .ZN(n3554) );
  AND2_X1 U3353 ( .A1(n3561), .A2(n3554), .ZN(n2858) );
  NAND2_X1 U33540 ( .A1(n4107), .A2(n3540), .ZN(n3557) );
  AND2_X1 U3355 ( .A1(n2858), .A2(n3557), .ZN(n3833) );
  NAND2_X1 U3356 ( .A1(n4104), .A2(n3892), .ZN(n3669) );
  AND2_X1 U3357 ( .A1(n3833), .A2(n3669), .ZN(n3630) );
  INV_X1 U3358 ( .A(n3630), .ZN(n3707) );
  OR2_X1 U3359 ( .A1(n4107), .A2(n3540), .ZN(n3558) );
  NAND2_X1 U3360 ( .A1(n3560), .A2(n3558), .ZN(n2857) );
  OR2_X1 U3361 ( .A1(n4105), .A2(n3881), .ZN(n3555) );
  INV_X1 U3362 ( .A(n3555), .ZN(n2856) );
  AOI21_X1 U3363 ( .B1(n2858), .B2(n2857), .A(n2856), .ZN(n3834) );
  OR2_X1 U3364 ( .A1(n4104), .A2(n3892), .ZN(n3670) );
  NAND2_X1 U3365 ( .A1(n3834), .A2(n3670), .ZN(n2859) );
  NAND2_X1 U3366 ( .A1(n2859), .A2(n3669), .ZN(n3710) );
  OR2_X1 U3367 ( .A1(n4103), .A2(n3808), .ZN(n3692) );
  AND2_X1 U3368 ( .A1(n4334), .A2(n3692), .ZN(n3715) );
  INV_X1 U3369 ( .A(n3715), .ZN(n2860) );
  NAND2_X1 U3370 ( .A1(n4101), .A2(n4347), .ZN(n3662) );
  AND2_X1 U3371 ( .A1(n2861), .A2(n3662), .ZN(n3635) );
  AND2_X1 U3372 ( .A1(n4103), .A2(n3808), .ZN(n3818) );
  NAND2_X1 U3373 ( .A1(n3818), .A2(n4334), .ZN(n2862) );
  NAND2_X1 U3374 ( .A1(n3635), .A2(n2862), .ZN(n3713) );
  INV_X1 U3375 ( .A(n3713), .ZN(n2863) );
  OR2_X1 U3376 ( .A1(n4101), .A2(n4347), .ZN(n4310) );
  OR2_X1 U3377 ( .A1(n4342), .A2(n4324), .ZN(n2864) );
  NAND2_X1 U3378 ( .A1(n4310), .A2(n2864), .ZN(n3717) );
  INV_X1 U3379 ( .A(n3717), .ZN(n2865) );
  NAND2_X1 U3380 ( .A1(n4311), .A2(n2865), .ZN(n4292) );
  NAND2_X1 U3381 ( .A1(n4316), .A2(n4301), .ZN(n3671) );
  NAND2_X1 U3382 ( .A1(n4342), .A2(n4324), .ZN(n4291) );
  AND2_X1 U3383 ( .A1(n3671), .A2(n4291), .ZN(n3716) );
  OR2_X1 U3384 ( .A1(n4316), .A2(n4301), .ZN(n4273) );
  OR2_X1 U3385 ( .A1(n4297), .A2(n4283), .ZN(n3691) );
  INV_X1 U3386 ( .A(n3652), .ZN(n3701) );
  NAND2_X1 U3387 ( .A1(n4297), .A2(n4283), .ZN(n3698) );
  NAND2_X1 U3388 ( .A1(n4278), .A2(n4265), .ZN(n3649) );
  INV_X1 U3389 ( .A(n4261), .ZN(n4253) );
  NAND2_X1 U3390 ( .A1(n4239), .A2(n2866), .ZN(n3702) );
  XNOR2_X1 U3391 ( .A(n2867), .B(n3695), .ZN(n2870) );
  INV_X1 U3392 ( .A(n2912), .ZN(n4449) );
  NAND2_X1 U3393 ( .A1(n4449), .A2(n3726), .ZN(n2869) );
  NAND2_X1 U3394 ( .A1(n4450), .A2(n4448), .ZN(n2868) );
  NAND2_X1 U3395 ( .A1(n2869), .A2(n2868), .ZN(n4821) );
  NAND2_X1 U3396 ( .A1(n2870), .A2(n4821), .ZN(n2875) );
  INV_X1 U3397 ( .A(n3006), .ZN(n2871) );
  NAND2_X1 U3398 ( .A1(n4449), .A2(n3127), .ZN(n4819) );
  NOR2_X1 U3399 ( .A1(n3658), .A2(n4819), .ZN(n2873) );
  AOI21_X1 U3400 ( .B1(n4256), .B2(n2260), .A(n2873), .ZN(n2874) );
  OAI211_X1 U3401 ( .C1(n3655), .C2(n4223), .A(n2875), .B(n2874), .ZN(n4231)
         );
  NAND2_X1 U3402 ( .A1(n2894), .A2(n2895), .ZN(n2879) );
  INV_X1 U3403 ( .A(IR_REG_24__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U3404 ( .A1(n2891), .A2(n2890), .ZN(n2884) );
  MUX2_X1 U3405 ( .A(n2891), .B(n2884), .S(B_REG_SCAN_IN), .Z(n2888) );
  INV_X1 U3406 ( .A(IR_REG_25__SCAN_IN), .ZN(n2885) );
  NAND2_X1 U3407 ( .A1(n2886), .A2(IR_REG_31__SCAN_IN), .ZN(n2887) );
  XNOR2_X1 U3408 ( .A(n2887), .B(IR_REG_26__SCAN_IN), .ZN(n2892) );
  INV_X1 U3409 ( .A(D_REG_1__SCAN_IN), .ZN(n2889) );
  NAND2_X1 U3410 ( .A1(n2936), .A2(n2889), .ZN(n3100) );
  INV_X1 U3411 ( .A(n2892), .ZN(n2909) );
  NAND2_X1 U3412 ( .A1(n2909), .A2(n2890), .ZN(n3003) );
  NAND2_X1 U3413 ( .A1(n3100), .A2(n3003), .ZN(n2908) );
  INV_X1 U3414 ( .A(n2890), .ZN(n2923) );
  INV_X1 U3415 ( .A(n2891), .ZN(n2893) );
  XNOR2_X1 U3416 ( .A(n2894), .B(n2895), .ZN(n3059) );
  AND2_X1 U3417 ( .A1(n3059), .A2(STATE_REG_SCAN_IN), .ZN(n2939) );
  NAND2_X1 U3418 ( .A1(n2912), .A2(n4828), .ZN(n2896) );
  NAND2_X1 U3419 ( .A1(n2896), .A2(n3006), .ZN(n3058) );
  AND2_X1 U3420 ( .A1(n3013), .A2(n3058), .ZN(n3102) );
  NOR4_X1 U3421 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2900) );
  NOR4_X1 U3422 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2899) );
  NOR4_X1 U3423 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2898) );
  NOR4_X1 U3424 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2897) );
  NAND4_X1 U3425 ( .A1(n2900), .A2(n2899), .A3(n2898), .A4(n2897), .ZN(n2906)
         );
  NOR2_X1 U3426 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_31__SCAN_IN), .ZN(n2904) );
  NOR4_X1 U3427 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2903) );
  NOR4_X1 U3428 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2902) );
  NOR4_X1 U3429 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2901) );
  NAND4_X1 U3430 ( .A1(n2904), .A2(n2903), .A3(n2902), .A4(n2901), .ZN(n2905)
         );
  OAI21_X1 U3431 ( .B1(n2906), .B2(n2905), .A(n2936), .ZN(n3004) );
  NAND2_X1 U3432 ( .A1(n4794), .A2(n3012), .ZN(n2907) );
  NAND4_X1 U3433 ( .A1(n2908), .A2(n3102), .A3(n3004), .A4(n2907), .ZN(n2915)
         );
  INV_X1 U3434 ( .A(D_REG_0__SCAN_IN), .ZN(n2941) );
  NAND2_X1 U3435 ( .A1(n2936), .A2(n2941), .ZN(n2910) );
  NAND2_X1 U3436 ( .A1(n2909), .A2(n2891), .ZN(n2938) );
  NAND2_X1 U3437 ( .A1(n2910), .A2(n2938), .ZN(n3101) );
  INV_X1 U3438 ( .A(n3101), .ZN(n3005) );
  INV_X2 U3439 ( .A(n4414), .ZN(n4849) );
  NAND2_X1 U3440 ( .A1(n3124), .A2(n2997), .ZN(n3171) );
  NAND2_X1 U3441 ( .A1(n3206), .A2(n3205), .ZN(n3208) );
  OAI21_X1 U3442 ( .B1(n4236), .B2(n3658), .A(n2268), .ZN(n4229) );
  NAND2_X1 U3443 ( .A1(n4849), .A2(n4406), .ZN(n4442) );
  NAND2_X1 U3444 ( .A1(n2914), .A2(n2913), .ZN(U3515) );
  INV_X1 U3445 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2917) );
  MUX2_X1 U3446 ( .A(n2917), .B(n2916), .S(n4411), .Z(n2919) );
  NAND2_X1 U3447 ( .A1(n4411), .A2(n4406), .ZN(n4396) );
  NAND2_X1 U3448 ( .A1(n2919), .A2(n2918), .ZN(U3547) );
  INV_X1 U3449 ( .A(n2939), .ZN(n3732) );
  OR2_X1 U3450 ( .A1(n2980), .A2(n3732), .ZN(n4117) );
  INV_X1 U3451 ( .A(n4117), .ZN(U4043) );
  INV_X1 U3452 ( .A(DATAI_21_), .ZN(n2921) );
  NAND2_X1 U3453 ( .A1(n3726), .A2(STATE_REG_SCAN_IN), .ZN(n2920) );
  OAI21_X1 U3454 ( .B1(STATE_REG_SCAN_IN), .B2(n2921), .A(n2920), .ZN(U3331)
         );
  INV_X1 U3455 ( .A(DATAI_15_), .ZN(n4482) );
  NAND2_X1 U3456 ( .A1(n4186), .A2(STATE_REG_SCAN_IN), .ZN(n2922) );
  OAI21_X1 U3457 ( .B1(STATE_REG_SCAN_IN), .B2(n4482), .A(n2922), .ZN(U3337)
         );
  INV_X1 U34580 ( .A(DATAI_25_), .ZN(n4557) );
  NAND2_X1 U34590 ( .A1(n2923), .A2(STATE_REG_SCAN_IN), .ZN(n2924) );
  OAI21_X1 U3460 ( .B1(STATE_REG_SCAN_IN), .B2(n4557), .A(n2924), .ZN(U3327)
         );
  INV_X1 U3461 ( .A(DATAI_29_), .ZN(n2927) );
  NAND2_X1 U3462 ( .A1(n2925), .A2(STATE_REG_SCAN_IN), .ZN(n2926) );
  OAI21_X1 U3463 ( .B1(STATE_REG_SCAN_IN), .B2(n2927), .A(n2926), .ZN(U3323)
         );
  INV_X1 U3464 ( .A(DATAI_24_), .ZN(n4565) );
  MUX2_X1 U3465 ( .A(n4565), .B(n2891), .S(STATE_REG_SCAN_IN), .Z(n2928) );
  INV_X1 U3466 ( .A(n2928), .ZN(U3328) );
  INV_X1 U34670 ( .A(n4204), .ZN(n4211) );
  NAND2_X1 U3468 ( .A1(n4211), .A2(STATE_REG_SCAN_IN), .ZN(n2929) );
  OAI21_X1 U34690 ( .B1(STATE_REG_SCAN_IN), .B2(n2737), .A(n2929), .ZN(U3335)
         );
  INV_X1 U3470 ( .A(DATAI_31_), .ZN(n2933) );
  OR4_X1 U34710 ( .A1(n2931), .A2(IR_REG_30__SCAN_IN), .A3(n2930), .A4(U3149), 
        .ZN(n2932) );
  OAI21_X1 U3472 ( .B1(STATE_REG_SCAN_IN), .B2(n2933), .A(n2932), .ZN(U3321)
         );
  MUX2_X1 U34730 ( .A(n4125), .B(n2550), .S(U3149), .Z(n2934) );
  INV_X1 U3474 ( .A(n2934), .ZN(U3351) );
  INV_X1 U34750 ( .A(DATAI_27_), .ZN(n4559) );
  NAND2_X1 U3476 ( .A1(n2951), .A2(STATE_REG_SCAN_IN), .ZN(n2935) );
  OAI21_X1 U34770 ( .B1(STATE_REG_SCAN_IN), .B2(n4559), .A(n2935), .ZN(U3325)
         );
  INV_X1 U3478 ( .A(n2936), .ZN(n2937) );
  INV_X1 U3480 ( .A(n2938), .ZN(n2940) );
  AOI22_X1 U34810 ( .A1(n2262), .A2(n2941), .B1(n2940), .B2(n2939), .ZN(U3458)
         );
  NAND2_X1 U34830 ( .A1(n4914), .A2(n3003), .ZN(n2942) );
  OAI21_X1 U3484 ( .B1(n4914), .B2(n2889), .A(n2942), .ZN(U3459) );
  AND2_X1 U34850 ( .A1(n3059), .A2(n3006), .ZN(n2944) );
  NOR2_X1 U3486 ( .A1(n3639), .A2(n2944), .ZN(n2950) );
  INV_X1 U34870 ( .A(n2950), .ZN(n2946) );
  OR2_X1 U3488 ( .A1(n3059), .A2(U3149), .ZN(n4455) );
  INV_X1 U34890 ( .A(n4455), .ZN(n2945) );
  OR2_X1 U3490 ( .A1(n3013), .A2(n2945), .ZN(n2949) );
  NOR2_X1 U34910 ( .A1(n4757), .A2(U4043), .ZN(U3148) );
  INV_X1 U3492 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4771) );
  AND2_X1 U34930 ( .A1(n2951), .A2(n4771), .ZN(n2947) );
  NOR2_X1 U3494 ( .A1(n4907), .A2(n2947), .ZN(n2988) );
  OAI21_X1 U34950 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2951), .A(n2988), .ZN(n2948) );
  MUX2_X1 U3496 ( .A(n2988), .B(n2948), .S(n2295), .Z(n2955) );
  AND2_X1 U34970 ( .A1(n2950), .A2(n2949), .ZN(n2963) );
  INV_X1 U3498 ( .A(n2963), .ZN(n2954) );
  AOI22_X1 U34990 ( .A1(n4757), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2953) );
  INV_X1 U3500 ( .A(n2951), .ZN(n3734) );
  AND2_X1 U35010 ( .A1(n2963), .A2(n3734), .ZN(n4744) );
  INV_X1 U3502 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2981) );
  NAND3_X1 U35030 ( .A1(n4744), .A2(IR_REG_0__SCAN_IN), .A3(n2981), .ZN(n2952)
         );
  OAI211_X1 U3504 ( .C1(n2955), .C2(n2954), .A(n2953), .B(n2952), .ZN(U3240)
         );
  NAND2_X1 U35050 ( .A1(n2963), .A2(n4907), .ZN(n4759) );
  INV_X1 U35060 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2956) );
  INV_X1 U35070 ( .A(n4137), .ZN(n2959) );
  NAND2_X1 U35080 ( .A1(n4121), .A2(REG1_REG_1__SCAN_IN), .ZN(n2958) );
  INV_X1 U35090 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4778) );
  NAND2_X1 U35100 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(
        n4126) );
  AOI21_X1 U35110 ( .B1(n4125), .B2(n4778), .A(n4126), .ZN(n2957) );
  NAND2_X1 U35120 ( .A1(n2958), .A2(n2957), .ZN(n4129) );
  NAND2_X1 U35130 ( .A1(n4129), .A2(n2958), .ZN(n4138) );
  INV_X1 U35140 ( .A(n4142), .ZN(n4454) );
  XOR2_X1 U35150 ( .A(REG1_REG_3__SCAN_IN), .B(n2976), .Z(n2967) );
  INV_X1 U35160 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2965) );
  NAND2_X1 U35170 ( .A1(n4124), .A2(n4123), .ZN(n4122) );
  NAND2_X1 U35180 ( .A1(n4121), .A2(REG2_REG_1__SCAN_IN), .ZN(n2960) );
  NAND2_X1 U35190 ( .A1(n4122), .A2(n2960), .ZN(n4135) );
  MUX2_X1 U35200 ( .A(n2961), .B(REG2_REG_2__SCAN_IN), .S(n4142), .Z(n4136) );
  NAND2_X1 U35210 ( .A1(n4135), .A2(n4136), .ZN(n4134) );
  XNOR2_X1 U35220 ( .A(n2970), .B(n4453), .ZN(n2964) );
  NOR2_X1 U35230 ( .A1(n4907), .A2(n3734), .ZN(n2962) );
  AND2_X1 U35240 ( .A1(n2963), .A2(n2962), .ZN(n4761) );
  INV_X1 U35250 ( .A(n4761), .ZN(n4739) );
  AOI211_X1 U35260 ( .C1(n2965), .C2(n2964), .A(n2972), .B(n4739), .ZN(n2966)
         );
  AOI21_X1 U35270 ( .B1(n4744), .B2(n2967), .A(n2966), .ZN(n2969) );
  NOR2_X1 U35280 ( .A1(STATE_REG_SCAN_IN), .A2(n2569), .ZN(n3064) );
  AOI21_X1 U35290 ( .B1(n4757), .B2(ADDR_REG_3__SCAN_IN), .A(n3064), .ZN(n2968) );
  OAI211_X1 U35300 ( .C1(n2338), .C2(n4759), .A(n2969), .B(n2968), .ZN(U3243)
         );
  AND2_X1 U35310 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3859) );
  OAI21_X1 U35320 ( .B1(REG2_REG_4__SCAN_IN), .B2(n2974), .A(n4761), .ZN(n2990) );
  XNOR2_X1 U35330 ( .A(REG1_REG_4__SCAN_IN), .B(n3232), .ZN(n2977) );
  NAND2_X1 U35340 ( .A1(n4744), .A2(n2977), .ZN(n2989) );
  INV_X1 U35350 ( .A(n2979), .ZN(n2978) );
  AND2_X2 U35360 ( .A1(n2978), .A2(n2980), .ZN(n3891) );
  NAND2_X1 U35370 ( .A1(n2993), .A2(n2983), .ZN(n2995) );
  NAND2_X1 U35380 ( .A1(n4120), .A2(n3431), .ZN(n2985) );
  AOI22_X1 U35390 ( .A1(n3126), .A2(n3891), .B1(n2982), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2984) );
  NAND2_X1 U35400 ( .A1(n2985), .A2(n2984), .ZN(n2994) );
  XOR2_X1 U35410 ( .A(n2995), .B(n2994), .Z(n3042) );
  NAND2_X1 U35420 ( .A1(n3042), .A2(n3734), .ZN(n2986) );
  INV_X1 U35430 ( .A(n4907), .ZN(n3011) );
  OAI211_X1 U35440 ( .C1(n4123), .C2(n3734), .A(n2986), .B(n3011), .ZN(n2987)
         );
  OAI211_X1 U35450 ( .C1(IR_REG_0__SCAN_IN), .C2(n2988), .A(n2987), .B(U4043), 
        .ZN(n4146) );
  OAI211_X1 U35460 ( .C1(n3245), .C2(n2990), .A(n2989), .B(n4146), .ZN(n2991)
         );
  AOI211_X1 U35470 ( .C1(n4757), .C2(ADDR_REG_4__SCAN_IN), .A(n3859), .B(n2991), .ZN(n2992) );
  OAI21_X1 U35480 ( .B1(n3243), .B2(n4759), .A(n2992), .ZN(U3244) );
  NAND2_X1 U35490 ( .A1(n4828), .A2(n4448), .ZN(n3733) );
  NAND2_X1 U35500 ( .A1(n2979), .A2(n3733), .ZN(n3054) );
  AOI22_X1 U35510 ( .A1(n2995), .A2(n2994), .B1(n2993), .B2(n3031), .ZN(n3027)
         );
  NAND2_X1 U35520 ( .A1(n2996), .A2(n3891), .ZN(n3000) );
  INV_X1 U35530 ( .A(n2997), .ZN(n2998) );
  NAND2_X1 U35540 ( .A1(n2998), .A2(n3051), .ZN(n2999) );
  NAND2_X1 U35550 ( .A1(n3000), .A2(n2999), .ZN(n3001) );
  XNOR2_X1 U35560 ( .A(n3001), .B(n3054), .ZN(n3024) );
  NAND2_X1 U35570 ( .A1(n2996), .A2(n3431), .ZN(n3002) );
  NAND2_X1 U35580 ( .A1(n3002), .A2(n2274), .ZN(n3023) );
  XNOR2_X1 U35590 ( .A(n3024), .B(n3023), .ZN(n3028) );
  XNOR2_X1 U35600 ( .A(n3027), .B(n3028), .ZN(n3022) );
  AND2_X1 U35610 ( .A1(n3004), .A2(n3003), .ZN(n3103) );
  NAND3_X1 U35620 ( .A1(n3005), .A2(n3103), .A3(n3100), .ZN(n3019) );
  INV_X1 U35630 ( .A(n3019), .ZN(n3009) );
  AOI21_X1 U35640 ( .B1(n4450), .B2(n3127), .A(n3006), .ZN(n3007) );
  AND2_X1 U35650 ( .A1(n4819), .A2(n3007), .ZN(n3018) );
  AND2_X1 U35660 ( .A1(n3018), .A2(n3013), .ZN(n3008) );
  NAND2_X1 U35670 ( .A1(n3009), .A2(n3008), .ZN(n4097) );
  NOR2_X1 U35680 ( .A1(n2979), .A2(n3733), .ZN(n3010) );
  NAND2_X1 U35690 ( .A1(n3010), .A2(n3013), .ZN(n3016) );
  NOR2_X1 U35700 ( .A1(n3019), .A2(n3016), .ZN(n3015) );
  AND2_X2 U35710 ( .A1(n3015), .A2(n3011), .ZN(n4090) );
  NAND2_X1 U35720 ( .A1(n3013), .A2(n4359), .ZN(n3014) );
  NAND3_X1 U35730 ( .A1(n4794), .A2(n3013), .A3(n3012), .ZN(n4875) );
  OAI21_X1 U35740 ( .B1(n3019), .B2(n3014), .A(n4875), .ZN(n4092) );
  AOI22_X1 U35750 ( .A1(n4090), .A2(n4120), .B1(n2998), .B2(n4893), .ZN(n3021)
         );
  AND2_X2 U35760 ( .A1(n3015), .A2(n4907), .ZN(n4089) );
  OAI21_X1 U35770 ( .B1(n4819), .B2(U3149), .A(n3016), .ZN(n3017) );
  NAND2_X1 U35780 ( .A1(n3019), .A2(n3017), .ZN(n3062) );
  NAND2_X1 U35790 ( .A1(n3019), .A2(n3018), .ZN(n3060) );
  NAND3_X1 U35800 ( .A1(n3062), .A2(n3060), .A3(n3102), .ZN(n3043) );
  AOI22_X1 U35810 ( .A1(n4089), .A2(n3034), .B1(n3043), .B2(
        REG3_REG_1__SCAN_IN), .ZN(n3020) );
  OAI211_X1 U3582 ( .C1(n3022), .C2(n4097), .A(n3021), .B(n3020), .ZN(U3219)
         );
  INV_X1 U3583 ( .A(n3024), .ZN(n3025) );
  OAI22_X1 U3584 ( .A1(n3028), .A2(n3027), .B1(n3026), .B2(n3025), .ZN(n3038)
         );
  NAND2_X1 U3585 ( .A1(n3034), .A2(n3891), .ZN(n3030) );
  NAND2_X1 U3586 ( .A1(n3172), .A2(n3051), .ZN(n3029) );
  NAND2_X1 U3587 ( .A1(n3030), .A2(n3029), .ZN(n3032) );
  XNOR2_X1 U3588 ( .A(n3032), .B(n3031), .ZN(n3036) );
  NOR2_X1 U3589 ( .A1(n3165), .A2(n3433), .ZN(n3033) );
  AOI21_X1 U3590 ( .B1(n3034), .B2(n3431), .A(n3033), .ZN(n3035) );
  NAND2_X1 U3591 ( .A1(n3036), .A2(n3035), .ZN(n3047) );
  OAI21_X1 U3592 ( .B1(n3036), .B2(n3035), .A(n3047), .ZN(n3037) );
  NOR2_X1 U3593 ( .A1(n3038), .A2(n3037), .ZN(n3049) );
  AOI21_X1 U3594 ( .B1(n3038), .B2(n3037), .A(n3049), .ZN(n3041) );
  AOI22_X1 U3595 ( .A1(n4090), .A2(n4118), .B1(n3172), .B2(n4893), .ZN(n3040)
         );
  AOI22_X1 U3596 ( .A1(n4089), .A2(n3050), .B1(n3043), .B2(REG3_REG_2__SCAN_IN), .ZN(n3039) );
  OAI211_X1 U3597 ( .C1(n3041), .C2(n4097), .A(n3040), .B(n3039), .ZN(U3234)
         );
  INV_X1 U3598 ( .A(n3042), .ZN(n3046) );
  AOI22_X1 U3599 ( .A1(n4089), .A2(n4118), .B1(n3126), .B2(n4893), .ZN(n3045)
         );
  NAND2_X1 U3600 ( .A1(n3043), .A2(REG3_REG_0__SCAN_IN), .ZN(n3044) );
  OAI211_X1 U3601 ( .C1(n3046), .C2(n4097), .A(n3045), .B(n3044), .ZN(U3229)
         );
  INV_X1 U3602 ( .A(n3047), .ZN(n3048) );
  NOR2_X1 U3603 ( .A1(n3049), .A2(n3048), .ZN(n3057) );
  AOI22_X1 U3604 ( .A1(n3050), .A2(n3947), .B1(n3891), .B2(n3199), .ZN(n3072)
         );
  NAND2_X1 U3605 ( .A1(n3050), .A2(n3891), .ZN(n3053) );
  NAND2_X1 U3606 ( .A1(n3199), .A2(n3946), .ZN(n3052) );
  NAND2_X1 U3607 ( .A1(n3053), .A2(n3052), .ZN(n3055) );
  XNOR2_X1 U3608 ( .A(n3055), .B(n3948), .ZN(n3074) );
  XOR2_X1 U3609 ( .A(n3072), .B(n3074), .Z(n3056) );
  AOI21_X1 U3610 ( .B1(n3057), .B2(n3056), .A(n3854), .ZN(n3069) );
  NAND4_X1 U3611 ( .A1(n3060), .A2(n2980), .A3(n3059), .A4(n3058), .ZN(n3061)
         );
  NAND2_X1 U3612 ( .A1(n3061), .A2(STATE_REG_SCAN_IN), .ZN(n3063) );
  AND2_X2 U3613 ( .A1(n3063), .A2(n3062), .ZN(n4903) );
  AOI22_X1 U3614 ( .A1(n4090), .A2(n3034), .B1(n4089), .B2(n4116), .ZN(n3066)
         );
  AOI21_X1 U3615 ( .B1(n4893), .B2(n3199), .A(n3064), .ZN(n3065) );
  OAI211_X1 U3616 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4903), .A(n3066), .B(n3065), 
        .ZN(n3067) );
  INV_X1 U3617 ( .A(n3067), .ZN(n3068) );
  OAI21_X1 U3618 ( .B1(n3069), .B2(n4097), .A(n3068), .ZN(U3215) );
  NOR2_X1 U3619 ( .A1(n3133), .A2(n3433), .ZN(n3070) );
  AOI21_X1 U3620 ( .B1(n4116), .B2(n3947), .A(n3070), .ZN(n3075) );
  INV_X1 U3621 ( .A(n3075), .ZN(n3078) );
  INV_X2 U3622 ( .A(n3924), .ZN(n3946) );
  AOI22_X1 U3623 ( .A1(n4116), .A2(n3891), .B1(n3946), .B2(n3860), .ZN(n3071)
         );
  XNOR2_X1 U3624 ( .A(n3071), .B(n3948), .ZN(n3076) );
  INV_X1 U3625 ( .A(n3076), .ZN(n3077) );
  INV_X1 U3626 ( .A(n3072), .ZN(n3073) );
  NOR2_X1 U3627 ( .A1(n3074), .A2(n3073), .ZN(n3853) );
  XNOR2_X1 U3628 ( .A(n3076), .B(n3075), .ZN(n3857) );
  NAND2_X1 U3629 ( .A1(n4115), .A2(n3899), .ZN(n3080) );
  NAND2_X1 U3630 ( .A1(n3153), .A2(n3946), .ZN(n3079) );
  NAND2_X1 U3631 ( .A1(n3080), .A2(n3079), .ZN(n3081) );
  XNOR2_X1 U3632 ( .A(n3081), .B(n3031), .ZN(n3083) );
  AOI22_X1 U3633 ( .A1(n4115), .A2(n3947), .B1(n3899), .B2(n3153), .ZN(n3082)
         );
  OR2_X1 U3634 ( .A1(n3083), .A2(n3082), .ZN(n3114) );
  INV_X1 U3635 ( .A(n3114), .ZN(n3084) );
  AND2_X1 U3636 ( .A1(n3083), .A2(n3082), .ZN(n3113) );
  NOR2_X1 U3637 ( .A1(n3084), .A2(n3113), .ZN(n3085) );
  XNOR2_X1 U3638 ( .A(n2289), .B(n3085), .ZN(n3089) );
  AOI22_X1 U3639 ( .A1(n4089), .A2(n4816), .B1(n4090), .B2(n4116), .ZN(n3087)
         );
  NOR2_X1 U3640 ( .A1(STATE_REG_SCAN_IN), .A2(n2590), .ZN(n4656) );
  AOI21_X1 U3641 ( .B1(n4893), .B2(n3153), .A(n4656), .ZN(n3086) );
  OAI211_X1 U3642 ( .C1(n4903), .C2(n3154), .A(n3087), .B(n3086), .ZN(n3088)
         );
  AOI21_X1 U3643 ( .B1(n3089), .B2(n4898), .A(n3088), .ZN(n3090) );
  INV_X1 U3644 ( .A(n3090), .ZN(U3224) );
  OAI21_X1 U3645 ( .B1(n3684), .B2(n3092), .A(n3091), .ZN(n4775) );
  OAI21_X1 U3646 ( .B1(n3094), .B2(n3602), .A(n3093), .ZN(n3098) );
  NAND2_X1 U3647 ( .A1(n4120), .A2(n2260), .ZN(n3096) );
  NAND2_X1 U3648 ( .A1(n3034), .A2(n2263), .ZN(n3095) );
  OAI211_X1 U3649 ( .C1(n4819), .C2(n2997), .A(n3096), .B(n3095), .ZN(n3097)
         );
  AOI21_X1 U3650 ( .B1(n3098), .B2(n4821), .A(n3097), .ZN(n3099) );
  OAI21_X1 U3651 ( .B1(n3842), .B2(n4775), .A(n3099), .ZN(n4777) );
  INV_X1 U3652 ( .A(n4777), .ZN(n3112) );
  NAND4_X1 U3653 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n3104)
         );
  INV_X1 U3654 ( .A(n4775), .ZN(n3110) );
  OR2_X1 U3655 ( .A1(n2979), .A2(n4828), .ZN(n3147) );
  INV_X1 U3656 ( .A(n3147), .ZN(n3105) );
  AND2_X1 U3657 ( .A1(n4328), .A2(n3105), .ZN(n4869) );
  AND2_X1 U3658 ( .A1(n4406), .A2(n4828), .ZN(n3106) );
  NAND2_X1 U3659 ( .A1(n4328), .A2(n3106), .ZN(n4871) );
  NAND2_X1 U3660 ( .A1(n2998), .A2(n3126), .ZN(n3107) );
  NAND2_X1 U3661 ( .A1(n3107), .A2(n3171), .ZN(n4773) );
  INV_X1 U3662 ( .A(n4875), .ZN(n4859) );
  AOI22_X1 U3663 ( .A1(n4858), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4859), .ZN(n3108) );
  OAI21_X1 U3664 ( .B1(n4871), .B2(n4773), .A(n3108), .ZN(n3109) );
  AOI21_X1 U3665 ( .B1(n3110), .B2(n4869), .A(n3109), .ZN(n3111) );
  OAI21_X1 U3666 ( .B1(n3112), .B2(n4858), .A(n3111), .ZN(U3289) );
  AOI22_X1 U3667 ( .A1(n4816), .A2(n3899), .B1(n3946), .B2(n3176), .ZN(n3115)
         );
  XNOR2_X1 U3668 ( .A(n3268), .B(n3269), .ZN(n3116) );
  XNOR2_X1 U3669 ( .A(n3271), .B(n3116), .ZN(n3122) );
  INV_X1 U3670 ( .A(n4802), .ZN(n3120) );
  AOI22_X1 U3671 ( .A1(n4089), .A2(n4114), .B1(n4090), .B2(n4115), .ZN(n3119)
         );
  NOR2_X1 U3672 ( .A1(STATE_REG_SCAN_IN), .A2(n3117), .ZN(n4666) );
  AOI21_X1 U3673 ( .B1(n4092), .B2(n3176), .A(n4666), .ZN(n3118) );
  OAI211_X1 U3674 ( .C1(n4903), .C2(n3120), .A(n3119), .B(n3118), .ZN(n3121)
         );
  AOI21_X1 U3675 ( .B1(n3122), .B2(n4898), .A(n3121), .ZN(n3123) );
  INV_X1 U3676 ( .A(n3123), .ZN(U3236) );
  NAND2_X1 U3677 ( .A1(n4120), .A2(n3124), .ZN(n3601) );
  NAND2_X1 U3678 ( .A1(n3125), .A2(n3601), .ZN(n4769) );
  AND2_X1 U3679 ( .A1(n3127), .A2(n3126), .ZN(n4768) );
  INV_X1 U3680 ( .A(n3842), .ZN(n3403) );
  OAI21_X1 U3681 ( .B1(n3403), .B2(n4821), .A(n4769), .ZN(n3128) );
  OAI21_X1 U3682 ( .B1(n2551), .B2(n3778), .A(n3128), .ZN(n4766) );
  AOI211_X1 U3683 ( .C1(n4794), .C2(n4769), .A(n4768), .B(n4766), .ZN(n4764)
         );
  NAND2_X1 U3684 ( .A1(n4844), .A2(REG1_REG_0__SCAN_IN), .ZN(n3129) );
  OAI21_X1 U3685 ( .B1(n4764), .B2(n4844), .A(n3129), .ZN(U3518) );
  INV_X1 U3686 ( .A(n3208), .ZN(n3130) );
  OAI211_X1 U3687 ( .C1(n3130), .C2(n3133), .A(n4406), .B(n3152), .ZN(n4791)
         );
  NOR2_X1 U3688 ( .A1(n4791), .A2(n4450), .ZN(n3141) );
  INV_X1 U3689 ( .A(n4821), .ZN(n4344) );
  XNOR2_X1 U3690 ( .A(n3131), .B(n3686), .ZN(n3140) );
  NAND2_X1 U3691 ( .A1(n3050), .A2(n2260), .ZN(n3132) );
  OAI21_X1 U3692 ( .B1(n4819), .B2(n3133), .A(n3132), .ZN(n3138) );
  NAND2_X1 U3693 ( .A1(n3134), .A2(n2432), .ZN(n3135) );
  NAND2_X1 U3694 ( .A1(n3136), .A2(n3135), .ZN(n3142) );
  NOR2_X1 U3695 ( .A1(n3142), .A2(n3842), .ZN(n3137) );
  AOI211_X1 U3696 ( .C1(n2263), .C2(n4115), .A(n3138), .B(n3137), .ZN(n3139)
         );
  OAI21_X1 U3697 ( .B1(n4344), .B2(n3140), .A(n3139), .ZN(n4792) );
  AOI211_X1 U3698 ( .C1(n4859), .C2(n3858), .A(n3141), .B(n4792), .ZN(n3144)
         );
  INV_X1 U3699 ( .A(n3142), .ZN(n4795) );
  AOI22_X1 U3700 ( .A1(n4795), .A2(n4869), .B1(REG2_REG_4__SCAN_IN), .B2(n4858), .ZN(n3143) );
  OAI21_X1 U3701 ( .B1(n3144), .B2(n4858), .A(n3143), .ZN(U3286) );
  INV_X1 U3702 ( .A(n3145), .ZN(n3612) );
  NAND2_X1 U3703 ( .A1(n3612), .A2(n3585), .ZN(n3677) );
  XOR2_X1 U3704 ( .A(n3146), .B(n3677), .Z(n3192) );
  INV_X1 U3705 ( .A(n3192), .ZN(n3160) );
  INV_X2 U3706 ( .A(n4858), .ZN(n4328) );
  NAND2_X1 U3707 ( .A1(n3842), .A2(n3147), .ZN(n4833) );
  NAND2_X1 U3708 ( .A1(n4328), .A2(n4833), .ZN(n4353) );
  XOR2_X1 U3709 ( .A(n3677), .B(n3148), .Z(n3151) );
  AOI22_X1 U3710 ( .A1(n4116), .A2(n2260), .B1(n3153), .B2(n4359), .ZN(n3150)
         );
  NAND2_X1 U3711 ( .A1(n4816), .A2(n2263), .ZN(n3149) );
  OAI211_X1 U3712 ( .C1(n3151), .C2(n4344), .A(n3150), .B(n3149), .ZN(n3191)
         );
  NAND2_X1 U3713 ( .A1(n3191), .A2(n4328), .ZN(n3159) );
  AOI21_X1 U3714 ( .B1(n3153), .B2(n3152), .A(n3183), .ZN(n3210) );
  NOR2_X1 U3715 ( .A1(n3154), .A2(n4875), .ZN(n3157) );
  INV_X1 U3716 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3155) );
  NOR2_X1 U3717 ( .A1(n4328), .A2(n3155), .ZN(n3156) );
  AOI211_X1 U3718 ( .C1(n3210), .C2(n4908), .A(n3157), .B(n3156), .ZN(n3158)
         );
  OAI211_X1 U3719 ( .C1(n3160), .C2(n4353), .A(n3159), .B(n3158), .ZN(U3285)
         );
  OAI21_X1 U3720 ( .B1(n3162), .B2(n3685), .A(n3161), .ZN(n4782) );
  NAND2_X1 U3721 ( .A1(n4118), .A2(n2260), .ZN(n3164) );
  NAND2_X1 U3722 ( .A1(n3050), .A2(n2263), .ZN(n3163) );
  OAI211_X1 U3723 ( .C1(n4819), .C2(n3165), .A(n3164), .B(n3163), .ZN(n3169)
         );
  XNOR2_X1 U3724 ( .A(n3166), .B(n3685), .ZN(n3167) );
  NOR2_X1 U3725 ( .A1(n3167), .A2(n4344), .ZN(n3168) );
  AOI211_X1 U3726 ( .C1(n3403), .C2(n4782), .A(n3169), .B(n3168), .ZN(n4785)
         );
  INV_X1 U3727 ( .A(n4785), .ZN(n3170) );
  AOI21_X1 U3728 ( .B1(n4794), .B2(n4782), .A(n3170), .ZN(n3214) );
  AOI21_X1 U3729 ( .B1(n3172), .B2(n3171), .A(n3206), .ZN(n4781) );
  INV_X1 U3730 ( .A(n4442), .ZN(n3307) );
  AOI22_X1 U3731 ( .A1(n4781), .A2(n3307), .B1(REG0_REG_2__SCAN_IN), .B2(n4414), .ZN(n3173) );
  OAI21_X1 U3732 ( .B1(n3214), .B2(n4414), .A(n3173), .ZN(U3471) );
  AND2_X1 U3733 ( .A1(n4811), .A2(n3613), .ZN(n3664) );
  XNOR2_X1 U3734 ( .A(n3174), .B(n3664), .ZN(n4805) );
  INV_X1 U3735 ( .A(n4805), .ZN(n3181) );
  XOR2_X1 U3736 ( .A(n3664), .B(n3175), .Z(n3179) );
  AOI22_X1 U3737 ( .A1(n4114), .A2(n2263), .B1(n3176), .B2(n4359), .ZN(n3178)
         );
  NAND2_X1 U3738 ( .A1(n4115), .A2(n2260), .ZN(n3177) );
  OAI211_X1 U3739 ( .C1(n3179), .C2(n4344), .A(n3178), .B(n3177), .ZN(n3180)
         );
  AOI21_X1 U3740 ( .B1(n3403), .B2(n4805), .A(n3180), .ZN(n4808) );
  OAI21_X1 U3741 ( .B1(n4774), .B2(n3181), .A(n4808), .ZN(n3189) );
  OAI21_X1 U3742 ( .B1(n3183), .B2(n3182), .A(n4825), .ZN(n4803) );
  INV_X1 U3743 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3184) );
  OAI22_X1 U3744 ( .A1(n4803), .A2(n4396), .B1(n4846), .B2(n3184), .ZN(n3185)
         );
  AOI21_X1 U3745 ( .B1(n3189), .B2(n4411), .A(n3185), .ZN(n3186) );
  INV_X1 U3746 ( .A(n3186), .ZN(U3524) );
  INV_X1 U3747 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3187) );
  OAI22_X1 U3748 ( .A1(n4803), .A2(n4442), .B1(n4849), .B2(n3187), .ZN(n3188)
         );
  AOI21_X1 U3749 ( .B1(n3189), .B2(n4849), .A(n3188), .ZN(n3190) );
  INV_X1 U3750 ( .A(n3190), .ZN(U3479) );
  AOI21_X1 U3751 ( .B1(n3192), .B2(n4840), .A(n3191), .ZN(n3212) );
  AOI22_X1 U3752 ( .A1(n3210), .A2(n3307), .B1(REG0_REG_5__SCAN_IN), .B2(n4414), .ZN(n3193) );
  OAI21_X1 U3753 ( .B1(n3212), .B2(n4414), .A(n3193), .ZN(U3477) );
  XNOR2_X1 U3754 ( .A(n3194), .B(n3683), .ZN(n4787) );
  INV_X1 U3755 ( .A(n3034), .ZN(n3202) );
  INV_X1 U3756 ( .A(n2260), .ZN(n4339) );
  OAI21_X1 U3757 ( .B1(n3197), .B2(n3196), .A(n3195), .ZN(n3198) );
  NAND2_X1 U3758 ( .A1(n3198), .A2(n4821), .ZN(n3201) );
  AOI22_X1 U3759 ( .A1(n4116), .A2(n2263), .B1(n4359), .B2(n3199), .ZN(n3200)
         );
  OAI211_X1 U3760 ( .C1(n3202), .C2(n4339), .A(n3201), .B(n3200), .ZN(n3203)
         );
  AOI21_X1 U3761 ( .B1(n3403), .B2(n4787), .A(n3203), .ZN(n4790) );
  INV_X1 U3762 ( .A(n4790), .ZN(n3204) );
  AOI21_X1 U3763 ( .B1(n4794), .B2(n4787), .A(n3204), .ZN(n3216) );
  OR2_X1 U3764 ( .A1(n3206), .A2(n3205), .ZN(n3207) );
  AND2_X1 U3765 ( .A1(n3208), .A2(n3207), .ZN(n4786) );
  AOI22_X1 U3766 ( .A1(n4786), .A2(n3307), .B1(REG0_REG_3__SCAN_IN), .B2(n4414), .ZN(n3209) );
  OAI21_X1 U3767 ( .B1(n3216), .B2(n4414), .A(n3209), .ZN(U3473) );
  INV_X1 U3768 ( .A(n4396), .ZN(n3303) );
  AOI22_X1 U3769 ( .A1(n3210), .A2(n3303), .B1(REG1_REG_5__SCAN_IN), .B2(n4844), .ZN(n3211) );
  OAI21_X1 U3770 ( .B1(n3212), .B2(n4844), .A(n3211), .ZN(U3523) );
  AOI22_X1 U3771 ( .A1(n4781), .A2(n3303), .B1(REG1_REG_2__SCAN_IN), .B2(n4844), .ZN(n3213) );
  OAI21_X1 U3772 ( .B1(n3214), .B2(n4844), .A(n3213), .ZN(U3520) );
  AOI22_X1 U3773 ( .A1(n4786), .A2(n3303), .B1(REG1_REG_3__SCAN_IN), .B2(n4844), .ZN(n3215) );
  OAI21_X1 U3774 ( .B1(n3216), .B2(n4844), .A(n3215), .ZN(U3521) );
  INV_X1 U3775 ( .A(n3619), .ZN(n3218) );
  AND2_X1 U3776 ( .A1(n3218), .A2(n3621), .ZN(n3663) );
  XNOR2_X1 U3777 ( .A(n3217), .B(n3663), .ZN(n3262) );
  INV_X1 U3778 ( .A(n3262), .ZN(n3228) );
  INV_X1 U3779 ( .A(n3301), .ZN(n3219) );
  AOI21_X1 U3780 ( .B1(n3319), .B2(n3219), .A(n3340), .ZN(n3264) );
  INV_X1 U3781 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3220) );
  OAI22_X1 U3782 ( .A1(n3322), .A2(n4875), .B1(n3220), .B2(n4328), .ZN(n3221)
         );
  AOI21_X1 U3783 ( .B1(n3264), .B2(n4908), .A(n3221), .ZN(n3227) );
  XNOR2_X1 U3784 ( .A(n3222), .B(n3663), .ZN(n3225) );
  AOI22_X1 U3785 ( .A1(n4814), .A2(n2260), .B1(n4359), .B2(n3319), .ZN(n3224)
         );
  NAND2_X1 U3786 ( .A1(n4112), .A2(n2263), .ZN(n3223) );
  OAI211_X1 U3787 ( .C1(n3225), .C2(n4344), .A(n3224), .B(n3223), .ZN(n3261)
         );
  NAND2_X1 U3788 ( .A1(n3261), .A2(n4328), .ZN(n3226) );
  OAI211_X1 U3789 ( .C1(n3228), .C2(n4353), .A(n3227), .B(n3226), .ZN(U3281)
         );
  INV_X1 U3790 ( .A(n4759), .ZN(n4182) );
  INV_X1 U3791 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4550) );
  NOR2_X1 U3792 ( .A1(STATE_REG_SCAN_IN), .A2(n4550), .ZN(n3318) );
  AOI21_X1 U3793 ( .B1(n4757), .B2(ADDR_REG_9__SCAN_IN), .A(n3318), .ZN(n3229)
         );
  INV_X1 U3794 ( .A(n3229), .ZN(n3242) );
  INV_X1 U3795 ( .A(n4673), .ZN(n4810) );
  INV_X1 U3796 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4845) );
  NOR2_X1 U3797 ( .A1(n4810), .A2(n4845), .ZN(n4679) );
  NAND2_X1 U3798 ( .A1(n3247), .A2(REG1_REG_5__SCAN_IN), .ZN(n3233) );
  INV_X1 U3799 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3230) );
  INV_X1 U3800 ( .A(n3247), .ZN(n4799) );
  AOI22_X1 U3801 ( .A1(n3247), .A2(REG1_REG_5__SCAN_IN), .B1(n3230), .B2(n4799), .ZN(n4660) );
  INV_X1 U3802 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U3803 ( .A1(n4660), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U3804 ( .A1(n3250), .A2(n3234), .ZN(n3235) );
  OAI22_X1 U3805 ( .A1(n4679), .A2(n4681), .B1(n4673), .B2(REG1_REG_7__SCAN_IN), .ZN(n3236) );
  NOR2_X1 U3806 ( .A1(n3254), .A2(n3236), .ZN(n3237) );
  INV_X1 U3807 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4687) );
  XNOR2_X1 U3808 ( .A(n3254), .B(n3236), .ZN(n4686) );
  NAND2_X1 U3809 ( .A1(n4452), .A2(REG1_REG_9__SCAN_IN), .ZN(n4156) );
  NOR2_X1 U3810 ( .A1(n4452), .A2(REG1_REG_9__SCAN_IN), .ZN(n4157) );
  INV_X1 U3811 ( .A(n4157), .ZN(n3238) );
  NAND2_X1 U3812 ( .A1(n4156), .A2(n3238), .ZN(n3240) );
  OAI21_X1 U3813 ( .B1(n4158), .B2(n3240), .A(n4744), .ZN(n3239) );
  AOI21_X1 U3814 ( .B1(n4158), .B2(n3240), .A(n3239), .ZN(n3241) );
  AOI211_X1 U3815 ( .C1(n4182), .C2(n4452), .A(n3242), .B(n3241), .ZN(n3260)
         );
  INV_X1 U3816 ( .A(n3244), .ZN(n3246) );
  NAND2_X1 U3817 ( .A1(n3247), .A2(REG2_REG_5__SCAN_IN), .ZN(n3248) );
  OAI21_X1 U3818 ( .B1(n3247), .B2(REG2_REG_5__SCAN_IN), .A(n3248), .ZN(n4654)
         );
  INV_X1 U3819 ( .A(n3250), .ZN(n4801) );
  NOR2_X1 U3820 ( .A1(n3251), .A2(n4801), .ZN(n3252) );
  INV_X1 U3821 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4665) );
  INV_X1 U3822 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U3823 ( .A1(n3253), .A2(n3255), .ZN(n3256) );
  NAND2_X1 U3824 ( .A1(n3256), .A2(n4690), .ZN(n3258) );
  MUX2_X1 U3825 ( .A(REG2_REG_9__SCAN_IN), .B(n3220), .S(n4452), .Z(n3257) );
  NAND2_X1 U3826 ( .A1(n3257), .A2(n3258), .ZN(n4147) );
  OAI211_X1 U3827 ( .C1(n3258), .C2(n3257), .A(n4761), .B(n4147), .ZN(n3259)
         );
  NAND2_X1 U3828 ( .A1(n3260), .A2(n3259), .ZN(U3249) );
  AOI21_X1 U3829 ( .B1(n3262), .B2(n4840), .A(n3261), .ZN(n3266) );
  AOI22_X1 U3830 ( .A1(n3264), .A2(n3303), .B1(REG1_REG_9__SCAN_IN), .B2(n4844), .ZN(n3263) );
  OAI21_X1 U3831 ( .B1(n3266), .B2(n4844), .A(n3263), .ZN(U3527) );
  AOI22_X1 U3832 ( .A1(n3264), .A2(n3307), .B1(REG0_REG_9__SCAN_IN), .B2(n4414), .ZN(n3265) );
  OAI21_X1 U3833 ( .B1(n3266), .B2(n4414), .A(n3265), .ZN(U3485) );
  AOI22_X1 U3834 ( .A1(n4114), .A2(n3899), .B1(n3946), .B2(n4824), .ZN(n3267)
         );
  XNOR2_X1 U3835 ( .A(n3267), .B(n3948), .ZN(n3277) );
  AOI22_X1 U3836 ( .A1(n4114), .A2(n3947), .B1(n3899), .B2(n4824), .ZN(n3278)
         );
  XNOR2_X1 U3837 ( .A(n3277), .B(n3278), .ZN(n3279) );
  XOR2_X1 U3838 ( .A(n3279), .B(n3280), .Z(n3275) );
  AOI22_X1 U3839 ( .A1(n4090), .A2(n4816), .B1(n4089), .B2(n4814), .ZN(n3273)
         );
  AND2_X1 U3840 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4677) );
  AOI21_X1 U3841 ( .B1(n4092), .B2(n4824), .A(n4677), .ZN(n3272) );
  OAI211_X1 U3842 ( .C1(n4903), .C2(n4838), .A(n3273), .B(n3272), .ZN(n3274)
         );
  AOI21_X1 U3843 ( .B1(n3275), .B2(n4898), .A(n3274), .ZN(n3276) );
  INV_X1 U3844 ( .A(n3276), .ZN(U3210) );
  NAND2_X1 U3845 ( .A1(n4814), .A2(n3899), .ZN(n3282) );
  NAND2_X1 U3846 ( .A1(n3302), .A2(n3946), .ZN(n3281) );
  NAND2_X1 U3847 ( .A1(n3282), .A2(n3281), .ZN(n3283) );
  XNOR2_X1 U3848 ( .A(n3283), .B(n3031), .ZN(n3285) );
  AOI22_X1 U3849 ( .A1(n4814), .A2(n3947), .B1(n3899), .B2(n3302), .ZN(n3284)
         );
  NOR2_X1 U3850 ( .A1(n3285), .A2(n3284), .ZN(n3314) );
  INV_X1 U3851 ( .A(n3314), .ZN(n3286) );
  NAND2_X1 U3852 ( .A1(n3285), .A2(n3284), .ZN(n3313) );
  NAND2_X1 U3853 ( .A1(n3286), .A2(n3313), .ZN(n3287) );
  XNOR2_X1 U3854 ( .A(n3315), .B(n3287), .ZN(n3292) );
  INV_X1 U3855 ( .A(n4851), .ZN(n3290) );
  AOI22_X1 U3856 ( .A1(n4089), .A2(n4113), .B1(n4090), .B2(n4114), .ZN(n3289)
         );
  INV_X1 U3857 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4613) );
  NOR2_X1 U3858 ( .A1(STATE_REG_SCAN_IN), .A2(n4613), .ZN(n4688) );
  AOI21_X1 U3859 ( .B1(n4893), .B2(n3302), .A(n4688), .ZN(n3288) );
  OAI211_X1 U3860 ( .C1(n4903), .C2(n3290), .A(n3289), .B(n3288), .ZN(n3291)
         );
  AOI21_X1 U3861 ( .B1(n3292), .B2(n4898), .A(n3291), .ZN(n3293) );
  INV_X1 U3862 ( .A(n3293), .ZN(U3218) );
  NAND2_X1 U3863 ( .A1(n3620), .A2(n3583), .ZN(n3674) );
  XOR2_X1 U3864 ( .A(n3674), .B(n3294), .Z(n4853) );
  XOR2_X1 U3865 ( .A(n3674), .B(n3295), .Z(n3298) );
  AOI22_X1 U3866 ( .A1(n4113), .A2(n2263), .B1(n3302), .B2(n4359), .ZN(n3297)
         );
  NAND2_X1 U3867 ( .A1(n4114), .A2(n2260), .ZN(n3296) );
  OAI211_X1 U3868 ( .C1(n3298), .C2(n4344), .A(n3297), .B(n3296), .ZN(n3299)
         );
  AOI21_X1 U3869 ( .B1(n4853), .B2(n3403), .A(n3299), .ZN(n4856) );
  INV_X1 U3870 ( .A(n4856), .ZN(n3300) );
  AOI21_X1 U3871 ( .B1(n4794), .B2(n4853), .A(n3300), .ZN(n3309) );
  AOI21_X1 U3872 ( .B1(n3302), .B2(n4826), .A(n3301), .ZN(n4852) );
  AOI22_X1 U3873 ( .A1(n4852), .A2(n3303), .B1(n4844), .B2(REG1_REG_8__SCAN_IN), .ZN(n3304) );
  OAI21_X1 U3874 ( .B1(n3309), .B2(n4844), .A(n3304), .ZN(U3526) );
  INV_X1 U3875 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3305) );
  NOR2_X1 U3876 ( .A1(n4849), .A2(n3305), .ZN(n3306) );
  AOI21_X1 U3877 ( .B1(n4852), .B2(n3307), .A(n3306), .ZN(n3308) );
  OAI21_X1 U3878 ( .B1(n3309), .B2(n4414), .A(n3308), .ZN(U3483) );
  NAND2_X1 U3879 ( .A1(n4113), .A2(n3899), .ZN(n3311) );
  NAND2_X1 U3880 ( .A1(n3319), .A2(n3946), .ZN(n3310) );
  NAND2_X1 U3881 ( .A1(n3311), .A2(n3310), .ZN(n3312) );
  XNOR2_X1 U3882 ( .A(n3312), .B(n3948), .ZN(n3354) );
  AOI22_X1 U3883 ( .A1(n4113), .A2(n3947), .B1(n3899), .B2(n3319), .ZN(n3355)
         );
  XNOR2_X1 U3884 ( .A(n3354), .B(n3355), .ZN(n3317) );
  OAI21_X1 U3885 ( .B1(n3315), .B2(n3314), .A(n3313), .ZN(n3316) );
  NAND2_X1 U3886 ( .A1(n3316), .A2(n3317), .ZN(n3980) );
  OAI21_X1 U3887 ( .B1(n3317), .B2(n3316), .A(n3980), .ZN(n3324) );
  AOI22_X1 U3888 ( .A1(n4090), .A2(n4814), .B1(n4089), .B2(n4112), .ZN(n3321)
         );
  AOI21_X1 U3889 ( .B1(n4092), .B2(n3319), .A(n3318), .ZN(n3320) );
  OAI211_X1 U3890 ( .C1(n4903), .C2(n3322), .A(n3321), .B(n3320), .ZN(n3323)
         );
  AOI21_X1 U3891 ( .B1(n3324), .B2(n4898), .A(n3323), .ZN(n3325) );
  INV_X1 U3892 ( .A(n3325), .ZN(U3228) );
  NAND2_X1 U3893 ( .A1(n3381), .A2(n3379), .ZN(n3676) );
  XNOR2_X1 U3894 ( .A(n3326), .B(n3676), .ZN(n3420) );
  INV_X1 U3895 ( .A(n3420), .ZN(n3338) );
  INV_X1 U3896 ( .A(n3327), .ZN(n3328) );
  AOI21_X1 U3897 ( .B1(n3405), .B2(n3329), .A(n3328), .ZN(n3382) );
  XOR2_X1 U3898 ( .A(n3676), .B(n3382), .Z(n3332) );
  AOI22_X1 U3899 ( .A1(n4111), .A2(n2260), .B1(n3436), .B2(n4359), .ZN(n3331)
         );
  NAND2_X1 U3900 ( .A1(n4109), .A2(n2263), .ZN(n3330) );
  OAI211_X1 U3901 ( .C1(n3332), .C2(n4344), .A(n3331), .B(n3330), .ZN(n3419)
         );
  AND2_X1 U3902 ( .A1(n3398), .A2(n3436), .ZN(n3333) );
  OR2_X1 U3903 ( .A1(n3333), .A2(n3390), .ZN(n3425) );
  AOI22_X1 U3904 ( .A1(n4858), .A2(REG2_REG_12__SCAN_IN), .B1(n3334), .B2(
        n4859), .ZN(n3335) );
  OAI21_X1 U3905 ( .B1(n3425), .B2(n4871), .A(n3335), .ZN(n3336) );
  AOI21_X1 U3906 ( .B1(n3419), .B2(n4328), .A(n3336), .ZN(n3337) );
  OAI21_X1 U3907 ( .B1(n3338), .B2(n4353), .A(n3337), .ZN(U3278) );
  OAI21_X1 U3908 ( .B1(n3340), .B2(n3339), .A(n3397), .ZN(n4861) );
  INV_X1 U3909 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U3910 ( .A1(n3592), .A2(n3588), .ZN(n3675) );
  XNOR2_X1 U3911 ( .A(n3341), .B(n3675), .ZN(n4863) );
  XNOR2_X1 U3912 ( .A(n3342), .B(n3675), .ZN(n3345) );
  AOI22_X1 U3913 ( .A1(n4111), .A2(n2263), .B1(n4359), .B2(n3985), .ZN(n3344)
         );
  NAND2_X1 U3914 ( .A1(n4113), .A2(n2260), .ZN(n3343) );
  OAI211_X1 U3915 ( .C1(n3345), .C2(n4344), .A(n3344), .B(n3343), .ZN(n3346)
         );
  AOI21_X1 U3916 ( .B1(n3403), .B2(n4863), .A(n3346), .ZN(n4866) );
  INV_X1 U3917 ( .A(n4866), .ZN(n3347) );
  AOI21_X1 U3918 ( .B1(n4794), .B2(n4863), .A(n3347), .ZN(n3350) );
  MUX2_X1 U3919 ( .A(n3348), .B(n3350), .S(n4411), .Z(n3349) );
  OAI21_X1 U3920 ( .B1(n4861), .B2(n4396), .A(n3349), .ZN(U3528) );
  INV_X1 U3921 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3351) );
  MUX2_X1 U3922 ( .A(n3351), .B(n3350), .S(n4849), .Z(n3352) );
  OAI21_X1 U3923 ( .B1(n4861), .B2(n4442), .A(n3352), .ZN(U3487) );
  AOI22_X1 U3924 ( .A1(n4112), .A2(n3947), .B1(n3899), .B2(n3985), .ZN(n3358)
         );
  AOI22_X1 U3925 ( .A1(n4112), .A2(n3899), .B1(n3946), .B2(n3985), .ZN(n3353)
         );
  XNOR2_X1 U3926 ( .A(n3353), .B(n3948), .ZN(n3359) );
  XOR2_X1 U3927 ( .A(n3358), .B(n3359), .Z(n3982) );
  INV_X1 U3928 ( .A(n3354), .ZN(n3356) );
  NAND2_X1 U3929 ( .A1(n3356), .A2(n3355), .ZN(n3979) );
  NAND2_X1 U3930 ( .A1(n3980), .A2(n3357), .ZN(n3981) );
  NAND2_X1 U3931 ( .A1(n3981), .A2(n3360), .ZN(n3426) );
  NAND2_X1 U3932 ( .A1(n4111), .A2(n3899), .ZN(n3362) );
  NAND2_X1 U3933 ( .A1(n3370), .A2(n3946), .ZN(n3361) );
  NAND2_X1 U3934 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  XNOR2_X1 U3935 ( .A(n3363), .B(n3948), .ZN(n3367) );
  NAND2_X1 U3936 ( .A1(n4111), .A2(n3947), .ZN(n3365) );
  NAND2_X1 U3937 ( .A1(n3370), .A2(n3899), .ZN(n3364) );
  NAND2_X1 U3938 ( .A1(n3365), .A2(n3364), .ZN(n3366) );
  NOR2_X1 U3939 ( .A1(n3367), .A2(n3366), .ZN(n3428) );
  INV_X1 U3940 ( .A(n3428), .ZN(n3368) );
  NAND2_X1 U3941 ( .A1(n3367), .A2(n3366), .ZN(n3427) );
  NAND2_X1 U3942 ( .A1(n3368), .A2(n3427), .ZN(n3369) );
  XNOR2_X1 U3943 ( .A(n3426), .B(n3369), .ZN(n3374) );
  AOI22_X1 U3944 ( .A1(n4090), .A2(n4112), .B1(n4089), .B2(n4110), .ZN(n3372)
         );
  AND2_X1 U3945 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4709) );
  AOI21_X1 U3946 ( .B1(n4092), .B2(n3370), .A(n4709), .ZN(n3371) );
  OAI211_X1 U3947 ( .C1(n4903), .C2(n4876), .A(n3372), .B(n3371), .ZN(n3373)
         );
  AOI21_X1 U3948 ( .B1(n3374), .B2(n4898), .A(n3373), .ZN(n3375) );
  INV_X1 U3949 ( .A(n3375), .ZN(U3233) );
  INV_X1 U3950 ( .A(n3443), .ZN(n3376) );
  OR2_X1 U3951 ( .A1(n3377), .A2(n3376), .ZN(n3668) );
  XNOR2_X1 U3952 ( .A(n3378), .B(n3668), .ZN(n3388) );
  INV_X1 U3953 ( .A(n3379), .ZN(n3380) );
  AOI21_X1 U3954 ( .B1(n3382), .B2(n3381), .A(n3380), .ZN(n3383) );
  XNOR2_X1 U3955 ( .A(n3383), .B(n3668), .ZN(n3386) );
  INV_X1 U3956 ( .A(n4110), .ZN(n3434) );
  AOI22_X1 U3957 ( .A1(n4886), .A2(n2263), .B1(n3509), .B2(n4359), .ZN(n3384)
         );
  OAI21_X1 U3958 ( .B1(n3434), .B2(n4339), .A(n3384), .ZN(n3385) );
  AOI21_X1 U3959 ( .B1(n3386), .B2(n4821), .A(n3385), .ZN(n3387) );
  OAI21_X1 U3960 ( .B1(n3388), .B2(n3842), .A(n3387), .ZN(n3460) );
  INV_X1 U3961 ( .A(n3460), .ZN(n3396) );
  INV_X1 U3962 ( .A(n3388), .ZN(n3461) );
  NOR2_X1 U3963 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  OR2_X1 U3964 ( .A1(n3453), .A2(n3391), .ZN(n3467) );
  AOI22_X1 U3965 ( .A1(n4858), .A2(REG2_REG_13__SCAN_IN), .B1(n3392), .B2(
        n4859), .ZN(n3393) );
  OAI21_X1 U3966 ( .B1(n3467), .B2(n4871), .A(n3393), .ZN(n3394) );
  AOI21_X1 U3967 ( .B1(n3461), .B2(n4869), .A(n3394), .ZN(n3395) );
  OAI21_X1 U3968 ( .B1(n3396), .B2(n4858), .A(n3395), .ZN(U3277) );
  INV_X1 U3969 ( .A(n3397), .ZN(n3399) );
  OAI21_X1 U3970 ( .B1(n3399), .B2(n3408), .A(n3398), .ZN(n4870) );
  NAND2_X1 U3971 ( .A1(n3400), .A2(n3404), .ZN(n3401) );
  NAND2_X1 U3972 ( .A1(n3402), .A2(n3401), .ZN(n4868) );
  NAND2_X1 U3973 ( .A1(n4868), .A2(n3403), .ZN(n3412) );
  XNOR2_X1 U3974 ( .A(n3405), .B(n3404), .ZN(n3410) );
  NAND2_X1 U3975 ( .A1(n4112), .A2(n2260), .ZN(n3407) );
  NAND2_X1 U3976 ( .A1(n4110), .A2(n2263), .ZN(n3406) );
  OAI211_X1 U3977 ( .C1(n4819), .C2(n3408), .A(n3407), .B(n3406), .ZN(n3409)
         );
  AOI21_X1 U3978 ( .B1(n3410), .B2(n4821), .A(n3409), .ZN(n3411) );
  AND2_X1 U3979 ( .A1(n3412), .A2(n3411), .ZN(n4880) );
  NAND2_X1 U3980 ( .A1(n4868), .A2(n4794), .ZN(n3413) );
  NAND2_X1 U3981 ( .A1(n4880), .A2(n3413), .ZN(n3416) );
  MUX2_X1 U3982 ( .A(REG1_REG_11__SCAN_IN), .B(n3416), .S(n4846), .Z(n3414) );
  INV_X1 U3983 ( .A(n3414), .ZN(n3415) );
  OAI21_X1 U3984 ( .B1(n4396), .B2(n4870), .A(n3415), .ZN(U3529) );
  MUX2_X1 U3985 ( .A(REG0_REG_11__SCAN_IN), .B(n3416), .S(n4849), .Z(n3417) );
  INV_X1 U3986 ( .A(n3417), .ZN(n3418) );
  OAI21_X1 U3987 ( .B1(n4870), .B2(n4442), .A(n3418), .ZN(U3489) );
  INV_X1 U3988 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3421) );
  AOI21_X1 U3989 ( .B1(n4840), .B2(n3420), .A(n3419), .ZN(n3423) );
  MUX2_X1 U3990 ( .A(n3421), .B(n3423), .S(n4849), .Z(n3422) );
  OAI21_X1 U3991 ( .B1(n3425), .B2(n4442), .A(n3422), .ZN(U3491) );
  INV_X1 U3992 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4718) );
  MUX2_X1 U3993 ( .A(n4718), .B(n3423), .S(n4411), .Z(n3424) );
  OAI21_X1 U3994 ( .B1(n3425), .B2(n4396), .A(n3424), .ZN(U3530) );
  INV_X1 U3995 ( .A(n3426), .ZN(n3429) );
  AOI22_X1 U3996 ( .A1(n4110), .A2(n3899), .B1(n3946), .B2(n3436), .ZN(n3430)
         );
  XOR2_X1 U3997 ( .A(n3948), .B(n3430), .Z(n3500) );
  INV_X1 U3998 ( .A(n3431), .ZN(n3926) );
  OAI22_X1 U3999 ( .A1(n3434), .A2(n3926), .B1(n3433), .B2(n3432), .ZN(n3501)
         );
  XNOR2_X1 U4000 ( .A(n3500), .B(n3501), .ZN(n3435) );
  XNOR2_X1 U4001 ( .A(n3502), .B(n3435), .ZN(n3441) );
  AOI22_X1 U4002 ( .A1(n4090), .A2(n4111), .B1(n4089), .B2(n4109), .ZN(n3438)
         );
  INV_X1 U4003 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4616) );
  NOR2_X1 U4004 ( .A1(STATE_REG_SCAN_IN), .A2(n4616), .ZN(n4719) );
  AOI21_X1 U4005 ( .B1(n4893), .B2(n3436), .A(n4719), .ZN(n3437) );
  OAI211_X1 U4006 ( .C1(n4903), .C2(n3439), .A(n3438), .B(n3437), .ZN(n3440)
         );
  AOI21_X1 U4007 ( .B1(n3441), .B2(n4898), .A(n3440), .ZN(n3442) );
  INV_X1 U4008 ( .A(n3442), .ZN(U3221) );
  AND2_X1 U4009 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  NAND2_X1 U4010 ( .A1(n3445), .A2(n3688), .ZN(n3484) );
  OAI21_X1 U4011 ( .B1(n3445), .B2(n3688), .A(n3484), .ZN(n3517) );
  INV_X1 U4012 ( .A(n3517), .ZN(n3459) );
  INV_X1 U4013 ( .A(n4108), .ZN(n3451) );
  OAI21_X1 U4014 ( .B1(n3446), .B2(n3706), .A(n3486), .ZN(n3447) );
  NAND2_X1 U4015 ( .A1(n3447), .A2(n4821), .ZN(n3450) );
  NOR2_X1 U4016 ( .A1(n3452), .A2(n4819), .ZN(n3448) );
  AOI21_X1 U4017 ( .B1(n4109), .B2(n2260), .A(n3448), .ZN(n3449) );
  OAI211_X1 U4018 ( .C1(n3451), .C2(n3778), .A(n3450), .B(n3449), .ZN(n3516)
         );
  OAI21_X1 U4019 ( .B1(n3453), .B2(n3452), .A(n3491), .ZN(n3523) );
  NOR2_X1 U4020 ( .A1(n3523), .A2(n4871), .ZN(n3457) );
  INV_X1 U4021 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3455) );
  INV_X1 U4022 ( .A(n3454), .ZN(n3531) );
  OAI22_X1 U4023 ( .A1(n4328), .A2(n3455), .B1(n3531), .B2(n4875), .ZN(n3456)
         );
  AOI211_X1 U4024 ( .C1(n3516), .C2(n4328), .A(n3457), .B(n3456), .ZN(n3458)
         );
  OAI21_X1 U4025 ( .B1(n3459), .B2(n4353), .A(n3458), .ZN(U3276) );
  INV_X1 U4026 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3462) );
  AOI21_X1 U4027 ( .B1(n4794), .B2(n3461), .A(n3460), .ZN(n3464) );
  MUX2_X1 U4028 ( .A(n3462), .B(n3464), .S(n4411), .Z(n3463) );
  OAI21_X1 U4029 ( .B1(n4396), .B2(n3467), .A(n3463), .ZN(U3531) );
  INV_X1 U4030 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3465) );
  MUX2_X1 U4031 ( .A(n3465), .B(n3464), .S(n4849), .Z(n3466) );
  OAI21_X1 U4032 ( .B1(n3467), .B2(n4442), .A(n3466), .ZN(U3493) );
  XNOR2_X1 U4033 ( .A(n3468), .B(n3475), .ZN(n3473) );
  NAND2_X1 U4034 ( .A1(n4107), .A2(n2263), .ZN(n3470) );
  NAND2_X1 U4035 ( .A1(n4108), .A2(n2260), .ZN(n3469) );
  OAI211_X1 U4036 ( .C1(n4819), .C2(n3471), .A(n3470), .B(n3469), .ZN(n3472)
         );
  AOI21_X1 U4037 ( .B1(n3473), .B2(n4821), .A(n3472), .ZN(n4409) );
  OAI21_X1 U4038 ( .B1(n3476), .B2(n3475), .A(n3474), .ZN(n4410) );
  OR2_X1 U4039 ( .A1(n4410), .A2(n4353), .ZN(n3482) );
  NAND2_X1 U4040 ( .A1(n3492), .A2(n4034), .ZN(n4405) );
  AND2_X1 U4041 ( .A1(n4405), .A2(n4908), .ZN(n3480) );
  INV_X1 U4042 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3478) );
  INV_X1 U40430 ( .A(n3477), .ZN(n4037) );
  OAI22_X1 U4044 ( .A1(n4328), .A2(n3478), .B1(n4037), .B2(n4875), .ZN(n3479)
         );
  AOI21_X1 U4045 ( .B1(n3480), .B2(n4407), .A(n3479), .ZN(n3481) );
  OAI211_X1 U4046 ( .C1(n4858), .C2(n4409), .A(n3482), .B(n3481), .ZN(U3274)
         );
  NAND2_X1 U4047 ( .A1(n3484), .A2(n3483), .ZN(n3485) );
  XNOR2_X1 U4048 ( .A(n3485), .B(n3687), .ZN(n3548) );
  INV_X1 U4049 ( .A(n3548), .ZN(n3499) );
  NAND2_X1 U4050 ( .A1(n3486), .A2(n3593), .ZN(n3487) );
  XNOR2_X1 U4051 ( .A(n3487), .B(n3687), .ZN(n3490) );
  AOI22_X1 U4052 ( .A1(n4886), .A2(n2260), .B1(n4359), .B2(n4894), .ZN(n3489)
         );
  NAND2_X1 U4053 ( .A1(n4885), .A2(n2263), .ZN(n3488) );
  OAI211_X1 U4054 ( .C1(n3490), .C2(n4344), .A(n3489), .B(n3488), .ZN(n3547)
         );
  INV_X1 U4055 ( .A(n3491), .ZN(n3494) );
  OAI21_X1 U4056 ( .B1(n3494), .B2(n3493), .A(n3492), .ZN(n3553) );
  AOI22_X1 U4057 ( .A1(n4858), .A2(REG2_REG_15__SCAN_IN), .B1(n3495), .B2(
        n4859), .ZN(n3496) );
  OAI21_X1 U4058 ( .B1(n3553), .B2(n4871), .A(n3496), .ZN(n3497) );
  AOI21_X1 U4059 ( .B1(n3547), .B2(n4328), .A(n3497), .ZN(n3498) );
  OAI21_X1 U4060 ( .B1(n3499), .B2(n4353), .A(n3498), .ZN(U3275) );
  NAND2_X1 U4061 ( .A1(n4109), .A2(n3899), .ZN(n3504) );
  NAND2_X1 U4062 ( .A1(n3509), .A2(n3946), .ZN(n3503) );
  NAND2_X1 U4063 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  XNOR2_X1 U4064 ( .A(n3505), .B(n3031), .ZN(n3507) );
  AOI22_X1 U4065 ( .A1(n4109), .A2(n3947), .B1(n3899), .B2(n3509), .ZN(n3506)
         );
  NAND2_X1 U4066 ( .A1(n3507), .A2(n3506), .ZN(n3524) );
  NAND2_X1 U4067 ( .A1(n2288), .A2(n3524), .ZN(n3508) );
  XNOR2_X1 U4068 ( .A(n3525), .B(n3508), .ZN(n3514) );
  AOI22_X1 U4069 ( .A1(n4089), .A2(n4886), .B1(n4090), .B2(n4110), .ZN(n3511)
         );
  INV_X1 U4070 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4548) );
  NOR2_X1 U4071 ( .A1(STATE_REG_SCAN_IN), .A2(n4548), .ZN(n4736) );
  AOI21_X1 U4072 ( .B1(n4092), .B2(n3509), .A(n4736), .ZN(n3510) );
  OAI211_X1 U4073 ( .C1(n4903), .C2(n3512), .A(n3511), .B(n3510), .ZN(n3513)
         );
  AOI21_X1 U4074 ( .B1(n3514), .B2(n4898), .A(n3513), .ZN(n3515) );
  INV_X1 U4075 ( .A(n3515), .ZN(U3231) );
  AOI21_X1 U4076 ( .B1(n3517), .B2(n4840), .A(n3516), .ZN(n3521) );
  INV_X1 U4077 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3518) );
  MUX2_X1 U4078 ( .A(n3521), .B(n3518), .S(n4414), .Z(n3519) );
  OAI21_X1 U4079 ( .B1(n3523), .B2(n4442), .A(n3519), .ZN(U3495) );
  INV_X1 U4080 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3520) );
  MUX2_X1 U4081 ( .A(n3521), .B(n3520), .S(n4844), .Z(n3522) );
  OAI21_X1 U4082 ( .B1(n4396), .B2(n3523), .A(n3522), .ZN(U3532) );
  AOI22_X1 U4083 ( .A1(n4886), .A2(n3947), .B1(n3899), .B2(n3528), .ZN(n3741)
         );
  AOI22_X1 U4084 ( .A1(n4886), .A2(n3899), .B1(n3946), .B2(n3528), .ZN(n3526)
         );
  XNOR2_X1 U4085 ( .A(n3526), .B(n3948), .ZN(n3739) );
  XOR2_X1 U4086 ( .A(n3741), .B(n3739), .Z(n3527) );
  XNOR2_X1 U4087 ( .A(n3742), .B(n3527), .ZN(n3533) );
  AOI22_X1 U4088 ( .A1(n4089), .A2(n4108), .B1(n4090), .B2(n4109), .ZN(n3530)
         );
  AND2_X1 U4089 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4166) );
  AOI21_X1 U4090 ( .B1(n4092), .B2(n3528), .A(n4166), .ZN(n3529) );
  OAI211_X1 U4091 ( .C1(n4903), .C2(n3531), .A(n3530), .B(n3529), .ZN(n3532)
         );
  AOI21_X1 U4092 ( .B1(n3533), .B2(n4898), .A(n3532), .ZN(n3534) );
  INV_X1 U4093 ( .A(n3534), .ZN(U3212) );
  NAND2_X1 U4094 ( .A1(n3558), .A2(n3557), .ZN(n3672) );
  XOR2_X1 U4095 ( .A(n3672), .B(n3535), .Z(n3575) );
  INV_X1 U4096 ( .A(n3575), .ZN(n3546) );
  INV_X1 U4097 ( .A(n4106), .ZN(n3996) );
  XNOR2_X1 U4098 ( .A(n3836), .B(n3672), .ZN(n3536) );
  NAND2_X1 U4099 ( .A1(n3536), .A2(n4821), .ZN(n3538) );
  AOI22_X1 U4100 ( .A1(n4885), .A2(n2260), .B1(n3769), .B2(n4359), .ZN(n3537)
         );
  OAI211_X1 U4101 ( .C1(n3996), .C2(n3778), .A(n3538), .B(n3537), .ZN(n3574)
         );
  INV_X1 U4102 ( .A(n4407), .ZN(n3541) );
  INV_X1 U4103 ( .A(n3777), .ZN(n3539) );
  OAI21_X1 U4104 ( .B1(n3541), .B2(n3540), .A(n3539), .ZN(n3581) );
  NOR2_X1 U4105 ( .A1(n3581), .A2(n4871), .ZN(n3544) );
  INV_X1 U4106 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3542) );
  OAI22_X1 U4107 ( .A1(n4328), .A2(n3542), .B1(n3772), .B2(n4875), .ZN(n3543)
         );
  AOI211_X1 U4108 ( .C1(n3574), .C2(n4328), .A(n3544), .B(n3543), .ZN(n3545)
         );
  OAI21_X1 U4109 ( .B1(n3546), .B2(n4353), .A(n3545), .ZN(U3273) );
  AOI21_X1 U4110 ( .B1(n3548), .B2(n4840), .A(n3547), .ZN(n3551) );
  INV_X1 U4111 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3549) );
  MUX2_X1 U4112 ( .A(n3551), .B(n3549), .S(n4414), .Z(n3550) );
  OAI21_X1 U4113 ( .B1(n3553), .B2(n4442), .A(n3550), .ZN(U3497) );
  INV_X1 U4114 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4171) );
  MUX2_X1 U4115 ( .A(n3551), .B(n4171), .S(n4844), .Z(n3552) );
  OAI21_X1 U4116 ( .B1(n4396), .B2(n3553), .A(n3552), .ZN(U3533) );
  NAND2_X1 U4117 ( .A1(n3555), .A2(n3554), .ZN(n3665) );
  XNOR2_X1 U4118 ( .A(n3556), .B(n3665), .ZN(n3794) );
  INV_X1 U4119 ( .A(n3794), .ZN(n3573) );
  INV_X1 U4120 ( .A(n3557), .ZN(n3559) );
  OAI21_X1 U4121 ( .B1(n3836), .B2(n3559), .A(n3558), .ZN(n3780) );
  INV_X1 U4122 ( .A(n3560), .ZN(n3562) );
  OAI21_X1 U4123 ( .B1(n3780), .B2(n3562), .A(n3561), .ZN(n3563) );
  XOR2_X1 U4124 ( .A(n3665), .B(n3563), .Z(n3566) );
  AOI22_X1 U4125 ( .A1(n4104), .A2(n2263), .B1(n4359), .B2(n3998), .ZN(n3565)
         );
  NAND2_X1 U4126 ( .A1(n4106), .A2(n2260), .ZN(n3564) );
  OAI211_X1 U4127 ( .C1(n3566), .C2(n4344), .A(n3565), .B(n3564), .ZN(n3793)
         );
  INV_X1 U4128 ( .A(n3776), .ZN(n3567) );
  OAI21_X1 U4129 ( .B1(n3567), .B2(n3881), .A(n2284), .ZN(n3800) );
  NOR2_X1 U4130 ( .A1(n3800), .A2(n4871), .ZN(n3571) );
  INV_X1 U4131 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3569) );
  OAI22_X1 U4132 ( .A1(n4328), .A2(n3569), .B1(n3568), .B2(n4875), .ZN(n3570)
         );
  AOI211_X1 U4133 ( .C1(n3793), .C2(n4328), .A(n3571), .B(n3570), .ZN(n3572)
         );
  OAI21_X1 U4134 ( .B1(n3573), .B2(n4353), .A(n3572), .ZN(U3271) );
  INV_X1 U4135 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3576) );
  AOI21_X1 U4136 ( .B1(n3575), .B2(n4840), .A(n3574), .ZN(n3578) );
  MUX2_X1 U4137 ( .A(n3576), .B(n3578), .S(n4846), .Z(n3577) );
  OAI21_X1 U4138 ( .B1(n4396), .B2(n3581), .A(n3577), .ZN(U3535) );
  INV_X1 U4139 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3579) );
  MUX2_X1 U4140 ( .A(n3579), .B(n3578), .S(n4849), .Z(n3580) );
  OAI21_X1 U4141 ( .B1(n3581), .B2(n4442), .A(n3580), .ZN(U3501) );
  INV_X1 U4142 ( .A(n3708), .ZN(n3632) );
  NAND2_X1 U4143 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  OR2_X1 U4144 ( .A1(n3619), .A2(n3584), .ZN(n3616) );
  INV_X1 U4145 ( .A(n3616), .ZN(n3587) );
  INV_X1 U4146 ( .A(n3585), .ZN(n3586) );
  NAND3_X1 U4147 ( .A1(n3587), .A2(n3586), .A3(n3613), .ZN(n3591) );
  AND2_X1 U4148 ( .A1(n3589), .A2(n3588), .ZN(n3623) );
  INV_X1 U4149 ( .A(n3623), .ZN(n3590) );
  AOI21_X1 U4150 ( .B1(n3592), .B2(n3591), .A(n3590), .ZN(n3596) );
  NAND2_X1 U4151 ( .A1(n3593), .A2(n3599), .ZN(n3705) );
  INV_X1 U4152 ( .A(n3594), .ZN(n3595) );
  NOR3_X1 U4153 ( .A1(n3596), .A2(n3705), .A3(n3595), .ZN(n3629) );
  NAND2_X1 U4154 ( .A1(n3598), .A2(n3597), .ZN(n3622) );
  NAND2_X1 U4155 ( .A1(n3622), .A2(n3599), .ZN(n3703) );
  INV_X1 U4156 ( .A(n3703), .ZN(n3628) );
  OAI211_X1 U4157 ( .C1(n3602), .C2(n3726), .A(n3601), .B(n3600), .ZN(n3605)
         );
  NAND3_X1 U4158 ( .A1(n3605), .A2(n3604), .A3(n3603), .ZN(n3608) );
  NAND3_X1 U4159 ( .A1(n3608), .A2(n3607), .A3(n3606), .ZN(n3611) );
  NAND3_X1 U4160 ( .A1(n3611), .A2(n3610), .A3(n3609), .ZN(n3615) );
  NAND4_X1 U4161 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3618)
         );
  AOI21_X1 U4162 ( .B1(n3618), .B2(n3617), .A(n3616), .ZN(n3626) );
  AOI21_X1 U4163 ( .B1(n3621), .B2(n3620), .A(n3619), .ZN(n3625) );
  INV_X1 U4164 ( .A(n3622), .ZN(n3624) );
  OAI211_X1 U4165 ( .C1(n3626), .C2(n3625), .A(n3624), .B(n3623), .ZN(n3627)
         );
  OAI21_X1 U4166 ( .B1(n3629), .B2(n3628), .A(n3627), .ZN(n3631) );
  OAI211_X1 U4167 ( .C1(n3632), .C2(n3631), .A(n3704), .B(n3630), .ZN(n3633)
         );
  OAI221_X1 U4168 ( .B1(n3818), .B2(n3710), .C1(n3818), .C2(n3633), .A(n3715), 
        .ZN(n3634) );
  AOI21_X1 U4169 ( .B1(n3635), .B2(n3634), .A(n3717), .ZN(n3653) );
  INV_X1 U4170 ( .A(n3716), .ZN(n3651) );
  INV_X1 U4171 ( .A(n3636), .ZN(n3637) );
  AOI21_X1 U4172 ( .B1(n4244), .B2(n3658), .A(n3637), .ZN(n3699) );
  INV_X1 U4173 ( .A(DATAI_30_), .ZN(n3638) );
  NOR2_X1 U4174 ( .A1(n3639), .A2(n3638), .ZN(n4360) );
  OR2_X1 U4175 ( .A1(n3655), .A2(n4360), .ZN(n3648) );
  NAND2_X1 U4176 ( .A1(n3640), .A2(REG1_REG_31__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4177 ( .A1(n3641), .A2(REG2_REG_31__SCAN_IN), .ZN(n3644) );
  NAND2_X1 U4178 ( .A1(n3642), .A2(REG0_REG_31__SCAN_IN), .ZN(n3643) );
  NAND3_X1 U4179 ( .A1(n3645), .A2(n3644), .A3(n3643), .ZN(n4099) );
  NAND2_X1 U4180 ( .A1(n3646), .A2(DATAI_31_), .ZN(n4222) );
  OR2_X1 U4181 ( .A1(n4099), .A2(n4222), .ZN(n3647) );
  AND2_X1 U4182 ( .A1(n3648), .A2(n3647), .ZN(n3654) );
  NAND4_X1 U4183 ( .A1(n3699), .A2(n3654), .A3(n3649), .A4(n3698), .ZN(n3650)
         );
  AOI221_X1 U4184 ( .B1(n3653), .B2(n3652), .C1(n3651), .C2(n3652), .A(n3650), 
        .ZN(n3661) );
  INV_X1 U4185 ( .A(n3654), .ZN(n3725) );
  NAND2_X1 U4186 ( .A1(n4099), .A2(n4222), .ZN(n3659) );
  INV_X1 U4187 ( .A(n3655), .ZN(n4100) );
  INV_X1 U4188 ( .A(n4360), .ZN(n3656) );
  OAI21_X1 U4189 ( .B1(n4100), .B2(n3656), .A(n3659), .ZN(n3667) );
  INV_X1 U4190 ( .A(n3667), .ZN(n3657) );
  OAI21_X1 U4191 ( .B1(n4244), .B2(n3658), .A(n3657), .ZN(n3700) );
  AOI21_X1 U4192 ( .B1(n3699), .B2(n3702), .A(n3700), .ZN(n3722) );
  AOI21_X1 U4193 ( .B1(n3725), .B2(n3659), .A(n3722), .ZN(n3660) );
  OR2_X1 U4194 ( .A1(n3661), .A2(n3660), .ZN(n3730) );
  AND2_X1 U4195 ( .A1(n4310), .A2(n3662), .ZN(n4338) );
  XNOR2_X1 U4196 ( .A(n4342), .B(n4315), .ZN(n4312) );
  NAND4_X1 U4197 ( .A1(n4338), .A2(n4312), .A3(n3664), .A4(n3663), .ZN(n3666)
         );
  NOR4_X1 U4198 ( .A1(n3725), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3682)
         );
  INV_X1 U4199 ( .A(n3668), .ZN(n3673) );
  NAND2_X1 U4200 ( .A1(n3670), .A2(n3669), .ZN(n3840) );
  NAND2_X1 U4201 ( .A1(n4273), .A2(n3671), .ZN(n4293) );
  NOR4_X1 U4202 ( .A1(n3673), .A2(n3840), .A3(n3672), .A4(n4293), .ZN(n3681)
         );
  NOR4_X1 U4203 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3680)
         );
  NOR4_X1 U4204 ( .A1(n2620), .A2(n3779), .A3(n4241), .A4(n3678), .ZN(n3679)
         );
  NAND4_X1 U4205 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n3697)
         );
  NOR4_X1 U4206 ( .A1(n3686), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(n3690)
         );
  NOR4_X1 U4207 ( .A1(n3688), .A2(n4335), .A3(n3687), .A4(n4769), .ZN(n3689)
         );
  NAND2_X1 U4208 ( .A1(n3690), .A2(n3689), .ZN(n3696) );
  NAND2_X1 U4209 ( .A1(n3698), .A2(n3691), .ZN(n4271) );
  INV_X1 U4210 ( .A(n4271), .ZN(n4276) );
  INV_X1 U4211 ( .A(n3692), .ZN(n3819) );
  NOR2_X1 U4212 ( .A1(n3819), .A2(n3818), .ZN(n3801) );
  NAND4_X1 U4213 ( .A1(n4261), .A2(n3693), .A3(n4276), .A4(n3801), .ZN(n3694)
         );
  NOR4_X1 U4214 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3728)
         );
  INV_X1 U4215 ( .A(n4222), .ZN(n4225) );
  INV_X1 U4216 ( .A(n4099), .ZN(n4224) );
  NAND3_X1 U4217 ( .A1(n4261), .A2(n3699), .A3(n3698), .ZN(n3721) );
  NOR3_X1 U4218 ( .A1(n3702), .A2(n3701), .A3(n3700), .ZN(n3720) );
  OAI211_X1 U4219 ( .C1(n3706), .C2(n3705), .A(n3704), .B(n3703), .ZN(n3709)
         );
  AOI21_X1 U4220 ( .B1(n3709), .B2(n3708), .A(n3707), .ZN(n3712) );
  INV_X1 U4221 ( .A(n3710), .ZN(n3711) );
  NOR2_X1 U4222 ( .A1(n3712), .A2(n3711), .ZN(n3714) );
  AOI21_X1 U4223 ( .B1(n3715), .B2(n3714), .A(n3713), .ZN(n3718) );
  OAI21_X1 U4224 ( .B1(n3718), .B2(n3717), .A(n3716), .ZN(n3719) );
  AOI22_X1 U4225 ( .A1(n3722), .A2(n3721), .B1(n3720), .B2(n3719), .ZN(n3723)
         );
  AOI21_X1 U4226 ( .B1(n4360), .B2(n4224), .A(n3723), .ZN(n3724) );
  AOI21_X1 U4227 ( .B1(n4225), .B2(n3725), .A(n3724), .ZN(n3727) );
  MUX2_X1 U4228 ( .A(n3728), .B(n3727), .S(n3726), .Z(n3729) );
  MUX2_X1 U4229 ( .A(n3730), .B(n3729), .S(n4449), .Z(n3731) );
  XNOR2_X1 U4230 ( .A(n3731), .B(n4450), .ZN(n3738) );
  NOR4_X1 U4231 ( .A1(n4907), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3735)
         );
  NAND2_X1 U4232 ( .A1(n3735), .A2(n3899), .ZN(n3736) );
  OAI211_X1 U4233 ( .C1(n4448), .C2(n4455), .A(n3736), .B(B_REG_SCAN_IN), .ZN(
        n3737) );
  OAI21_X1 U4234 ( .B1(n3738), .B2(n4455), .A(n3737), .ZN(U3239) );
  AOI21_X1 U4235 ( .B1(n3742), .B2(n3741), .A(n3739), .ZN(n3740) );
  INV_X1 U4236 ( .A(n3740), .ZN(n3743) );
  NAND2_X1 U4237 ( .A1(n4108), .A2(n3899), .ZN(n3745) );
  NAND2_X1 U4238 ( .A1(n4894), .A2(n3946), .ZN(n3744) );
  NAND2_X1 U4239 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  XNOR2_X1 U4240 ( .A(n3746), .B(n3031), .ZN(n4896) );
  NAND2_X1 U4241 ( .A1(n4108), .A2(n3947), .ZN(n3748) );
  NAND2_X1 U4242 ( .A1(n4894), .A2(n3899), .ZN(n3747) );
  AND2_X1 U4243 ( .A1(n3748), .A2(n3747), .ZN(n4895) );
  NAND2_X1 U4244 ( .A1(n4885), .A2(n3899), .ZN(n3750) );
  NAND2_X1 U4245 ( .A1(n4034), .A2(n3946), .ZN(n3749) );
  NAND2_X1 U4246 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  XNOR2_X1 U4247 ( .A(n3751), .B(n3948), .ZN(n3754) );
  NAND2_X1 U4248 ( .A1(n4885), .A2(n3947), .ZN(n3753) );
  NAND2_X1 U4249 ( .A1(n4034), .A2(n3899), .ZN(n3752) );
  NAND2_X1 U4250 ( .A1(n3753), .A2(n3752), .ZN(n3755) );
  NAND2_X1 U4251 ( .A1(n3754), .A2(n3755), .ZN(n4031) );
  OAI21_X1 U4252 ( .B1(n4896), .B2(n4895), .A(n4031), .ZN(n3760) );
  NAND3_X1 U4253 ( .A1(n4031), .A2(n4895), .A3(n4896), .ZN(n3758) );
  INV_X1 U4254 ( .A(n3754), .ZN(n3757) );
  INV_X1 U4255 ( .A(n3755), .ZN(n3756) );
  NAND2_X1 U4256 ( .A1(n3757), .A2(n3756), .ZN(n4030) );
  NAND2_X1 U4257 ( .A1(n4107), .A2(n3899), .ZN(n3762) );
  NAND2_X1 U4258 ( .A1(n3769), .A2(n3946), .ZN(n3761) );
  NAND2_X1 U4259 ( .A1(n3762), .A2(n3761), .ZN(n3763) );
  XNOR2_X1 U4260 ( .A(n3763), .B(n3948), .ZN(n3767) );
  NAND2_X1 U4261 ( .A1(n4107), .A2(n3947), .ZN(n3765) );
  NAND2_X1 U4262 ( .A1(n3769), .A2(n3899), .ZN(n3764) );
  NAND2_X1 U4263 ( .A1(n3765), .A2(n3764), .ZN(n3766) );
  NOR2_X1 U4264 ( .A1(n3767), .A2(n3766), .ZN(n3866) );
  NAND2_X1 U4265 ( .A1(n3767), .A2(n3766), .ZN(n3867) );
  NOR2_X1 U4266 ( .A1(n3866), .A2(n2363), .ZN(n3768) );
  XNOR2_X1 U4267 ( .A(n3868), .B(n3768), .ZN(n3774) );
  AOI22_X1 U4268 ( .A1(n4090), .A2(n4885), .B1(n4089), .B2(n4106), .ZN(n3771)
         );
  INV_X1 U4269 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4626) );
  NOR2_X1 U4270 ( .A1(STATE_REG_SCAN_IN), .A2(n4626), .ZN(n4202) );
  AOI21_X1 U4271 ( .B1(n4893), .B2(n3769), .A(n4202), .ZN(n3770) );
  OAI211_X1 U4272 ( .C1(n4903), .C2(n3772), .A(n3771), .B(n3770), .ZN(n3773)
         );
  AOI21_X1 U4273 ( .B1(n3774), .B2(n4898), .A(n3773), .ZN(n3775) );
  INV_X1 U4274 ( .A(n3775), .ZN(U3225) );
  OAI211_X1 U4275 ( .C1(n3777), .C2(n3872), .A(n3776), .B(n4406), .ZN(n4402)
         );
  INV_X1 U4276 ( .A(n4105), .ZN(n3839) );
  OAI22_X1 U4277 ( .A1(n3839), .A2(n3778), .B1(n3872), .B2(n4819), .ZN(n3783)
         );
  XNOR2_X1 U4278 ( .A(n3780), .B(n3779), .ZN(n3781) );
  NOR2_X1 U4279 ( .A1(n3781), .A2(n4344), .ZN(n3782) );
  AOI211_X1 U4280 ( .C1(n2260), .C2(n4107), .A(n3783), .B(n3782), .ZN(n4403)
         );
  OAI21_X1 U4281 ( .B1(n4450), .B2(n4402), .A(n4403), .ZN(n3791) );
  INV_X1 U4282 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4208) );
  INV_X1 U4283 ( .A(n3784), .ZN(n4080) );
  OAI22_X1 U4284 ( .A1(n4328), .A2(n4208), .B1(n4080), .B2(n4875), .ZN(n3790)
         );
  INV_X1 U4285 ( .A(n3785), .ZN(n3786) );
  AOI21_X1 U4286 ( .B1(n3788), .B2(n3787), .A(n3786), .ZN(n4404) );
  NOR2_X1 U4287 ( .A1(n4404), .A2(n4353), .ZN(n3789) );
  AOI211_X1 U4288 ( .C1(n4328), .C2(n3791), .A(n3790), .B(n3789), .ZN(n3792)
         );
  INV_X1 U4289 ( .A(n3792), .ZN(U3272) );
  INV_X1 U4290 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3795) );
  AOI21_X1 U4291 ( .B1(n3794), .B2(n4840), .A(n3793), .ZN(n3797) );
  MUX2_X1 U4292 ( .A(n3795), .B(n3797), .S(n4411), .Z(n3796) );
  OAI21_X1 U4293 ( .B1(n4396), .B2(n3800), .A(n3796), .ZN(U3537) );
  INV_X1 U4294 ( .A(REG0_REG_19__SCAN_IN), .ZN(n3798) );
  MUX2_X1 U4295 ( .A(n3798), .B(n3797), .S(n4849), .Z(n3799) );
  OAI21_X1 U4296 ( .B1(n3800), .B2(n4442), .A(n3799), .ZN(U3505) );
  XOR2_X1 U4297 ( .A(n3801), .B(n3815), .Z(n4393) );
  INV_X1 U4298 ( .A(n4393), .ZN(n3812) );
  XNOR2_X1 U4299 ( .A(n3821), .B(n3801), .ZN(n3802) );
  NAND2_X1 U4300 ( .A1(n3802), .A2(n4821), .ZN(n3804) );
  AOI22_X1 U4301 ( .A1(n4102), .A2(n2263), .B1(n4359), .B2(n4010), .ZN(n3803)
         );
  OAI211_X1 U4302 ( .C1(n3995), .C2(n4339), .A(n3804), .B(n3803), .ZN(n4392)
         );
  INV_X1 U4303 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3806) );
  INV_X1 U4304 ( .A(n3805), .ZN(n4013) );
  OAI22_X1 U4305 ( .A1(n4328), .A2(n3806), .B1(n4013), .B2(n4875), .ZN(n3810)
         );
  INV_X1 U4306 ( .A(n3827), .ZN(n3807) );
  OAI21_X1 U4307 ( .B1(n3846), .B2(n3808), .A(n3807), .ZN(n4443) );
  NOR2_X1 U4308 ( .A1(n4443), .A2(n4871), .ZN(n3809) );
  AOI211_X1 U4309 ( .C1(n4392), .C2(n4328), .A(n3810), .B(n3809), .ZN(n3811)
         );
  OAI21_X1 U4310 ( .B1(n3812), .B2(n4353), .A(n3811), .ZN(U3269) );
  OAI21_X1 U4311 ( .B1(n3815), .B2(n3814), .A(n3813), .ZN(n3817) );
  AND2_X1 U4312 ( .A1(n3817), .A2(n4335), .ZN(n4332) );
  INV_X1 U4313 ( .A(n4332), .ZN(n3816) );
  OAI21_X1 U4314 ( .B1(n3817), .B2(n4335), .A(n3816), .ZN(n4391) );
  INV_X1 U4315 ( .A(n3818), .ZN(n3820) );
  AOI21_X1 U4316 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n4336) );
  XNOR2_X1 U4317 ( .A(n4336), .B(n4335), .ZN(n3825) );
  NAND2_X1 U4318 ( .A1(n4101), .A2(n2263), .ZN(n3823) );
  NAND2_X1 U4319 ( .A1(n4103), .A2(n2260), .ZN(n3822) );
  OAI211_X1 U4320 ( .C1(n4819), .C2(n4064), .A(n3823), .B(n3822), .ZN(n3824)
         );
  AOI21_X1 U4321 ( .B1(n3825), .B2(n4821), .A(n3824), .ZN(n4390) );
  INV_X1 U4322 ( .A(n4390), .ZN(n3831) );
  INV_X1 U4323 ( .A(n3826), .ZN(n4068) );
  OR2_X1 U4324 ( .A1(n3827), .A2(n4064), .ZN(n4388) );
  NAND3_X1 U4325 ( .A1(n4388), .A2(n4387), .A3(n4908), .ZN(n3829) );
  NAND2_X1 U4326 ( .A1(n4858), .A2(REG2_REG_22__SCAN_IN), .ZN(n3828) );
  OAI211_X1 U4327 ( .C1(n4875), .C2(n4068), .A(n3829), .B(n3828), .ZN(n3830)
         );
  AOI21_X1 U4328 ( .B1(n3831), .B2(n4328), .A(n3830), .ZN(n3832) );
  OAI21_X1 U4329 ( .B1(n4391), .B2(n4353), .A(n3832), .ZN(U3268) );
  INV_X1 U4330 ( .A(n3833), .ZN(n3835) );
  OAI21_X1 U4331 ( .B1(n3836), .B2(n3835), .A(n3834), .ZN(n3837) );
  XOR2_X1 U4332 ( .A(n3840), .B(n3837), .Z(n3845) );
  AOI22_X1 U4333 ( .A1(n4103), .A2(n2263), .B1(n4053), .B2(n4359), .ZN(n3838)
         );
  OAI21_X1 U4334 ( .B1(n3839), .B2(n4339), .A(n3838), .ZN(n3844) );
  XNOR2_X1 U4335 ( .A(n3841), .B(n3840), .ZN(n4401) );
  NOR2_X1 U4336 ( .A1(n4401), .A2(n3842), .ZN(n3843) );
  AOI211_X1 U4337 ( .C1(n3845), .C2(n4821), .A(n3844), .B(n3843), .ZN(n4400)
         );
  INV_X1 U4338 ( .A(n4401), .ZN(n3851) );
  INV_X1 U4339 ( .A(n3846), .ZN(n4398) );
  NAND2_X1 U4340 ( .A1(n2284), .A2(n4053), .ZN(n4397) );
  AND3_X1 U4341 ( .A1(n4398), .A2(n4908), .A3(n4397), .ZN(n3850) );
  INV_X1 U4342 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3848) );
  INV_X1 U4343 ( .A(n3847), .ZN(n4056) );
  OAI22_X1 U4344 ( .A1(n4328), .A2(n3848), .B1(n4056), .B2(n4875), .ZN(n3849)
         );
  AOI211_X1 U4345 ( .C1(n3851), .C2(n4869), .A(n3850), .B(n3849), .ZN(n3852)
         );
  OAI21_X1 U4346 ( .B1(n4400), .B2(n4858), .A(n3852), .ZN(U3270) );
  OR2_X1 U4347 ( .A1(n3854), .A2(n3853), .ZN(n3856) );
  AOI211_X1 U4348 ( .C1(n3857), .C2(n3856), .A(n4097), .B(n3855), .ZN(n3865)
         );
  INV_X1 U4349 ( .A(n3858), .ZN(n3863) );
  AOI22_X1 U4350 ( .A1(n4090), .A2(n3050), .B1(n4089), .B2(n4115), .ZN(n3862)
         );
  AOI21_X1 U4351 ( .B1(n4893), .B2(n3860), .A(n3859), .ZN(n3861) );
  OAI211_X1 U4352 ( .C1(n4903), .C2(n3863), .A(n3862), .B(n3861), .ZN(n3864)
         );
  OR2_X1 U4353 ( .A1(n3865), .A2(n3864), .ZN(U3227) );
  NAND2_X1 U4354 ( .A1(n4106), .A2(n3899), .ZN(n3870) );
  NAND2_X1 U4355 ( .A1(n4077), .A2(n3946), .ZN(n3869) );
  NAND2_X1 U4356 ( .A1(n3870), .A2(n3869), .ZN(n3871) );
  XNOR2_X1 U4357 ( .A(n3871), .B(n3031), .ZN(n4074) );
  NOR2_X1 U4358 ( .A1(n3872), .A2(n3433), .ZN(n3873) );
  AOI21_X1 U4359 ( .B1(n4106), .B2(n3947), .A(n3873), .ZN(n4073) );
  INV_X1 U4360 ( .A(n4074), .ZN(n3875) );
  INV_X1 U4361 ( .A(n4073), .ZN(n3874) );
  NAND2_X1 U4362 ( .A1(n3875), .A2(n3874), .ZN(n3876) );
  NAND2_X1 U4363 ( .A1(n3877), .A2(n3876), .ZN(n3991) );
  INV_X1 U4364 ( .A(n3991), .ZN(n3886) );
  NAND2_X1 U4365 ( .A1(n4105), .A2(n3899), .ZN(n3879) );
  NAND2_X1 U4366 ( .A1(n3998), .A2(n3946), .ZN(n3878) );
  NAND2_X1 U4367 ( .A1(n3879), .A2(n3878), .ZN(n3880) );
  XNOR2_X1 U4368 ( .A(n3880), .B(n3031), .ZN(n3884) );
  NOR2_X1 U4369 ( .A1(n3881), .A2(n3433), .ZN(n3882) );
  AOI21_X1 U4370 ( .B1(n4105), .B2(n3947), .A(n3882), .ZN(n3883) );
  NAND2_X1 U4371 ( .A1(n3884), .A2(n3883), .ZN(n3887) );
  OAI21_X1 U4372 ( .B1(n3884), .B2(n3883), .A(n3887), .ZN(n3994) );
  NAND2_X1 U4373 ( .A1(n3886), .A2(n3885), .ZN(n3992) );
  NAND2_X1 U4374 ( .A1(n4104), .A2(n3899), .ZN(n3889) );
  NAND2_X1 U4375 ( .A1(n4053), .A2(n3946), .ZN(n3888) );
  NAND2_X1 U4376 ( .A1(n3889), .A2(n3888), .ZN(n3890) );
  XNOR2_X1 U4377 ( .A(n3890), .B(n3031), .ZN(n3903) );
  INV_X1 U4378 ( .A(n3903), .ZN(n3895) );
  NOR2_X1 U4379 ( .A1(n3433), .A2(n3892), .ZN(n3893) );
  AOI21_X1 U4380 ( .B1(n4104), .B2(n3947), .A(n3893), .ZN(n3902) );
  INV_X1 U4381 ( .A(n3902), .ZN(n3894) );
  NAND2_X1 U4382 ( .A1(n3895), .A2(n3894), .ZN(n4051) );
  NAND2_X1 U4383 ( .A1(n4103), .A2(n3899), .ZN(n3897) );
  NAND2_X1 U4384 ( .A1(n4010), .A2(n3946), .ZN(n3896) );
  NAND2_X1 U4385 ( .A1(n3897), .A2(n3896), .ZN(n3898) );
  XNOR2_X1 U4386 ( .A(n3898), .B(n3948), .ZN(n4007) );
  NAND2_X1 U4387 ( .A1(n4103), .A2(n3947), .ZN(n3901) );
  NAND2_X1 U4388 ( .A1(n4010), .A2(n3899), .ZN(n3900) );
  NAND2_X1 U4389 ( .A1(n3901), .A2(n3900), .ZN(n4006) );
  NAND2_X1 U4390 ( .A1(n3903), .A2(n3902), .ZN(n4050) );
  OAI21_X1 U4391 ( .B1(n4007), .B2(n4006), .A(n4050), .ZN(n3904) );
  AOI21_X1 U4392 ( .B1(n4004), .B2(n4051), .A(n3904), .ZN(n3908) );
  INV_X1 U4393 ( .A(n4007), .ZN(n3906) );
  INV_X1 U4394 ( .A(n4006), .ZN(n3905) );
  NOR2_X1 U4395 ( .A1(n3906), .A2(n3905), .ZN(n3907) );
  NOR2_X1 U4396 ( .A1(n3908), .A2(n3907), .ZN(n4060) );
  OAI22_X1 U4397 ( .A1(n4340), .A2(n3433), .B1(n3924), .B2(n4064), .ZN(n3909)
         );
  XNOR2_X1 U4398 ( .A(n3909), .B(n3948), .ZN(n3914) );
  OAI22_X1 U4399 ( .A1(n4340), .A2(n3926), .B1(n3433), .B2(n4064), .ZN(n3913)
         );
  XNOR2_X1 U4400 ( .A(n3914), .B(n3913), .ZN(n4063) );
  NAND2_X1 U4401 ( .A1(n4060), .A2(n3910), .ZN(n3968) );
  NOR2_X1 U4402 ( .A1(n3433), .A2(n4347), .ZN(n3911) );
  AOI21_X1 U4403 ( .B1(n4101), .B2(n3947), .A(n3911), .ZN(n3917) );
  OAI22_X1 U4404 ( .A1(n4319), .A2(n3433), .B1(n3924), .B2(n4347), .ZN(n3912)
         );
  XNOR2_X1 U4405 ( .A(n3912), .B(n3948), .ZN(n3916) );
  XOR2_X1 U4406 ( .A(n3917), .B(n3916), .Z(n3969) );
  NOR2_X1 U4407 ( .A1(n3914), .A2(n3913), .ZN(n3970) );
  NOR2_X1 U4408 ( .A1(n3969), .A2(n3970), .ZN(n3915) );
  INV_X1 U4409 ( .A(n3916), .ZN(n3918) );
  OR2_X1 U4410 ( .A1(n3918), .A2(n3917), .ZN(n3922) );
  NAND2_X1 U4411 ( .A1(n4342), .A2(n3899), .ZN(n3920) );
  NAND2_X1 U4412 ( .A1(n4315), .A2(n3946), .ZN(n3919) );
  NAND2_X1 U4413 ( .A1(n3920), .A2(n3919), .ZN(n3921) );
  XNOR2_X1 U4414 ( .A(n3921), .B(n3031), .ZN(n3923) );
  OAI22_X1 U4415 ( .A1(n4300), .A2(n3926), .B1(n3433), .B2(n4324), .ZN(n4042)
         );
  OAI22_X1 U4416 ( .A1(n3927), .A2(n3433), .B1(n3924), .B2(n4301), .ZN(n3925)
         );
  NAND2_X1 U4417 ( .A1(n3928), .A2(n4018), .ZN(n3931) );
  INV_X1 U4418 ( .A(n4017), .ZN(n3929) );
  NAND2_X1 U4419 ( .A1(n3929), .A2(n2282), .ZN(n3930) );
  NAND2_X1 U4420 ( .A1(n3931), .A2(n3930), .ZN(n4087) );
  NAND2_X1 U4421 ( .A1(n4297), .A2(n3899), .ZN(n3933) );
  NAND2_X1 U4422 ( .A1(n4091), .A2(n3946), .ZN(n3932) );
  NAND2_X1 U4423 ( .A1(n3933), .A2(n3932), .ZN(n3934) );
  XNOR2_X1 U4424 ( .A(n3934), .B(n3031), .ZN(n3937) );
  NOR2_X1 U4425 ( .A1(n3433), .A2(n4283), .ZN(n3935) );
  AOI21_X1 U4426 ( .B1(n4297), .B2(n3947), .A(n3935), .ZN(n3936) );
  NOR2_X1 U4427 ( .A1(n3937), .A2(n3936), .ZN(n4085) );
  NAND2_X1 U4428 ( .A1(n3937), .A2(n3936), .ZN(n4084) );
  NAND2_X1 U4429 ( .A1(n4278), .A2(n3899), .ZN(n3939) );
  NAND2_X1 U4430 ( .A1(n4255), .A2(n3946), .ZN(n3938) );
  NAND2_X1 U4431 ( .A1(n3939), .A2(n3938), .ZN(n3940) );
  XNOR2_X1 U4432 ( .A(n3940), .B(n3948), .ZN(n3944) );
  NAND2_X1 U4433 ( .A1(n4278), .A2(n3947), .ZN(n3942) );
  NAND2_X1 U4434 ( .A1(n4255), .A2(n3899), .ZN(n3941) );
  NAND2_X1 U4435 ( .A1(n3942), .A2(n3941), .ZN(n3943) );
  NAND2_X1 U4436 ( .A1(n3944), .A2(n3943), .ZN(n3945) );
  OAI21_X1 U4437 ( .B1(n3944), .B2(n3943), .A(n3945), .ZN(n3959) );
  AOI22_X1 U4438 ( .A1(n4256), .A2(n3899), .B1(n3946), .B2(n4243), .ZN(n3951)
         );
  AOI22_X1 U4439 ( .A1(n4256), .A2(n3947), .B1(n3899), .B2(n4243), .ZN(n3949)
         );
  XNOR2_X1 U4440 ( .A(n3949), .B(n3948), .ZN(n3950) );
  INV_X1 U4441 ( .A(n4235), .ZN(n3955) );
  AOI22_X1 U4442 ( .A1(n4089), .A2(n4244), .B1(n4090), .B2(n4278), .ZN(n3954)
         );
  AOI22_X1 U4443 ( .A1(n4893), .A2(n4243), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3953) );
  OAI211_X1 U4444 ( .C1(n4903), .C2(n3955), .A(n3954), .B(n3953), .ZN(n3956)
         );
  INV_X1 U4445 ( .A(n3956), .ZN(n3957) );
  OAI21_X1 U4446 ( .B1(n3958), .B2(n4097), .A(n3957), .ZN(U3217) );
  AOI21_X1 U4447 ( .B1(n3960), .B2(n3959), .A(n4097), .ZN(n3966) );
  INV_X1 U4448 ( .A(n4260), .ZN(n3963) );
  AOI22_X1 U4449 ( .A1(n4089), .A2(n4256), .B1(n4090), .B2(n4297), .ZN(n3962)
         );
  AOI22_X1 U4450 ( .A1(n4893), .A2(n4255), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3961) );
  OAI211_X1 U4451 ( .C1(n4903), .C2(n3963), .A(n3962), .B(n3961), .ZN(n3964)
         );
  AOI21_X1 U4452 ( .B1(n3966), .B2(n3965), .A(n3964), .ZN(n3967) );
  INV_X1 U4453 ( .A(n3967), .ZN(U3211) );
  INV_X1 U4454 ( .A(n3968), .ZN(n4061) );
  OAI21_X1 U4455 ( .B1(n4061), .B2(n3970), .A(n3969), .ZN(n3972) );
  NAND3_X1 U4456 ( .A1(n3972), .A2(n4898), .A3(n3971), .ZN(n3978) );
  AOI22_X1 U4457 ( .A1(n4893), .A2(n3973), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3977) );
  AOI22_X1 U4458 ( .A1(n4089), .A2(n4342), .B1(n4090), .B2(n4102), .ZN(n3976)
         );
  INV_X1 U4459 ( .A(n4349), .ZN(n3974) );
  OR2_X1 U4460 ( .A1(n4903), .A2(n3974), .ZN(n3975) );
  NAND4_X1 U4461 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(U3213)
         );
  AND2_X1 U4462 ( .A1(n3980), .A2(n3979), .ZN(n3983) );
  OAI211_X1 U4463 ( .C1(n3983), .C2(n3982), .A(n4898), .B(n3981), .ZN(n3990)
         );
  NOR2_X1 U4464 ( .A1(STATE_REG_SCAN_IN), .A2(n3984), .ZN(n4702) );
  AOI21_X1 U4465 ( .B1(n4092), .B2(n3985), .A(n4702), .ZN(n3989) );
  AOI22_X1 U4466 ( .A1(n4090), .A2(n4113), .B1(n4089), .B2(n4111), .ZN(n3988)
         );
  INV_X1 U4467 ( .A(n4860), .ZN(n3986) );
  OR2_X1 U4468 ( .A1(n4903), .A2(n3986), .ZN(n3987) );
  NAND4_X1 U4469 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(U3214)
         );
  INV_X1 U4470 ( .A(n3992), .ZN(n3993) );
  AOI21_X1 U4471 ( .B1(n3991), .B2(n3994), .A(n3993), .ZN(n4003) );
  INV_X1 U4472 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4610) );
  NOR2_X1 U4473 ( .A1(STATE_REG_SCAN_IN), .A2(n4610), .ZN(n4756) );
  INV_X1 U4474 ( .A(n4090), .ZN(n4888) );
  INV_X1 U4475 ( .A(n4089), .ZN(n4889) );
  OAI22_X1 U4476 ( .A1(n3996), .A2(n4888), .B1(n4889), .B2(n3995), .ZN(n3997)
         );
  AOI211_X1 U4477 ( .C1(n3998), .C2(n4893), .A(n4756), .B(n3997), .ZN(n4002)
         );
  INV_X1 U4478 ( .A(n4903), .ZN(n4000) );
  NAND2_X1 U4479 ( .A1(n4000), .A2(n3999), .ZN(n4001) );
  OAI211_X1 U4480 ( .C1(n4003), .C2(n4097), .A(n4002), .B(n4001), .ZN(U3216)
         );
  INV_X1 U4481 ( .A(n4050), .ZN(n4005) );
  OAI21_X1 U4482 ( .B1(n4004), .B2(n4005), .A(n4051), .ZN(n4009) );
  XNOR2_X1 U4483 ( .A(n4007), .B(n4006), .ZN(n4008) );
  XNOR2_X1 U4484 ( .A(n4009), .B(n4008), .ZN(n4015) );
  AOI22_X1 U4485 ( .A1(n4090), .A2(n4104), .B1(n4089), .B2(n4102), .ZN(n4012)
         );
  AOI22_X1 U4486 ( .A1(n4092), .A2(n4010), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n4011) );
  OAI211_X1 U4487 ( .C1(n4903), .C2(n4013), .A(n4012), .B(n4011), .ZN(n4014)
         );
  AOI21_X1 U4488 ( .B1(n4015), .B2(n4898), .A(n4014), .ZN(n4016) );
  INV_X1 U4489 ( .A(n4016), .ZN(U3220) );
  XNOR2_X1 U4490 ( .A(n2282), .B(n4018), .ZN(n4019) );
  XNOR2_X1 U4491 ( .A(n4017), .B(n4019), .ZN(n4025) );
  INV_X1 U4492 ( .A(n4304), .ZN(n4022) );
  AOI22_X1 U4493 ( .A1(n4090), .A2(n4342), .B1(n4089), .B2(n4297), .ZN(n4021)
         );
  AOI22_X1 U4494 ( .A1(n4893), .A2(n4296), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n4020) );
  OAI211_X1 U4495 ( .C1(n4903), .C2(n4022), .A(n4021), .B(n4020), .ZN(n4023)
         );
  INV_X1 U4496 ( .A(n4023), .ZN(n4024) );
  OAI21_X1 U4497 ( .B1(n4025), .B2(n4097), .A(n4024), .ZN(U3222) );
  INV_X1 U4498 ( .A(n4895), .ZN(n4027) );
  NOR2_X1 U4499 ( .A1(n4026), .A2(n4027), .ZN(n4029) );
  INV_X1 U4500 ( .A(n4026), .ZN(n4028) );
  OAI22_X1 U4501 ( .A1(n4029), .A2(n4896), .B1(n4028), .B2(n4895), .ZN(n4033)
         );
  NAND2_X1 U4502 ( .A1(n4031), .A2(n4030), .ZN(n4032) );
  XNOR2_X1 U4503 ( .A(n4033), .B(n4032), .ZN(n4039) );
  AOI22_X1 U4504 ( .A1(n4090), .A2(n4108), .B1(n4089), .B2(n4107), .ZN(n4036)
         );
  NOR2_X1 U4505 ( .A1(STATE_REG_SCAN_IN), .A2(n4624), .ZN(n4743) );
  AOI21_X1 U4506 ( .B1(n4893), .B2(n4034), .A(n4743), .ZN(n4035) );
  OAI211_X1 U4507 ( .C1(n4903), .C2(n4037), .A(n4036), .B(n4035), .ZN(n4038)
         );
  AOI21_X1 U4508 ( .B1(n4039), .B2(n4898), .A(n4038), .ZN(n4040) );
  INV_X1 U4509 ( .A(n4040), .ZN(U3223) );
  NOR2_X1 U4510 ( .A1(n2271), .A2(n4041), .ZN(n4043) );
  XNOR2_X1 U4511 ( .A(n4043), .B(n4042), .ZN(n4049) );
  INV_X1 U4512 ( .A(n4044), .ZN(n4320) );
  AOI22_X1 U4513 ( .A1(n4090), .A2(n4101), .B1(n4089), .B2(n4316), .ZN(n4046)
         );
  AOI22_X1 U4514 ( .A1(n4893), .A2(n4315), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n4045) );
  OAI211_X1 U4515 ( .C1(n4903), .C2(n4320), .A(n4046), .B(n4045), .ZN(n4047)
         );
  INV_X1 U4516 ( .A(n4047), .ZN(n4048) );
  OAI21_X1 U4517 ( .B1(n4049), .B2(n4097), .A(n4048), .ZN(U3226) );
  NAND2_X1 U4518 ( .A1(n4051), .A2(n4050), .ZN(n4052) );
  XOR2_X1 U4519 ( .A(n4052), .B(n4004), .Z(n4058) );
  AOI22_X1 U4520 ( .A1(n4089), .A2(n4103), .B1(n4090), .B2(n4105), .ZN(n4055)
         );
  AOI22_X1 U4521 ( .A1(n4092), .A2(n4053), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n4054) );
  OAI211_X1 U4522 ( .C1(n4903), .C2(n4056), .A(n4055), .B(n4054), .ZN(n4057)
         );
  AOI21_X1 U4523 ( .B1(n4058), .B2(n4898), .A(n4057), .ZN(n4059) );
  INV_X1 U4524 ( .A(n4059), .ZN(U3230) );
  AOI21_X1 U4525 ( .B1(n4063), .B2(n4062), .A(n4061), .ZN(n4071) );
  AOI22_X1 U4526 ( .A1(n4089), .A2(n4101), .B1(n4090), .B2(n4103), .ZN(n4067)
         );
  INV_X1 U4527 ( .A(n4064), .ZN(n4065) );
  AOI22_X1 U4528 ( .A1(n4893), .A2(n4065), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n4066) );
  OAI211_X1 U4529 ( .C1(n4903), .C2(n4068), .A(n4067), .B(n4066), .ZN(n4069)
         );
  INV_X1 U4530 ( .A(n4069), .ZN(n4070) );
  OAI21_X1 U4531 ( .B1(n4071), .B2(n4097), .A(n4070), .ZN(U3232) );
  XNOR2_X1 U4532 ( .A(n4074), .B(n4073), .ZN(n4075) );
  XNOR2_X1 U4533 ( .A(n4072), .B(n4075), .ZN(n4082) );
  AOI22_X1 U4534 ( .A1(n4090), .A2(n4107), .B1(n4089), .B2(n4105), .ZN(n4079)
         );
  NOR2_X1 U4535 ( .A1(STATE_REG_SCAN_IN), .A2(n4076), .ZN(n4215) );
  AOI21_X1 U4536 ( .B1(n4092), .B2(n4077), .A(n4215), .ZN(n4078) );
  OAI211_X1 U4537 ( .C1(n4903), .C2(n4080), .A(n4079), .B(n4078), .ZN(n4081)
         );
  AOI21_X1 U4538 ( .B1(n4082), .B2(n4898), .A(n4081), .ZN(n4083) );
  INV_X1 U4539 ( .A(n4083), .ZN(U3235) );
  NOR2_X1 U4540 ( .A1(n4085), .A2(n2374), .ZN(n4086) );
  XNOR2_X1 U4541 ( .A(n4087), .B(n4086), .ZN(n4098) );
  INV_X1 U4542 ( .A(n4088), .ZN(n4286) );
  AOI22_X1 U4543 ( .A1(n4090), .A2(n4316), .B1(n4089), .B2(n4278), .ZN(n4094)
         );
  AOI22_X1 U4544 ( .A1(n4092), .A2(n4091), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4093) );
  OAI211_X1 U4545 ( .C1(n4903), .C2(n4286), .A(n4094), .B(n4093), .ZN(n4095)
         );
  INV_X1 U4546 ( .A(n4095), .ZN(n4096) );
  OAI21_X1 U4547 ( .B1(n4098), .B2(n4097), .A(n4096), .ZN(U3237) );
  MUX2_X1 U4548 ( .A(DATAO_REG_31__SCAN_IN), .B(n4099), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4549 ( .A(DATAO_REG_30__SCAN_IN), .B(n4100), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4550 ( .A(n4244), .B(DATAO_REG_29__SCAN_IN), .S(n4117), .Z(U3579)
         );
  MUX2_X1 U4551 ( .A(n4256), .B(DATAO_REG_28__SCAN_IN), .S(n4117), .Z(U3578)
         );
  MUX2_X1 U4552 ( .A(n4278), .B(DATAO_REG_27__SCAN_IN), .S(n4117), .Z(U3577)
         );
  MUX2_X1 U4553 ( .A(n4297), .B(DATAO_REG_26__SCAN_IN), .S(n4117), .Z(U3576)
         );
  INV_X1 U4554 ( .A(U4043), .ZN(n4119) );
  MUX2_X1 U4555 ( .A(n4316), .B(DATAO_REG_25__SCAN_IN), .S(n4119), .Z(U3575)
         );
  MUX2_X1 U4556 ( .A(n4342), .B(DATAO_REG_24__SCAN_IN), .S(n4119), .Z(U3574)
         );
  MUX2_X1 U4557 ( .A(n4101), .B(DATAO_REG_23__SCAN_IN), .S(n4117), .Z(U3573)
         );
  MUX2_X1 U4558 ( .A(n4102), .B(DATAO_REG_22__SCAN_IN), .S(n4119), .Z(U3572)
         );
  MUX2_X1 U4559 ( .A(n4103), .B(DATAO_REG_21__SCAN_IN), .S(n4117), .Z(U3571)
         );
  MUX2_X1 U4560 ( .A(n4104), .B(DATAO_REG_20__SCAN_IN), .S(n4117), .Z(U3570)
         );
  MUX2_X1 U4561 ( .A(n4105), .B(DATAO_REG_19__SCAN_IN), .S(n4119), .Z(U3569)
         );
  MUX2_X1 U4562 ( .A(n4106), .B(DATAO_REG_18__SCAN_IN), .S(n4117), .Z(U3568)
         );
  MUX2_X1 U4563 ( .A(n4107), .B(DATAO_REG_17__SCAN_IN), .S(n4117), .Z(U3567)
         );
  MUX2_X1 U4564 ( .A(n4885), .B(DATAO_REG_16__SCAN_IN), .S(n4119), .Z(U3566)
         );
  MUX2_X1 U4565 ( .A(n4108), .B(DATAO_REG_15__SCAN_IN), .S(n4117), .Z(U3565)
         );
  MUX2_X1 U4566 ( .A(n4886), .B(DATAO_REG_14__SCAN_IN), .S(n4117), .Z(U3564)
         );
  MUX2_X1 U4567 ( .A(n4109), .B(DATAO_REG_13__SCAN_IN), .S(n4119), .Z(U3563)
         );
  MUX2_X1 U4568 ( .A(n4110), .B(DATAO_REG_12__SCAN_IN), .S(n4117), .Z(U3562)
         );
  MUX2_X1 U4569 ( .A(n4111), .B(DATAO_REG_11__SCAN_IN), .S(n4117), .Z(U3561)
         );
  MUX2_X1 U4570 ( .A(n4112), .B(DATAO_REG_10__SCAN_IN), .S(n4119), .Z(U3560)
         );
  MUX2_X1 U4571 ( .A(n4113), .B(DATAO_REG_9__SCAN_IN), .S(n4119), .Z(U3559) );
  MUX2_X1 U4572 ( .A(n4814), .B(DATAO_REG_8__SCAN_IN), .S(n4117), .Z(U3558) );
  MUX2_X1 U4573 ( .A(n4114), .B(DATAO_REG_7__SCAN_IN), .S(n4119), .Z(U3557) );
  MUX2_X1 U4574 ( .A(n4816), .B(DATAO_REG_6__SCAN_IN), .S(n4117), .Z(U3556) );
  MUX2_X1 U4575 ( .A(n4115), .B(DATAO_REG_5__SCAN_IN), .S(n4117), .Z(U3555) );
  MUX2_X1 U4576 ( .A(n4116), .B(DATAO_REG_4__SCAN_IN), .S(n4117), .Z(U3554) );
  MUX2_X1 U4577 ( .A(n3050), .B(DATAO_REG_3__SCAN_IN), .S(n4117), .Z(U3553) );
  MUX2_X1 U4578 ( .A(n3034), .B(DATAO_REG_2__SCAN_IN), .S(n4119), .Z(U3552) );
  MUX2_X1 U4579 ( .A(n4118), .B(DATAO_REG_1__SCAN_IN), .S(n4119), .Z(U3551) );
  MUX2_X1 U4580 ( .A(n4120), .B(DATAO_REG_0__SCAN_IN), .S(n4119), .Z(U3550) );
  NAND2_X1 U4581 ( .A1(n4182), .A2(n4121), .ZN(n4133) );
  AOI22_X1 U4582 ( .A1(n4757), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4132) );
  OAI211_X1 U4583 ( .C1(n4124), .C2(n4123), .A(n4761), .B(n4122), .ZN(n4131)
         );
  MUX2_X1 U4584 ( .A(REG1_REG_1__SCAN_IN), .B(n4778), .S(n4125), .Z(n4127) );
  NAND2_X1 U4585 ( .A1(n4127), .A2(n4126), .ZN(n4128) );
  NAND3_X1 U4586 ( .A1(n4744), .A2(n4129), .A3(n4128), .ZN(n4130) );
  NAND4_X1 U4587 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(U3241)
         );
  AOI22_X1 U4588 ( .A1(n4757), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4145) );
  OAI211_X1 U4589 ( .C1(n4136), .C2(n4135), .A(n4761), .B(n4134), .ZN(n4141)
         );
  XNOR2_X1 U4590 ( .A(n4138), .B(n4137), .ZN(n4139) );
  NAND2_X1 U4591 ( .A1(n4744), .A2(n4139), .ZN(n4140) );
  AND2_X1 U4592 ( .A1(n4141), .A2(n4140), .ZN(n4144) );
  OR2_X1 U4593 ( .A1(n4759), .A2(n4142), .ZN(n4143) );
  NAND4_X1 U4594 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(U3242)
         );
  NAND2_X1 U4595 ( .A1(n4705), .A2(REG2_REG_11__SCAN_IN), .ZN(n4151) );
  INV_X1 U4596 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4874) );
  AOI22_X1 U4597 ( .A1(n4705), .A2(REG2_REG_11__SCAN_IN), .B1(n4874), .B2(
        n4867), .ZN(n4713) );
  NAND2_X1 U4598 ( .A1(n4452), .A2(REG2_REG_9__SCAN_IN), .ZN(n4148) );
  NAND2_X1 U4599 ( .A1(n4694), .A2(n4149), .ZN(n4150) );
  NAND2_X1 U4600 ( .A1(n4713), .A2(n4712), .ZN(n4711) );
  NAND2_X1 U4601 ( .A1(n4161), .A2(n4152), .ZN(n4153) );
  NAND2_X1 U4602 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4722), .ZN(n4721) );
  INV_X1 U4603 ( .A(n4164), .ZN(n4884) );
  INV_X1 U4604 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4731) );
  NOR2_X1 U4605 ( .A1(n4884), .A2(n4731), .ZN(n4730) );
  OAI22_X1 U4606 ( .A1(n4732), .A2(n4730), .B1(n4164), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n4154) );
  NOR2_X2 U4607 ( .A1(n4154), .A2(n4172), .ZN(n4177) );
  AOI211_X1 U4608 ( .C1(n3455), .C2(n4155), .A(n4176), .B(n4739), .ZN(n4170)
         );
  OAI21_X1 U4609 ( .B1(n4158), .B2(n4157), .A(n4156), .ZN(n4159) );
  NAND2_X1 U4610 ( .A1(n4694), .A2(n4159), .ZN(n4160) );
  XOR2_X1 U4611 ( .A(n4159), .B(n4694), .Z(n4698) );
  NAND2_X1 U4612 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4698), .ZN(n4697) );
  INV_X1 U4613 ( .A(n4161), .ZN(n4882) );
  NOR2_X1 U4614 ( .A1(n4162), .A2(n4882), .ZN(n4163) );
  NAND2_X1 U4615 ( .A1(n4164), .A2(REG1_REG_13__SCAN_IN), .ZN(n4725) );
  NOR2_X1 U4616 ( .A1(n4164), .A2(REG1_REG_13__SCAN_IN), .ZN(n4726) );
  AOI21_X1 U4617 ( .B1(n4728), .B2(n4725), .A(n4726), .ZN(n4173) );
  XNOR2_X1 U4618 ( .A(n4173), .B(n4172), .ZN(n4165) );
  NAND2_X1 U4619 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4165), .ZN(n4174) );
  OAI211_X1 U4620 ( .C1(n4165), .C2(REG1_REG_14__SCAN_IN), .A(n4744), .B(n4174), .ZN(n4168) );
  AOI21_X1 U4621 ( .B1(n4757), .B2(ADDR_REG_14__SCAN_IN), .A(n4166), .ZN(n4167) );
  OAI211_X1 U4622 ( .C1(n4759), .C2(n4172), .A(n4168), .B(n4167), .ZN(n4169)
         );
  OR2_X1 U4623 ( .A1(n4170), .A2(n4169), .ZN(U3254) );
  INV_X1 U4624 ( .A(n4744), .ZN(n4762) );
  XNOR2_X1 U4625 ( .A(n4186), .B(n4171), .ZN(n4188) );
  INV_X1 U4626 ( .A(n4172), .ZN(n4451) );
  NAND2_X1 U4627 ( .A1(n4451), .A2(n4173), .ZN(n4175) );
  NAND2_X1 U4628 ( .A1(n4175), .A2(n4174), .ZN(n4187) );
  XNOR2_X1 U4629 ( .A(n4188), .B(n4187), .ZN(n4185) );
  AND2_X1 U4630 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4892) );
  NAND2_X1 U4631 ( .A1(n4186), .A2(REG2_REG_15__SCAN_IN), .ZN(n4195) );
  OAI21_X1 U4632 ( .B1(n4186), .B2(REG2_REG_15__SCAN_IN), .A(n4195), .ZN(n4179) );
  OR2_X2 U4633 ( .A1(n4180), .A2(n4179), .ZN(n4196) );
  INV_X1 U4634 ( .A(n4196), .ZN(n4178) );
  AOI211_X1 U4635 ( .C1(n4180), .C2(n4179), .A(n4178), .B(n4739), .ZN(n4181)
         );
  AOI211_X1 U4636 ( .C1(n4757), .C2(ADDR_REG_15__SCAN_IN), .A(n4892), .B(n4181), .ZN(n4184) );
  NAND2_X1 U4637 ( .A1(n4182), .A2(n4186), .ZN(n4183) );
  OAI211_X1 U4638 ( .C1(n4762), .C2(n4185), .A(n4184), .B(n4183), .ZN(U3255)
         );
  AOI22_X1 U4639 ( .A1(n4188), .A2(n4187), .B1(REG1_REG_15__SCAN_IN), .B2(
        n4186), .ZN(n4189) );
  INV_X1 U4640 ( .A(n4189), .ZN(n4191) );
  NOR2_X1 U4641 ( .A1(n4190), .A2(n4191), .ZN(n4192) );
  NOR2_X1 U4642 ( .A1(n4211), .A2(REG1_REG_17__SCAN_IN), .ZN(n4217) );
  INV_X1 U4643 ( .A(n4217), .ZN(n4193) );
  OAI21_X1 U4644 ( .B1(n4204), .B2(n3576), .A(n4193), .ZN(n4194) );
  AOI21_X1 U4645 ( .B1(n2272), .B2(n4194), .A(n4216), .ZN(n4207) );
  XNOR2_X1 U4646 ( .A(n4204), .B(REG2_REG_17__SCAN_IN), .ZN(n4200) );
  NAND2_X1 U4647 ( .A1(n4197), .A2(n4905), .ZN(n4198) );
  NAND2_X1 U4648 ( .A1(n4199), .A2(n4200), .ZN(n4210) );
  AOI221_X1 U4649 ( .B1(n4200), .B2(n4210), .C1(n4199), .C2(n4210), .A(n4739), 
        .ZN(n4201) );
  OR2_X1 U4650 ( .A1(n4202), .A2(n4201), .ZN(n4203) );
  AOI21_X1 U4651 ( .B1(n4757), .B2(ADDR_REG_17__SCAN_IN), .A(n4203), .ZN(n4206) );
  OR2_X1 U4652 ( .A1(n4759), .A2(n4204), .ZN(n4205) );
  OAI211_X1 U4653 ( .C1(n4207), .C2(n4762), .A(n4206), .B(n4205), .ZN(U3257)
         );
  INV_X1 U4654 ( .A(n4221), .ZN(n4754) );
  NOR2_X1 U4655 ( .A1(n4754), .A2(n4208), .ZN(n4209) );
  AOI21_X1 U4656 ( .B1(n4208), .B2(n4754), .A(n4209), .ZN(n4213) );
  OAI21_X1 U4657 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4211), .A(n4210), .ZN(n4212) );
  AOI211_X1 U4658 ( .C1(n4213), .C2(n4212), .A(n4753), .B(n4739), .ZN(n4214)
         );
  AOI211_X1 U4659 ( .C1(n4757), .C2(ADDR_REG_18__SCAN_IN), .A(n4215), .B(n4214), .ZN(n4220) );
  XNOR2_X1 U4660 ( .A(n4754), .B(REG1_REG_18__SCAN_IN), .ZN(n4749) );
  NOR2_X1 U4661 ( .A1(n4217), .A2(n4216), .ZN(n4750) );
  XNOR2_X1 U4662 ( .A(n4749), .B(n4750), .ZN(n4218) );
  NAND2_X1 U4663 ( .A1(n4744), .A2(n4218), .ZN(n4219) );
  OAI211_X1 U4664 ( .C1(n4221), .C2(n4759), .A(n4220), .B(n4219), .ZN(U3258)
         );
  XNOR2_X1 U4665 ( .A(n4357), .B(n4222), .ZN(n4416) );
  NOR2_X1 U4666 ( .A1(n4224), .A2(n4223), .ZN(n4358) );
  AOI21_X1 U4667 ( .B1(n4225), .B2(n4359), .A(n4358), .ZN(n4412) );
  NOR2_X1 U4668 ( .A1(n4412), .A2(n4858), .ZN(n4226) );
  AOI21_X1 U4669 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4858), .A(n4226), .ZN(n4227) );
  OAI21_X1 U4670 ( .B1(n4416), .B2(n4871), .A(n4227), .ZN(U3260) );
  OAI22_X1 U4671 ( .A1(n4229), .A2(n4871), .B1(n4228), .B2(n4875), .ZN(n4230)
         );
  OAI21_X1 U4672 ( .B1(n4231), .B2(n4230), .A(n4328), .ZN(n4233) );
  NAND2_X1 U4673 ( .A1(n4858), .A2(REG2_REG_29__SCAN_IN), .ZN(n4232) );
  OAI211_X1 U4674 ( .C1(n2275), .C2(n4353), .A(n4233), .B(n4232), .ZN(U3354)
         );
  XNOR2_X1 U4675 ( .A(n4234), .B(n4241), .ZN(n4365) );
  AOI22_X1 U4676 ( .A1(n4858), .A2(REG2_REG_28__SCAN_IN), .B1(n4235), .B2(
        n4859), .ZN(n4251) );
  INV_X1 U4677 ( .A(n4236), .ZN(n4237) );
  OAI211_X1 U4678 ( .C1(n2299), .C2(n4238), .A(n4237), .B(n4406), .ZN(n4363)
         );
  INV_X1 U4679 ( .A(n4239), .ZN(n4240) );
  NOR2_X1 U4680 ( .A1(n4252), .A2(n4240), .ZN(n4242) );
  XNOR2_X1 U4681 ( .A(n4242), .B(n4241), .ZN(n4248) );
  AOI22_X1 U4682 ( .A1(n4244), .A2(n2263), .B1(n4243), .B2(n4359), .ZN(n4245)
         );
  OAI21_X1 U4683 ( .B1(n4246), .B2(n4339), .A(n4245), .ZN(n4247) );
  AOI21_X1 U4684 ( .B1(n4248), .B2(n4821), .A(n4247), .ZN(n4364) );
  OAI21_X1 U4685 ( .B1(n4450), .B2(n4363), .A(n4364), .ZN(n4249) );
  NAND2_X1 U4686 ( .A1(n4249), .A2(n4328), .ZN(n4250) );
  OAI211_X1 U4687 ( .C1(n4365), .C2(n4353), .A(n4251), .B(n4250), .ZN(U3262)
         );
  AOI21_X1 U4688 ( .B1(n4254), .B2(n4253), .A(n4252), .ZN(n4259) );
  AOI22_X1 U4689 ( .A1(n4256), .A2(n2263), .B1(n4255), .B2(n4359), .ZN(n4258)
         );
  NAND2_X1 U4690 ( .A1(n4297), .A2(n2260), .ZN(n4257) );
  OAI211_X1 U4691 ( .C1(n4259), .C2(n4344), .A(n4258), .B(n4257), .ZN(n4366)
         );
  AOI21_X1 U4692 ( .B1(n4260), .B2(n4859), .A(n4366), .ZN(n4270) );
  XNOR2_X1 U4693 ( .A(n4262), .B(n4261), .ZN(n4367) );
  INV_X1 U4694 ( .A(n4353), .ZN(n4263) );
  NAND2_X1 U4695 ( .A1(n4367), .A2(n4263), .ZN(n4269) );
  INV_X1 U4696 ( .A(n4370), .ZN(n4266) );
  OAI21_X1 U4697 ( .B1(n4266), .B2(n4265), .A(n4264), .ZN(n4424) );
  INV_X1 U4698 ( .A(n4424), .ZN(n4267) );
  AOI22_X1 U4699 ( .A1(n4267), .A2(n4908), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4858), .ZN(n4268) );
  OAI211_X1 U4700 ( .C1(n4858), .C2(n4270), .A(n4269), .B(n4268), .ZN(U3263)
         );
  XNOR2_X1 U4701 ( .A(n4272), .B(n4271), .ZN(n4374) );
  INV_X1 U4702 ( .A(n4273), .ZN(n4274) );
  OR2_X1 U4703 ( .A1(n4275), .A2(n4274), .ZN(n4277) );
  XNOR2_X1 U4704 ( .A(n4277), .B(n4276), .ZN(n4282) );
  NAND2_X1 U4705 ( .A1(n4316), .A2(n2260), .ZN(n4280) );
  NAND2_X1 U4706 ( .A1(n4278), .A2(n2263), .ZN(n4279) );
  OAI211_X1 U4707 ( .C1(n4819), .C2(n4283), .A(n4280), .B(n4279), .ZN(n4281)
         );
  AOI21_X1 U4708 ( .B1(n4282), .B2(n4821), .A(n4281), .ZN(n4373) );
  INV_X1 U4709 ( .A(n4373), .ZN(n4288) );
  OR2_X1 U4710 ( .A1(n4303), .A2(n4283), .ZN(n4371) );
  NAND3_X1 U4711 ( .A1(n4371), .A2(n4370), .A3(n4908), .ZN(n4285) );
  NAND2_X1 U4712 ( .A1(n4858), .A2(REG2_REG_26__SCAN_IN), .ZN(n4284) );
  OAI211_X1 U4713 ( .C1(n4875), .C2(n4286), .A(n4285), .B(n4284), .ZN(n4287)
         );
  AOI21_X1 U4714 ( .B1(n4288), .B2(n4328), .A(n4287), .ZN(n4289) );
  OAI21_X1 U4715 ( .B1(n4374), .B2(n4353), .A(n4289), .ZN(U3264) );
  XOR2_X1 U4716 ( .A(n4293), .B(n4290), .Z(n4376) );
  INV_X1 U4717 ( .A(n4376), .ZN(n4308) );
  NAND2_X1 U4718 ( .A1(n4292), .A2(n4291), .ZN(n4294) );
  XNOR2_X1 U4719 ( .A(n4294), .B(n4293), .ZN(n4295) );
  NAND2_X1 U4720 ( .A1(n4295), .A2(n4821), .ZN(n4299) );
  AOI22_X1 U4721 ( .A1(n4297), .A2(n2263), .B1(n4359), .B2(n4296), .ZN(n4298)
         );
  OAI211_X1 U4722 ( .C1(n4300), .C2(n4339), .A(n4299), .B(n4298), .ZN(n4375)
         );
  NOR2_X1 U4723 ( .A1(n4322), .A2(n4301), .ZN(n4302) );
  OR2_X1 U4724 ( .A1(n4303), .A2(n4302), .ZN(n4429) );
  AOI22_X1 U4725 ( .A1(n4858), .A2(REG2_REG_25__SCAN_IN), .B1(n4304), .B2(
        n4859), .ZN(n4305) );
  OAI21_X1 U4726 ( .B1(n4429), .B2(n4871), .A(n4305), .ZN(n4306) );
  AOI21_X1 U4727 ( .B1(n4375), .B2(n4328), .A(n4306), .ZN(n4307) );
  OAI21_X1 U4728 ( .B1(n4308), .B2(n4353), .A(n4307), .ZN(U3265) );
  XNOR2_X1 U4729 ( .A(n4309), .B(n4312), .ZN(n4380) );
  INV_X1 U4730 ( .A(n4380), .ZN(n4330) );
  NAND2_X1 U4731 ( .A1(n4311), .A2(n4310), .ZN(n4313) );
  XNOR2_X1 U4732 ( .A(n4313), .B(n4312), .ZN(n4314) );
  NAND2_X1 U4733 ( .A1(n4314), .A2(n4821), .ZN(n4318) );
  AOI22_X1 U4734 ( .A1(n4316), .A2(n2263), .B1(n4359), .B2(n4315), .ZN(n4317)
         );
  OAI211_X1 U4735 ( .C1(n4319), .C2(n4339), .A(n4318), .B(n4317), .ZN(n4379)
         );
  INV_X1 U4736 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4321) );
  OAI22_X1 U4737 ( .A1(n4328), .A2(n4321), .B1(n4320), .B2(n4875), .ZN(n4327)
         );
  INV_X1 U4738 ( .A(n4346), .ZN(n4325) );
  INV_X1 U4739 ( .A(n4322), .ZN(n4323) );
  OAI21_X1 U4740 ( .B1(n4325), .B2(n4324), .A(n4323), .ZN(n4433) );
  NOR2_X1 U4741 ( .A1(n4433), .A2(n4871), .ZN(n4326) );
  AOI211_X1 U4742 ( .C1(n4328), .C2(n4379), .A(n4327), .B(n4326), .ZN(n4329)
         );
  OAI21_X1 U4743 ( .B1(n4330), .B2(n4353), .A(n4329), .ZN(U3266) );
  NOR2_X1 U4744 ( .A1(n4332), .A2(n4331), .ZN(n4333) );
  XOR2_X1 U4745 ( .A(n4338), .B(n4333), .Z(n4384) );
  INV_X1 U4746 ( .A(n4384), .ZN(n4354) );
  OAI21_X1 U4747 ( .B1(n4336), .B2(n4335), .A(n4334), .ZN(n4337) );
  XOR2_X1 U4748 ( .A(n4338), .B(n4337), .Z(n4345) );
  OAI22_X1 U4749 ( .A1(n4340), .A2(n4339), .B1(n4819), .B2(n4347), .ZN(n4341)
         );
  AOI21_X1 U4750 ( .B1(n2263), .B2(n4342), .A(n4341), .ZN(n4343) );
  OAI21_X1 U4751 ( .B1(n4345), .B2(n4344), .A(n4343), .ZN(n4383) );
  INV_X1 U4752 ( .A(n4387), .ZN(n4348) );
  OAI21_X1 U4753 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(n4437) );
  AOI22_X1 U4754 ( .A1(n4858), .A2(REG2_REG_23__SCAN_IN), .B1(n4349), .B2(
        n4859), .ZN(n4350) );
  OAI21_X1 U4755 ( .B1(n4437), .B2(n4871), .A(n4350), .ZN(n4351) );
  AOI21_X1 U4756 ( .B1(n4383), .B2(n4328), .A(n4351), .ZN(n4352) );
  OAI21_X1 U4757 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(U3267) );
  NOR2_X1 U4758 ( .A1(n4412), .A2(n4844), .ZN(n4355) );
  AOI21_X1 U4759 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4844), .A(n4355), .ZN(n4356) );
  OAI21_X1 U4760 ( .B1(n4416), .B2(n4396), .A(n4356), .ZN(U3549) );
  AOI21_X1 U4761 ( .B1(n4360), .B2(n2268), .A(n4357), .ZN(n4909) );
  INV_X1 U4762 ( .A(n4909), .ZN(n4419) );
  INV_X1 U4763 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4361) );
  AOI21_X1 U4764 ( .B1(n4360), .B2(n4359), .A(n4358), .ZN(n4911) );
  MUX2_X1 U4765 ( .A(n4361), .B(n4911), .S(n4411), .Z(n4362) );
  OAI21_X1 U4766 ( .B1(n4419), .B2(n4396), .A(n4362), .ZN(U3548) );
  OAI211_X1 U4767 ( .C1(n4365), .C2(n2466), .A(n4364), .B(n4363), .ZN(n4420)
         );
  MUX2_X1 U4768 ( .A(REG1_REG_28__SCAN_IN), .B(n4420), .S(n4411), .Z(U3546) );
  INV_X1 U4769 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4368) );
  AOI21_X1 U4770 ( .B1(n4367), .B2(n4840), .A(n4366), .ZN(n4421) );
  MUX2_X1 U4771 ( .A(n4368), .B(n4421), .S(n4411), .Z(n4369) );
  OAI21_X1 U4772 ( .B1(n4396), .B2(n4424), .A(n4369), .ZN(U3545) );
  NAND3_X1 U4773 ( .A1(n4371), .A2(n4406), .A3(n4370), .ZN(n4372) );
  OAI211_X1 U4774 ( .C1(n4374), .C2(n2466), .A(n4373), .B(n4372), .ZN(n4425)
         );
  MUX2_X1 U4775 ( .A(REG1_REG_26__SCAN_IN), .B(n4425), .S(n4411), .Z(U3544) );
  INV_X1 U4776 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4377) );
  AOI21_X1 U4777 ( .B1(n4376), .B2(n4840), .A(n4375), .ZN(n4426) );
  MUX2_X1 U4778 ( .A(n4377), .B(n4426), .S(n4846), .Z(n4378) );
  OAI21_X1 U4779 ( .B1(n4396), .B2(n4429), .A(n4378), .ZN(U3543) );
  INV_X1 U4780 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4381) );
  AOI21_X1 U4781 ( .B1(n4380), .B2(n4840), .A(n4379), .ZN(n4430) );
  MUX2_X1 U4782 ( .A(n4381), .B(n4430), .S(n4411), .Z(n4382) );
  OAI21_X1 U4783 ( .B1(n4396), .B2(n4433), .A(n4382), .ZN(U3542) );
  INV_X1 U4784 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4385) );
  AOI21_X1 U4785 ( .B1(n4384), .B2(n4840), .A(n4383), .ZN(n4434) );
  MUX2_X1 U4786 ( .A(n4385), .B(n4434), .S(n4846), .Z(n4386) );
  OAI21_X1 U4787 ( .B1(n4396), .B2(n4437), .A(n4386), .ZN(U3541) );
  NAND3_X1 U4788 ( .A1(n4388), .A2(n4406), .A3(n4387), .ZN(n4389) );
  OAI211_X1 U4789 ( .C1(n4391), .C2(n2466), .A(n4390), .B(n4389), .ZN(n4438)
         );
  MUX2_X1 U4790 ( .A(REG1_REG_22__SCAN_IN), .B(n4438), .S(n4846), .Z(U3540) );
  INV_X1 U4791 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4394) );
  AOI21_X1 U4792 ( .B1(n4393), .B2(n4840), .A(n4392), .ZN(n4439) );
  MUX2_X1 U4793 ( .A(n4394), .B(n4439), .S(n4411), .Z(n4395) );
  OAI21_X1 U4794 ( .B1(n4396), .B2(n4443), .A(n4395), .ZN(U3539) );
  NAND3_X1 U4795 ( .A1(n4398), .A2(n4397), .A3(n4406), .ZN(n4399) );
  OAI211_X1 U4796 ( .C1(n4401), .C2(n4774), .A(n4400), .B(n4399), .ZN(n4444)
         );
  MUX2_X1 U4797 ( .A(REG1_REG_20__SCAN_IN), .B(n4444), .S(n4846), .Z(U3538) );
  OAI211_X1 U4798 ( .C1(n4404), .C2(n2466), .A(n4403), .B(n4402), .ZN(n4445)
         );
  MUX2_X1 U4799 ( .A(REG1_REG_18__SCAN_IN), .B(n4445), .S(n4411), .Z(U3536) );
  NAND3_X1 U4800 ( .A1(n4407), .A2(n4406), .A3(n4405), .ZN(n4408) );
  OAI211_X1 U4801 ( .C1(n4410), .C2(n2466), .A(n4409), .B(n4408), .ZN(n4446)
         );
  MUX2_X1 U4802 ( .A(REG1_REG_16__SCAN_IN), .B(n4446), .S(n4411), .Z(U3534) );
  NOR2_X1 U4803 ( .A1(n4412), .A2(n4414), .ZN(n4413) );
  AOI21_X1 U4804 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4414), .A(n4413), .ZN(n4415) );
  OAI21_X1 U4805 ( .B1(n4416), .B2(n4442), .A(n4415), .ZN(U3517) );
  INV_X1 U4806 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4417) );
  MUX2_X1 U4807 ( .A(n4417), .B(n4911), .S(n4849), .Z(n4418) );
  OAI21_X1 U4808 ( .B1(n4419), .B2(n4442), .A(n4418), .ZN(U3516) );
  MUX2_X1 U4809 ( .A(REG0_REG_28__SCAN_IN), .B(n4420), .S(n4849), .Z(U3514) );
  INV_X1 U4810 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4422) );
  MUX2_X1 U4811 ( .A(n4422), .B(n4421), .S(n4849), .Z(n4423) );
  OAI21_X1 U4812 ( .B1(n4424), .B2(n4442), .A(n4423), .ZN(U3513) );
  MUX2_X1 U4813 ( .A(REG0_REG_26__SCAN_IN), .B(n4425), .S(n4849), .Z(U3512) );
  INV_X1 U4814 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4427) );
  MUX2_X1 U4815 ( .A(n4427), .B(n4426), .S(n4849), .Z(n4428) );
  OAI21_X1 U4816 ( .B1(n4429), .B2(n4442), .A(n4428), .ZN(U3511) );
  INV_X1 U4817 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4431) );
  MUX2_X1 U4818 ( .A(n4431), .B(n4430), .S(n4849), .Z(n4432) );
  OAI21_X1 U4819 ( .B1(n4433), .B2(n4442), .A(n4432), .ZN(U3510) );
  INV_X1 U4820 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4435) );
  MUX2_X1 U4821 ( .A(n4435), .B(n4434), .S(n4849), .Z(n4436) );
  OAI21_X1 U4822 ( .B1(n4437), .B2(n4442), .A(n4436), .ZN(U3509) );
  MUX2_X1 U4823 ( .A(REG0_REG_22__SCAN_IN), .B(n4438), .S(n4849), .Z(U3508) );
  INV_X1 U4824 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4440) );
  MUX2_X1 U4825 ( .A(n4440), .B(n4439), .S(n4849), .Z(n4441) );
  OAI21_X1 U4826 ( .B1(n4443), .B2(n4442), .A(n4441), .ZN(U3507) );
  MUX2_X1 U4827 ( .A(REG0_REG_20__SCAN_IN), .B(n4444), .S(n4849), .Z(U3506) );
  MUX2_X1 U4828 ( .A(REG0_REG_18__SCAN_IN), .B(n4445), .S(n4849), .Z(U3503) );
  MUX2_X1 U4829 ( .A(REG0_REG_16__SCAN_IN), .B(n4446), .S(n4849), .Z(U3499) );
  MUX2_X1 U4830 ( .A(n4447), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4831 ( .A(n2892), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4832 ( .A(DATAI_22_), .B(n4448), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4833 ( .A(n4449), .B(DATAI_20_), .S(U3149), .Z(U3332) );
  MUX2_X1 U4834 ( .A(n4450), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4835 ( .A(DATAI_18_), .B(n4754), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U4836 ( .A(DATAI_14_), .B(n4451), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U4837 ( .A(n4452), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4838 ( .A(n2973), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U4839 ( .A(n4453), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4840 ( .A(n4454), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U4841 ( .A(DATAI_23_), .ZN(n4474) );
  OAI21_X1 U4842 ( .B1(STATE_REG_SCAN_IN), .B2(n4474), .A(n4455), .ZN(U3329)
         );
  AND2_X1 U4843 ( .A1(D_REG_2__SCAN_IN), .A2(n2262), .ZN(U3320) );
  AND2_X1 U4844 ( .A1(D_REG_3__SCAN_IN), .A2(n2262), .ZN(U3319) );
  AND2_X1 U4845 ( .A1(D_REG_4__SCAN_IN), .A2(n2262), .ZN(U3318) );
  AND2_X1 U4846 ( .A1(D_REG_5__SCAN_IN), .A2(n2262), .ZN(U3317) );
  AND2_X1 U4847 ( .A1(D_REG_7__SCAN_IN), .A2(n2262), .ZN(U3315) );
  AND2_X1 U4848 ( .A1(D_REG_8__SCAN_IN), .A2(n2262), .ZN(U3314) );
  AND2_X1 U4849 ( .A1(D_REG_9__SCAN_IN), .A2(n2262), .ZN(U3313) );
  AND2_X1 U4850 ( .A1(D_REG_10__SCAN_IN), .A2(n2262), .ZN(U3312) );
  AND2_X1 U4851 ( .A1(D_REG_11__SCAN_IN), .A2(n2262), .ZN(U3311) );
  AND2_X1 U4852 ( .A1(D_REG_12__SCAN_IN), .A2(n2262), .ZN(U3310) );
  AND2_X1 U4853 ( .A1(D_REG_13__SCAN_IN), .A2(n2262), .ZN(U3309) );
  AND2_X1 U4854 ( .A1(D_REG_14__SCAN_IN), .A2(n2262), .ZN(U3308) );
  AND2_X1 U4855 ( .A1(D_REG_15__SCAN_IN), .A2(n2262), .ZN(U3307) );
  AND2_X1 U4856 ( .A1(D_REG_16__SCAN_IN), .A2(n2262), .ZN(U3306) );
  AND2_X1 U4857 ( .A1(D_REG_17__SCAN_IN), .A2(n2262), .ZN(U3305) );
  AND2_X1 U4858 ( .A1(D_REG_18__SCAN_IN), .A2(n2262), .ZN(U3304) );
  AND2_X1 U4859 ( .A1(D_REG_19__SCAN_IN), .A2(n2262), .ZN(U3303) );
  AND2_X1 U4860 ( .A1(D_REG_20__SCAN_IN), .A2(n2262), .ZN(U3302) );
  AND2_X1 U4861 ( .A1(D_REG_21__SCAN_IN), .A2(n2262), .ZN(U3301) );
  AND2_X1 U4862 ( .A1(D_REG_22__SCAN_IN), .A2(n2262), .ZN(U3300) );
  AND2_X1 U4863 ( .A1(D_REG_23__SCAN_IN), .A2(n2262), .ZN(U3299) );
  AND2_X1 U4864 ( .A1(D_REG_24__SCAN_IN), .A2(n2262), .ZN(U3298) );
  AND2_X1 U4865 ( .A1(D_REG_25__SCAN_IN), .A2(n2262), .ZN(U3297) );
  AND2_X1 U4866 ( .A1(D_REG_26__SCAN_IN), .A2(n2262), .ZN(U3296) );
  AND2_X1 U4867 ( .A1(D_REG_27__SCAN_IN), .A2(n2262), .ZN(U3295) );
  AND2_X1 U4868 ( .A1(D_REG_28__SCAN_IN), .A2(n2262), .ZN(U3294) );
  AND2_X1 U4869 ( .A1(D_REG_29__SCAN_IN), .A2(n2262), .ZN(U3293) );
  AND2_X1 U4870 ( .A1(D_REG_30__SCAN_IN), .A2(n2262), .ZN(U3292) );
  AND2_X1 U4871 ( .A1(D_REG_31__SCAN_IN), .A2(n2262), .ZN(U3291) );
  NAND2_X1 U4872 ( .A1(n2262), .A2(D_REG_6__SCAN_IN), .ZN(n4653) );
  INV_X1 U4873 ( .A(keyinput_121), .ZN(n4536) );
  AOI22_X1 U4874 ( .A1(n4548), .A2(keyinput_118), .B1(n2295), .B2(keyinput_119), .ZN(n4457) );
  OAI221_X1 U4875 ( .B1(n4548), .B2(keyinput_118), .C1(n2295), .C2(
        keyinput_119), .A(n4457), .ZN(n4534) );
  OAI22_X1 U4876 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_110), .B1(
        REG3_REG_25__SCAN_IN), .B2(keyinput_109), .ZN(n4458) );
  AOI221_X1 U4877 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_110), .C1(
        keyinput_109), .C2(REG3_REG_25__SCAN_IN), .A(n4458), .ZN(n4527) );
  INV_X1 U4878 ( .A(keyinput_103), .ZN(n4514) );
  INV_X1 U4879 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4602) );
  INV_X1 U4880 ( .A(keyinput_99), .ZN(n4508) );
  OAI22_X1 U4881 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_96), .B1(keyinput_95), 
        .B2(DATAI_0_), .ZN(n4459) );
  AOI221_X1 U4882 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_96), .C1(DATAI_0_), 
        .C2(keyinput_95), .A(n4459), .ZN(n4506) );
  AOI22_X1 U4883 ( .A1(DATAI_5_), .A2(keyinput_90), .B1(DATAI_6_), .B2(
        keyinput_89), .ZN(n4460) );
  OAI221_X1 U4884 ( .B1(DATAI_5_), .B2(keyinput_90), .C1(DATAI_6_), .C2(
        keyinput_89), .A(n4460), .ZN(n4501) );
  INV_X1 U4885 ( .A(keyinput_82), .ZN(n4488) );
  INV_X1 U4886 ( .A(DATAI_13_), .ZN(n4883) );
  OAI22_X1 U4887 ( .A1(n4462), .A2(keyinput_77), .B1(keyinput_76), .B2(
        DATAI_19_), .ZN(n4461) );
  AOI221_X1 U4888 ( .B1(n4462), .B2(keyinput_77), .C1(DATAI_19_), .C2(
        keyinput_76), .A(n4461), .ZN(n4486) );
  INV_X1 U4889 ( .A(keyinput_71), .ZN(n4472) );
  XOR2_X1 U4890 ( .A(DATAI_29_), .B(keyinput_66), .Z(n4470) );
  AOI22_X1 U4891 ( .A1(DATAI_31_), .A2(keyinput_64), .B1(DATAI_30_), .B2(
        keyinput_65), .ZN(n4463) );
  OAI221_X1 U4892 ( .B1(DATAI_31_), .B2(keyinput_64), .C1(DATAI_30_), .C2(
        keyinput_65), .A(n4463), .ZN(n4469) );
  INV_X1 U4893 ( .A(DATAI_26_), .ZN(n4465) );
  AOI22_X1 U4894 ( .A1(n4559), .A2(keyinput_68), .B1(keyinput_69), .B2(n4465), 
        .ZN(n4464) );
  OAI221_X1 U4895 ( .B1(n4559), .B2(keyinput_68), .C1(n4465), .C2(keyinput_69), 
        .A(n4464), .ZN(n4468) );
  AOI22_X1 U4896 ( .A1(DATAI_25_), .A2(keyinput_70), .B1(DATAI_28_), .B2(
        keyinput_67), .ZN(n4466) );
  OAI221_X1 U4897 ( .B1(DATAI_25_), .B2(keyinput_70), .C1(DATAI_28_), .C2(
        keyinput_67), .A(n4466), .ZN(n4467) );
  AOI211_X1 U4898 ( .C1(n4470), .C2(n4469), .A(n4468), .B(n4467), .ZN(n4471)
         );
  AOI221_X1 U4899 ( .B1(DATAI_24_), .B2(n4472), .C1(n4565), .C2(keyinput_71), 
        .A(n4471), .ZN(n4478) );
  INV_X1 U4900 ( .A(DATAI_22_), .ZN(n4568) );
  AOI22_X1 U4901 ( .A1(n4474), .A2(keyinput_72), .B1(keyinput_73), .B2(n4568), 
        .ZN(n4473) );
  OAI221_X1 U4902 ( .B1(n4474), .B2(keyinput_72), .C1(n4568), .C2(keyinput_73), 
        .A(n4473), .ZN(n4477) );
  OAI22_X1 U4903 ( .A1(DATAI_21_), .A2(keyinput_74), .B1(keyinput_75), .B2(
        DATAI_20_), .ZN(n4475) );
  AOI221_X1 U4904 ( .B1(DATAI_21_), .B2(keyinput_74), .C1(DATAI_20_), .C2(
        keyinput_75), .A(n4475), .ZN(n4476) );
  OAI21_X1 U4905 ( .B1(n4478), .B2(n4477), .A(n4476), .ZN(n4485) );
  AOI22_X1 U4906 ( .A1(n2737), .A2(keyinput_78), .B1(keyinput_81), .B2(n4480), 
        .ZN(n4479) );
  OAI221_X1 U4907 ( .B1(n2737), .B2(keyinput_78), .C1(n4480), .C2(keyinput_81), 
        .A(n4479), .ZN(n4484) );
  AOI22_X1 U4908 ( .A1(DATAI_16_), .A2(keyinput_79), .B1(n4482), .B2(
        keyinput_80), .ZN(n4481) );
  OAI221_X1 U4909 ( .B1(DATAI_16_), .B2(keyinput_79), .C1(n4482), .C2(
        keyinput_80), .A(n4481), .ZN(n4483) );
  AOI211_X1 U4910 ( .C1(n4486), .C2(n4485), .A(n4484), .B(n4483), .ZN(n4487)
         );
  AOI221_X1 U4911 ( .B1(DATAI_13_), .B2(n4488), .C1(n4883), .C2(keyinput_82), 
        .A(n4487), .ZN(n4495) );
  INV_X1 U4912 ( .A(DATAI_12_), .ZN(n4881) );
  AOI22_X1 U4913 ( .A1(DATAI_11_), .A2(keyinput_84), .B1(n4881), .B2(
        keyinput_83), .ZN(n4489) );
  OAI221_X1 U4914 ( .B1(DATAI_11_), .B2(keyinput_84), .C1(n4881), .C2(
        keyinput_83), .A(n4489), .ZN(n4494) );
  OAI22_X1 U4915 ( .A1(DATAI_10_), .A2(keyinput_85), .B1(DATAI_9_), .B2(
        keyinput_86), .ZN(n4490) );
  AOI221_X1 U4916 ( .B1(DATAI_10_), .B2(keyinput_85), .C1(keyinput_86), .C2(
        DATAI_9_), .A(n4490), .ZN(n4493) );
  INV_X1 U4917 ( .A(DATAI_8_), .ZN(n4850) );
  INV_X1 U4918 ( .A(DATAI_7_), .ZN(n4809) );
  OAI22_X1 U4919 ( .A1(n4850), .A2(keyinput_87), .B1(n4809), .B2(keyinput_88), 
        .ZN(n4491) );
  AOI221_X1 U4920 ( .B1(n4850), .B2(keyinput_87), .C1(keyinput_88), .C2(n4809), 
        .A(n4491), .ZN(n4492) );
  OAI211_X1 U4921 ( .C1(n4495), .C2(n4494), .A(n4493), .B(n4492), .ZN(n4500)
         );
  INV_X1 U4922 ( .A(DATAI_3_), .ZN(n4591) );
  OAI22_X1 U4923 ( .A1(n4591), .A2(keyinput_92), .B1(keyinput_94), .B2(
        DATAI_1_), .ZN(n4496) );
  AOI221_X1 U4924 ( .B1(n4591), .B2(keyinput_92), .C1(DATAI_1_), .C2(
        keyinput_94), .A(n4496), .ZN(n4499) );
  OAI22_X1 U4925 ( .A1(DATAI_4_), .A2(keyinput_91), .B1(DATAI_2_), .B2(
        keyinput_93), .ZN(n4497) );
  AOI221_X1 U4926 ( .B1(DATAI_4_), .B2(keyinput_91), .C1(keyinput_93), .C2(
        DATAI_2_), .A(n4497), .ZN(n4498) );
  OAI211_X1 U4927 ( .C1(n4501), .C2(n4500), .A(n4499), .B(n4498), .ZN(n4505)
         );
  AOI22_X1 U4928 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_97), .B1(n4503), 
        .B2(keyinput_98), .ZN(n4502) );
  OAI221_X1 U4929 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_97), .C1(n4503), 
        .C2(keyinput_98), .A(n4502), .ZN(n4504) );
  AOI21_X1 U4930 ( .B1(n4506), .B2(n4505), .A(n4504), .ZN(n4507) );
  AOI221_X1 U4931 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_99), .C1(n4602), 
        .C2(n4508), .A(n4507), .ZN(n4511) );
  AOI22_X1 U4932 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_101), .B1(n2569), 
        .B2(keyinput_102), .ZN(n4509) );
  OAI221_X1 U4933 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_101), .C1(n2569), 
        .C2(keyinput_102), .A(n4509), .ZN(n4510) );
  AOI211_X1 U4934 ( .C1(n4608), .C2(keyinput_100), .A(n4511), .B(n4510), .ZN(
        n4512) );
  OAI21_X1 U4935 ( .B1(n4608), .B2(keyinput_100), .A(n4512), .ZN(n4513) );
  OAI221_X1 U4936 ( .B1(REG3_REG_19__SCAN_IN), .B2(n4514), .C1(n4610), .C2(
        keyinput_103), .A(n4513), .ZN(n4520) );
  OAI22_X1 U4937 ( .A1(n2802), .A2(keyinput_104), .B1(REG3_REG_21__SCAN_IN), 
        .B2(keyinput_107), .ZN(n4515) );
  AOI221_X1 U4938 ( .B1(n2802), .B2(keyinput_104), .C1(keyinput_107), .C2(
        REG3_REG_21__SCAN_IN), .A(n4515), .ZN(n4519) );
  XOR2_X1 U4939 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_106), .Z(n4518) );
  OAI22_X1 U4940 ( .A1(n4616), .A2(keyinput_108), .B1(keyinput_105), .B2(
        REG3_REG_8__SCAN_IN), .ZN(n4516) );
  AOI221_X1 U4941 ( .B1(n4616), .B2(keyinput_108), .C1(REG3_REG_8__SCAN_IN), 
        .C2(keyinput_105), .A(n4516), .ZN(n4517) );
  NAND4_X1 U4942 ( .A1(n4520), .A2(n4519), .A3(n4518), .A4(n4517), .ZN(n4526)
         );
  AOI22_X1 U4943 ( .A1(n4626), .A2(keyinput_112), .B1(n2590), .B2(keyinput_111), .ZN(n4521) );
  OAI221_X1 U4944 ( .B1(n4626), .B2(keyinput_112), .C1(n2590), .C2(
        keyinput_111), .A(n4521), .ZN(n4525) );
  AOI22_X1 U4945 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_114), .B1(n4523), 
        .B2(keyinput_113), .ZN(n4522) );
  OAI221_X1 U4946 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_114), .C1(n4523), 
        .C2(keyinput_113), .A(n4522), .ZN(n4524) );
  AOI211_X1 U4947 ( .C1(n4527), .C2(n4526), .A(n4525), .B(n4524), .ZN(n4531)
         );
  OAI22_X1 U4948 ( .A1(n4635), .A2(keyinput_117), .B1(keyinput_116), .B2(
        REG3_REG_0__SCAN_IN), .ZN(n4528) );
  AOI221_X1 U4949 ( .B1(n4635), .B2(keyinput_117), .C1(REG3_REG_0__SCAN_IN), 
        .C2(keyinput_116), .A(n4528), .ZN(n4529) );
  OAI21_X1 U4950 ( .B1(keyinput_115), .B2(REG3_REG_9__SCAN_IN), .A(n4529), 
        .ZN(n4530) );
  AOI211_X1 U4951 ( .C1(keyinput_115), .C2(REG3_REG_9__SCAN_IN), .A(n4531), 
        .B(n4530), .ZN(n4533) );
  NAND2_X1 U4952 ( .A1(n2405), .A2(keyinput_120), .ZN(n4532) );
  OAI221_X1 U4953 ( .B1(n4534), .B2(n4533), .C1(n2405), .C2(keyinput_120), .A(
        n4532), .ZN(n4535) );
  OAI221_X1 U4954 ( .B1(IR_REG_2__SCAN_IN), .B2(n4536), .C1(n2565), .C2(
        keyinput_121), .A(n4535), .ZN(n4540) );
  XNOR2_X1 U4955 ( .A(n4537), .B(keyinput_123), .ZN(n4539) );
  XNOR2_X1 U4956 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n4538) );
  NAND3_X1 U4957 ( .A1(n4540), .A2(n4539), .A3(n4538), .ZN(n4542) );
  XNOR2_X1 U4958 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_124), .ZN(n4541) );
  NAND2_X1 U4959 ( .A1(n4542), .A2(n4541), .ZN(n4545) );
  OAI22_X1 U4960 ( .A1(n2642), .A2(keyinput_125), .B1(keyinput_127), .B2(
        IR_REG_8__SCAN_IN), .ZN(n4543) );
  AOI221_X1 U4961 ( .B1(n2642), .B2(keyinput_125), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_127), .A(n4543), .ZN(n4544) );
  OAI211_X1 U4962 ( .C1(IR_REG_7__SCAN_IN), .C2(keyinput_126), .A(n4545), .B(
        n4544), .ZN(n4546) );
  AOI21_X1 U4963 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_126), .A(n4546), .ZN(
        n4651) );
  INV_X1 U4964 ( .A(keyinput_57), .ZN(n4640) );
  AOI22_X1 U4965 ( .A1(n4548), .A2(keyinput_54), .B1(n2295), .B2(keyinput_55), 
        .ZN(n4547) );
  OAI221_X1 U4966 ( .B1(n4548), .B2(keyinput_54), .C1(n2295), .C2(keyinput_55), 
        .A(n4547), .ZN(n4637) );
  OAI22_X1 U4967 ( .A1(n4550), .A2(keyinput_51), .B1(REG3_REG_0__SCAN_IN), 
        .B2(keyinput_52), .ZN(n4549) );
  AOI221_X1 U4968 ( .B1(n4550), .B2(keyinput_51), .C1(keyinput_52), .C2(
        REG3_REG_0__SCAN_IN), .A(n4549), .ZN(n4633) );
  INV_X1 U4969 ( .A(keyinput_39), .ZN(n4611) );
  INV_X1 U4970 ( .A(keyinput_35), .ZN(n4603) );
  OAI22_X1 U4971 ( .A1(U3149), .A2(keyinput_32), .B1(keyinput_31), .B2(
        DATAI_0_), .ZN(n4551) );
  AOI221_X1 U4972 ( .B1(U3149), .B2(keyinput_32), .C1(DATAI_0_), .C2(
        keyinput_31), .A(n4551), .ZN(n4600) );
  AOI22_X1 U4973 ( .A1(DATAI_6_), .A2(keyinput_25), .B1(DATAI_7_), .B2(
        keyinput_24), .ZN(n4552) );
  OAI221_X1 U4974 ( .B1(DATAI_6_), .B2(keyinput_25), .C1(DATAI_7_), .C2(
        keyinput_24), .A(n4552), .ZN(n4596) );
  INV_X1 U4975 ( .A(keyinput_18), .ZN(n4581) );
  INV_X1 U4976 ( .A(DATAI_19_), .ZN(n4554) );
  OAI22_X1 U4977 ( .A1(n4554), .A2(keyinput_12), .B1(keyinput_13), .B2(
        DATAI_18_), .ZN(n4553) );
  AOI221_X1 U4978 ( .B1(n4554), .B2(keyinput_12), .C1(DATAI_18_), .C2(
        keyinput_13), .A(n4553), .ZN(n4579) );
  INV_X1 U4979 ( .A(keyinput_7), .ZN(n4566) );
  XNOR2_X1 U4980 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n4563) );
  AOI22_X1 U4981 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(DATAI_30_), .B2(
        keyinput_1), .ZN(n4555) );
  OAI221_X1 U4982 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(DATAI_30_), .C2(
        keyinput_1), .A(n4555), .ZN(n4562) );
  INV_X1 U4983 ( .A(DATAI_28_), .ZN(n4906) );
  AOI22_X1 U4984 ( .A1(n4906), .A2(keyinput_3), .B1(keyinput_6), .B2(n4557), 
        .ZN(n4556) );
  OAI221_X1 U4985 ( .B1(n4906), .B2(keyinput_3), .C1(n4557), .C2(keyinput_6), 
        .A(n4556), .ZN(n4561) );
  AOI22_X1 U4986 ( .A1(DATAI_26_), .A2(keyinput_5), .B1(n4559), .B2(keyinput_4), .ZN(n4558) );
  OAI221_X1 U4987 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(n4559), .C2(
        keyinput_4), .A(n4558), .ZN(n4560) );
  AOI211_X1 U4988 ( .C1(n4563), .C2(n4562), .A(n4561), .B(n4560), .ZN(n4564)
         );
  AOI221_X1 U4989 ( .B1(DATAI_24_), .B2(n4566), .C1(n4565), .C2(keyinput_7), 
        .A(n4564), .ZN(n4573) );
  AOI22_X1 U4990 ( .A1(DATAI_23_), .A2(keyinput_8), .B1(n4568), .B2(keyinput_9), .ZN(n4567) );
  OAI221_X1 U4991 ( .B1(DATAI_23_), .B2(keyinput_8), .C1(n4568), .C2(
        keyinput_9), .A(n4567), .ZN(n4572) );
  INV_X1 U4992 ( .A(DATAI_20_), .ZN(n4570) );
  OAI22_X1 U4993 ( .A1(n4570), .A2(keyinput_11), .B1(keyinput_10), .B2(
        DATAI_21_), .ZN(n4569) );
  AOI221_X1 U4994 ( .B1(n4570), .B2(keyinput_11), .C1(DATAI_21_), .C2(
        keyinput_10), .A(n4569), .ZN(n4571) );
  OAI21_X1 U4995 ( .B1(n4573), .B2(n4572), .A(n4571), .ZN(n4578) );
  AOI22_X1 U4996 ( .A1(n4904), .A2(keyinput_15), .B1(n2737), .B2(keyinput_14), 
        .ZN(n4574) );
  OAI221_X1 U4997 ( .B1(n4904), .B2(keyinput_15), .C1(n2737), .C2(keyinput_14), 
        .A(n4574), .ZN(n4577) );
  AOI22_X1 U4998 ( .A1(DATAI_14_), .A2(keyinput_17), .B1(DATAI_15_), .B2(
        keyinput_16), .ZN(n4575) );
  OAI221_X1 U4999 ( .B1(DATAI_14_), .B2(keyinput_17), .C1(DATAI_15_), .C2(
        keyinput_16), .A(n4575), .ZN(n4576) );
  AOI211_X1 U5000 ( .C1(n4579), .C2(n4578), .A(n4577), .B(n4576), .ZN(n4580)
         );
  AOI221_X1 U5001 ( .B1(DATAI_13_), .B2(keyinput_18), .C1(n4883), .C2(n4581), 
        .A(n4580), .ZN(n4589) );
  AOI22_X1 U5002 ( .A1(n2670), .A2(keyinput_20), .B1(n4881), .B2(keyinput_19), 
        .ZN(n4582) );
  OAI221_X1 U5003 ( .B1(n2670), .B2(keyinput_20), .C1(n4881), .C2(keyinput_19), 
        .A(n4582), .ZN(n4588) );
  OAI22_X1 U5004 ( .A1(DATAI_10_), .A2(keyinput_21), .B1(DATAI_5_), .B2(
        keyinput_26), .ZN(n4583) );
  AOI221_X1 U5005 ( .B1(DATAI_10_), .B2(keyinput_21), .C1(keyinput_26), .C2(
        DATAI_5_), .A(n4583), .ZN(n4587) );
  INV_X1 U5006 ( .A(DATAI_9_), .ZN(n4585) );
  OAI22_X1 U5007 ( .A1(n4585), .A2(keyinput_22), .B1(n4850), .B2(keyinput_23), 
        .ZN(n4584) );
  AOI221_X1 U5008 ( .B1(n4585), .B2(keyinput_22), .C1(keyinput_23), .C2(n4850), 
        .A(n4584), .ZN(n4586) );
  OAI211_X1 U5009 ( .C1(n4589), .C2(n4588), .A(n4587), .B(n4586), .ZN(n4595)
         );
  OAI22_X1 U5010 ( .A1(n4591), .A2(keyinput_28), .B1(keyinput_30), .B2(
        DATAI_1_), .ZN(n4590) );
  AOI221_X1 U5011 ( .B1(n4591), .B2(keyinput_28), .C1(DATAI_1_), .C2(
        keyinput_30), .A(n4590), .ZN(n4594) );
  OAI22_X1 U5012 ( .A1(DATAI_4_), .A2(keyinput_27), .B1(DATAI_2_), .B2(
        keyinput_29), .ZN(n4592) );
  AOI221_X1 U5013 ( .B1(DATAI_4_), .B2(keyinput_27), .C1(keyinput_29), .C2(
        DATAI_2_), .A(n4592), .ZN(n4593) );
  OAI211_X1 U5014 ( .C1(n4596), .C2(n4595), .A(n4594), .B(n4593), .ZN(n4599)
         );
  AOI22_X1 U5015 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_34), .B1(
        REG3_REG_7__SCAN_IN), .B2(keyinput_33), .ZN(n4597) );
  OAI221_X1 U5016 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_34), .C1(
        REG3_REG_7__SCAN_IN), .C2(keyinput_33), .A(n4597), .ZN(n4598) );
  AOI21_X1 U5017 ( .B1(n4600), .B2(n4599), .A(n4598), .ZN(n4601) );
  AOI221_X1 U5018 ( .B1(REG3_REG_14__SCAN_IN), .B2(n4603), .C1(n4602), .C2(
        keyinput_35), .A(n4601), .ZN(n4607) );
  OAI22_X1 U5019 ( .A1(n2569), .A2(keyinput_38), .B1(REG3_REG_10__SCAN_IN), 
        .B2(keyinput_37), .ZN(n4604) );
  AOI221_X1 U5020 ( .B1(n2569), .B2(keyinput_38), .C1(keyinput_37), .C2(
        REG3_REG_10__SCAN_IN), .A(n4604), .ZN(n4605) );
  OAI21_X1 U5021 ( .B1(keyinput_36), .B2(n4608), .A(n4605), .ZN(n4606) );
  AOI211_X1 U5022 ( .C1(keyinput_36), .C2(n4608), .A(n4607), .B(n4606), .ZN(
        n4609) );
  AOI221_X1 U5023 ( .B1(REG3_REG_19__SCAN_IN), .B2(n4611), .C1(n4610), .C2(
        keyinput_39), .A(n4609), .ZN(n4622) );
  AOI22_X1 U5024 ( .A1(n2775), .A2(keyinput_43), .B1(n4613), .B2(keyinput_41), 
        .ZN(n4612) );
  OAI221_X1 U5025 ( .B1(n2775), .B2(keyinput_43), .C1(n4613), .C2(keyinput_41), 
        .A(n4612), .ZN(n4614) );
  INV_X1 U5026 ( .A(n4614), .ZN(n4620) );
  INV_X1 U5027 ( .A(keyinput_40), .ZN(n4615) );
  XNOR2_X1 U5028 ( .A(n4615), .B(REG3_REG_28__SCAN_IN), .ZN(n4619) );
  XOR2_X1 U5029 ( .A(keyinput_44), .B(n4616), .Z(n4618) );
  XNOR2_X1 U5030 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .ZN(n4617) );
  NAND4_X1 U5031 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n4621)
         );
  NOR2_X1 U5032 ( .A1(n4622), .A2(n4621), .ZN(n4631) );
  AOI22_X1 U5033 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_45), .B1(n4624), 
        .B2(keyinput_46), .ZN(n4623) );
  OAI221_X1 U5034 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_45), .C1(n4624), 
        .C2(keyinput_46), .A(n4623), .ZN(n4630) );
  OAI22_X1 U5035 ( .A1(n2590), .A2(keyinput_47), .B1(n4626), .B2(keyinput_48), 
        .ZN(n4625) );
  AOI221_X1 U5036 ( .B1(n2590), .B2(keyinput_47), .C1(keyinput_48), .C2(n4626), 
        .A(n4625), .ZN(n4629) );
  OAI22_X1 U5037 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_50), .B1(keyinput_49), .B2(REG3_REG_24__SCAN_IN), .ZN(n4627) );
  AOI221_X1 U5038 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_50), .C1(
        REG3_REG_24__SCAN_IN), .C2(keyinput_49), .A(n4627), .ZN(n4628) );
  OAI211_X1 U5039 ( .C1(n4631), .C2(n4630), .A(n4629), .B(n4628), .ZN(n4632)
         );
  OAI211_X1 U5040 ( .C1(n4635), .C2(keyinput_53), .A(n4633), .B(n4632), .ZN(
        n4634) );
  AOI21_X1 U5041 ( .B1(n4635), .B2(keyinput_53), .A(n4634), .ZN(n4636) );
  OAI22_X1 U5042 ( .A1(keyinput_56), .A2(n2405), .B1(n4637), .B2(n4636), .ZN(
        n4638) );
  AOI21_X1 U5043 ( .B1(keyinput_56), .B2(n2405), .A(n4638), .ZN(n4639) );
  AOI221_X1 U5044 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_57), .C1(n2565), .C2(
        n4640), .A(n4639), .ZN(n4645) );
  XNOR2_X1 U5045 ( .A(n4641), .B(keyinput_58), .ZN(n4643) );
  XNOR2_X1 U5046 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_59), .ZN(n4642) );
  NAND2_X1 U5047 ( .A1(n4643), .A2(n4642), .ZN(n4644) );
  OAI22_X1 U5048 ( .A1(n4645), .A2(n4644), .B1(IR_REG_5__SCAN_IN), .B2(
        keyinput_60), .ZN(n4646) );
  AOI21_X1 U5049 ( .B1(keyinput_60), .B2(IR_REG_5__SCAN_IN), .A(n4646), .ZN(
        n4650) );
  XNOR2_X1 U5050 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .ZN(n4649) );
  AOI22_X1 U5051 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_62), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_61), .ZN(n4647) );
  OAI221_X1 U5052 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_62), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_61), .A(n4647), .ZN(n4648) );
  NOR4_X1 U5053 ( .A1(n4651), .A2(n4650), .A3(n4649), .A4(n4648), .ZN(n4652)
         );
  XNOR2_X1 U5054 ( .A(n4653), .B(n4652), .ZN(U3316) );
  AOI211_X1 U5055 ( .C1(n4655), .C2(n4654), .A(n2290), .B(n4739), .ZN(n4657)
         );
  AOI211_X1 U5056 ( .C1(n4757), .C2(ADDR_REG_5__SCAN_IN), .A(n4657), .B(n4656), 
        .ZN(n4662) );
  OAI211_X1 U5057 ( .C1(n4660), .C2(n4659), .A(n4744), .B(n4658), .ZN(n4661)
         );
  OAI211_X1 U5058 ( .C1(n4759), .C2(n4799), .A(n4662), .B(n4661), .ZN(U3245)
         );
  AOI211_X1 U5059 ( .C1(n4665), .C2(n4664), .A(n4663), .B(n4739), .ZN(n4667)
         );
  AOI211_X1 U5060 ( .C1(n4757), .C2(ADDR_REG_6__SCAN_IN), .A(n4667), .B(n4666), 
        .ZN(n4671) );
  OAI211_X1 U5061 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4669), .A(n4744), .B(n4668), 
        .ZN(n4670) );
  OAI211_X1 U5062 ( .C1(n4759), .C2(n4801), .A(n4671), .B(n4670), .ZN(U3246)
         );
  AOI22_X1 U5063 ( .A1(n4673), .A2(n4672), .B1(REG2_REG_7__SCAN_IN), .B2(n4810), .ZN(n4675) );
  OAI21_X1 U5064 ( .B1(n4676), .B2(n4675), .A(n4761), .ZN(n4674) );
  AOI21_X1 U5065 ( .B1(n4676), .B2(n4675), .A(n4674), .ZN(n4678) );
  AOI211_X1 U5066 ( .C1(n4757), .C2(ADDR_REG_7__SCAN_IN), .A(n4678), .B(n4677), 
        .ZN(n4684) );
  AOI21_X1 U5067 ( .B1(n4810), .B2(n4845), .A(n4679), .ZN(n4682) );
  AOI21_X1 U5068 ( .B1(n4682), .B2(n4681), .A(n4762), .ZN(n4680) );
  OAI21_X1 U5069 ( .B1(n4682), .B2(n4681), .A(n4680), .ZN(n4683) );
  OAI211_X1 U5070 ( .C1(n4759), .C2(n4810), .A(n4684), .B(n4683), .ZN(U3247)
         );
  AOI211_X1 U5071 ( .C1(n4687), .C2(n4686), .A(n4685), .B(n4762), .ZN(n4689)
         );
  AOI211_X1 U5072 ( .C1(n4757), .C2(ADDR_REG_8__SCAN_IN), .A(n4689), .B(n4688), 
        .ZN(n4693) );
  OAI211_X1 U5073 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4691), .A(n4761), .B(n4690), 
        .ZN(n4692) );
  OAI211_X1 U5074 ( .C1(n4759), .C2(n3254), .A(n4693), .B(n4692), .ZN(U3248)
         );
  OAI211_X1 U5075 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4696), .A(n4761), .B(n4695), .ZN(n4700) );
  OAI211_X1 U5076 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4698), .A(n4744), .B(n4697), .ZN(n4699) );
  OAI211_X1 U5077 ( .C1(n4759), .C2(n2422), .A(n4700), .B(n4699), .ZN(n4701)
         );
  AOI211_X1 U5078 ( .C1(n4757), .C2(ADDR_REG_10__SCAN_IN), .A(n4702), .B(n4701), .ZN(n4703) );
  INV_X1 U5079 ( .A(n4703), .ZN(U3250) );
  INV_X1 U5080 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5081 ( .A1(n4705), .A2(REG1_REG_11__SCAN_IN), .B1(n4704), .B2(
        n4867), .ZN(n4708) );
  OAI21_X1 U5082 ( .B1(n4708), .B2(n4707), .A(n4744), .ZN(n4706) );
  AOI21_X1 U5083 ( .B1(n4708), .B2(n4707), .A(n4706), .ZN(n4710) );
  AOI211_X1 U5084 ( .C1(n4757), .C2(ADDR_REG_11__SCAN_IN), .A(n4710), .B(n4709), .ZN(n4715) );
  OAI211_X1 U5085 ( .C1(n4713), .C2(n4712), .A(n4761), .B(n4711), .ZN(n4714)
         );
  OAI211_X1 U5086 ( .C1(n4759), .C2(n4867), .A(n4715), .B(n4714), .ZN(U3251)
         );
  AOI211_X1 U5087 ( .C1(n4718), .C2(n4717), .A(n4716), .B(n4762), .ZN(n4720)
         );
  AOI211_X1 U5088 ( .C1(n4757), .C2(ADDR_REG_12__SCAN_IN), .A(n4720), .B(n4719), .ZN(n4724) );
  OAI211_X1 U5089 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4722), .A(n4761), .B(n4721), .ZN(n4723) );
  OAI211_X1 U5090 ( .C1(n4759), .C2(n4882), .A(n4724), .B(n4723), .ZN(U3252)
         );
  INV_X1 U5091 ( .A(n4725), .ZN(n4727) );
  NOR2_X1 U5092 ( .A1(n4727), .A2(n4726), .ZN(n4729) );
  XOR2_X1 U5093 ( .A(n4729), .B(n4728), .Z(n4738) );
  AOI21_X1 U5094 ( .B1(n4884), .B2(n4731), .A(n4730), .ZN(n4733) );
  XNOR2_X1 U5095 ( .A(n4733), .B(n4732), .ZN(n4734) );
  OAI22_X1 U5096 ( .A1(n4884), .A2(n4759), .B1(n4739), .B2(n4734), .ZN(n4735)
         );
  AOI211_X1 U5097 ( .C1(n4757), .C2(ADDR_REG_13__SCAN_IN), .A(n4736), .B(n4735), .ZN(n4737) );
  OAI21_X1 U5098 ( .B1(n4738), .B2(n4762), .A(n4737), .ZN(U3253) );
  AOI221_X1 U5099 ( .B1(n4741), .B2(n4740), .C1(n3478), .C2(n4740), .A(n4739), 
        .ZN(n4742) );
  AOI211_X1 U5100 ( .C1(n4757), .C2(ADDR_REG_16__SCAN_IN), .A(n4743), .B(n4742), .ZN(n4748) );
  OAI221_X1 U5101 ( .B1(n4746), .B2(REG1_REG_16__SCAN_IN), .C1(n4746), .C2(
        n4745), .A(n4744), .ZN(n4747) );
  OAI211_X1 U5102 ( .C1(n4759), .C2(n4905), .A(n4748), .B(n4747), .ZN(U3256)
         );
  INV_X1 U5103 ( .A(n4749), .ZN(n4751) );
  MUX2_X1 U5104 ( .A(REG1_REG_19__SCAN_IN), .B(n3795), .S(n4828), .Z(n4752) );
  MUX2_X1 U5105 ( .A(REG2_REG_19__SCAN_IN), .B(n3569), .S(n4828), .Z(n4755) );
  AOI21_X1 U5106 ( .B1(n4757), .B2(ADDR_REG_19__SCAN_IN), .A(n4756), .ZN(n4758) );
  OAI21_X1 U5107 ( .B1(n4828), .B2(n4759), .A(n4758), .ZN(n4760) );
  AOI22_X1 U5108 ( .A1(STATE_REG_SCAN_IN), .A2(n2295), .B1(n2296), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5109 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5110 ( .A1(n4849), .A2(n4764), .B1(n4763), .B2(n4414), .ZN(U3467)
         );
  INV_X1 U5111 ( .A(n4765), .ZN(n4767) );
  AOI21_X1 U5112 ( .B1(n4768), .B2(n4767), .A(n4766), .ZN(n4772) );
  AOI22_X1 U5113 ( .A1(n4769), .A2(n4869), .B1(REG3_REG_0__SCAN_IN), .B2(n4859), .ZN(n4770) );
  OAI221_X1 U5114 ( .B1(n4858), .B2(n4772), .C1(n4328), .C2(n4771), .A(n4770), 
        .ZN(U3290) );
  OAI22_X1 U5115 ( .A1(n4775), .A2(n4774), .B1(n4823), .B2(n4773), .ZN(n4776)
         );
  NOR2_X1 U5116 ( .A1(n4777), .A2(n4776), .ZN(n4780) );
  AOI22_X1 U5117 ( .A1(n4846), .A2(n4780), .B1(n4778), .B2(n4844), .ZN(U3519)
         );
  INV_X1 U5118 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4779) );
  AOI22_X1 U5119 ( .A1(n4849), .A2(n4780), .B1(n4779), .B2(n4414), .ZN(U3469)
         );
  AOI22_X1 U5120 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4858), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4859), .ZN(n4784) );
  AOI22_X1 U5121 ( .A1(n4782), .A2(n4869), .B1(n4908), .B2(n4781), .ZN(n4783)
         );
  OAI211_X1 U5122 ( .C1(n4858), .C2(n4785), .A(n4784), .B(n4783), .ZN(U3288)
         );
  AOI22_X1 U5123 ( .A1(n4858), .A2(REG2_REG_3__SCAN_IN), .B1(n4859), .B2(n2569), .ZN(n4789) );
  AOI22_X1 U5124 ( .A1(n4787), .A2(n4869), .B1(n4908), .B2(n4786), .ZN(n4788)
         );
  OAI211_X1 U5125 ( .C1(n4858), .C2(n4790), .A(n4789), .B(n4788), .ZN(U3287)
         );
  INV_X1 U5126 ( .A(n4791), .ZN(n4793) );
  AOI211_X1 U5127 ( .C1(n4795), .C2(n4794), .A(n4793), .B(n4792), .ZN(n4797)
         );
  AOI22_X1 U5128 ( .A1(n4846), .A2(n4797), .B1(n3231), .B2(n4844), .ZN(U3522)
         );
  INV_X1 U5129 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4796) );
  AOI22_X1 U5130 ( .A1(n4849), .A2(n4797), .B1(n4796), .B2(n4414), .ZN(U3475)
         );
  INV_X1 U5131 ( .A(DATAI_5_), .ZN(n4798) );
  AOI22_X1 U5132 ( .A1(STATE_REG_SCAN_IN), .A2(n4799), .B1(n4798), .B2(U3149), 
        .ZN(U3347) );
  INV_X1 U5133 ( .A(DATAI_6_), .ZN(n4800) );
  AOI22_X1 U5134 ( .A1(STATE_REG_SCAN_IN), .A2(n4801), .B1(n4800), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5135 ( .A1(n4802), .A2(n4859), .B1(REG2_REG_6__SCAN_IN), .B2(n4858), .ZN(n4807) );
  INV_X1 U5136 ( .A(n4803), .ZN(n4804) );
  AOI22_X1 U5137 ( .A1(n4805), .A2(n4869), .B1(n4908), .B2(n4804), .ZN(n4806)
         );
  OAI211_X1 U5138 ( .C1(n4858), .C2(n4808), .A(n4807), .B(n4806), .ZN(U3284)
         );
  AOI22_X1 U5139 ( .A1(STATE_REG_SCAN_IN), .A2(n4810), .B1(n4809), .B2(U3149), 
        .ZN(U3345) );
  NAND2_X1 U5140 ( .A1(n4812), .A2(n4811), .ZN(n4813) );
  XNOR2_X1 U5141 ( .A(n4813), .B(n4830), .ZN(n4822) );
  NAND2_X1 U5142 ( .A1(n4814), .A2(n2263), .ZN(n4818) );
  NAND2_X1 U5143 ( .A1(n4816), .A2(n2260), .ZN(n4817) );
  OAI211_X1 U5144 ( .C1(n4819), .C2(n2292), .A(n4818), .B(n4817), .ZN(n4820)
         );
  AOI21_X1 U5145 ( .B1(n4822), .B2(n4821), .A(n4820), .ZN(n4842) );
  AOI21_X1 U5146 ( .B1(n4825), .B2(n4824), .A(n4823), .ZN(n4827) );
  AND2_X1 U5147 ( .A1(n4827), .A2(n4826), .ZN(n4839) );
  AOI21_X1 U5148 ( .B1(n4839), .B2(n4828), .A(n4858), .ZN(n4835) );
  NAND2_X1 U5149 ( .A1(n4829), .A2(n4830), .ZN(n4831) );
  AND2_X1 U5150 ( .A1(n4832), .A2(n4831), .ZN(n4841) );
  NAND2_X1 U5151 ( .A1(n4841), .A2(n4833), .ZN(n4834) );
  NAND3_X1 U5152 ( .A1(n4842), .A2(n4835), .A3(n4834), .ZN(n4836) );
  OAI21_X1 U5153 ( .B1(REG2_REG_7__SCAN_IN), .B2(n4328), .A(n4836), .ZN(n4837)
         );
  OAI21_X1 U5154 ( .B1(n4838), .B2(n4875), .A(n4837), .ZN(U3283) );
  AOI21_X1 U5155 ( .B1(n4841), .B2(n4840), .A(n4839), .ZN(n4843) );
  AND2_X1 U5156 ( .A1(n4843), .A2(n4842), .ZN(n4848) );
  AOI22_X1 U5157 ( .A1(n4846), .A2(n4848), .B1(n4845), .B2(n4844), .ZN(U3525)
         );
  INV_X1 U5158 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4847) );
  AOI22_X1 U5159 ( .A1(n4849), .A2(n4848), .B1(n4847), .B2(n4414), .ZN(U3481)
         );
  AOI22_X1 U5160 ( .A1(STATE_REG_SCAN_IN), .A2(n3254), .B1(n4850), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5161 ( .A1(n4851), .A2(n4859), .B1(REG2_REG_8__SCAN_IN), .B2(n4858), .ZN(n4855) );
  AOI22_X1 U5162 ( .A1(n4853), .A2(n4869), .B1(n4908), .B2(n4852), .ZN(n4854)
         );
  OAI211_X1 U5163 ( .C1(n4858), .C2(n4856), .A(n4855), .B(n4854), .ZN(U3282)
         );
  INV_X1 U5164 ( .A(DATAI_10_), .ZN(n4857) );
  AOI22_X1 U5165 ( .A1(STATE_REG_SCAN_IN), .A2(n2422), .B1(n4857), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5166 ( .A1(n4860), .A2(n4859), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4858), .ZN(n4865) );
  INV_X1 U5167 ( .A(n4861), .ZN(n4862) );
  AOI22_X1 U5168 ( .A1(n4863), .A2(n4869), .B1(n4908), .B2(n4862), .ZN(n4864)
         );
  OAI211_X1 U5169 ( .C1(n4858), .C2(n4866), .A(n4865), .B(n4864), .ZN(U3280)
         );
  AOI22_X1 U5170 ( .A1(STATE_REG_SCAN_IN), .A2(n4867), .B1(n2670), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5171 ( .A(n4868), .ZN(n4873) );
  INV_X1 U5172 ( .A(n4869), .ZN(n4872) );
  OAI22_X1 U5173 ( .A1(n4873), .A2(n4872), .B1(n4871), .B2(n4870), .ZN(n4878)
         );
  OAI22_X1 U5174 ( .A1(n4876), .A2(n4875), .B1(n4874), .B2(n4328), .ZN(n4877)
         );
  NOR2_X1 U5175 ( .A1(n4878), .A2(n4877), .ZN(n4879) );
  OAI21_X1 U5176 ( .B1(n4880), .B2(n4858), .A(n4879), .ZN(U3279) );
  AOI22_X1 U5177 ( .A1(STATE_REG_SCAN_IN), .A2(n4882), .B1(n4881), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5178 ( .A1(STATE_REG_SCAN_IN), .A2(n4884), .B1(n4883), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5179 ( .A(n4885), .ZN(n4890) );
  INV_X1 U5180 ( .A(n4886), .ZN(n4887) );
  OAI22_X1 U5181 ( .A1(n4890), .A2(n4889), .B1(n4888), .B2(n4887), .ZN(n4891)
         );
  AOI211_X1 U5182 ( .C1(n4894), .C2(n4893), .A(n4892), .B(n4891), .ZN(n4901)
         );
  XNOR2_X1 U5183 ( .A(n4896), .B(n4895), .ZN(n4897) );
  XNOR2_X1 U5184 ( .A(n4026), .B(n4897), .ZN(n4899) );
  NAND2_X1 U5185 ( .A1(n4899), .A2(n4898), .ZN(n4900) );
  OAI211_X1 U5186 ( .C1(n4903), .C2(n4902), .A(n4901), .B(n4900), .ZN(U3238)
         );
  AOI22_X1 U5187 ( .A1(STATE_REG_SCAN_IN), .A2(n4905), .B1(n4904), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5188 ( .A1(STATE_REG_SCAN_IN), .A2(n4907), .B1(n4906), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5189 ( .A1(n4909), .A2(n4908), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4858), .ZN(n4910) );
  OAI21_X1 U5190 ( .B1(n4858), .B2(n4911), .A(n4910), .ZN(U3261) );
  NAND2_X1 U2297 ( .A1(n2980), .A2(n2979), .ZN(n3924) );
  OAI22_X1 U2301 ( .A1(n3245), .A2(n2417), .B1(n2418), .B2(n3249), .ZN(n3251)
         );
  CLKBUF_X1 U2306 ( .A(n2558), .Z(n2684) );
  XNOR2_X1 U2331 ( .A(n3251), .B(n4801), .ZN(n4664) );
  BUF_X4 U2773 ( .A(n2566), .Z(n3639) );
  AND2_X1 U2774 ( .A1(n2937), .A2(n3013), .ZN(n4914) );
  CLKBUF_X1 U2881 ( .A(n4846), .Z(n4411) );
endmodule

