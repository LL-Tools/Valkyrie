

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4268, n4269, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010;

  OAI21_X1 U4774 ( .B1(n8550), .B2(n4835), .A(n4281), .ZN(n6367) );
  OR2_X1 U4775 ( .A1(n6276), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6286) );
  OAI22_X1 U4776 ( .A1(n6690), .A2(n6689), .B1(n6702), .B2(n5683), .ZN(n6656)
         );
  INV_X1 U4777 ( .A(n5817), .ZN(n5885) );
  NAND4_X2 U4778 ( .A1(n4903), .A2(n4902), .A3(n4901), .A4(n4900), .ZN(n5732)
         );
  AND2_X1 U4780 ( .A1(n9389), .A2(n4898), .ZN(n4966) );
  NAND2_X1 U4781 ( .A1(n8153), .A2(n8152), .ZN(n6834) );
  NAND2_X1 U4782 ( .A1(n5982), .A2(n5981), .ZN(n6101) );
  AOI21_X1 U4783 ( .B1(n7600), .B2(n7595), .A(n7596), .ZN(n7563) );
  INV_X1 U4784 ( .A(n5791), .ZN(n5908) );
  OR2_X1 U4785 ( .A1(n9157), .A2(n6441), .ZN(n7795) );
  INV_X1 U4786 ( .A(n4941), .ZN(n6008) );
  INV_X1 U4787 ( .A(n6183), .ZN(n6199) );
  OAI22_X1 U4788 ( .A1(n6656), .A2(n6657), .B1(n5684), .B2(n6546), .ZN(n9845)
         );
  NAND2_X1 U4789 ( .A1(n8190), .A2(n8182), .ZN(n8321) );
  INV_X1 U4790 ( .A(n8278), .ZN(n8301) );
  INV_X1 U4791 ( .A(n6922), .ZN(n6881) );
  AND2_X1 U4792 ( .A1(n6320), .A2(n6319), .ZN(n6588) );
  OR2_X1 U4793 ( .A1(n8883), .A2(n8886), .ZN(n8884) );
  AND2_X1 U4795 ( .A1(n4899), .A2(n4898), .ZN(n5001) );
  OAI21_X1 U4796 ( .B1(n7195), .B2(n7777), .A(n5478), .ZN(n7249) );
  NAND2_X2 U4797 ( .A1(n5640), .A2(n5641), .ZN(n5989) );
  OAI21_X1 U4798 ( .B1(n8005), .B2(n8555), .A(n7974), .ZN(n8080) );
  AND2_X1 U4799 ( .A1(n6293), .A2(n6292), .ZN(n8508) );
  OAI21_X1 U4800 ( .B1(n4293), .B2(n9934), .A(n6435), .ZN(n4578) );
  NAND2_X1 U4801 ( .A1(n6367), .A2(n8310), .ZN(n8515) );
  AND2_X1 U4802 ( .A1(n8875), .A2(n5934), .ZN(n6480) );
  XNOR2_X1 U4803 ( .A(n6450), .B(n6453), .ZN(n7903) );
  INV_X1 U4804 ( .A(n6929), .ZN(n6758) );
  NOR2_X2 U4805 ( .A1(n5564), .A2(n5509), .ZN(n5531) );
  NAND2_X2 U4806 ( .A1(n5515), .A2(n5514), .ZN(n5528) );
  AND4_X4 U4807 ( .A1(n5997), .A2(n5996), .A3(n5995), .A4(n5994), .ZN(n6929)
         );
  NOR2_X2 U4808 ( .A1(n6173), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6185) );
  XNOR2_X2 U4809 ( .A(n5732), .B(n9683), .ZN(n6903) );
  OR2_X2 U4810 ( .A1(n5078), .A2(n9617), .ZN(n7648) );
  NAND4_X2 U4811 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n8985)
         );
  NAND2_X1 U4812 ( .A1(n5982), .A2(n5981), .ZN(n4268) );
  OAI211_X2 U4813 ( .C1(n5236), .C2(n4390), .A(n4387), .B(n4385), .ZN(n7928)
         );
  XNOR2_X1 U4814 ( .A(n8685), .B(n8508), .ZN(n8497) );
  INV_X1 U4815 ( .A(n8985), .ZN(n6441) );
  NAND4_X1 U4816 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n8393)
         );
  INV_X1 U4817 ( .A(n6870), .ZN(n9879) );
  INV_X2 U4818 ( .A(n5287), .ZN(n5340) );
  INV_X2 U4820 ( .A(n5989), .ZN(n6204) );
  AOI21_X1 U4822 ( .B1(n8515), .B2(n4826), .A(n4824), .ZN(n4823) );
  NOR2_X1 U4823 ( .A1(n8853), .A2(n8764), .ZN(n8769) );
  OAI21_X1 U4824 ( .B1(n8497), .B2(n4825), .A(n8270), .ZN(n4824) );
  AOI21_X1 U4825 ( .B1(n8578), .B2(n8563), .A(n8564), .ZN(n8562) );
  NOR2_X1 U4826 ( .A1(n8497), .A2(n4829), .ZN(n4826) );
  XNOR2_X1 U4827 ( .A(n7722), .B(n7721), .ZN(n7724) );
  NAND2_X1 U4828 ( .A1(n6411), .A2(n6410), .ZN(n7722) );
  OR2_X1 U4829 ( .A1(n8265), .A2(n8264), .ZN(n8341) );
  NAND2_X1 U4830 ( .A1(n7617), .A2(n7616), .ZN(n4651) );
  NAND2_X1 U4831 ( .A1(n7454), .A2(n4649), .ZN(n7515) );
  NAND2_X1 U4832 ( .A1(n4849), .A2(n4847), .ZN(n7323) );
  OAI22_X1 U4833 ( .A1(n7249), .A2(n5479), .B1(n9768), .B2(n8892), .ZN(n7345)
         );
  AND2_X1 U4834 ( .A1(n7453), .A2(n7457), .ZN(n4649) );
  XNOR2_X1 U4835 ( .A(n7452), .B(n8197), .ZN(n7413) );
  NAND2_X1 U4836 ( .A1(n7182), .A2(n4873), .ZN(n7263) );
  NAND2_X1 U4837 ( .A1(n6073), .A2(n6072), .ZN(n7273) );
  NAND2_X1 U4838 ( .A1(n5080), .A2(n7772), .ZN(n7842) );
  AOI21_X1 U4839 ( .B1(n6517), .B2(n6495), .A(n6494), .ZN(n6493) );
  OAI21_X1 U4840 ( .B1(n6777), .B2(n6515), .A(n6514), .ZN(n6517) );
  NOR2_X1 U4841 ( .A1(n6286), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6297) );
  AOI21_X1 U4842 ( .B1(n6725), .B2(n6718), .A(n6717), .ZN(n6720) );
  AOI21_X1 U4843 ( .B1(n4654), .B2(n7057), .A(n4319), .ZN(n4652) );
  NAND2_X1 U4844 ( .A1(n4683), .A2(n5179), .ZN(n5197) );
  NAND2_X1 U4845 ( .A1(n8192), .A2(n8183), .ZN(n8322) );
  AND2_X1 U4846 ( .A1(n8178), .A2(n8175), .ZN(n8318) );
  NAND2_X2 U4847 ( .A1(n6396), .A2(n8618), .ZN(n8608) );
  NAND2_X1 U4848 ( .A1(n6057), .A2(n6043), .ZN(n8316) );
  NAND2_X1 U4849 ( .A1(n5042), .A2(n5041), .ZN(n5078) );
  OR2_X1 U4850 ( .A1(n9619), .A2(n7045), .ZN(n7643) );
  NAND2_X1 U4851 ( .A1(n6758), .A2(n6013), .ZN(n8153) );
  INV_X1 U4852 ( .A(n7283), .ZN(n8391) );
  NAND2_X1 U4853 ( .A1(n4328), .A2(n4583), .ZN(n6922) );
  OAI21_X1 U4854 ( .B1(n5950), .B2(n5958), .A(n9104), .ZN(n8894) );
  AND4_X1 U4855 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n7283)
         );
  NAND4_X1 U4856 ( .A1(n4988), .A2(n4987), .A3(n4986), .A4(n4985), .ZN(n9653)
         );
  AND3_X2 U4857 ( .A1(n6001), .A2(n6000), .A3(n5999), .ZN(n6865) );
  OR2_X1 U4858 ( .A1(n4268), .A2(n5993), .ZN(n5994) );
  INV_X2 U4859 ( .A(n4377), .ZN(n5937) );
  CLKBUF_X2 U4860 ( .A(n6017), .Z(n4271) );
  INV_X1 U4861 ( .A(n5980), .ZN(n5981) );
  OR2_X1 U4862 ( .A1(n8742), .A2(n5974), .ZN(n5975) );
  XNOR2_X1 U4863 ( .A(n5978), .B(n5977), .ZN(n5980) );
  XNOR2_X1 U4864 ( .A(n5522), .B(n5517), .ZN(n7448) );
  AOI21_X1 U4865 ( .B1(n4714), .B2(n5103), .A(n4713), .ZN(n4712) );
  NAND2_X2 U4866 ( .A1(n4927), .A2(n6008), .ZN(n7751) );
  NAND2_X1 U4867 ( .A1(n4897), .A2(n4896), .ZN(n9396) );
  XNOR2_X1 U4868 ( .A(n4893), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4899) );
  XNOR2_X1 U4869 ( .A(n5536), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6858) );
  NAND2_X1 U4870 ( .A1(n4896), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U4871 ( .A1(n5417), .A2(n6458), .ZN(n4927) );
  XNOR2_X1 U4872 ( .A(n6306), .B(n6305), .ZN(n8303) );
  XNOR2_X1 U4873 ( .A(n4906), .B(n4905), .ZN(n5417) );
  OAI21_X1 U4874 ( .B1(n5633), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6306) );
  OR2_X1 U4875 ( .A1(n6135), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6144) );
  INV_X2 U4876 ( .A(n8748), .ZN(n7936) );
  NAND2_X1 U4877 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U4878 ( .A1(n4860), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U4879 ( .A1(n4662), .A2(n4660), .ZN(n4941) );
  AND3_X1 U4880 ( .A1(n4781), .A2(n5405), .A3(n5413), .ZN(n4889) );
  INV_X4 U4881 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U4882 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4421) );
  NOR2_X1 U4883 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4422) );
  INV_X1 U4884 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5405) );
  INV_X1 U4885 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5413) );
  INV_X4 U4886 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4887 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n6985) );
  NOR2_X2 U4888 ( .A1(n7372), .A2(n7371), .ZN(n9142) );
  NAND2_X1 U4889 ( .A1(n5989), .A2(n6008), .ZN(n6082) );
  NAND2_X4 U4890 ( .A1(n5982), .A2(n5980), .ZN(n6077) );
  XNOR2_X1 U4892 ( .A(n5580), .B(n5579), .ZN(n6532) );
  NAND2_X1 U4893 ( .A1(n5979), .A2(n5981), .ZN(n6017) );
  XNOR2_X2 U4894 ( .A(n5975), .B(n8743), .ZN(n5979) );
  AOI21_X1 U4895 ( .B1(n4430), .B2(n4877), .A(n8301), .ZN(n4429) );
  INV_X1 U4896 ( .A(n4431), .ZN(n4430) );
  AOI21_X1 U4897 ( .B1(n4434), .B2(n4436), .A(n8498), .ZN(n4431) );
  OR2_X1 U4898 ( .A1(n6414), .A2(n8030), .ZN(n8349) );
  NAND2_X1 U4900 ( .A1(n4927), .A2(n7725), .ZN(n5071) );
  OAI21_X1 U4901 ( .B1(n5265), .B2(n5264), .A(n5263), .ZN(n5281) );
  NOR2_X1 U4902 ( .A1(n4973), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n4608) );
  NAND3_X1 U4903 ( .A1(n6320), .A2(n5527), .A3(n5526), .ZN(n6747) );
  NOR2_X1 U4904 ( .A1(n5485), .A2(n4818), .ZN(n4816) );
  AND2_X1 U4905 ( .A1(n9199), .A2(n8901), .ZN(n5485) );
  INV_X1 U4906 ( .A(n5015), .ZN(n6560) );
  INV_X1 U4907 ( .A(n7751), .ZN(n5256) );
  NOR2_X1 U4908 ( .A1(n4904), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4894) );
  AND2_X1 U4909 ( .A1(n7358), .A2(n6110), .ZN(n6124) );
  OR2_X1 U4910 ( .A1(n6112), .A2(n8322), .ZN(n6127) );
  NOR2_X1 U4911 ( .A1(n4569), .A2(n6294), .ZN(n4568) );
  INV_X1 U4912 ( .A(n4571), .ZN(n4569) );
  OR2_X1 U4913 ( .A1(n6465), .A2(n6449), .ZN(n7796) );
  INV_X1 U4914 ( .A(n5327), .ZN(n4487) );
  INV_X1 U4915 ( .A(n5179), .ZN(n4682) );
  OR2_X1 U4916 ( .A1(n8679), .A2(n8285), .ZN(n8354) );
  INV_X1 U4917 ( .A(n4439), .ZN(n4436) );
  NOR2_X1 U4918 ( .A1(n8274), .A2(n8344), .ZN(n4439) );
  NAND2_X1 U4919 ( .A1(n6786), .A2(n5600), .ZN(n5603) );
  AOI21_X1 U4920 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n6772), .A(n8442), .ZN(
        n5671) );
  OR2_X1 U4921 ( .A1(n8702), .A2(n8519), .ZN(n6261) );
  OR2_X1 U4922 ( .A1(n8702), .A2(n8541), .ZN(n8310) );
  OR2_X1 U4923 ( .A1(n8719), .A2(n7957), .ZN(n8246) );
  NAND2_X1 U4924 ( .A1(n4859), .A2(n4858), .ZN(n5509) );
  AND2_X1 U4925 ( .A1(n4422), .A2(n4421), .ZN(n4859) );
  AND2_X1 U4926 ( .A1(n4349), .A2(n4863), .ZN(n4770) );
  NAND2_X1 U4927 ( .A1(n7928), .A2(n7146), .ZN(n5943) );
  AOI21_X1 U4928 ( .B1(n4789), .B2(n4787), .A(n4314), .ZN(n4786) );
  INV_X1 U4929 ( .A(n4790), .ZN(n4787) );
  INV_X1 U4930 ( .A(n4789), .ZN(n4788) );
  NAND2_X1 U4931 ( .A1(n9173), .A2(n9036), .ZN(n4794) );
  OR2_X1 U4932 ( .A1(n7086), .A2(n7400), .ZN(n7848) );
  CLKBUF_X1 U4933 ( .A(n4946), .Z(n7834) );
  AND2_X1 U4934 ( .A1(n5435), .A2(n9381), .ZN(n6470) );
  NAND2_X1 U4935 ( .A1(n4464), .A2(n5347), .ZN(n5361) );
  AND2_X1 U4936 ( .A1(n5362), .A2(n5351), .ZN(n5360) );
  AND2_X1 U4937 ( .A1(n5270), .A2(n5269), .ZN(n5280) );
  OAI21_X1 U4938 ( .B1(n5250), .B2(n5249), .A(n5248), .ZN(n5265) );
  AND2_X1 U4939 ( .A1(n5232), .A2(n5218), .ZN(n5230) );
  AOI21_X1 U4940 ( .B1(n4712), .B2(n4710), .A(n4324), .ZN(n4709) );
  NOR2_X1 U4941 ( .A1(n4884), .A2(n4973), .ZN(n5128) );
  NOR2_X1 U4942 ( .A1(n5125), .A2(n4715), .ZN(n4714) );
  INV_X1 U4943 ( .A(n5102), .ZN(n4715) );
  OAI21_X1 U4944 ( .B1(n4941), .B2(n4911), .A(n4910), .ZN(n4939) );
  AND2_X1 U4945 ( .A1(n7137), .A2(n7135), .ZN(n4654) );
  AND2_X1 U4946 ( .A1(n7975), .A2(n8541), .ZN(n7976) );
  NAND2_X1 U4947 ( .A1(n4646), .A2(n4645), .ZN(n7970) );
  NOR2_X1 U4948 ( .A1(n4647), .A2(n4341), .ZN(n4645) );
  INV_X1 U4949 ( .A(n6101), .ZN(n6307) );
  NAND2_X1 U4950 ( .A1(n4733), .A2(n4752), .ZN(n4732) );
  XNOR2_X1 U4951 ( .A(n5990), .B(n5671), .ZN(n8459) );
  NOR2_X1 U4952 ( .A1(n5534), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U4953 ( .A1(n6418), .A2(n6417), .ZN(n8351) );
  AND2_X1 U4954 ( .A1(n6297), .A2(n8027), .ZN(n8487) );
  OR2_X1 U4955 ( .A1(n8291), .A2(n6021), .ZN(n6022) );
  NAND2_X1 U4956 ( .A1(n6321), .A2(n6593), .ZN(n6862) );
  NAND2_X1 U4957 ( .A1(n6757), .A2(n8301), .ZN(n8607) );
  OR2_X1 U4958 ( .A1(n8661), .A2(n8606), .ZN(n8575) );
  NOR2_X1 U4959 ( .A1(n7543), .A2(n4559), .ZN(n4558) );
  INV_X1 U4960 ( .A(n6170), .ZN(n4559) );
  NOR2_X1 U4961 ( .A1(n6745), .A2(n6376), .ZN(n6762) );
  INV_X1 U4962 ( .A(n9861), .ZN(n9872) );
  AND2_X1 U4963 ( .A1(n6747), .A2(n6595), .ZN(n6752) );
  CLKBUF_X1 U4964 ( .A(n5531), .Z(n5558) );
  INV_X1 U4965 ( .A(n4766), .ZN(n4765) );
  INV_X1 U4966 ( .A(n9048), .ZN(n8798) );
  NAND2_X1 U4967 ( .A1(n4394), .A2(n4400), .ZN(n5836) );
  OR2_X1 U4968 ( .A1(n5830), .A2(n4337), .ZN(n4394) );
  NAND2_X1 U4969 ( .A1(n4967), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4902) );
  AND2_X1 U4970 ( .A1(n4899), .A2(n9396), .ZN(n4951) );
  AND2_X1 U4971 ( .A1(n9464), .A2(n9465), .ZN(n9462) );
  NAND2_X1 U4972 ( .A1(n8280), .A2(n5318), .ZN(n4484) );
  NOR2_X1 U4973 ( .A1(n6465), .A2(n4526), .ZN(n4525) );
  INV_X1 U4974 ( .A(n4527), .ZN(n4526) );
  OR2_X1 U4975 ( .A1(n9025), .A2(n9173), .ZN(n9011) );
  NOR2_X1 U4976 ( .A1(n9060), .A2(n7700), .ZN(n9045) );
  OR2_X1 U4977 ( .A1(n9204), .A2(n9125), .ZN(n5483) );
  OR2_X1 U4978 ( .A1(n7201), .A2(n8906), .ZN(n5478) );
  NAND2_X1 U4979 ( .A1(n5131), .A2(n5130), .ZN(n7100) );
  INV_X1 U4980 ( .A(n8912), .ZN(n6956) );
  INV_X2 U4981 ( .A(n6008), .ZN(n7746) );
  NAND2_X1 U4982 ( .A1(n4607), .A2(n4297), .ZN(n4904) );
  NOR2_X1 U4983 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4891) );
  NAND2_X1 U4984 ( .A1(n5235), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U4985 ( .A1(n5368), .A2(n5367), .ZN(n9168) );
  NOR2_X1 U4986 ( .A1(n7641), .A2(n4600), .ZN(n4599) );
  INV_X1 U4987 ( .A(n7840), .ZN(n4600) );
  MUX2_X1 U4988 ( .A(n8161), .B(n8160), .S(n8278), .Z(n8162) );
  AND2_X1 U4989 ( .A1(n8164), .A2(n8316), .ZN(n4460) );
  NAND2_X1 U4990 ( .A1(n4604), .A2(n4601), .ZN(n7654) );
  NAND2_X1 U4991 ( .A1(n4603), .A2(n4602), .ZN(n4601) );
  OR2_X1 U4992 ( .A1(n8203), .A2(n4445), .ZN(n4443) );
  NAND2_X1 U4993 ( .A1(n7667), .A2(n7666), .ZN(n4585) );
  NAND2_X1 U4994 ( .A1(n4589), .A2(n4586), .ZN(n7667) );
  OAI21_X1 U4995 ( .B1(n4588), .B2(n4587), .A(n7888), .ZN(n4586) );
  INV_X1 U4996 ( .A(n4590), .ZN(n4589) );
  INV_X1 U4997 ( .A(n7852), .ZN(n4587) );
  AOI22_X1 U4998 ( .A1(n4450), .A2(n4275), .B1(n4451), .B2(n4316), .ZN(n8248)
         );
  NAND2_X1 U4999 ( .A1(n8235), .A2(n4453), .ZN(n4450) );
  NAND2_X1 U5000 ( .A1(n7708), .A2(n7707), .ZN(n4618) );
  MUX2_X1 U5001 ( .A(n8252), .B(n8251), .S(n8301), .Z(n8258) );
  NOR2_X1 U5002 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4880) );
  INV_X1 U5003 ( .A(n4435), .ZN(n4434) );
  OAI21_X1 U5004 ( .B1(n4436), .B2(n8276), .A(n4326), .ZN(n4435) );
  NAND2_X1 U5005 ( .A1(n4433), .A2(n8301), .ZN(n4432) );
  NAND2_X1 U5006 ( .A1(n4876), .A2(n8286), .ZN(n4433) );
  OR2_X1 U5007 ( .A1(n6109), .A2(n8321), .ZN(n6123) );
  AND2_X1 U5008 ( .A1(n8303), .A2(n7067), .ZN(n6369) );
  AND2_X1 U5009 ( .A1(n5743), .A2(n6907), .ZN(n4370) );
  NAND2_X1 U5010 ( .A1(n4375), .A2(n4377), .ZN(n4373) );
  AND2_X1 U5011 ( .A1(n9643), .A2(n7645), .ZN(n4796) );
  INV_X1 U5012 ( .A(n5471), .ZN(n4799) );
  NOR2_X1 U5013 ( .A1(n8895), .A2(n5177), .ZN(n4539) );
  INV_X1 U5014 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5160) );
  NOR2_X1 U5015 ( .A1(n4711), .A2(n4707), .ZN(n4706) );
  INV_X1 U5016 ( .A(n5082), .ZN(n4707) );
  NAND2_X1 U5017 ( .A1(n4712), .A2(n5138), .ZN(n4711) );
  NAND2_X1 U5018 ( .A1(n5108), .A2(n5107), .ZN(n5124) );
  INV_X1 U5019 ( .A(n5050), .ZN(n4466) );
  OAI21_X1 U5020 ( .B1(n9818), .B2(n5577), .A(n5578), .ZN(n9810) );
  NAND2_X1 U5021 ( .A1(n4743), .A2(n4742), .ZN(n5666) );
  NAND2_X1 U5022 ( .A1(n6600), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4742) );
  NOR2_X1 U5023 ( .A1(n8405), .A2(n4352), .ZN(n5669) );
  NOR2_X1 U5024 ( .A1(n6130), .A2(n7332), .ZN(n6131) );
  NOR2_X1 U5025 ( .A1(n4567), .A2(n4563), .ZN(n4562) );
  INV_X1 U5026 ( .A(n4866), .ZN(n4563) );
  INV_X1 U5027 ( .A(n4568), .ZN(n4567) );
  NAND2_X1 U5028 ( .A1(n4568), .A2(n4566), .ZN(n4565) );
  INV_X1 U5029 ( .A(n4574), .ZN(n4566) );
  NAND2_X1 U5030 ( .A1(n4831), .A2(n8267), .ZN(n4830) );
  INV_X1 U5031 ( .A(n8266), .ZN(n4831) );
  OR2_X1 U5032 ( .A1(n8696), .A2(n8531), .ZN(n8267) );
  NAND2_X1 U5033 ( .A1(n6362), .A2(n4841), .ZN(n4840) );
  NOR2_X1 U5034 ( .A1(n8616), .A2(n4842), .ZN(n4841) );
  NAND3_X1 U5035 ( .A1(n4856), .A2(n4540), .A3(n5592), .ZN(n4853) );
  INV_X1 U5036 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U5037 ( .A1(n4380), .A2(n4379), .ZN(n5858) );
  AOI21_X1 U5038 ( .B1(n4381), .B2(n4382), .A(n4347), .ZN(n4379) );
  NOR2_X1 U5039 ( .A1(n5785), .A2(n4778), .ZN(n4777) );
  INV_X1 U5040 ( .A(n7069), .ZN(n4778) );
  NAND2_X1 U5041 ( .A1(n8754), .A2(n4402), .ZN(n4401) );
  INV_X1 U5042 ( .A(n5829), .ZN(n4402) );
  INV_X1 U5043 ( .A(n7821), .ZN(n4632) );
  INV_X1 U5044 ( .A(n7741), .ZN(n4633) );
  NOR2_X1 U5045 ( .A1(n9563), .A2(n4508), .ZN(n8936) );
  AND2_X1 U5046 ( .A1(n9568), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4508) );
  NOR2_X1 U5047 ( .A1(n9164), .A2(n9157), .ZN(n4527) );
  NAND2_X1 U5048 ( .A1(n4702), .A2(n4700), .ZN(n5416) );
  NAND2_X1 U5049 ( .A1(n4701), .A2(n7798), .ZN(n4700) );
  INV_X1 U5050 ( .A(n4703), .ZN(n4701) );
  INV_X1 U5051 ( .A(n9017), .ZN(n4699) );
  NOR2_X1 U5052 ( .A1(n9033), .A2(n4698), .ZN(n4697) );
  OR2_X1 U5053 ( .A1(n9173), .A2(n5491), .ZN(n7803) );
  NOR2_X1 U5054 ( .A1(n9188), .A2(n9194), .ZN(n4532) );
  NAND2_X1 U5055 ( .A1(n8814), .A2(n4539), .ZN(n4538) );
  NAND2_X1 U5056 ( .A1(n9219), .A2(n8903), .ZN(n4814) );
  OR2_X1 U5057 ( .A1(n9219), .A2(n9143), .ZN(n7858) );
  NOR2_X1 U5058 ( .A1(n8895), .A2(n8904), .ZN(n4810) );
  NAND2_X1 U5059 ( .A1(n9743), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U5060 ( .A1(n7098), .A2(n5500), .ZN(n7254) );
  AND2_X1 U5061 ( .A1(n5942), .A2(n5456), .ZN(n6471) );
  OAI21_X1 U5062 ( .B1(n7724), .B2(SI_29_), .A(n7723), .ZN(n7743) );
  NAND2_X1 U5063 ( .A1(n4820), .A2(n4514), .ZN(n4819) );
  NOR2_X1 U5064 ( .A1(n4821), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4820) );
  INV_X1 U5065 ( .A(n4890), .ZN(n4514) );
  NAND2_X1 U5066 ( .A1(n4463), .A2(n5362), .ZN(n5376) );
  AND2_X1 U5067 ( .A1(n5377), .A2(n5366), .ZN(n5375) );
  NAND2_X1 U5068 ( .A1(n5408), .A2(n5407), .ZN(n5429) );
  AOI21_X1 U5069 ( .B1(n4488), .B2(n4491), .A(n4487), .ZN(n4486) );
  AND2_X1 U5070 ( .A1(n5347), .A2(n5334), .ZN(n5345) );
  INV_X1 U5071 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5450) );
  INV_X1 U5072 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U5073 ( .A1(n4474), .A2(n4472), .ZN(n5250) );
  AOI21_X1 U5074 ( .B1(n4476), .B2(n4479), .A(n4473), .ZN(n4472) );
  INV_X1 U5075 ( .A(n5232), .ZN(n4473) );
  OR2_X1 U5076 ( .A1(n5051), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5085) );
  NOR2_X2 U5077 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4936) );
  XNOR2_X1 U5078 ( .A(n4939), .B(SI_1_), .ZN(n4937) );
  INV_X1 U5079 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4661) );
  INV_X1 U5080 ( .A(n8387), .ZN(n7516) );
  INV_X1 U5081 ( .A(n4654), .ZN(n4653) );
  INV_X1 U5082 ( .A(n7303), .ZN(n7916) );
  AND2_X1 U5083 ( .A1(n4298), .A2(n7954), .ZN(n4648) );
  NAND2_X1 U5084 ( .A1(n7938), .A2(n7992), .ZN(n7995) );
  OAI21_X1 U5085 ( .B1(n8351), .B2(n8350), .A(n8357), .ZN(n4852) );
  AND2_X1 U5086 ( .A1(n8353), .A2(n4877), .ZN(n8357) );
  OR2_X1 U5087 ( .A1(n8358), .A2(n4851), .ZN(n4850) );
  NOR2_X1 U5088 ( .A1(n8305), .A2(n4345), .ZN(n4851) );
  NOR2_X1 U5089 ( .A1(n8290), .A2(n8289), .ZN(n8364) );
  NAND2_X1 U5090 ( .A1(n4426), .A2(n4423), .ZN(n8290) );
  AOI21_X1 U5091 ( .B1(n8275), .B2(n8276), .A(n4436), .ZN(n8288) );
  NAND3_X1 U5092 ( .A1(n5549), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n5547) );
  AND4_X1 U5093 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n7282)
         );
  OR2_X1 U5094 ( .A1(n4271), .A2(n9273), .ZN(n6091) );
  OR2_X1 U5095 ( .A1(n5584), .A2(n6546), .ZN(n5585) );
  INV_X1 U5096 ( .A(n4731), .ZN(n4730) );
  NAND2_X1 U5097 ( .A1(n9848), .A2(n5651), .ZN(n5652) );
  NAND2_X1 U5098 ( .A1(n4748), .A2(n4747), .ZN(n4746) );
  OR2_X1 U5099 ( .A1(n5603), .A2(n6552), .ZN(n5604) );
  NAND2_X1 U5100 ( .A1(n5656), .A2(n6552), .ZN(n6499) );
  OR2_X1 U5101 ( .A1(n7607), .A2(n7606), .ZN(n4743) );
  AOI21_X1 U5102 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6600), .A(n7593), .ZN(
        n5619) );
  XNOR2_X1 U5103 ( .A(n5669), .B(n8417), .ZN(n8425) );
  NOR2_X1 U5104 ( .A1(n8425), .A2(n8424), .ZN(n8423) );
  AOI21_X1 U5105 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6653), .A(n8395), .ZN(
        n5622) );
  NOR2_X1 U5106 ( .A1(n5628), .A2(n8451), .ZN(n8481) );
  OR2_X1 U5107 ( .A1(n8668), .A2(n8074), .ZN(n8593) );
  AOI21_X1 U5108 ( .B1(n4545), .B2(n4544), .A(n4315), .ZN(n4543) );
  INV_X1 U5109 ( .A(n4550), .ZN(n4544) );
  AND4_X1 U5110 ( .A1(n5988), .A2(n5987), .A3(n5986), .A4(n5985), .ZN(n8604)
         );
  NOR2_X1 U5111 ( .A1(n4552), .A2(n4551), .ZN(n4550) );
  INV_X1 U5112 ( .A(n8621), .ZN(n4551) );
  NAND2_X1 U5113 ( .A1(n8622), .A2(n4549), .ZN(n4548) );
  INV_X1 U5114 ( .A(n4552), .ZN(n4549) );
  OR2_X1 U5115 ( .A1(n8053), .A2(n8139), .ZN(n8231) );
  NAND2_X1 U5116 ( .A1(n7324), .A2(n6150), .ZN(n7437) );
  NAND2_X1 U5117 ( .A1(n7210), .A2(n8327), .ZN(n4849) );
  NAND3_X1 U5118 ( .A1(n4556), .A2(n4554), .A3(n4557), .ZN(n7324) );
  NOR2_X1 U5119 ( .A1(n8209), .A2(n4555), .ZN(n4554) );
  OAI211_X1 U5120 ( .C1(n6391), .C2(n6390), .A(n6389), .B(n6388), .ZN(n6396)
         );
  NOR2_X1 U5121 ( .A1(n4313), .A2(n4572), .ZN(n4571) );
  NOR2_X1 U5122 ( .A1(n6283), .A2(n4573), .ZN(n4572) );
  NAND2_X1 U5123 ( .A1(n6272), .A2(n6273), .ZN(n4573) );
  NOR2_X1 U5124 ( .A1(n6283), .A2(n4575), .ZN(n4574) );
  INV_X1 U5125 ( .A(n6272), .ZN(n4575) );
  OR2_X1 U5126 ( .A1(n8696), .A2(n8381), .ZN(n6272) );
  INV_X1 U5127 ( .A(n8267), .ZN(n4832) );
  INV_X1 U5128 ( .A(n8341), .ZN(n8505) );
  AND2_X1 U5129 ( .A1(n6264), .A2(n6263), .ZN(n7977) );
  NAND2_X1 U5130 ( .A1(n4834), .A2(n8255), .ZN(n4833) );
  AND2_X1 U5131 ( .A1(n8310), .A2(n8309), .ZN(n8529) );
  OR2_X1 U5132 ( .A1(n8713), .A2(n8567), .ZN(n6239) );
  INV_X1 U5133 ( .A(n9858), .ZN(n8605) );
  OR2_X1 U5134 ( .A1(n8713), .A2(n8542), .ZN(n8253) );
  NAND2_X1 U5135 ( .A1(n8550), .A2(n8254), .ZN(n4837) );
  OAI21_X1 U5136 ( .B1(n8562), .B2(n8552), .A(n8551), .ZN(n8554) );
  NAND2_X1 U5137 ( .A1(n4840), .A2(n8234), .ZN(n8598) );
  AND2_X1 U5138 ( .A1(n8236), .A2(n8234), .ZN(n8622) );
  AND2_X1 U5139 ( .A1(n8231), .A2(n8230), .ZN(n8335) );
  NAND2_X1 U5140 ( .A1(n7524), .A2(n6169), .ZN(n4560) );
  NAND2_X1 U5141 ( .A1(n6358), .A2(n8219), .ZN(n7545) );
  INV_X1 U5142 ( .A(n8607), .ZN(n9859) );
  AND2_X1 U5143 ( .A1(n6871), .A2(n8301), .ZN(n9858) );
  NAND2_X1 U5144 ( .A1(n4582), .A2(n4581), .ZN(n5976) );
  NOR2_X1 U5145 ( .A1(n4872), .A2(n4843), .ZN(n4581) );
  INV_X1 U5146 ( .A(n5528), .ZN(n4582) );
  NAND2_X1 U5147 ( .A1(n4844), .A2(n5973), .ZN(n4843) );
  XNOR2_X1 U5148 ( .A(n5542), .B(n5973), .ZN(n5640) );
  NAND2_X1 U5149 ( .A1(n4290), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5542) );
  AND2_X1 U5150 ( .A1(n5521), .A2(n5520), .ZN(n6320) );
  INV_X1 U5151 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4462) );
  INV_X1 U5152 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5565) );
  NOR2_X1 U5153 ( .A1(n5611), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5569) );
  INV_X1 U5154 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5592) );
  INV_X1 U5155 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5579) );
  XNOR2_X1 U5156 ( .A(n5797), .B(n5795), .ZN(n7184) );
  INV_X1 U5157 ( .A(n5796), .ZN(n5795) );
  INV_X1 U5158 ( .A(n4764), .ZN(n4763) );
  OAI21_X1 U5159 ( .B1(n4287), .B2(n4765), .A(n7396), .ZN(n4764) );
  NAND2_X1 U5160 ( .A1(n4273), .A2(n4310), .ZN(n4766) );
  INV_X1 U5161 ( .A(n5900), .ZN(n5901) );
  OAI21_X1 U5162 ( .B1(n5899), .B2(n5898), .A(n5897), .ZN(n5900) );
  NAND2_X1 U5163 ( .A1(n8822), .A2(n8824), .ZN(n8823) );
  NAND2_X1 U5164 ( .A1(n7184), .A2(n7183), .ZN(n7182) );
  AOI21_X1 U5165 ( .B1(n4769), .B2(n4404), .A(n4403), .ZN(n8763) );
  NOR2_X1 U5166 ( .A1(n4283), .A2(n4771), .ZN(n4404) );
  INV_X1 U5167 ( .A(n8761), .ZN(n4403) );
  INV_X1 U5168 ( .A(n5895), .ZN(n8762) );
  OAI21_X1 U5169 ( .B1(n8822), .B2(n5906), .A(n4772), .ZN(n8871) );
  INV_X1 U5170 ( .A(n4773), .ZN(n4772) );
  OAI21_X1 U5171 ( .B1(n8824), .B2(n5906), .A(n8795), .ZN(n4773) );
  OR2_X1 U5172 ( .A1(n4337), .A2(n5835), .ZN(n4399) );
  OR2_X1 U5173 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  NOR2_X1 U5174 ( .A1(n4401), .A2(n5835), .ZN(n4396) );
  AND2_X1 U5175 ( .A1(n4401), .A2(n5835), .ZN(n4400) );
  NAND2_X1 U5176 ( .A1(n5429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U5177 ( .A1(n5455), .A2(n5454), .ZN(n5730) );
  AND2_X1 U5178 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  AND2_X1 U5179 ( .A1(n6621), .A2(n4418), .ZN(n9468) );
  OR2_X1 U5180 ( .A1(n6618), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4418) );
  NOR2_X1 U5181 ( .A1(n9462), .A2(n4296), .ZN(n9426) );
  OR2_X1 U5182 ( .A1(n9426), .A2(n9427), .ZN(n4502) );
  OR2_X1 U5183 ( .A1(n9506), .A2(n9507), .ZN(n4413) );
  OR2_X1 U5184 ( .A1(n9502), .A2(n9503), .ZN(n4506) );
  NAND2_X1 U5185 ( .A1(n4413), .A2(n4412), .ZN(n4411) );
  NAND2_X1 U5186 ( .A1(n6630), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4412) );
  AND2_X1 U5187 ( .A1(n4411), .A2(n4410), .ZN(n9520) );
  INV_X1 U5188 ( .A(n9522), .ZN(n4410) );
  AND2_X1 U5189 ( .A1(n4506), .A2(n4505), .ZN(n9517) );
  NAND2_X1 U5190 ( .A1(n6630), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4505) );
  OR2_X1 U5191 ( .A1(n9517), .A2(n9518), .ZN(n4504) );
  NOR2_X1 U5192 ( .A1(n9401), .A2(n4511), .ZN(n9533) );
  AND2_X1 U5193 ( .A1(n9406), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4511) );
  AOI21_X1 U5194 ( .B1(n9406), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9398), .ZN(
        n9537) );
  AOI21_X1 U5195 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9568), .A(n9560), .ZN(
        n8927) );
  NAND2_X1 U5196 ( .A1(n8929), .A2(n4406), .ZN(n8954) );
  INV_X1 U5197 ( .A(n8932), .ZN(n4406) );
  OR2_X1 U5198 ( .A1(n8941), .A2(n8940), .ZN(n8948) );
  NAND2_X1 U5199 ( .A1(n5416), .A2(n7761), .ZN(n5415) );
  NOR2_X1 U5200 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  INV_X1 U5201 ( .A(n5490), .ZN(n4791) );
  INV_X1 U5202 ( .A(n4794), .ZN(n4792) );
  NAND2_X1 U5203 ( .A1(n4329), .A2(n4794), .ZN(n4789) );
  OR2_X1 U5204 ( .A1(n9188), .A2(n9047), .ZN(n5487) );
  AND3_X1 U5205 ( .A1(n4673), .A2(n4671), .A3(n4672), .ZN(n9060) );
  OR2_X1 U5206 ( .A1(n9120), .A2(n9144), .ZN(n4867) );
  AOI21_X1 U5207 ( .B1(n4813), .B2(n4804), .A(n4802), .ZN(n9116) );
  AND2_X1 U5208 ( .A1(n4807), .A2(n5480), .ZN(n4804) );
  OAI21_X1 U5209 ( .B1(n4805), .B2(n4803), .A(n4320), .ZN(n4802) );
  INV_X1 U5210 ( .A(n5480), .ZN(n4803) );
  NAND2_X1 U5211 ( .A1(n4806), .A2(n4814), .ZN(n4805) );
  INV_X1 U5212 ( .A(n4809), .ZN(n4806) );
  AND2_X1 U5213 ( .A1(n4812), .A2(n4814), .ZN(n4807) );
  NAND2_X1 U5214 ( .A1(n4687), .A2(n4686), .ZN(n7372) );
  NAND2_X1 U5215 ( .A1(n4692), .A2(n7669), .ZN(n4686) );
  NAND3_X1 U5216 ( .A1(n4689), .A2(n7669), .A3(n4688), .ZN(n4687) );
  NAND2_X1 U5217 ( .A1(n7671), .A2(n7858), .ZN(n7371) );
  NOR2_X1 U5218 ( .A1(n7782), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U5219 ( .A1(n4813), .A2(n4812), .ZN(n4811) );
  INV_X1 U5220 ( .A(n4810), .ZN(n4808) );
  INV_X1 U5221 ( .A(n7371), .ZN(n7782) );
  NOR2_X1 U5222 ( .A1(n9769), .A2(n7928), .ZN(n6469) );
  AOI21_X1 U5223 ( .B1(n7091), .B2(n7093), .A(n4317), .ZN(n7195) );
  OAI21_X1 U5224 ( .B1(n7077), .B2(n7776), .A(n4795), .ZN(n7091) );
  OR2_X1 U5225 ( .A1(n7086), .A2(n8907), .ZN(n4795) );
  AND2_X1 U5226 ( .A1(n7776), .A2(n7655), .ZN(n5122) );
  NAND2_X1 U5227 ( .A1(n5090), .A2(n5089), .ZN(n5476) );
  NOR2_X1 U5228 ( .A1(n9631), .A2(n4522), .ZN(n7085) );
  OR2_X1 U5229 ( .A1(n9630), .A2(n7181), .ZN(n9631) );
  NAND2_X1 U5230 ( .A1(n4999), .A2(n7840), .ZN(n7639) );
  NOR2_X1 U5231 ( .A1(n4625), .A2(n4965), .ZN(n4622) );
  INV_X1 U5232 ( .A(n4947), .ZN(n4625) );
  NAND2_X1 U5233 ( .A1(n5461), .A2(n7838), .ZN(n7764) );
  OR2_X1 U5234 ( .A1(n7823), .A2(n9473), .ZN(n9616) );
  INV_X1 U5235 ( .A(n9655), .ZN(n9138) );
  OR2_X1 U5236 ( .A1(n5727), .A2(n7928), .ZN(n6905) );
  INV_X1 U5237 ( .A(n9616), .ZN(n9652) );
  INV_X1 U5238 ( .A(n9769), .ZN(n9666) );
  NAND2_X1 U5239 ( .A1(n5283), .A2(n5282), .ZN(n9199) );
  NAND2_X1 U5240 ( .A1(n7757), .A2(n5494), .ZN(n9655) );
  NAND2_X1 U5241 ( .A1(n5433), .A2(n5453), .ZN(n9379) );
  XNOR2_X1 U5242 ( .A(n7743), .B(n7742), .ZN(n8280) );
  XNOR2_X1 U5243 ( .A(n6407), .B(n6406), .ZN(n7591) );
  NAND2_X1 U5244 ( .A1(n4494), .A2(n5296), .ZN(n5313) );
  NAND2_X1 U5245 ( .A1(n5271), .A2(n4495), .ZN(n4494) );
  AND3_X1 U5246 ( .A1(n5128), .A2(n4336), .A3(n4779), .ZN(n5411) );
  NAND2_X1 U5247 ( .A1(n4885), .A2(n4781), .ZN(n4780) );
  AND2_X1 U5248 ( .A1(n5405), .A2(n5404), .ZN(n4386) );
  NAND2_X1 U5249 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4389), .ZN(n4388) );
  NAND2_X1 U5250 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n4389) );
  NAND2_X1 U5251 ( .A1(n5219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U5252 ( .A1(n4405), .A2(n4782), .ZN(n5219) );
  INV_X1 U5253 ( .A(n5143), .ZN(n4405) );
  NAND2_X1 U5254 ( .A1(n4475), .A2(n4480), .ZN(n5231) );
  NAND2_X1 U5255 ( .A1(n5197), .A2(n4482), .ZN(n4475) );
  OAI21_X1 U5256 ( .B1(n5197), .B2(n5196), .A(n5195), .ZN(n5213) );
  OAI211_X1 U5257 ( .C1(n5159), .C2(n4680), .A(n4677), .B(n4676), .ZN(n6675)
         );
  AOI21_X1 U5258 ( .B1(n4679), .B2(n4681), .A(n4292), .ZN(n4676) );
  INV_X1 U5259 ( .A(n4681), .ZN(n4680) );
  INV_X1 U5260 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5165) );
  XNOR2_X1 U5261 ( .A(n5181), .B(n5180), .ZN(n6651) );
  NAND2_X1 U5262 ( .A1(n4708), .A2(n4712), .ZN(n5142) );
  NAND2_X1 U5263 ( .A1(n5104), .A2(n4714), .ZN(n4708) );
  INV_X4 U5264 ( .A(n6008), .ZN(n7725) );
  XNOR2_X1 U5265 ( .A(n5025), .B(SI_6_), .ZN(n5023) );
  NAND2_X1 U5266 ( .A1(n5010), .A2(n5009), .ZN(n5014) );
  AND2_X1 U5267 ( .A1(n5072), .A2(n5020), .ZN(n6633) );
  INV_X1 U5268 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U5269 ( .A1(n7136), .A2(n4654), .ZN(n7238) );
  NAND2_X1 U5270 ( .A1(n4638), .A2(n4641), .ZN(n4634) );
  AOI21_X1 U5271 ( .B1(n4640), .B2(n4638), .A(n4637), .ZN(n4636) );
  NAND2_X1 U5272 ( .A1(n7983), .A2(n7984), .ZN(n8023) );
  INV_X1 U5273 ( .A(n8519), .ZN(n8541) );
  AOI21_X1 U5274 ( .B1(n8080), .B2(n8081), .A(n7976), .ZN(n8046) );
  OR2_X1 U5275 ( .A1(n6017), .A2(n9813), .ZN(n5997) );
  AND4_X1 U5276 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n8606)
         );
  AND2_X1 U5277 ( .A1(n6766), .A2(n6765), .ZN(n8132) );
  INV_X1 U5278 ( .A(n7067), .ZN(n8368) );
  XNOR2_X1 U5279 ( .A(n5619), .B(n7561), .ZN(n7559) );
  OR2_X1 U5280 ( .A1(n7559), .A2(n7560), .ZN(n4728) );
  OAI21_X1 U5281 ( .B1(n7559), .B2(n4726), .A(n4725), .ZN(n8395) );
  NAND2_X1 U5282 ( .A1(n4729), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4726) );
  NAND2_X1 U5283 ( .A1(n5620), .A2(n4729), .ZN(n4725) );
  INV_X1 U5284 ( .A(n8396), .ZN(n4729) );
  NOR2_X1 U5285 ( .A1(n8486), .A2(n8485), .ZN(n4740) );
  NAND2_X1 U5286 ( .A1(n5558), .A2(n4461), .ZN(n5629) );
  AOI21_X1 U5287 ( .B1(n4276), .B2(n9827), .A(n4365), .ZN(n5724) );
  NOR2_X1 U5288 ( .A1(n8469), .A2(n5674), .ZN(n5675) );
  AND2_X1 U5289 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  NAND2_X1 U5290 ( .A1(n6432), .A2(n6431), .ZN(n6433) );
  NOR2_X1 U5291 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  OR2_X1 U5292 ( .A1(n6764), .A2(n6743), .ZN(n6381) );
  INV_X1 U5293 ( .A(n7201), .ZN(n5500) );
  AND2_X1 U5294 ( .A1(n5963), .A2(n5952), .ZN(n8876) );
  AND2_X1 U5295 ( .A1(n5965), .A2(n5417), .ZN(n8887) );
  INV_X1 U5296 ( .A(n7146), .ZN(n7895) );
  NAND4_X1 U5297 ( .A1(n4972), .A2(n4971), .A3(n4970), .A4(n4969), .ZN(n8912)
         );
  NAND3_X1 U5298 ( .A1(n4954), .A2(n4953), .A3(n4952), .ZN(n5754) );
  OR2_X1 U5299 ( .A1(n5287), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4952) );
  AND2_X1 U5300 ( .A1(n4950), .A2(n4949), .ZN(n4954) );
  NAND4_X1 U5301 ( .A1(n4935), .A2(n4934), .A3(n4933), .A4(n4932), .ZN(n6911)
         );
  NAND2_X1 U5302 ( .A1(n4966), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4934) );
  NAND2_X1 U5303 ( .A1(n4966), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4903) );
  OR2_X1 U5304 ( .A1(n6641), .A2(n9473), .ZN(n9543) );
  NAND2_X1 U5305 ( .A1(n9589), .A2(n9590), .ZN(n9588) );
  NAND2_X1 U5306 ( .A1(n8948), .A2(n4509), .ZN(n9585) );
  AND2_X1 U5307 ( .A1(n9587), .A2(n8947), .ZN(n4509) );
  XNOR2_X1 U5308 ( .A(n4415), .B(n4414), .ZN(n8960) );
  INV_X1 U5309 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n4414) );
  NAND2_X1 U5310 ( .A1(n9607), .A2(n8957), .ZN(n4415) );
  AOI21_X1 U5311 ( .B1(n9383), .B2(n5318), .A(n7752), .ZN(n9154) );
  NAND2_X1 U5312 ( .A1(n8998), .A2(n4525), .ZN(n8976) );
  INV_X1 U5313 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4892) );
  NOR2_X1 U5314 ( .A1(n4606), .A2(n4594), .ZN(n4593) );
  NAND2_X1 U5315 ( .A1(n4599), .A2(n7753), .ZN(n4594) );
  OAI211_X1 U5316 ( .C1(n4999), .C2(n4598), .A(n7642), .B(n4591), .ZN(n4603)
         );
  NAND2_X1 U5317 ( .A1(n4592), .A2(n7768), .ZN(n4591) );
  INV_X1 U5318 ( .A(n4599), .ZN(n4592) );
  AND2_X1 U5319 ( .A1(n4458), .A2(n4459), .ZN(n8169) );
  AOI21_X1 U5320 ( .B1(n8162), .B2(n4460), .A(n4325), .ZN(n4459) );
  AOI21_X1 U5321 ( .B1(n7651), .B2(n7658), .A(n7888), .ZN(n4590) );
  OAI211_X1 U5322 ( .C1(n7650), .C2(n7649), .A(n7656), .B(n7852), .ZN(n7651)
         );
  NOR2_X1 U5323 ( .A1(n7660), .A2(n7659), .ZN(n4588) );
  AND2_X1 U5324 ( .A1(n4441), .A2(n4334), .ZN(n4440) );
  NAND2_X1 U5325 ( .A1(n7672), .A2(n7671), .ZN(n4629) );
  AOI21_X1 U5326 ( .B1(n4585), .B2(n4688), .A(n4584), .ZN(n7670) );
  NAND2_X1 U5327 ( .A1(n7661), .A2(n7859), .ZN(n4584) );
  NAND2_X1 U5328 ( .A1(n4626), .A2(n9130), .ZN(n7682) );
  NAND2_X1 U5329 ( .A1(n4628), .A2(n4627), .ZN(n4626) );
  AOI21_X1 U5330 ( .B1(n7673), .B2(n7753), .A(n7676), .ZN(n4627) );
  NAND2_X1 U5331 ( .A1(n4629), .A2(n7888), .ZN(n4628) );
  AND2_X1 U5332 ( .A1(n8243), .A2(n4457), .ZN(n4453) );
  AND2_X1 U5333 ( .A1(n8575), .A2(n8593), .ZN(n4457) );
  NAND2_X1 U5334 ( .A1(n4456), .A2(n8278), .ZN(n4455) );
  INV_X1 U5335 ( .A(n8240), .ZN(n4456) );
  OR2_X1 U5336 ( .A1(n8241), .A2(n8301), .ZN(n4452) );
  OAI21_X1 U5337 ( .B1(n8248), .B2(n8247), .A(n4454), .ZN(n8250) );
  AND2_X1 U5338 ( .A1(n8246), .A2(n8245), .ZN(n4454) );
  INV_X1 U5339 ( .A(n7711), .ZN(n4615) );
  NAND2_X1 U5340 ( .A1(n4618), .A2(n4617), .ZN(n4616) );
  NAND2_X1 U5341 ( .A1(n8310), .A2(n4836), .ZN(n4448) );
  INV_X1 U5342 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5507) );
  INV_X1 U5343 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U5344 ( .A1(n7715), .A2(n7803), .ZN(n4614) );
  OR2_X1 U5345 ( .A1(n4611), .A2(n7713), .ZN(n4610) );
  NOR2_X1 U5346 ( .A1(n7717), .A2(n4612), .ZN(n4611) );
  INV_X1 U5347 ( .A(n7714), .ZN(n4612) );
  NOR2_X1 U5348 ( .A1(n7717), .A2(n7712), .ZN(n4613) );
  AOI21_X1 U5349 ( .B1(n4480), .B2(n4478), .A(n4477), .ZN(n4476) );
  INV_X1 U5350 ( .A(n5230), .ZN(n4477) );
  INV_X1 U5351 ( .A(n4482), .ZN(n4478) );
  INV_X1 U5352 ( .A(n4480), .ZN(n4479) );
  NOR2_X1 U5353 ( .A1(n5180), .A2(n4685), .ZN(n4684) );
  INV_X1 U5354 ( .A(n5158), .ZN(n4685) );
  NAND2_X1 U5355 ( .A1(n5162), .A2(n5161), .ZN(n5179) );
  NOR2_X1 U5356 ( .A1(n4714), .A2(n5141), .ZN(n4710) );
  NOR2_X1 U5357 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4882) );
  NOR2_X1 U5358 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4881) );
  INV_X1 U5359 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4663) );
  INV_X1 U5360 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4664) );
  AOI21_X1 U5361 ( .B1(n4429), .B2(n4425), .A(n4424), .ZN(n4423) );
  NAND2_X1 U5362 ( .A1(n4434), .A2(n4877), .ZN(n4425) );
  NOR2_X1 U5363 ( .A1(n4309), .A2(n4432), .ZN(n4424) );
  OAI21_X1 U5364 ( .B1(n4429), .B2(n4428), .A(n4427), .ZN(n4426) );
  NOR2_X1 U5365 ( .A1(n4432), .A2(n4436), .ZN(n4428) );
  INV_X1 U5366 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U5367 ( .A1(n4368), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9816) );
  INV_X1 U5368 ( .A(n9814), .ZN(n4368) );
  NAND2_X1 U5369 ( .A1(n4732), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5370 ( .A1(n4828), .A2(n4286), .ZN(n4825) );
  OR2_X1 U5371 ( .A1(n6163), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6173) );
  NOR2_X1 U5372 ( .A1(n9920), .A2(n8387), .ZN(n4555) );
  AND2_X1 U5373 ( .A1(n6122), .A2(n7272), .ZN(n6132) );
  AND2_X1 U5374 ( .A1(n7334), .A2(n8202), .ZN(n6122) );
  NAND2_X1 U5375 ( .A1(n6128), .A2(n6127), .ZN(n7336) );
  NOR2_X1 U5376 ( .A1(n6126), .A2(n6125), .ZN(n6128) );
  INV_X1 U5377 ( .A(n6123), .ZN(n6126) );
  AND2_X1 U5378 ( .A1(n8323), .A2(n6113), .ZN(n7334) );
  AND2_X1 U5379 ( .A1(n6123), .A2(n6127), .ZN(n6113) );
  NAND2_X1 U5380 ( .A1(n7916), .A2(n6111), .ZN(n8192) );
  INV_X1 U5381 ( .A(n6862), .ZN(n6391) );
  INV_X1 U5382 ( .A(n8518), .ZN(n7979) );
  AND2_X1 U5383 ( .A1(n6179), .A2(n7544), .ZN(n8333) );
  NAND2_X1 U5384 ( .A1(n5516), .A2(n4846), .ZN(n4845) );
  INV_X1 U5385 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5516) );
  INV_X1 U5386 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U5387 ( .A1(n5549), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5519) );
  INV_X1 U5388 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5510) );
  OR2_X1 U5389 ( .A1(n5606), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5611) );
  INV_X1 U5390 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4657) );
  INV_X1 U5391 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5506) );
  OAI211_X1 U5392 ( .C1(n4376), .C2(n5746), .A(n4374), .B(n4371), .ZN(n5736)
         );
  NAND2_X1 U5393 ( .A1(n4377), .A2(n5731), .ZN(n4376) );
  NAND2_X1 U5394 ( .A1(n5746), .A2(n4370), .ZN(n4374) );
  NOR2_X1 U5395 ( .A1(n4771), .A2(n4283), .ZN(n4768) );
  NAND2_X1 U5396 ( .A1(n5321), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U5397 ( .A1(n5337), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5354) );
  INV_X1 U5398 ( .A(n5339), .ZN(n5337) );
  NOR2_X1 U5399 ( .A1(n7804), .A2(n4670), .ZN(n4675) );
  NOR2_X1 U5400 ( .A1(n7683), .A2(n9109), .ZN(n4670) );
  INV_X1 U5401 ( .A(n5322), .ZN(n5321) );
  OR2_X1 U5402 ( .A1(n5223), .A2(n5222), .ZN(n5241) );
  NAND2_X1 U5403 ( .A1(n7781), .A2(n7661), .ZN(n4692) );
  INV_X1 U5404 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5170) );
  INV_X1 U5405 ( .A(n7779), .ZN(n5178) );
  INV_X1 U5406 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5147) );
  OR2_X1 U5407 ( .A1(n5148), .A2(n5147), .ZN(n5171) );
  INV_X1 U5408 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5091) );
  AOI21_X1 U5409 ( .B1(n7645), .B2(n4799), .A(n4312), .ZN(n4798) );
  NAND2_X1 U5410 ( .A1(n9683), .A2(n6671), .ZN(n4517) );
  INV_X1 U5411 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9238) );
  INV_X1 U5412 ( .A(SI_15_), .ZN(n9300) );
  NOR2_X1 U5413 ( .A1(n9100), .A2(n9199), .ZN(n9091) );
  NOR2_X1 U5414 ( .A1(n7254), .A2(n4537), .ZN(n7375) );
  INV_X1 U5415 ( .A(n4539), .ZN(n4537) );
  NAND2_X1 U5416 ( .A1(n4272), .A2(n4516), .ZN(n9664) );
  NOR2_X1 U5417 ( .A1(n7834), .A2(n4517), .ZN(n6822) );
  CLKBUF_X1 U5418 ( .A(n4929), .Z(n6907) );
  AND2_X1 U5419 ( .A1(n7744), .A2(n7729), .ZN(n7742) );
  NAND2_X1 U5420 ( .A1(n5376), .A2(n5375), .ZN(n5378) );
  AND2_X1 U5421 ( .A1(n5392), .A2(n5382), .ZN(n5390) );
  NOR2_X1 U5422 ( .A1(n5312), .A2(n4493), .ZN(n4492) );
  INV_X1 U5423 ( .A(n5296), .ZN(n4493) );
  NOR2_X1 U5424 ( .A1(n5297), .A2(n4496), .ZN(n4495) );
  INV_X1 U5425 ( .A(n5270), .ZN(n4496) );
  INV_X1 U5426 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5406) );
  AND2_X1 U5427 ( .A1(n4483), .A2(n5195), .ZN(n4482) );
  INV_X1 U5428 ( .A(n5212), .ZN(n4483) );
  AOI21_X1 U5429 ( .B1(n5196), .B2(n4482), .A(n4481), .ZN(n4480) );
  INV_X1 U5430 ( .A(n5211), .ZN(n4481) );
  NOR2_X1 U5431 ( .A1(n4679), .A2(n5196), .ZN(n4678) );
  INV_X1 U5432 ( .A(n4684), .ZN(n4679) );
  NOR2_X1 U5433 ( .A1(n5193), .A2(n4682), .ZN(n4681) );
  INV_X1 U5434 ( .A(n4884), .ZN(n4609) );
  INV_X1 U5435 ( .A(n5124), .ZN(n4713) );
  NAND2_X1 U5436 ( .A1(n5083), .A2(n5082), .ZN(n5104) );
  OAI211_X1 U5437 ( .C1(n4470), .C2(n4469), .A(n5034), .B(n4468), .ZN(n5081)
         );
  INV_X1 U5438 ( .A(n4469), .ZN(n4465) );
  NAND2_X1 U5439 ( .A1(n4466), .A2(n5029), .ZN(n4469) );
  OR3_X1 U5440 ( .A1(n5039), .A2(P1_IR_REG_7__SCAN_IN), .A3(
        P1_IR_REG_6__SCAN_IN), .ZN(n5051) );
  NOR2_X1 U5441 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4369) );
  INV_X1 U5442 ( .A(n8125), .ZN(n4637) );
  INV_X1 U5443 ( .A(n8385), .ZN(n7999) );
  INV_X1 U5444 ( .A(n6992), .ZN(n6885) );
  NAND2_X1 U5445 ( .A1(n4651), .A2(n4650), .ZN(n7937) );
  AND2_X1 U5446 ( .A1(n7624), .A2(n7620), .ZN(n4650) );
  INV_X1 U5447 ( .A(n8388), .ZN(n8197) );
  OR2_X1 U5448 ( .A1(n6197), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6208) );
  INV_X1 U5449 ( .A(n7978), .ZN(n4642) );
  AND2_X1 U5450 ( .A1(n8300), .A2(n8299), .ZN(n8490) );
  AND3_X1 U5451 ( .A1(n6231), .A2(n6230), .A3(n6229), .ZN(n7957) );
  NAND4_X1 U5452 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n7303)
         );
  OR2_X1 U5453 ( .A1(n9810), .A2(n9809), .ZN(n9812) );
  NAND2_X1 U5454 ( .A1(n9816), .A2(n5646), .ZN(n6692) );
  NAND2_X1 U5455 ( .A1(n9812), .A2(n5578), .ZN(n6695) );
  NAND2_X1 U5456 ( .A1(n4735), .A2(n9832), .ZN(n9837) );
  NAND2_X1 U5457 ( .A1(n4736), .A2(n9833), .ZN(n4735) );
  NAND2_X1 U5458 ( .A1(n4737), .A2(n5585), .ZN(n9835) );
  NOR2_X1 U5459 ( .A1(n4734), .A2(n9869), .ZN(n4737) );
  INV_X1 U5460 ( .A(n9833), .ZN(n4734) );
  NAND2_X1 U5461 ( .A1(n4753), .A2(n6781), .ZN(n6710) );
  NAND2_X1 U5462 ( .A1(n4752), .A2(n9941), .ZN(n4751) );
  NAND2_X1 U5463 ( .A1(n4364), .A2(n6781), .ZN(n6783) );
  NAND2_X1 U5464 ( .A1(n4746), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4745) );
  AND2_X1 U5465 ( .A1(n7116), .A2(n5614), .ZN(n7221) );
  AND2_X1 U5466 ( .A1(n7109), .A2(n5660), .ZN(n7218) );
  NOR2_X1 U5467 ( .A1(n7218), .A2(n7217), .ZN(n7216) );
  AOI21_X1 U5468 ( .B1(n7509), .B2(n5702), .A(n7497), .ZN(n7600) );
  INV_X1 U5469 ( .A(n5666), .ZN(n5665) );
  NOR2_X1 U5470 ( .A1(n8423), .A2(n5670), .ZN(n8444) );
  NOR2_X1 U5471 ( .A1(n8444), .A2(n8443), .ZN(n8442) );
  INV_X1 U5472 ( .A(n8434), .ZN(n4719) );
  NOR2_X1 U5473 ( .A1(n8433), .A2(n5626), .ZN(n5627) );
  NAND2_X1 U5474 ( .A1(n4756), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U5475 ( .A1(n5672), .A2(n4756), .ZN(n4754) );
  INV_X1 U5476 ( .A(n8470), .ZN(n4756) );
  OR2_X1 U5477 ( .A1(n5723), .A2(n4366), .ZN(n4365) );
  NAND2_X1 U5478 ( .A1(n5720), .A2(n8015), .ZN(n4366) );
  NAND2_X1 U5479 ( .A1(n6227), .A2(n6226), .ZN(n6234) );
  AND2_X1 U5480 ( .A1(n6218), .A2(n6217), .ZN(n6227) );
  NOR2_X1 U5481 ( .A1(n4335), .A2(n4839), .ZN(n4838) );
  INV_X1 U5482 ( .A(n8234), .ZN(n4839) );
  NAND2_X1 U5483 ( .A1(n6187), .A2(n5983), .ZN(n6197) );
  AND2_X1 U5484 ( .A1(n6185), .A2(n6184), .ZN(n6187) );
  AND2_X1 U5485 ( .A1(n8215), .A2(n8214), .ZN(n8328) );
  NOR2_X1 U5486 ( .A1(n8330), .A2(n4848), .ZN(n4847) );
  INV_X1 U5487 ( .A(n8206), .ZN(n4848) );
  INV_X1 U5488 ( .A(n4555), .ZN(n4553) );
  AND2_X1 U5489 ( .A1(n8207), .A2(n8206), .ZN(n8327) );
  NAND2_X1 U5490 ( .A1(n9908), .A2(n7303), .ZN(n8183) );
  INV_X1 U5491 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U5492 ( .A1(n6099), .A2(n7111), .ZN(n6116) );
  INV_X1 U5493 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6086) );
  AND2_X1 U5494 ( .A1(n6087), .A2(n6086), .ZN(n6099) );
  AND4_X1 U5495 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n7172)
         );
  AND2_X1 U5496 ( .A1(n8171), .A2(n8176), .ZN(n8319) );
  NAND2_X1 U5497 ( .A1(n6370), .A2(n6756), .ZN(n7364) );
  INV_X1 U5498 ( .A(n8151), .ZN(n6344) );
  NAND2_X1 U5499 ( .A1(n4561), .A2(n4564), .ZN(n6405) );
  AND2_X1 U5500 ( .A1(n4565), .A2(n4576), .ZN(n4564) );
  NAND2_X1 U5501 ( .A1(n8271), .A2(n8508), .ZN(n4576) );
  NOR2_X1 U5502 ( .A1(n8508), .A2(n8605), .ZN(n6314) );
  AND2_X1 U5503 ( .A1(n8246), .A2(n8249), .ZN(n8564) );
  AND2_X1 U5504 ( .A1(n6216), .A2(n6215), .ZN(n7955) );
  INV_X1 U5505 ( .A(n8333), .ZN(n8221) );
  INV_X1 U5506 ( .A(n8329), .ZN(n8217) );
  NAND2_X1 U5507 ( .A1(n8361), .A2(n8359), .ZN(n9913) );
  OR2_X1 U5508 ( .A1(n8278), .A2(n6860), .ZN(n6756) );
  INV_X1 U5509 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5514) );
  CLKBUF_X1 U5510 ( .A(n5528), .Z(n5539) );
  INV_X1 U5511 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6305) );
  INV_X1 U5512 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U5513 ( .A1(n5558), .A2(n5560), .ZN(n5562) );
  INV_X1 U5514 ( .A(n5582), .ZN(n4855) );
  NOR2_X1 U5515 ( .A1(n5582), .A2(n4854), .ZN(n5586) );
  INV_X1 U5516 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U5517 ( .A1(n5830), .A2(n5829), .ZN(n5833) );
  OR2_X1 U5518 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  AND2_X1 U5519 ( .A1(n5887), .A2(n5886), .ZN(n8766) );
  NAND2_X1 U5520 ( .A1(n4776), .A2(n4774), .ZN(n5797) );
  AOI21_X1 U5521 ( .B1(n4777), .B2(n6948), .A(n4775), .ZN(n4774) );
  INV_X1 U5522 ( .A(n4362), .ZN(n4775) );
  AOI22_X1 U5523 ( .A1(n5939), .A2(n6908), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5956), .ZN(n5741) );
  AOI21_X1 U5524 ( .B1(n4763), .B2(n4765), .A(n5820), .ZN(n4761) );
  NAND2_X1 U5525 ( .A1(n7263), .A2(n7262), .ZN(n4767) );
  NAND2_X1 U5526 ( .A1(n4758), .A2(n4757), .ZN(n4879) );
  NAND2_X1 U5527 ( .A1(n4284), .A2(n4355), .ZN(n4381) );
  OR2_X1 U5528 ( .A1(n8806), .A2(n4384), .ZN(n4383) );
  NAND2_X1 U5529 ( .A1(n5843), .A2(n4355), .ZN(n4382) );
  AND3_X1 U5530 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5002) );
  NOR2_X1 U5531 ( .A1(n5354), .A2(n8797), .ZN(n5369) );
  NOR2_X1 U5532 ( .A1(n5951), .A2(n7896), .ZN(n5963) );
  INV_X1 U5533 ( .A(n7755), .ZN(n4500) );
  OAI21_X1 U5534 ( .B1(n7737), .B2(n7792), .A(n4305), .ZN(n4499) );
  MUX2_X1 U5535 ( .A(n7821), .B(n7754), .S(n7753), .Z(n7755) );
  INV_X1 U5536 ( .A(n4966), .ZN(n5000) );
  INV_X1 U5537 ( .A(n5001), .ZN(n5287) );
  AND2_X1 U5538 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8917) );
  AOI21_X1 U5539 ( .B1(n6624), .B2(P1_REG1_REG_3__SCAN_IN), .A(n9429), .ZN(
        n9491) );
  NAND2_X1 U5540 ( .A1(n6624), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4501) );
  NOR2_X1 U5541 ( .A1(n9520), .A2(n4409), .ZN(n9415) );
  AND2_X1 U5542 ( .A1(n6633), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4409) );
  AND2_X1 U5543 ( .A1(n4504), .A2(n4503), .ZN(n9412) );
  NAND2_X1 U5544 ( .A1(n6633), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4503) );
  NOR2_X1 U5545 ( .A1(n9410), .A2(n4513), .ZN(n9441) );
  AND2_X1 U5546 ( .A1(n6635), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4513) );
  NOR2_X1 U5547 ( .A1(n9444), .A2(n4417), .ZN(n6638) );
  AND2_X1 U5548 ( .A1(n6637), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4417) );
  NOR2_X1 U5549 ( .A1(n9441), .A2(n9442), .ZN(n9440) );
  NAND2_X1 U5550 ( .A1(n6638), .A2(n6639), .ZN(n6845) );
  NOR2_X1 U5551 ( .A1(n9536), .A2(n4408), .ZN(n6849) );
  AND2_X1 U5552 ( .A1(n9531), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4408) );
  NOR2_X1 U5553 ( .A1(n9533), .A2(n9534), .ZN(n9532) );
  NAND2_X1 U5554 ( .A1(n6849), .A2(n6848), .ZN(n8924) );
  NOR2_X1 U5555 ( .A1(n9551), .A2(n4353), .ZN(n9565) );
  NOR2_X1 U5556 ( .A1(n9565), .A2(n9564), .ZN(n9563) );
  XNOR2_X1 U5557 ( .A(n8936), .B(n8937), .ZN(n9578) );
  OR2_X1 U5558 ( .A1(n6641), .A2(n9476), .ZN(n9575) );
  AND2_X1 U5559 ( .A1(n8998), .A2(n4279), .ZN(n8975) );
  NOR2_X1 U5560 ( .A1(n7762), .A2(n4704), .ZN(n4703) );
  AOI21_X1 U5561 ( .B1(n4786), .B2(n4788), .A(n4346), .ZN(n4784) );
  INV_X1 U5562 ( .A(n7762), .ZN(n8984) );
  NOR2_X1 U5563 ( .A1(n9168), .A2(n9011), .ZN(n8998) );
  NAND2_X1 U5564 ( .A1(n9044), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5565 ( .A1(n4699), .A2(n4697), .ZN(n4695) );
  NAND2_X1 U5566 ( .A1(n4699), .A2(n7710), .ZN(n4694) );
  NAND2_X1 U5567 ( .A1(n9091), .A2(n4528), .ZN(n9025) );
  NOR2_X1 U5568 ( .A1(n9178), .A2(n4530), .ZN(n4528) );
  NAND2_X1 U5569 ( .A1(n4675), .A2(n7683), .ZN(n4672) );
  NAND2_X1 U5570 ( .A1(n9091), .A2(n9082), .ZN(n9075) );
  NAND2_X1 U5571 ( .A1(n9091), .A2(n4532), .ZN(n9054) );
  AOI21_X1 U5572 ( .B1(n9110), .B2(n9109), .A(n7683), .ZN(n9087) );
  NOR2_X1 U5573 ( .A1(n9133), .A2(n9208), .ZN(n9117) );
  AND2_X1 U5574 ( .A1(n7681), .A2(n7680), .ZN(n9122) );
  NOR3_X1 U5575 ( .A1(n9142), .A2(n9141), .A3(n9140), .ZN(n9139) );
  NAND2_X1 U5576 ( .A1(n4536), .A2(n9137), .ZN(n4535) );
  INV_X1 U5577 ( .A(n4538), .ZN(n4536) );
  NOR2_X1 U5578 ( .A1(n7254), .A2(n4538), .ZN(n9132) );
  NOR2_X1 U5579 ( .A1(n5171), .A2(n5170), .ZN(n5187) );
  AND2_X1 U5580 ( .A1(n5187), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5205) );
  INV_X1 U5581 ( .A(n4692), .ZN(n4690) );
  NAND2_X1 U5582 ( .A1(n7661), .A2(n7663), .ZN(n7779) );
  AND2_X1 U5583 ( .A1(n7666), .A2(n7662), .ZN(n7777) );
  NAND2_X1 U5584 ( .A1(n9749), .A2(n4521), .ZN(n4520) );
  NOR2_X1 U5585 ( .A1(n4522), .A2(n7100), .ZN(n4521) );
  INV_X1 U5586 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5115) );
  NOR2_X1 U5587 ( .A1(n5116), .A2(n5115), .ZN(n5132) );
  OR2_X1 U5588 ( .A1(n5092), .A2(n5091), .ZN(n5116) );
  NAND2_X1 U5589 ( .A1(n5114), .A2(n5113), .ZN(n7086) );
  NAND2_X1 U5590 ( .A1(n4519), .A2(n4518), .ZN(n7097) );
  NOR2_X1 U5591 ( .A1(n7086), .A2(n4522), .ZN(n4518) );
  INV_X1 U5592 ( .A(n9631), .ZN(n4519) );
  AOI21_X1 U5593 ( .B1(n6996), .B2(n6997), .A(n5477), .ZN(n7077) );
  AND2_X1 U5594 ( .A1(n7848), .A2(n7656), .ZN(n7776) );
  INV_X1 U5595 ( .A(n6997), .ZN(n7773) );
  INV_X1 U5596 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5043) );
  OR2_X1 U5597 ( .A1(n5056), .A2(n5043), .ZN(n5092) );
  INV_X1 U5598 ( .A(n9637), .ZN(n9619) );
  AND2_X1 U5599 ( .A1(n9646), .A2(n9714), .ZN(n9644) );
  NAND2_X1 U5600 ( .A1(n4515), .A2(n4272), .ZN(n9665) );
  NOR2_X1 U5601 ( .A1(n4517), .A2(n5762), .ZN(n4515) );
  NOR2_X1 U5602 ( .A1(n9665), .A2(n6961), .ZN(n9646) );
  AOI21_X1 U5603 ( .B1(n5464), .B2(n4623), .A(n4620), .ZN(n4619) );
  OAI211_X1 U5604 ( .C1(n5015), .C2(n9471), .A(n4944), .B(n4943), .ZN(n4946)
         );
  OR2_X1 U5605 ( .A1(n7751), .A2(n6534), .ZN(n4943) );
  NOR2_X1 U5606 ( .A1(n5740), .A2(n6671), .ZN(n6910) );
  NAND2_X1 U5607 ( .A1(n5353), .A2(n5352), .ZN(n9173) );
  NAND2_X1 U5608 ( .A1(n5258), .A2(n5257), .ZN(n9204) );
  NAND2_X1 U5609 ( .A1(n5204), .A2(n5203), .ZN(n9219) );
  OR2_X1 U5610 ( .A1(n6802), .A2(n7895), .ZN(n9769) );
  OR2_X1 U5611 ( .A1(n7886), .A2(n6802), .ZN(n9767) );
  NAND2_X1 U5612 ( .A1(n7235), .A2(n7837), .ZN(n6802) );
  NAND2_X1 U5613 ( .A1(n9622), .A2(n9680), .ZN(n9773) );
  AND2_X1 U5614 ( .A1(n6472), .A2(n6471), .ZN(n6487) );
  INV_X1 U5615 ( .A(n7896), .ZN(n9380) );
  XNOR2_X1 U5616 ( .A(n4908), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6458) );
  XNOR2_X1 U5617 ( .A(n5391), .B(n5390), .ZN(n7540) );
  XNOR2_X1 U5618 ( .A(n5432), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5453) );
  XNOR2_X1 U5619 ( .A(n5430), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5455) );
  OAI21_X1 U5620 ( .B1(n5429), .B2(n5428), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5430) );
  AND2_X1 U5621 ( .A1(n5329), .A2(n5317), .ZN(n5327) );
  AOI21_X1 U5622 ( .B1(n4490), .B2(n4492), .A(n4489), .ZN(n4488) );
  INV_X1 U5623 ( .A(n5311), .ZN(n4489) );
  INV_X1 U5624 ( .A(n4495), .ZN(n4490) );
  INV_X1 U5625 ( .A(n4492), .ZN(n4491) );
  XNOR2_X1 U5626 ( .A(n5451), .B(n5450), .ZN(n6562) );
  XNOR2_X1 U5627 ( .A(n5410), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5495) );
  INV_X1 U5628 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4822) );
  INV_X1 U5629 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5183) );
  XNOR2_X1 U5630 ( .A(n5126), .B(n5125), .ZN(n6583) );
  OAI21_X1 U5631 ( .B1(n5104), .B2(n5103), .A(n5102), .ZN(n5126) );
  XNOR2_X1 U5632 ( .A(n5081), .B(n4289), .ZN(n6566) );
  NAND2_X1 U5633 ( .A1(n4467), .A2(n5029), .ZN(n5049) );
  NAND2_X1 U5634 ( .A1(n4470), .A2(n4471), .ZN(n4467) );
  INV_X1 U5635 ( .A(n5013), .ZN(n4669) );
  OAI21_X1 U5636 ( .B1(n4497), .B2(n4937), .A(n4940), .ZN(n4958) );
  XNOR2_X1 U5637 ( .A(n4419), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U5638 ( .A1(n4420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4419) );
  AND4_X1 U5639 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n7919)
         );
  AND3_X1 U5640 ( .A1(n6047), .A2(n6046), .A3(n6045), .ZN(n6942) );
  INV_X1 U5641 ( .A(n7971), .ZN(n7972) );
  OAI22_X1 U5642 ( .A1(n7914), .A2(n7240), .B1(n7282), .B2(n7912), .ZN(n7407)
         );
  NAND2_X1 U5643 ( .A1(n4651), .A2(n7620), .ZN(n7626) );
  AND2_X1 U5644 ( .A1(n4646), .A2(n7967), .ZN(n8104) );
  NAND2_X1 U5645 ( .A1(n7454), .A2(n7453), .ZN(n7455) );
  INV_X1 U5646 ( .A(n8132), .ZN(n8116) );
  NAND2_X1 U5647 ( .A1(n7059), .A2(n7058), .ZN(n7136) );
  INV_X1 U5648 ( .A(n8095), .ZN(n8136) );
  NAND2_X1 U5649 ( .A1(n6759), .A2(n8618), .ZN(n8129) );
  NAND2_X1 U5650 ( .A1(n4635), .A2(n4638), .ZN(n8124) );
  NAND2_X1 U5651 ( .A1(n8080), .A2(n4639), .ZN(n4635) );
  INV_X1 U5652 ( .A(n8129), .ZN(n8145) );
  NOR2_X1 U5653 ( .A1(n8133), .A2(n4644), .ZN(n4643) );
  INV_X1 U5654 ( .A(n7941), .ZN(n4644) );
  NAND2_X1 U5655 ( .A1(n7995), .A2(n7941), .ZN(n8134) );
  INV_X1 U5656 ( .A(n8075), .ZN(n8141) );
  AOI21_X1 U5657 ( .B1(n4852), .B2(n4302), .A(n4850), .ZN(n8366) );
  NAND2_X1 U5658 ( .A1(n6260), .A2(n6259), .ZN(n8519) );
  INV_X1 U5659 ( .A(n7957), .ZN(n8581) );
  AOI22_X1 U5660 ( .A1(n6183), .A2(P2_REG0_REG_2__SCAN_IN), .B1(n6420), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n4583) );
  OR2_X2 U5661 ( .A1(n6747), .A2(n5530), .ZN(n8474) );
  OR2_X1 U5662 ( .A1(P2_U3150), .A2(n5719), .ZN(n9831) );
  NAND2_X1 U5663 ( .A1(n4732), .A2(n6787), .ZN(n6707) );
  OAI22_X1 U5664 ( .A1(n6706), .A2(n6705), .B1(n4752), .B2(n5687), .ZN(n6779)
         );
  NAND2_X1 U5665 ( .A1(n4744), .A2(n6499), .ZN(n6520) );
  INV_X1 U5666 ( .A(n4745), .ZN(n4744) );
  NAND2_X1 U5667 ( .A1(n4746), .A2(n6499), .ZN(n6518) );
  NAND2_X1 U5668 ( .A1(n5605), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6524) );
  AOI21_X1 U5669 ( .B1(n6094), .B2(n5698), .A(n7106), .ZN(n7215) );
  INV_X1 U5670 ( .A(n4723), .ZN(n7503) );
  OR2_X1 U5671 ( .A1(n7504), .A2(n7505), .ZN(n4723) );
  INV_X1 U5672 ( .A(n5617), .ZN(n4722) );
  INV_X1 U5673 ( .A(n4743), .ZN(n7605) );
  OAI21_X1 U5674 ( .B1(n7504), .B2(n4721), .A(n4720), .ZN(n7593) );
  NAND2_X1 U5675 ( .A1(n4724), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U5676 ( .A1(n5617), .A2(n4724), .ZN(n4720) );
  INV_X1 U5677 ( .A(n7594), .ZN(n4724) );
  INV_X1 U5678 ( .A(n5620), .ZN(n4727) );
  XNOR2_X1 U5679 ( .A(n5622), .B(n8417), .ZN(n8415) );
  NOR2_X1 U5680 ( .A1(n8415), .A2(n8416), .ZN(n8414) );
  NAND2_X1 U5681 ( .A1(n4718), .A2(n4716), .ZN(n8433) );
  NAND2_X1 U5682 ( .A1(n5623), .A2(n4719), .ZN(n4718) );
  OR2_X1 U5683 ( .A1(n8415), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U5684 ( .A1(n4719), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U5685 ( .A1(n6275), .A2(n6274), .ZN(n8512) );
  OR2_X1 U5686 ( .A1(n8595), .A2(n8594), .ZN(n8663) );
  NAND2_X1 U5687 ( .A1(n6207), .A2(n6206), .ZN(n8661) );
  OAI21_X1 U5688 ( .B1(n8623), .B2(n4546), .A(n4543), .ZN(n8588) );
  NAND2_X1 U5689 ( .A1(n4547), .A2(n4548), .ZN(n8601) );
  NAND2_X1 U5690 ( .A1(n8623), .A2(n4550), .ZN(n4547) );
  NAND2_X1 U5691 ( .A1(n6196), .A2(n6195), .ZN(n8668) );
  NAND2_X1 U5692 ( .A1(n6142), .A2(n6141), .ZN(n9930) );
  OR2_X1 U5693 ( .A1(n9913), .A2(n6393), .ZN(n7441) );
  INV_X1 U5694 ( .A(n9865), .ZN(n8618) );
  INV_X1 U5695 ( .A(n8615), .ZN(n9867) );
  INV_X1 U5696 ( .A(n9913), .ZN(n9931) );
  AND3_X1 U5697 ( .A1(n6752), .A2(n9931), .A3(n6393), .ZN(n9865) );
  AND2_X1 U5698 ( .A1(n6329), .A2(n6328), .ZN(n6342) );
  NAND2_X1 U5699 ( .A1(n8283), .A2(n8282), .ZN(n8679) );
  NAND2_X1 U5700 ( .A1(n4570), .A2(n4571), .ZN(n8496) );
  NAND2_X1 U5701 ( .A1(n8516), .A2(n4574), .ZN(n4570) );
  OAI21_X1 U5702 ( .B1(n8515), .B2(n4286), .A(n4828), .ZN(n8495) );
  OAI21_X1 U5703 ( .B1(n8516), .B2(n6273), .A(n6272), .ZN(n8506) );
  INV_X1 U5704 ( .A(n4827), .ZN(n8504) );
  AOI21_X1 U5705 ( .B1(n8515), .B2(n8266), .A(n4832), .ZN(n4827) );
  INV_X1 U5706 ( .A(n7977), .ZN(n8696) );
  NAND2_X1 U5707 ( .A1(n6252), .A2(n6251), .ZN(n8702) );
  NAND2_X1 U5708 ( .A1(n4837), .A2(n4834), .ZN(n8526) );
  NAND2_X1 U5709 ( .A1(n4837), .A2(n8253), .ZN(n8537) );
  NAND2_X1 U5710 ( .A1(n6233), .A2(n6232), .ZN(n8713) );
  NAND2_X1 U5711 ( .A1(n6225), .A2(n6224), .ZN(n8719) );
  INV_X1 U5712 ( .A(n7955), .ZN(n8726) );
  AOI21_X1 U5713 ( .B1(n8623), .B2(n8621), .A(n8622), .ZN(n8629) );
  NAND2_X1 U5714 ( .A1(n6182), .A2(n6181), .ZN(n8053) );
  AND2_X1 U5715 ( .A1(n7579), .A2(n7578), .ZN(n7587) );
  NAND2_X1 U5716 ( .A1(n6172), .A2(n6171), .ZN(n8225) );
  NAND2_X1 U5717 ( .A1(n6162), .A2(n6161), .ZN(n7990) );
  INV_X1 U5718 ( .A(n8736), .ZN(n8725) );
  OR2_X1 U5719 ( .A1(n9934), .A2(n9913), .ZN(n8736) );
  NAND2_X1 U5720 ( .A1(n6752), .A2(n6589), .ZN(n6597) );
  INV_X1 U5721 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5977) );
  INV_X1 U5722 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7382) );
  INV_X1 U5723 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9297) );
  INV_X1 U5724 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7161) );
  INV_X1 U5725 ( .A(n6858), .ZN(n8361) );
  INV_X1 U5726 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9349) );
  INV_X1 U5727 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7068) );
  XNOR2_X1 U5728 ( .A(n5635), .B(n5634), .ZN(n7067) );
  INV_X1 U5729 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6919) );
  INV_X1 U5730 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6775) );
  INV_X1 U5731 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6655) );
  INV_X1 U5732 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5566) );
  INV_X1 U5733 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6580) );
  INV_X1 U5734 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6567) );
  INV_X1 U5735 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6559) );
  INV_X1 U5736 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5601) );
  OR2_X1 U5737 ( .A1(n5598), .A2(n5597), .ZN(n6543) );
  OR2_X1 U5738 ( .A1(n5644), .A2(n5974), .ZN(n5580) );
  NAND2_X1 U5739 ( .A1(n5576), .A2(n5575), .ZN(n9818) );
  INV_X1 U5740 ( .A(n9047), .ZN(n9074) );
  AND2_X1 U5741 ( .A1(n8763), .A2(n8762), .ZN(n8764) );
  NAND2_X1 U5742 ( .A1(n5395), .A2(n5394), .ZN(n9157) );
  OAI21_X1 U5743 ( .B1(n7263), .B2(n4765), .A(n4763), .ZN(n7395) );
  NAND2_X1 U5744 ( .A1(n4762), .A2(n4766), .ZN(n7397) );
  NAND2_X1 U5745 ( .A1(n7263), .A2(n4287), .ZN(n4762) );
  NAND2_X1 U5746 ( .A1(n8823), .A2(n5907), .ZN(n8794) );
  INV_X1 U5747 ( .A(n8904), .ZN(n8809) );
  INV_X1 U5748 ( .A(n8889), .ZN(n8846) );
  NAND2_X1 U5749 ( .A1(n8805), .A2(n5843), .ZN(n8817) );
  NAND2_X1 U5750 ( .A1(n5221), .A2(n5220), .ZN(n9213) );
  NOR2_X1 U5751 ( .A1(n6678), .A2(n4871), .ZN(n8835) );
  NAND2_X1 U5752 ( .A1(n5304), .A2(n5303), .ZN(n9188) );
  INV_X1 U5753 ( .A(n8887), .ZN(n8867) );
  NAND2_X1 U5754 ( .A1(n4378), .A2(n4381), .ZN(n8861) );
  OR2_X1 U5755 ( .A1(n8804), .A2(n4382), .ZN(n4378) );
  NOR2_X1 U5756 ( .A1(n6947), .A2(n6948), .ZN(n6946) );
  AND2_X1 U5757 ( .A1(n5965), .A2(n9473), .ZN(n8878) );
  OAI21_X1 U5758 ( .B1(n8874), .B2(n8873), .A(n8872), .ZN(n8877) );
  INV_X1 U5759 ( .A(n8905), .ZN(n8892) );
  INV_X1 U5760 ( .A(n8878), .ZN(n8891) );
  AOI21_X1 U5761 ( .B1(n4400), .B2(n4337), .A(n4396), .ZN(n4395) );
  NAND2_X1 U5762 ( .A1(n5830), .A2(n4400), .ZN(n4397) );
  OR2_X1 U5763 ( .A1(n5830), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U5764 ( .A1(n6675), .A2(n5318), .ZN(n5186) );
  AOI211_X1 U5765 ( .C1(n7891), .C2(n9027), .A(n7890), .B(n7889), .ZN(n7892)
         );
  OAI21_X1 U5766 ( .B1(n7758), .B2(n4631), .A(n4630), .ZN(n7889) );
  NAND2_X1 U5767 ( .A1(n4631), .A2(n7888), .ZN(n4630) );
  OR2_X1 U5768 ( .A1(n6492), .A2(n5956), .ZN(n7896) );
  XNOR2_X1 U5769 ( .A(n5448), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7898) );
  INV_X1 U5770 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9480) );
  INV_X1 U5771 ( .A(n4502), .ZN(n9425) );
  INV_X1 U5772 ( .A(n4413), .ZN(n9505) );
  INV_X1 U5773 ( .A(n4506), .ZN(n9501) );
  INV_X1 U5774 ( .A(n4411), .ZN(n9521) );
  INV_X1 U5775 ( .A(n4504), .ZN(n9516) );
  NOR2_X1 U5776 ( .A1(n9440), .A2(n4512), .ZN(n6616) );
  AND2_X1 U5777 ( .A1(n6637), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5778 ( .A1(n6616), .A2(n6617), .ZN(n6840) );
  NOR2_X1 U5779 ( .A1(n9400), .A2(n9399), .ZN(n9398) );
  NAND2_X1 U5780 ( .A1(n6845), .A2(n4416), .ZN(n9400) );
  OR2_X1 U5781 ( .A1(n6846), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4416) );
  NOR2_X1 U5782 ( .A1(n9532), .A2(n4510), .ZN(n6842) );
  AND2_X1 U5783 ( .A1(n9531), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5784 ( .A1(n6842), .A2(n6843), .ZN(n8933) );
  NOR2_X1 U5785 ( .A1(n9549), .A2(n9550), .ZN(n9548) );
  NAND2_X1 U5786 ( .A1(n8924), .A2(n4407), .ZN(n9549) );
  NAND2_X1 U5787 ( .A1(n6854), .A2(n9796), .ZN(n4407) );
  AOI21_X1 U5788 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9556), .A(n9548), .ZN(
        n9561) );
  INV_X1 U5789 ( .A(n8929), .ZN(n8931) );
  NAND2_X1 U5790 ( .A1(n8954), .A2(n4361), .ZN(n9589) );
  AND2_X1 U5791 ( .A1(n8948), .A2(n8947), .ZN(n9586) );
  OR2_X1 U5792 ( .A1(n9604), .A2(n9603), .ZN(n9607) );
  NAND2_X1 U5793 ( .A1(n9585), .A2(n4363), .ZN(n9599) );
  AND2_X1 U5794 ( .A1(n9585), .A2(n8950), .ZN(n9601) );
  OAI21_X1 U5795 ( .B1(n8960), .B2(n9602), .A(n9543), .ZN(n8958) );
  AOI21_X1 U5796 ( .B1(n6464), .B2(n9655), .A(n6463), .ZN(n7911) );
  NAND2_X1 U5797 ( .A1(n6462), .A2(n6461), .ZN(n6463) );
  OR2_X1 U5798 ( .A1(n9161), .A2(n9152), .ZN(n5505) );
  AOI21_X1 U5799 ( .B1(n5426), .B2(n5425), .A(n5424), .ZN(n9160) );
  INV_X1 U5800 ( .A(n5423), .ZN(n5424) );
  AND2_X1 U5801 ( .A1(n5415), .A2(n9655), .ZN(n5426) );
  NAND2_X1 U5802 ( .A1(n4785), .A2(n4789), .ZN(n8997) );
  NAND2_X1 U5803 ( .A1(n9024), .A2(n4790), .ZN(n4785) );
  AND2_X1 U5804 ( .A1(n4793), .A2(n4295), .ZN(n9010) );
  NAND2_X1 U5805 ( .A1(n9024), .A2(n5490), .ZN(n4793) );
  AND2_X1 U5806 ( .A1(n4815), .A2(n4278), .ZN(n9069) );
  NAND2_X1 U5807 ( .A1(n5484), .A2(n4817), .ZN(n9085) );
  NAND2_X1 U5808 ( .A1(n4801), .A2(n4805), .ZN(n9131) );
  NAND2_X1 U5809 ( .A1(n4813), .A2(n4807), .ZN(n4801) );
  NAND2_X1 U5810 ( .A1(n4811), .A2(n4808), .ZN(n7369) );
  INV_X1 U5811 ( .A(n5177), .ZN(n9768) );
  NAND2_X1 U5812 ( .A1(n9380), .A2(n6469), .ZN(n9104) );
  NAND2_X1 U5813 ( .A1(n5146), .A2(n5145), .ZN(n7201) );
  NOR2_X1 U5814 ( .A1(n9631), .A2(n5078), .ZN(n7002) );
  NAND2_X1 U5815 ( .A1(n9642), .A2(n9643), .ZN(n4800) );
  OR2_X1 U5816 ( .A1(n5501), .A2(n9027), .ZN(n8982) );
  NAND2_X1 U5817 ( .A1(n4624), .A2(n7838), .ZN(n9650) );
  NAND2_X1 U5818 ( .A1(n4622), .A2(n4948), .ZN(n4624) );
  INV_X1 U5819 ( .A(n5755), .ZN(n9695) );
  NAND2_X1 U5820 ( .A1(n4948), .A2(n4947), .ZN(n6809) );
  INV_X1 U5821 ( .A(n9113), .ZN(n9673) );
  INV_X1 U5822 ( .A(n9152), .ZN(n9670) );
  AND2_X2 U5823 ( .A1(n6487), .A2(n6486), .ZN(n9803) );
  AND2_X2 U5824 ( .A1(n6487), .A2(n6473), .ZN(n9777) );
  AND2_X1 U5825 ( .A1(n9380), .A2(n9379), .ZN(n9678) );
  XNOR2_X1 U5826 ( .A(n7749), .B(n7748), .ZN(n9383) );
  MUX2_X1 U5827 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4895), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n4897) );
  OR2_X1 U5828 ( .A1(n4894), .A2(n9384), .ZN(n4895) );
  INV_X1 U5829 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4905) );
  CLKBUF_X1 U5830 ( .A(n6458), .Z(n9474) );
  INV_X1 U5831 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9228) );
  INV_X1 U5832 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7392) );
  XNOR2_X1 U5833 ( .A(n5328), .B(n5327), .ZN(n7297) );
  OAI21_X1 U5834 ( .B1(n5271), .B2(n4491), .A(n4488), .ZN(n5328) );
  INV_X1 U5835 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7233) );
  INV_X1 U5836 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7169) );
  INV_X1 U5837 ( .A(n5495), .ZN(n7837) );
  XNOR2_X1 U5838 ( .A(n5414), .B(n5413), .ZN(n7146) );
  INV_X1 U5839 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9350) );
  INV_X1 U5840 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7926) );
  OAI21_X1 U5841 ( .B1(n5404), .B2(P1_IR_REG_31__SCAN_IN), .A(n4388), .ZN(
        n4387) );
  NAND2_X1 U5842 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n4390) );
  NAND2_X1 U5843 ( .A1(n5236), .A2(n5405), .ZN(n5255) );
  INV_X1 U5844 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9274) );
  AND2_X1 U5845 ( .A1(n5182), .A2(n5167), .ZN(n9568) );
  AND2_X1 U5846 ( .A1(n5111), .A2(n5088), .ZN(n9406) );
  INV_X1 U5847 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6571) );
  INV_X1 U5848 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U5849 ( .A1(n5014), .A2(n5013), .ZN(n5024) );
  XNOR2_X1 U5850 ( .A(n4915), .B(n4914), .ZN(n6619) );
  NAND2_X1 U5851 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4914) );
  AND4_X1 U5852 ( .A1(n7572), .A2(n7571), .A3(n7570), .A4(n7569), .ZN(n7573)
         );
  INV_X1 U5853 ( .A(n4728), .ZN(n7558) );
  NAND2_X1 U5854 ( .A1(n8483), .A2(n8484), .ZN(n4738) );
  NOR2_X1 U5855 ( .A1(n8482), .A2(n4740), .ZN(n4739) );
  NAND2_X1 U5856 ( .A1(n4367), .A2(n4307), .ZN(P2_U3201) );
  INV_X1 U5857 ( .A(n5726), .ZN(n4367) );
  AND2_X1 U5858 ( .A1(n4579), .A2(n4580), .ZN(n7934) );
  OAI21_X1 U5859 ( .B1(n6400), .B2(n8615), .A(n6399), .ZN(n6401) );
  NOR2_X1 U5860 ( .A1(n6438), .A2(n4864), .ZN(n6439) );
  OAI21_X1 U5861 ( .B1(n4579), .B2(n9934), .A(n4577), .ZN(P2_U3456) );
  INV_X1 U5862 ( .A(n4578), .ZN(n4577) );
  NOR2_X1 U5863 ( .A1(n6434), .A2(n4870), .ZN(n6435) );
  MUX2_X1 U5864 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9225), .S(n9777), .Z(n9365)
         );
  NAND2_X1 U5865 ( .A1(n6858), .A2(n8373), .ZN(n8278) );
  NAND2_X1 U5866 ( .A1(n6448), .A2(n6447), .ZN(n6465) );
  INV_X1 U5867 ( .A(n5791), .ZN(n5912) );
  AND2_X1 U5868 ( .A1(n4769), .A2(n5869), .ZN(n8784) );
  AND2_X1 U5869 ( .A1(n9689), .A2(n9695), .ZN(n4272) );
  INV_X1 U5870 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5404) );
  NOR2_X1 U5871 ( .A1(n5814), .A2(n5813), .ZN(n4273) );
  AND4_X1 U5872 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5533), .ZN(n4274)
         );
  OAI22_X1 U5873 ( .A1(n8080), .A2(n4634), .B1(n4636), .B2(n7981), .ZN(n7983)
         );
  NAND2_X1 U5874 ( .A1(n8804), .A2(n8806), .ZN(n8805) );
  OAI21_X1 U5875 ( .B1(n4819), .B2(n5143), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5432) );
  NAND2_X1 U5876 ( .A1(n5336), .A2(n5335), .ZN(n9178) );
  AND2_X1 U5877 ( .A1(n4455), .A2(n4452), .ZN(n4275) );
  INV_X1 U5878 ( .A(n8305), .ZN(n8678) );
  NAND2_X1 U5879 ( .A1(n8293), .A2(n8292), .ZN(n8305) );
  XOR2_X1 U5880 ( .A(n5718), .B(n5717), .Z(n4276) );
  OR2_X1 U5881 ( .A1(n8895), .A2(n8809), .ZN(n7859) );
  AND2_X1 U5882 ( .A1(n8481), .A2(n8480), .ZN(n4277) );
  AOI21_X1 U5883 ( .B1(n4639), .B2(n7976), .A(n4327), .ZN(n4638) );
  NAND2_X1 U5884 ( .A1(n9096), .A2(n9112), .ZN(n4278) );
  AND2_X1 U5885 ( .A1(n4525), .A2(n4524), .ZN(n4279) );
  AND2_X1 U5886 ( .A1(n4545), .A2(n8313), .ZN(n4280) );
  AND2_X1 U5887 ( .A1(n8259), .A2(n4833), .ZN(n4281) );
  NOR2_X1 U5888 ( .A1(n4358), .A2(n6131), .ZN(n4282) );
  NAND2_X1 U5889 ( .A1(n8785), .A2(n5888), .ZN(n4283) );
  INV_X1 U5890 ( .A(n5843), .ZN(n4384) );
  OR2_X1 U5891 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  NAND2_X1 U5892 ( .A1(n4383), .A2(n8815), .ZN(n4284) );
  OR2_X1 U5893 ( .A1(n6396), .A2(n7441), .ZN(n8620) );
  INV_X1 U5894 ( .A(n8620), .ZN(n9864) );
  NAND2_X1 U5895 ( .A1(n5729), .A2(n5730), .ZN(n5743) );
  INV_X1 U5896 ( .A(n5193), .ZN(n5196) );
  AND2_X1 U5897 ( .A1(n5026), .A2(SI_6_), .ZN(n4285) );
  INV_X1 U5898 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U5899 ( .A1(n4936), .A2(n4369), .ZN(n4973) );
  OR2_X1 U5900 ( .A1(n8265), .A2(n4832), .ZN(n4286) );
  INV_X2 U5901 ( .A(n5000), .ZN(n7731) );
  OR2_X1 U5902 ( .A1(n9178), .A2(n8798), .ZN(n7799) );
  AND2_X1 U5903 ( .A1(n4273), .A2(n7262), .ZN(n4287) );
  NAND2_X1 U5904 ( .A1(n8895), .A2(n8809), .ZN(n7669) );
  NAND2_X1 U5905 ( .A1(n4548), .A2(n4301), .ZN(n4546) );
  OR2_X1 U5906 ( .A1(n9164), .A2(n5493), .ZN(n7798) );
  NAND2_X1 U5907 ( .A1(n5803), .A2(n5802), .ZN(n4288) );
  AND2_X1 U5908 ( .A1(n5082), .A2(n5038), .ZN(n4289) );
  INV_X1 U5909 ( .A(n8531), .ZN(n8381) );
  AND2_X1 U5910 ( .A1(n6271), .A2(n6270), .ZN(n8531) );
  OR3_X1 U5911 ( .A1(n5528), .A2(n4872), .A3(n4845), .ZN(n4290) );
  AND2_X1 U5912 ( .A1(n8213), .A2(n8328), .ZN(n4291) );
  INV_X1 U5913 ( .A(n7870), .ZN(n4704) );
  AND2_X1 U5914 ( .A1(n5193), .A2(n4682), .ZN(n4292) );
  AND2_X1 U5915 ( .A1(n4580), .A2(n6433), .ZN(n4293) );
  NAND2_X1 U5916 ( .A1(n8115), .A2(n7954), .ZN(n8011) );
  INV_X1 U5917 ( .A(n7887), .ZN(n4631) );
  XNOR2_X1 U5918 ( .A(n8763), .B(n8762), .ZN(n8852) );
  NOR2_X1 U5919 ( .A1(n5582), .A2(n4853), .ZN(n5595) );
  AND2_X1 U5920 ( .A1(n4502), .A2(n4501), .ZN(n4294) );
  NAND2_X1 U5921 ( .A1(n9030), .A2(n8798), .ZN(n4295) );
  AND2_X1 U5922 ( .A1(n6618), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4296) );
  AND3_X1 U5923 ( .A1(n4609), .A2(n4608), .A3(n4891), .ZN(n4297) );
  INV_X1 U5924 ( .A(n5138), .ZN(n5141) );
  NOR2_X1 U5925 ( .A1(n8099), .A2(n8102), .ZN(n4298) );
  NAND2_X1 U5926 ( .A1(n9920), .A2(n8387), .ZN(n4299) );
  OR2_X1 U5927 ( .A1(n9194), .A2(n9059), .ZN(n4300) );
  OR2_X1 U5928 ( .A1(n8668), .A2(n8625), .ZN(n4301) );
  NOR2_X1 U5929 ( .A1(n8356), .A2(n8355), .ZN(n4302) );
  NAND2_X1 U5930 ( .A1(n5273), .A2(n5272), .ZN(n9194) );
  AND2_X1 U5931 ( .A1(n9002), .A2(n7870), .ZN(n4303) );
  NOR2_X1 U5932 ( .A1(n8457), .A2(n5672), .ZN(n4304) );
  NAND2_X1 U5933 ( .A1(n5384), .A2(n5383), .ZN(n9164) );
  AND3_X1 U5934 ( .A1(n6042), .A2(n6041), .A3(n6040), .ZN(n9890) );
  AND3_X1 U5935 ( .A1(n4633), .A2(n4632), .A3(n7820), .ZN(n4305) );
  NAND2_X1 U5936 ( .A1(n5186), .A2(n5185), .ZN(n8895) );
  AND2_X1 U5937 ( .A1(n5495), .A2(n7146), .ZN(n5498) );
  AND2_X1 U5938 ( .A1(n4696), .A2(n7799), .ZN(n4306) );
  AND4_X1 U5939 ( .A1(n6039), .A2(n6038), .A3(n6037), .A4(n6036), .ZN(n8165)
         );
  NAND2_X1 U5940 ( .A1(n5643), .A2(n5642), .ZN(n4307) );
  AND2_X1 U5941 ( .A1(n4862), .A2(n6024), .ZN(n4308) );
  INV_X1 U5942 ( .A(n8344), .ZN(n8277) );
  NAND2_X1 U5943 ( .A1(n8349), .A2(n8284), .ZN(n8344) );
  AND2_X1 U5944 ( .A1(n4434), .A2(n4876), .ZN(n4309) );
  NAND2_X1 U5945 ( .A1(n5815), .A2(n4288), .ZN(n4310) );
  AND2_X1 U5946 ( .A1(n4443), .A2(n4291), .ZN(n4311) );
  INV_X1 U5947 ( .A(n4829), .ZN(n4828) );
  OAI21_X1 U5948 ( .B1(n8265), .B2(n4830), .A(n8147), .ZN(n4829) );
  INV_X1 U5949 ( .A(n4606), .ZN(n4605) );
  NOR2_X1 U5950 ( .A1(n9637), .A2(n7045), .ZN(n4312) );
  NOR2_X1 U5951 ( .A1(n8690), .A2(n7979), .ZN(n4313) );
  INV_X1 U5952 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4781) );
  NOR2_X1 U5953 ( .A1(n7637), .A2(n9001), .ZN(n4314) );
  NOR2_X1 U5954 ( .A1(n8123), .A2(n8074), .ZN(n4315) );
  AND2_X1 U5955 ( .A1(n4455), .A2(n8278), .ZN(n4316) );
  AND2_X1 U5956 ( .A1(n9757), .A2(n7489), .ZN(n4317) );
  AND2_X1 U5957 ( .A1(n9002), .A2(n4703), .ZN(n4318) );
  NAND2_X1 U5958 ( .A1(n5858), .A2(n4863), .ZN(n8776) );
  AND2_X1 U5959 ( .A1(n7237), .A2(n7919), .ZN(n4319) );
  NAND2_X1 U5960 ( .A1(n9137), .A2(n7374), .ZN(n4320) );
  OR2_X1 U5961 ( .A1(n5528), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n4321) );
  OR3_X1 U5962 ( .A1(n5143), .A2(n4890), .A3(n4821), .ZN(n4322) );
  INV_X1 U5963 ( .A(n4530), .ZN(n4529) );
  NAND2_X1 U5964 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  INV_X1 U5965 ( .A(n8498), .ZN(n4438) );
  INV_X1 U5966 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5560) );
  INV_X1 U5967 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U5968 ( .A1(n8661), .A2(n8582), .ZN(n4323) );
  AND2_X1 U5969 ( .A1(n5140), .A2(SI_12_), .ZN(n4324) );
  NAND2_X1 U5970 ( .A1(n8176), .A2(n8167), .ZN(n4325) );
  XNOR2_X1 U5971 ( .A(n7970), .B(n7971), .ZN(n8005) );
  OR2_X1 U5972 ( .A1(n8344), .A2(n8279), .ZN(n4326) );
  INV_X1 U5973 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U5974 ( .A1(n5644), .A2(n5579), .ZN(n5582) );
  AND2_X1 U5975 ( .A1(n4642), .A2(n8531), .ZN(n4327) );
  AND2_X1 U5976 ( .A1(n6019), .A2(n6020), .ZN(n4328) );
  INV_X1 U5977 ( .A(n7891), .ZN(n4498) );
  NAND2_X1 U5978 ( .A1(n5492), .A2(n4295), .ZN(n4329) );
  INV_X1 U5979 ( .A(n4546), .ZN(n4545) );
  AND2_X1 U5980 ( .A1(n7798), .A2(n9003), .ZN(n4330) );
  AND2_X1 U5981 ( .A1(n7646), .A2(n7652), .ZN(n4331) );
  NOR2_X1 U5982 ( .A1(n8081), .A2(n7976), .ZN(n4332) );
  NAND2_X1 U5983 ( .A1(n8871), .A2(n5920), .ZN(n8875) );
  OAI21_X1 U5984 ( .B1(n4543), .B2(n8594), .A(n4323), .ZN(n4542) );
  AND2_X1 U5985 ( .A1(n4278), .A2(n4300), .ZN(n4333) );
  NAND2_X1 U5986 ( .A1(n6896), .A2(n6033), .ZN(n8164) );
  AND2_X1 U5987 ( .A1(n8217), .A2(n8216), .ZN(n4334) );
  OR2_X1 U5988 ( .A1(n8602), .A2(n8313), .ZN(n4335) );
  INV_X1 U5989 ( .A(n4835), .ZN(n4834) );
  NAND2_X1 U5990 ( .A1(n4836), .A2(n8253), .ZN(n4835) );
  AND3_X1 U5991 ( .A1(n5406), .A2(n5405), .A3(n5404), .ZN(n4336) );
  INV_X1 U5992 ( .A(n6552), .ZN(n4747) );
  NAND2_X1 U5993 ( .A1(n5498), .A2(n5730), .ZN(n5791) );
  NAND2_X1 U5994 ( .A1(n6296), .A2(n6295), .ZN(n8286) );
  INV_X1 U5995 ( .A(n8286), .ZN(n4437) );
  AND2_X1 U5996 ( .A1(n4767), .A2(n4288), .ZN(n7422) );
  INV_X1 U5997 ( .A(n9033), .ZN(n4617) );
  AND2_X1 U5998 ( .A1(n5832), .A2(n5829), .ZN(n4337) );
  NAND2_X1 U5999 ( .A1(n5320), .A2(n5319), .ZN(n9183) );
  INV_X1 U6000 ( .A(n9183), .ZN(n4531) );
  NAND2_X1 U6001 ( .A1(n4484), .A2(n7730), .ZN(n8978) );
  INV_X1 U6002 ( .A(n8978), .ZN(n4524) );
  OR2_X1 U6003 ( .A1(n7250), .A2(n7665), .ZN(n4691) );
  XNOR2_X1 U6004 ( .A(n7724), .B(SI_29_), .ZN(n8750) );
  AND2_X1 U6005 ( .A1(n8707), .A2(n8555), .ZN(n8312) );
  INV_X1 U6006 ( .A(n8312), .ZN(n4836) );
  INV_X1 U6007 ( .A(n4946), .ZN(n9689) );
  OAI211_X1 U6008 ( .C1(n5943), .C2(n7898), .A(n5730), .B(n6905), .ZN(n5817)
         );
  INV_X1 U6009 ( .A(n7768), .ZN(n4598) );
  INV_X1 U6010 ( .A(n8271), .ZN(n8685) );
  AND2_X1 U6011 ( .A1(n6285), .A2(n6284), .ZN(n8271) );
  NAND2_X1 U6012 ( .A1(n4560), .A2(n6170), .ZN(n7546) );
  NAND2_X1 U6013 ( .A1(n7796), .A2(n7818), .ZN(n7792) );
  INV_X1 U6014 ( .A(n7792), .ZN(n6453) );
  NAND2_X1 U6015 ( .A1(n5239), .A2(n5238), .ZN(n9208) );
  NAND2_X1 U6016 ( .A1(n7413), .A2(n7412), .ZN(n7454) );
  NAND2_X1 U6017 ( .A1(n4609), .A2(n4608), .ZN(n5143) );
  INV_X1 U6018 ( .A(n8546), .ZN(n8707) );
  NAND2_X1 U6019 ( .A1(n6241), .A2(n6240), .ZN(n8546) );
  INV_X1 U6020 ( .A(n8754), .ZN(n5832) );
  AND2_X1 U6021 ( .A1(n4691), .A2(n4690), .ZN(n4338) );
  AND2_X1 U6022 ( .A1(n4849), .A2(n8206), .ZN(n4339) );
  NOR2_X1 U6023 ( .A1(n8414), .A2(n5623), .ZN(n4340) );
  NAND2_X1 U6024 ( .A1(n9091), .A2(n4529), .ZN(n4533) );
  AND2_X1 U6025 ( .A1(n7969), .A2(n8567), .ZN(n4341) );
  AND2_X1 U6026 ( .A1(n4728), .A2(n4727), .ZN(n4342) );
  INV_X1 U6027 ( .A(n4818), .ZN(n4817) );
  AND2_X1 U6028 ( .A1(n4811), .A2(n4809), .ZN(n4343) );
  AND3_X1 U6029 ( .A1(n5831), .A2(n5833), .A3(n5832), .ZN(n4344) );
  OR2_X1 U6030 ( .A1(n8490), .A2(n8360), .ZN(n4345) );
  NOR2_X1 U6031 ( .A1(n9168), .A2(n9020), .ZN(n4346) );
  NOR2_X1 U6032 ( .A1(n8863), .A2(n5856), .ZN(n4347) );
  OR2_X1 U6033 ( .A1(n5143), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n4348) );
  INV_X1 U6034 ( .A(n7981), .ZN(n4641) );
  INV_X1 U6035 ( .A(n5869), .ZN(n4771) );
  INV_X1 U6036 ( .A(n4640), .ZN(n4639) );
  OR2_X1 U6037 ( .A1(n8047), .A2(n4332), .ZN(n4640) );
  INV_X1 U6038 ( .A(n7807), .ZN(n4674) );
  NOR2_X1 U6039 ( .A1(n8777), .A2(n5868), .ZN(n4349) );
  OR2_X1 U6040 ( .A1(n5143), .A2(n4821), .ZN(n4350) );
  INV_X1 U6041 ( .A(n7967), .ZN(n4647) );
  AND2_X1 U6042 ( .A1(n6382), .A2(n6381), .ZN(n9934) );
  OR2_X1 U6043 ( .A1(n7254), .A2(n5177), .ZN(n4351) );
  OR2_X1 U6044 ( .A1(n7898), .A2(n7928), .ZN(n7888) );
  AND2_X1 U6045 ( .A1(n6653), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4352) );
  AND2_X1 U6046 ( .A1(n9556), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4353) );
  NAND2_X1 U6047 ( .A1(n5475), .A2(n5474), .ZN(n6996) );
  NAND2_X1 U6048 ( .A1(n4797), .A2(n4798), .ZN(n9620) );
  NAND2_X1 U6049 ( .A1(n4800), .A2(n5471), .ZN(n7034) );
  NAND2_X1 U6050 ( .A1(n8833), .A2(n5766), .ZN(n6735) );
  NAND2_X1 U6051 ( .A1(n6025), .A2(n6024), .ZN(n9857) );
  INV_X1 U6052 ( .A(n6869), .ZN(n6863) );
  NOR2_X1 U6053 ( .A1(n6946), .A2(n5785), .ZN(n4354) );
  OR2_X1 U6054 ( .A1(n5850), .A2(n5849), .ZN(n4355) );
  INV_X1 U6055 ( .A(n6320), .ZN(n6325) );
  AND3_X1 U6056 ( .A1(n4557), .A2(n4556), .A3(n4553), .ZN(n4356) );
  NOR2_X1 U6057 ( .A1(n7254), .A2(n4535), .ZN(n4534) );
  AND2_X1 U6058 ( .A1(n4723), .A2(n4722), .ZN(n4357) );
  AND2_X1 U6059 ( .A1(n6132), .A2(n7273), .ZN(n4358) );
  NOR2_X1 U6060 ( .A1(n4520), .A2(n9631), .ZN(n7098) );
  AND2_X1 U6061 ( .A1(n7859), .A2(n7669), .ZN(n7781) );
  INV_X1 U6062 ( .A(n7781), .ZN(n4812) );
  AND2_X1 U6063 ( .A1(n7136), .A2(n7135), .ZN(n4359) );
  INV_X1 U6064 ( .A(n9844), .ZN(n9827) );
  AND2_X1 U6065 ( .A1(n4730), .A2(n6787), .ZN(n4360) );
  AND2_X1 U6066 ( .A1(n6097), .A2(n6096), .ZN(n9908) );
  AND2_X2 U6067 ( .A1(n6342), .A2(n6389), .ZN(n9952) );
  OR2_X1 U6068 ( .A1(n8955), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4361) );
  INV_X1 U6069 ( .A(n5078), .ZN(n4523) );
  INV_X1 U6070 ( .A(n8608), .ZN(n9870) );
  INV_X1 U6071 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4846) );
  OR2_X1 U6072 ( .A1(n5790), .A2(n5789), .ZN(n4362) );
  NAND2_X1 U6073 ( .A1(n9683), .A2(n6671), .ZN(n6906) );
  INV_X1 U6074 ( .A(n4517), .ZN(n4516) );
  AND2_X1 U6075 ( .A1(n9600), .A2(n8950), .ZN(n4363) );
  AND2_X1 U6076 ( .A1(n4753), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4364) );
  INV_X1 U6077 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5061) );
  NOR2_X1 U6078 ( .A1(n5976), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U6079 ( .A1(n5652), .A2(n6538), .ZN(n6781) );
  OR2_X1 U6080 ( .A1(n5652), .A2(n6538), .ZN(n4753) );
  NAND2_X1 U6081 ( .A1(n5594), .A2(n6538), .ZN(n6787) );
  NAND2_X1 U6082 ( .A1(n6538), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4750) );
  INV_X1 U6083 ( .A(n6538), .ZN(n4752) );
  NAND2_X1 U6084 ( .A1(n4655), .A2(n4658), .ZN(n5564) );
  NOR2_X2 U6085 ( .A1(n5528), .A2(n4845), .ZN(n4659) );
  XNOR2_X1 U6086 ( .A(n5666), .B(n6649), .ZN(n7567) );
  INV_X1 U6087 ( .A(n5656), .ZN(n4748) );
  NOR2_X1 U6088 ( .A1(n7495), .A2(n5663), .ZN(n7607) );
  NAND2_X1 U6089 ( .A1(n4373), .A2(n4372), .ZN(n4371) );
  NAND2_X1 U6090 ( .A1(n5731), .A2(n5743), .ZN(n4372) );
  INV_X1 U6091 ( .A(n5743), .ZN(n4377) );
  NAND2_X1 U6092 ( .A1(n9683), .A2(n5731), .ZN(n4375) );
  NOR2_X1 U6093 ( .A1(n5736), .A2(n5735), .ZN(n5745) );
  NAND2_X1 U6094 ( .A1(n8804), .A2(n4381), .ZN(n4380) );
  NAND2_X1 U6095 ( .A1(n5236), .A2(n4386), .ZN(n4385) );
  OAI21_X1 U6096 ( .B1(n8835), .B2(n4393), .A(n4391), .ZN(n5777) );
  INV_X1 U6097 ( .A(n4392), .ZN(n4391) );
  OAI21_X1 U6098 ( .B1(n8834), .B2(n4393), .A(n5774), .ZN(n4392) );
  INV_X1 U6099 ( .A(n5766), .ZN(n4393) );
  NAND2_X1 U6100 ( .A1(n8835), .A2(n8834), .ZN(n8833) );
  NAND3_X1 U6101 ( .A1(n4398), .A2(n4397), .A3(n4395), .ZN(n8883) );
  NAND2_X1 U6102 ( .A1(n6618), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6621) );
  INV_X1 U6103 ( .A(n4936), .ZN(n4420) );
  INV_X1 U6104 ( .A(n8275), .ZN(n4427) );
  NAND2_X1 U6105 ( .A1(n4442), .A2(n4440), .ZN(n8223) );
  NAND3_X1 U6106 ( .A1(n4443), .A2(n4444), .A3(n4291), .ZN(n4441) );
  NAND2_X1 U6107 ( .A1(n8205), .A2(n4311), .ZN(n4442) );
  OR2_X1 U6108 ( .A1(n4445), .A2(n8204), .ZN(n4444) );
  NAND2_X1 U6109 ( .A1(n8208), .A2(n8209), .ZN(n4445) );
  NAND2_X1 U6110 ( .A1(n8263), .A2(n4446), .ZN(n8269) );
  NAND2_X1 U6111 ( .A1(n4447), .A2(n8278), .ZN(n4446) );
  OAI21_X1 U6112 ( .B1(n4449), .B2(n4448), .A(n8309), .ZN(n4447) );
  NOR2_X1 U6113 ( .A1(n8260), .A2(n8311), .ZN(n4449) );
  NAND2_X1 U6114 ( .A1(n8239), .A2(n8238), .ZN(n4451) );
  NAND2_X1 U6115 ( .A1(n8163), .A2(n4460), .ZN(n4458) );
  OAI21_X1 U6116 ( .B1(n8163), .B2(n8162), .A(n8316), .ZN(n8174) );
  NAND3_X1 U6117 ( .A1(n5558), .A2(n4461), .A3(n4462), .ZN(n5633) );
  NAND2_X1 U6118 ( .A1(n5361), .A2(n5360), .ZN(n4463) );
  NAND2_X1 U6119 ( .A1(n5346), .A2(n5345), .ZN(n4464) );
  NAND2_X1 U6120 ( .A1(n4465), .A2(n4667), .ZN(n4468) );
  INV_X1 U6121 ( .A(n4667), .ZN(n4471) );
  NAND2_X1 U6122 ( .A1(n4668), .A2(n5014), .ZN(n4470) );
  NAND2_X1 U6123 ( .A1(n5197), .A2(n4476), .ZN(n4474) );
  NAND2_X1 U6124 ( .A1(n5271), .A2(n4488), .ZN(n4485) );
  NAND2_X1 U6125 ( .A1(n4485), .A2(n4486), .ZN(n5330) );
  NAND2_X1 U6126 ( .A1(n5271), .A2(n5270), .ZN(n5298) );
  INV_X1 U6127 ( .A(n4938), .ZN(n4497) );
  NAND3_X1 U6128 ( .A1(n4500), .A2(n4499), .A3(n4498), .ZN(n7758) );
  NAND3_X1 U6129 ( .A1(n9480), .A2(n4915), .A3(n4507), .ZN(n4955) );
  MUX2_X1 U6130 ( .A(n9397), .B(P1_IR_REG_0__SCAN_IN), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  MUX2_X1 U6131 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9397), .S(n4927), .Z(n6908) );
  AND2_X1 U6132 ( .A1(n8998), .A2(n4527), .ZN(n8967) );
  NAND2_X1 U6133 ( .A1(n8998), .A2(n8994), .ZN(n8988) );
  INV_X1 U6134 ( .A(n4533), .ZN(n9041) );
  INV_X1 U6135 ( .A(n4534), .ZN(n9133) );
  NAND2_X1 U6136 ( .A1(n4856), .A2(n4540), .ZN(n4854) );
  NAND2_X1 U6137 ( .A1(n4855), .A2(n4540), .ZN(n5587) );
  XNOR2_X1 U6138 ( .A(n5583), .B(n4540), .ZN(n6546) );
  INV_X1 U6139 ( .A(n8623), .ZN(n4541) );
  AOI21_X1 U6140 ( .B1(n4541), .B2(n4280), .A(n4542), .ZN(n8580) );
  AND2_X1 U6141 ( .A1(n8067), .A2(n8382), .ZN(n4552) );
  NAND2_X1 U6142 ( .A1(n6131), .A2(n4299), .ZN(n4557) );
  NAND3_X1 U6143 ( .A1(n6132), .A2(n7273), .A3(n4299), .ZN(n4556) );
  NAND2_X1 U6144 ( .A1(n4560), .A2(n4558), .ZN(n6180) );
  NAND2_X1 U6145 ( .A1(n6262), .A2(n4866), .ZN(n8516) );
  NAND2_X1 U6146 ( .A1(n6262), .A2(n4562), .ZN(n4561) );
  NAND2_X1 U6147 ( .A1(n6429), .A2(n9861), .ZN(n4579) );
  NAND2_X1 U6148 ( .A1(n4579), .A2(n4293), .ZN(n6436) );
  INV_X1 U6149 ( .A(n6428), .ZN(n4580) );
  NAND2_X1 U6150 ( .A1(n6025), .A2(n4308), .ZN(n7125) );
  NAND2_X1 U6151 ( .A1(n6055), .A2(n7125), .ZN(n7126) );
  INV_X2 U6152 ( .A(n6017), .ZN(n6420) );
  AOI22_X1 U6153 ( .A1(n4595), .A2(n7753), .B1(n4999), .B2(n4593), .ZN(n4604)
         );
  NAND3_X1 U6154 ( .A1(n4597), .A2(n4596), .A3(n4331), .ZN(n4595) );
  NAND2_X1 U6155 ( .A1(n4605), .A2(n7645), .ZN(n4596) );
  NAND2_X1 U6156 ( .A1(n4605), .A2(n4598), .ZN(n4597) );
  NOR2_X1 U6157 ( .A1(n4874), .A2(n7753), .ZN(n4602) );
  NAND2_X1 U6158 ( .A1(n7644), .A2(n7643), .ZN(n4606) );
  INV_X1 U6159 ( .A(n4819), .ZN(n4607) );
  AOI21_X1 U6160 ( .B1(n4614), .B2(n4613), .A(n4610), .ZN(n7720) );
  AND2_X1 U6161 ( .A1(n4616), .A2(n4615), .ZN(n7715) );
  INV_X1 U6162 ( .A(n7839), .ZN(n4620) );
  NAND2_X1 U6163 ( .A1(n4621), .A2(n4619), .ZN(n6954) );
  NAND3_X1 U6164 ( .A1(n4622), .A2(n4948), .A3(n5464), .ZN(n4621) );
  INV_X1 U6165 ( .A(n7838), .ZN(n4623) );
  AOI21_X1 U6166 ( .B1(n7682), .B2(n7864), .A(n7868), .ZN(n7684) );
  NOR3_X1 U6167 ( .A1(n7684), .A2(n7690), .A3(n7683), .ZN(n7685) );
  AOI21_X1 U6168 ( .B1(n7694), .B2(n7693), .A(n7692), .ZN(n7699) );
  MUX2_X1 U6169 ( .A(n7686), .B(n7685), .S(n7888), .Z(n7694) );
  OAI21_X1 U6170 ( .B1(n7654), .B2(n7653), .A(n7652), .ZN(n7657) );
  NAND2_X1 U6171 ( .A1(n4931), .A2(n4930), .ZN(n6817) );
  OAI211_X1 U6172 ( .C1(n7699), .C2(n7698), .A(n9046), .B(n7786), .ZN(n7708)
         );
  AOI21_X1 U6173 ( .B1(n8539), .B2(n6250), .A(n6249), .ZN(n8528) );
  INV_X1 U6174 ( .A(n4656), .ZN(n4655) );
  NAND4_X2 U6175 ( .A1(n4924), .A2(n4923), .A3(n4922), .A4(n4921), .ZN(n5740)
         );
  NAND2_X1 U6176 ( .A1(n7995), .A2(n4643), .ZN(n8055) );
  NAND2_X1 U6177 ( .A1(n8115), .A2(n4648), .ZN(n4646) );
  OAI21_X2 U6178 ( .B1(n7059), .B2(n4653), .A(n4652), .ZN(n7914) );
  INV_X1 U6179 ( .A(n4853), .ZN(n4658) );
  NOR2_X2 U6180 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5644) );
  NAND4_X1 U6181 ( .A1(n5579), .A2(n5506), .A3(n9239), .A4(n4657), .ZN(n4656)
         );
  INV_X1 U6182 ( .A(n4659), .ZN(n5524) );
  NAND2_X1 U6183 ( .A1(n4659), .A2(n5517), .ZN(n5549) );
  NAND3_X1 U6184 ( .A1(n4661), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4660) );
  NAND3_X1 U6185 ( .A1(n6985), .A2(n4664), .A3(n4663), .ZN(n4662) );
  OAI21_X1 U6186 ( .B1(n5014), .B2(n4666), .A(n4665), .ZN(n5069) );
  AOI21_X1 U6187 ( .B1(n4669), .B2(n5023), .A(n4285), .ZN(n4665) );
  INV_X1 U6188 ( .A(n5023), .ZN(n4666) );
  OAI21_X1 U6189 ( .B1(n5023), .B2(n4285), .A(n5070), .ZN(n4667) );
  NOR2_X1 U6190 ( .A1(n4285), .A2(n4669), .ZN(n4668) );
  NOR2_X1 U6191 ( .A1(n9062), .A2(n4674), .ZN(n4671) );
  NAND2_X1 U6192 ( .A1(n9110), .A2(n4675), .ZN(n4673) );
  NAND3_X1 U6193 ( .A1(n4673), .A2(n4672), .A3(n7807), .ZN(n9061) );
  NAND2_X1 U6194 ( .A1(n5159), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U6195 ( .A1(n5159), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U6196 ( .A1(n5159), .A2(n5158), .ZN(n5181) );
  INV_X1 U6197 ( .A(n7665), .ZN(n4688) );
  INV_X1 U6198 ( .A(n7250), .ZN(n4689) );
  INV_X1 U6199 ( .A(n9044), .ZN(n4693) );
  OAI21_X1 U6200 ( .B1(n4693), .B2(n4695), .A(n4694), .ZN(n9016) );
  NAND2_X1 U6201 ( .A1(n9044), .A2(n7704), .ZN(n9032) );
  INV_X1 U6202 ( .A(n4696), .ZN(n9031) );
  INV_X1 U6203 ( .A(n7704), .ZN(n4698) );
  NAND2_X1 U6204 ( .A1(n9004), .A2(n4330), .ZN(n4702) );
  NAND2_X1 U6205 ( .A1(n9004), .A2(n9003), .ZN(n9002) );
  NAND2_X1 U6206 ( .A1(n5083), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U6207 ( .A1(n4705), .A2(n4709), .ZN(n5156) );
  XNOR2_X1 U6208 ( .A(n5616), .B(n7509), .ZN(n7504) );
  NAND2_X1 U6209 ( .A1(n4731), .A2(n6787), .ZN(n5599) );
  INV_X1 U6210 ( .A(n5594), .ZN(n4733) );
  NAND2_X1 U6211 ( .A1(n5585), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U6212 ( .A1(n5585), .A2(n9833), .ZN(n6660) );
  NAND3_X1 U6213 ( .A1(n4741), .A2(n4739), .A3(n4738), .ZN(P2_U3200) );
  OAI21_X1 U6214 ( .B1(n8479), .B2(n4277), .A(n5642), .ZN(n4741) );
  NAND2_X1 U6215 ( .A1(n4745), .A2(n6499), .ZN(n5657) );
  NAND2_X1 U6216 ( .A1(n4749), .A2(n4750), .ZN(n5654) );
  NAND2_X1 U6217 ( .A1(n5652), .A2(n4751), .ZN(n4749) );
  OAI21_X1 U6218 ( .B1(n8459), .B2(n4755), .A(n4754), .ZN(n8469) );
  NOR2_X1 U6219 ( .A1(n8459), .A2(n8458), .ZN(n8457) );
  INV_X1 U6220 ( .A(n4759), .ZN(n4757) );
  XNOR2_X1 U6221 ( .A(n5749), .B(n4377), .ZN(n4759) );
  INV_X1 U6222 ( .A(n5751), .ZN(n4758) );
  NAND2_X1 U6223 ( .A1(n5751), .A2(n4759), .ZN(n5752) );
  NAND2_X1 U6224 ( .A1(n7263), .A2(n4763), .ZN(n4760) );
  NAND2_X1 U6225 ( .A1(n4760), .A2(n4761), .ZN(n7468) );
  NAND2_X1 U6226 ( .A1(n5858), .A2(n4770), .ZN(n4769) );
  NAND2_X1 U6227 ( .A1(n4769), .A2(n4768), .ZN(n5894) );
  NAND2_X1 U6228 ( .A1(n6947), .A2(n4777), .ZN(n4776) );
  NOR2_X1 U6229 ( .A1(n4821), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4782) );
  NOR2_X1 U6230 ( .A1(n4821), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U6231 ( .A1(n5831), .A2(n5833), .ZN(n8753) );
  NAND2_X1 U6232 ( .A1(n4783), .A2(n4784), .ZN(n8983) );
  NAND2_X1 U6233 ( .A1(n9024), .A2(n4786), .ZN(n4783) );
  NAND2_X1 U6234 ( .A1(n9642), .A2(n4796), .ZN(n4797) );
  INV_X1 U6235 ( .A(n7345), .ZN(n4813) );
  NAND2_X1 U6236 ( .A1(n4815), .A2(n4333), .ZN(n5486) );
  NAND2_X1 U6237 ( .A1(n5484), .A2(n4816), .ZN(n4815) );
  NOR2_X1 U6238 ( .A1(n9103), .A2(n9089), .ZN(n4818) );
  INV_X1 U6239 ( .A(n6834), .ZN(n6345) );
  NAND2_X1 U6240 ( .A1(n6929), .A2(n6865), .ZN(n8152) );
  NAND2_X1 U6241 ( .A1(n6344), .A2(n6345), .ZN(n6833) );
  INV_X1 U6242 ( .A(n4823), .ZN(n6416) );
  NAND2_X1 U6243 ( .A1(n4840), .A2(n4838), .ZN(n8574) );
  NAND2_X1 U6244 ( .A1(n6362), .A2(n8231), .ZN(n8617) );
  INV_X1 U6245 ( .A(n8231), .ZN(n4842) );
  INV_X1 U6246 ( .A(n4845), .ZN(n4844) );
  NOR2_X1 U6247 ( .A1(n8852), .A2(n8854), .ZN(n8853) );
  NAND2_X2 U6248 ( .A1(n5743), .A2(n5817), .ZN(n5746) );
  NAND2_X1 U6249 ( .A1(n5947), .A2(n4869), .ZN(n5972) );
  OAI21_X1 U6250 ( .B1(n6480), .B2(n6479), .A(n8876), .ZN(n6485) );
  NAND2_X1 U6251 ( .A1(n5409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5410) );
  AND2_X1 U6252 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  INV_X1 U6253 ( .A(n9396), .ZN(n4898) );
  INV_X2 U6254 ( .A(n5071), .ZN(n5318) );
  XNOR2_X1 U6255 ( .A(n6870), .B(n6863), .ZN(n6880) );
  AND2_X1 U6256 ( .A1(n7273), .A2(n7272), .ZN(n7335) );
  NAND2_X1 U6257 ( .A1(n4904), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4906) );
  INV_X1 U6258 ( .A(n5754), .ZN(n6820) );
  CLKBUF_X1 U6259 ( .A(n5640), .Z(n8370) );
  AND2_X1 U6260 ( .A1(n8574), .A2(n8573), .ZN(n8662) );
  INV_X1 U6262 ( .A(n6430), .ZN(n6432) );
  NOR2_X1 U6263 ( .A1(n6099), .A2(n6088), .ZN(n4857) );
  INV_X1 U6264 ( .A(n9822), .ZN(n5642) );
  AND2_X1 U6265 ( .A1(n5508), .A2(n5507), .ZN(n4858) );
  AND2_X1 U6266 ( .A1(n5165), .A2(n5183), .ZN(n4860) );
  OR2_X1 U6267 ( .A1(n5730), .A2(n6574), .ZN(n4861) );
  OR2_X1 U6268 ( .A1(n8393), .A2(n6033), .ZN(n4862) );
  OR2_X1 U6269 ( .A1(n5857), .A2(n8862), .ZN(n4863) );
  AND2_X1 U6270 ( .A1(n9950), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4864) );
  OR2_X1 U6271 ( .A1(n9160), .A2(n9658), .ZN(n4865) );
  OR2_X1 U6272 ( .A1(n8646), .A2(n8541), .ZN(n4866) );
  OR2_X1 U6273 ( .A1(n9082), .A2(n9090), .ZN(n4868) );
  AND2_X1 U6274 ( .A1(n5946), .A2(n5945), .ZN(n4869) );
  AND2_X1 U6275 ( .A1(n9934), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4870) );
  INV_X1 U6276 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5127) );
  INV_X1 U6277 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4911) );
  AND2_X1 U6278 ( .A1(n5761), .A2(n5760), .ZN(n4871) );
  OR2_X1 U6279 ( .A1(n5548), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4872) );
  OR2_X1 U6280 ( .A1(n5797), .A2(n5796), .ZN(n4873) );
  NAND2_X1 U6281 ( .A1(n7646), .A2(n7009), .ZN(n4874) );
  AND2_X1 U6282 ( .A1(n8363), .A2(n8362), .ZN(n4875) );
  INV_X1 U6283 ( .A(n8165), .ZN(n6877) );
  AND2_X1 U6284 ( .A1(n8354), .A2(n8349), .ZN(n4876) );
  AND2_X1 U6285 ( .A1(n8307), .A2(n8284), .ZN(n4877) );
  AND2_X1 U6286 ( .A1(n5505), .A2(n5504), .ZN(n4878) );
  OR2_X1 U6287 ( .A1(n6380), .A2(n8373), .ZN(n9915) );
  INV_X1 U6288 ( .A(n9915), .ZN(n6431) );
  NAND2_X1 U6289 ( .A1(n8171), .A2(n8178), .ZN(n8168) );
  NOR3_X1 U6290 ( .A1(n8186), .A2(n8323), .A3(n8194), .ZN(n8205) );
  AND2_X1 U6291 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  NAND2_X1 U6292 ( .A1(n8262), .A2(n8301), .ZN(n8263) );
  OAI211_X1 U6293 ( .C1(n8269), .C2(n8517), .A(n8505), .B(n8268), .ZN(n8275)
         );
  NOR2_X1 U6294 ( .A1(n8546), .A2(n8555), .ZN(n6249) );
  OR2_X1 U6295 ( .A1(n5891), .A2(n8787), .ZN(n8761) );
  NAND2_X1 U6296 ( .A1(n7880), .A2(n8972), .ZN(n7820) );
  NAND2_X1 U6297 ( .A1(n5178), .A2(n7662), .ZN(n7665) );
  INV_X1 U6298 ( .A(n6619), .ZN(n4916) );
  NAND2_X1 U6299 ( .A1(n6407), .A2(n6406), .ZN(n6411) );
  INV_X1 U6300 ( .A(n7970), .ZN(n7973) );
  NAND2_X1 U6301 ( .A1(n6507), .A2(n5610), .ZN(n5613) );
  NAND2_X1 U6302 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  NOR2_X1 U6303 ( .A1(n5286), .A2(n8789), .ZN(n5305) );
  INV_X1 U6304 ( .A(n5409), .ZN(n5408) );
  NAND2_X1 U6305 ( .A1(n4941), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4910) );
  AND2_X1 U6306 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  NAND2_X1 U6307 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  INV_X1 U6308 ( .A(n7625), .ZN(n7624) );
  INV_X1 U6309 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6048) );
  INV_X1 U6310 ( .A(n6077), .ZN(n6419) );
  NAND2_X1 U6311 ( .A1(n5584), .A2(n6546), .ZN(n9833) );
  INV_X1 U6312 ( .A(n5625), .ZN(n5626) );
  AND2_X1 U6313 ( .A1(n9839), .A2(n8368), .ZN(n5723) );
  NAND2_X1 U6314 ( .A1(n9870), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6397) );
  OR2_X1 U6315 ( .A1(n6116), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6135) );
  NOR2_X1 U6316 ( .A1(n6075), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6087) );
  NOR2_X1 U6317 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6049) );
  AND2_X1 U6318 ( .A1(n5944), .A2(n8876), .ZN(n5945) );
  INV_X1 U6319 ( .A(n5791), .ZN(n5939) );
  NOR2_X1 U6320 ( .A1(n9277), .A2(n5385), .ZN(n5398) );
  OR2_X1 U6321 ( .A1(n5284), .A2(n8845), .ZN(n5286) );
  NAND2_X1 U6322 ( .A1(n5205), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5223) );
  NOR2_X1 U6323 ( .A1(n5062), .A2(n5061), .ZN(n5064) );
  NOR2_X1 U6324 ( .A1(n5416), .A2(n7761), .ZN(n6452) );
  INV_X1 U6325 ( .A(n7098), .ZN(n7198) );
  NAND2_X1 U6326 ( .A1(n5216), .A2(n5215), .ZN(n5232) );
  INV_X1 U6327 ( .A(n8625), .ZN(n8074) );
  OR2_X1 U6328 ( .A1(n8487), .A2(n6298), .ZN(n8028) );
  NAND2_X1 U6329 ( .A1(n5603), .A2(n6552), .ZN(n6504) );
  OR2_X1 U6330 ( .A1(n6242), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6253) );
  OR2_X1 U6331 ( .A1(n6234), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6242) );
  INV_X1 U6332 ( .A(n8622), .ZN(n8616) );
  INV_X1 U6333 ( .A(n8318), .ZN(n6072) );
  OR2_X1 U6334 ( .A1(n8490), .A2(n8489), .ZN(n8676) );
  NAND2_X1 U6335 ( .A1(n8574), .A2(n6363), .ZN(n6364) );
  NAND2_X1 U6336 ( .A1(n7323), .A2(n8212), .ZN(n7443) );
  INV_X1 U6337 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8743) );
  INV_X1 U6338 ( .A(n7474), .ZN(n7489) );
  AND2_X1 U6339 ( .A1(n5963), .A2(n6801), .ZN(n5965) );
  INV_X1 U6340 ( .A(n5730), .ZN(n5956) );
  AND2_X1 U6341 ( .A1(n5399), .A2(n5418), .ZN(n5964) );
  NOR2_X1 U6342 ( .A1(n5241), .A2(n5240), .ZN(n5259) );
  INV_X1 U6343 ( .A(n6465), .ZN(n8968) );
  AND2_X1 U6344 ( .A1(n7911), .A2(n6466), .ZN(n6467) );
  AOI22_X1 U6345 ( .A1(n8983), .A2(n7762), .B1(n5493), .B2(n8994), .ZN(n6444)
         );
  INV_X1 U6346 ( .A(n9767), .ZN(n9734) );
  INV_X1 U6347 ( .A(n5781), .ZN(n9714) );
  OR2_X1 U6348 ( .A1(n5497), .A2(n6801), .ZN(n9622) );
  XNOR2_X1 U6349 ( .A(n5194), .B(n9300), .ZN(n5193) );
  NAND2_X1 U6350 ( .A1(n6012), .A2(n4913), .ZN(n4938) );
  INV_X1 U6351 ( .A(n8555), .ZN(n8532) );
  INV_X1 U6352 ( .A(n8138), .ZN(n8092) );
  OR2_X1 U6353 ( .A1(n6063), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6075) );
  INV_X1 U6354 ( .A(n8359), .ZN(n8373) );
  AND3_X1 U6355 ( .A1(n6238), .A2(n6237), .A3(n6236), .ZN(n8542) );
  AND4_X1 U6356 ( .A1(n6192), .A2(n6191), .A3(n6190), .A4(n6189), .ZN(n8139)
         );
  INV_X1 U6357 ( .A(n9831), .ZN(n9841) );
  INV_X1 U6358 ( .A(n9890), .ZN(n8166) );
  NAND2_X1 U6359 ( .A1(n8355), .A2(n6377), .ZN(n9861) );
  INV_X1 U6360 ( .A(n8672), .ZN(n8658) );
  AND2_X1 U6361 ( .A1(n6375), .A2(n6341), .ZN(n6389) );
  AND2_X1 U6362 ( .A1(n7527), .A2(n7526), .ZN(n7534) );
  AND2_X1 U6363 ( .A1(n7308), .A2(n7281), .ZN(n9906) );
  NAND2_X1 U6364 ( .A1(n7364), .A2(n9915), .ZN(n9921) );
  XNOR2_X1 U6365 ( .A(n5529), .B(n4846), .ZN(n6746) );
  INV_X1 U6366 ( .A(n9602), .ZN(n9591) );
  INV_X1 U6367 ( .A(n9575), .ZN(n9598) );
  INV_X1 U6368 ( .A(n7928), .ZN(n9027) );
  AND2_X1 U6369 ( .A1(n7705), .A2(n7704), .ZN(n9046) );
  AND2_X1 U6370 ( .A1(n7688), .A2(n7867), .ZN(n9109) );
  INV_X1 U6371 ( .A(n8982), .ZN(n9669) );
  INV_X1 U6372 ( .A(n9618), .ZN(n9651) );
  INV_X1 U6373 ( .A(n9660), .ZN(n7202) );
  AND2_X1 U6374 ( .A1(n5434), .A2(n9382), .ZN(n6486) );
  INV_X1 U6375 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6474) );
  INV_X1 U6376 ( .A(n9773), .ZN(n9222) );
  INV_X1 U6377 ( .A(n6486), .ZN(n6473) );
  XNOR2_X1 U6378 ( .A(n5112), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9531) );
  INV_X1 U6379 ( .A(n6085), .ZN(n9903) );
  AND2_X1 U6380 ( .A1(n8300), .A2(n6311), .ZN(n8030) );
  INV_X1 U6381 ( .A(n8542), .ZN(n8567) );
  INV_X1 U6382 ( .A(n8139), .ZN(n8626) );
  NAND2_X1 U6383 ( .A1(P2_U3893), .A2(n8370), .ZN(n9844) );
  AND4_X1 U6384 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n8431)
         );
  NAND2_X1 U6385 ( .A1(n8608), .A2(n6395), .ZN(n8615) );
  NAND2_X1 U6386 ( .A1(n9952), .A2(n9931), .ZN(n8672) );
  NAND2_X1 U6387 ( .A1(n9952), .A2(n9921), .ZN(n8673) );
  INV_X1 U6388 ( .A(n9952), .ZN(n9950) );
  OR2_X1 U6389 ( .A1(n9934), .A2(n9926), .ZN(n8738) );
  INV_X2 U6390 ( .A(n9934), .ZN(n9932) );
  AND2_X1 U6391 ( .A1(n6746), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6595) );
  INV_X1 U6392 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7300) );
  INV_X1 U6393 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6774) );
  INV_X1 U6394 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6554) );
  INV_X1 U6395 ( .A(n9204), .ZN(n9103) );
  INV_X1 U6396 ( .A(n7100), .ZN(n9757) );
  INV_X1 U6397 ( .A(n9178), .ZN(n9030) );
  INV_X1 U6398 ( .A(n8894), .ZN(n8851) );
  INV_X1 U6399 ( .A(n8876), .ZN(n8897) );
  NAND4_X1 U6400 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n9020)
         );
  OR2_X1 U6401 ( .A1(n6641), .A2(n6640), .ZN(n9602) );
  INV_X1 U6402 ( .A(n9486), .ZN(n9613) );
  OR2_X1 U6403 ( .A1(n9658), .A2(n5499), .ZN(n9152) );
  INV_X2 U6404 ( .A(n9113), .ZN(n9658) );
  NAND2_X1 U6405 ( .A1(n5501), .A2(n9104), .ZN(n9113) );
  INV_X1 U6406 ( .A(n9803), .ZN(n9800) );
  OR2_X1 U6407 ( .A1(n9777), .A2(n6474), .ZN(n6475) );
  INV_X1 U6408 ( .A(n9777), .ZN(n9775) );
  INV_X1 U6409 ( .A(n9678), .ZN(n9679) );
  INV_X1 U6410 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7296) );
  INV_X1 U6411 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6605) );
  INV_X1 U6412 ( .A(n9386), .ZN(n9392) );
  INV_X1 U6413 ( .A(n8474), .ZN(P2_U3893) );
  INV_X1 U6414 ( .A(n8913), .ZN(P1_U3973) );
  NAND2_X1 U6415 ( .A1(n4865), .A2(n4878), .ZN(P1_U3265) );
  NOR2_X1 U6416 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4883) );
  NAND4_X1 U6417 ( .A1(n4883), .A2(n4882), .A3(n4881), .A4(n4880), .ZN(n4884)
         );
  NOR2_X1 U6418 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4888) );
  NOR2_X1 U6419 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4887) );
  NOR2_X1 U6420 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4886) );
  NAND4_X1 U6421 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n4890)
         );
  NAND2_X1 U6422 ( .A1(n4894), .A2(n4892), .ZN(n4896) );
  INV_X1 U6423 ( .A(n4899), .ZN(n9389) );
  AND2_X2 U6424 ( .A1(n9389), .A2(n9396), .ZN(n4967) );
  NAND2_X1 U6425 ( .A1(n4951), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U6426 ( .A1(n5001), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U6427 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n4907) );
  NAND2_X1 U6428 ( .A1(n5432), .A2(n4907), .ZN(n4908) );
  INV_X1 U6429 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4909) );
  OR2_X1 U6430 ( .A1(n7751), .A2(n4909), .ZN(n4920) );
  AND2_X1 U6431 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4912) );
  NAND2_X1 U6432 ( .A1(n6008), .A2(n4912), .ZN(n6012) );
  AND2_X1 U6433 ( .A1(n4941), .A2(SI_0_), .ZN(n4926) );
  NAND2_X1 U6434 ( .A1(n4926), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4913) );
  XNOR2_X1 U6435 ( .A(n4937), .B(n4938), .ZN(n5998) );
  INV_X1 U6436 ( .A(n5998), .ZN(n6536) );
  OR2_X1 U6437 ( .A1(n5071), .A2(n6536), .ZN(n4919) );
  INV_X1 U6438 ( .A(n5015), .ZN(n4917) );
  INV_X1 U6439 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4915) );
  NAND2_X1 U6440 ( .A1(n4917), .A2(n4916), .ZN(n4918) );
  NAND3_X1 U6441 ( .A1(n4920), .A2(n4919), .A3(n4918), .ZN(n4929) );
  INV_X2 U6442 ( .A(n4929), .ZN(n9683) );
  INV_X1 U6443 ( .A(n6903), .ZN(n4928) );
  NAND2_X1 U6444 ( .A1(n4966), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U6445 ( .A1(n4967), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U6446 ( .A1(n5001), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U6447 ( .A1(n4951), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4921) );
  INV_X1 U6448 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4925) );
  XNOR2_X1 U6449 ( .A(n4926), .B(n4925), .ZN(n9397) );
  INV_X1 U6450 ( .A(n6908), .ZN(n6671) );
  NAND2_X1 U6451 ( .A1(n4928), .A2(n6910), .ZN(n4931) );
  INV_X1 U6452 ( .A(n5732), .ZN(n6819) );
  NAND2_X1 U6453 ( .A1(n6819), .A2(n6907), .ZN(n4930) );
  NAND2_X1 U6454 ( .A1(n4967), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U6455 ( .A1(n4951), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6456 ( .A1(n5001), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4932) );
  INV_X1 U6457 ( .A(n6618), .ZN(n9471) );
  NAND2_X1 U6458 ( .A1(n4939), .A2(SI_1_), .ZN(n4940) );
  MUX2_X1 U6459 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4941), .Z(n4959) );
  INV_X1 U6460 ( .A(SI_2_), .ZN(n4942) );
  XNOR2_X1 U6461 ( .A(n4959), .B(n4942), .ZN(n4957) );
  XNOR2_X1 U6462 ( .A(n4958), .B(n4957), .ZN(n6535) );
  OR2_X1 U6463 ( .A1(n5071), .A2(n6535), .ZN(n4944) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6534) );
  XNOR2_X1 U6465 ( .A(n6911), .B(n9689), .ZN(n7763) );
  INV_X1 U6466 ( .A(n7763), .ZN(n4945) );
  NAND2_X1 U6467 ( .A1(n6817), .A2(n4945), .ZN(n4948) );
  INV_X1 U6468 ( .A(n6911), .ZN(n7835) );
  NAND2_X1 U6469 ( .A1(n7835), .A2(n7834), .ZN(n4947) );
  NAND2_X1 U6470 ( .A1(n4967), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n4950) );
  NAND2_X1 U6471 ( .A1(n4966), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U6472 ( .A1(n7732), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U6473 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4955), .ZN(n4956) );
  XNOR2_X1 U6474 ( .A(n4956), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6624) );
  INV_X1 U6475 ( .A(n6624), .ZN(n9435) );
  NAND2_X1 U6476 ( .A1(n4958), .A2(n4957), .ZN(n4961) );
  NAND2_X1 U6477 ( .A1(n4959), .A2(SI_2_), .ZN(n4960) );
  NAND2_X1 U6478 ( .A1(n4961), .A2(n4960), .ZN(n4977) );
  INV_X1 U6479 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6548) );
  INV_X1 U6480 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6533) );
  MUX2_X1 U6481 ( .A(n6548), .B(n6533), .S(n7746), .Z(n4978) );
  XNOR2_X1 U6482 ( .A(n4978), .B(SI_3_), .ZN(n4962) );
  XNOR2_X1 U6483 ( .A(n4977), .B(n4962), .ZN(n6547) );
  OR2_X1 U6484 ( .A1(n5071), .A2(n6547), .ZN(n4964) );
  OR2_X1 U6485 ( .A1(n7751), .A2(n6533), .ZN(n4963) );
  OAI211_X1 U6486 ( .C1(n5015), .C2(n9435), .A(n4964), .B(n4963), .ZN(n5755)
         );
  NAND2_X1 U6487 ( .A1(n6820), .A2(n5755), .ZN(n5461) );
  INV_X1 U6488 ( .A(n5461), .ZN(n4965) );
  NAND2_X1 U6489 ( .A1(n5754), .A2(n9695), .ZN(n7838) );
  NAND2_X1 U6490 ( .A1(n4966), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U6491 ( .A1(n4967), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4971) );
  INV_X1 U6492 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n4968) );
  XNOR2_X1 U6493 ( .A(n4968), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U6494 ( .A1(n5001), .A2(n9657), .ZN(n4970) );
  NAND2_X1 U6495 ( .A1(n7732), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U6496 ( .A1(n4973), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4974) );
  XNOR2_X1 U6497 ( .A(n4974), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6627) );
  INV_X1 U6498 ( .A(n6627), .ZN(n9496) );
  INV_X1 U6499 ( .A(SI_3_), .ZN(n4975) );
  NAND2_X1 U6500 ( .A1(n4978), .A2(n4975), .ZN(n4976) );
  NAND2_X1 U6501 ( .A1(n4977), .A2(n4976), .ZN(n4981) );
  INV_X1 U6502 ( .A(n4978), .ZN(n4979) );
  NAND2_X1 U6503 ( .A1(n4979), .A2(SI_3_), .ZN(n4980) );
  NAND2_X1 U6504 ( .A1(n4981), .A2(n4980), .ZN(n4991) );
  INV_X1 U6505 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6550) );
  INV_X1 U6506 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6537) );
  MUX2_X1 U6507 ( .A(n6550), .B(n6537), .S(n7746), .Z(n4992) );
  XNOR2_X1 U6508 ( .A(n4992), .B(SI_4_), .ZN(n4990) );
  XNOR2_X1 U6509 ( .A(n4991), .B(n4990), .ZN(n6549) );
  OR2_X1 U6510 ( .A1(n5071), .A2(n6549), .ZN(n4983) );
  OR2_X1 U6511 ( .A1(n7751), .A2(n6537), .ZN(n4982) );
  OAI211_X1 U6512 ( .C1(n5015), .C2(n9496), .A(n4983), .B(n4982), .ZN(n5762)
         );
  NAND2_X1 U6513 ( .A1(n6956), .A2(n5762), .ZN(n5464) );
  INV_X1 U6514 ( .A(n5762), .ZN(n9701) );
  NAND2_X1 U6515 ( .A1(n8912), .A2(n9701), .ZN(n7839) );
  NAND2_X1 U6516 ( .A1(n4967), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6517 ( .A1(n7731), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4987) );
  AOI21_X1 U6518 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n4984) );
  NOR2_X1 U6519 ( .A1(n4984), .A2(n5002), .ZN(n6962) );
  NAND2_X1 U6520 ( .A1(n5340), .A2(n6962), .ZN(n4986) );
  NAND2_X1 U6521 ( .A1(n7732), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4985) );
  INV_X1 U6522 ( .A(n9653), .ZN(n5468) );
  NOR2_X1 U6523 ( .A1(n4973), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5017) );
  OR2_X1 U6524 ( .A1(n5017), .A2(n9384), .ZN(n4989) );
  XNOR2_X1 U6525 ( .A(n4989), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6630) );
  INV_X1 U6526 ( .A(n6630), .ZN(n9511) );
  NAND2_X1 U6527 ( .A1(n4991), .A2(n4990), .ZN(n4995) );
  INV_X1 U6528 ( .A(n4992), .ZN(n4993) );
  NAND2_X1 U6529 ( .A1(n4993), .A2(SI_4_), .ZN(n4994) );
  NAND2_X1 U6530 ( .A1(n4995), .A2(n4994), .ZN(n5010) );
  INV_X1 U6531 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6539) );
  INV_X1 U6532 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6540) );
  MUX2_X1 U6533 ( .A(n6539), .B(n6540), .S(n7746), .Z(n5011) );
  XNOR2_X1 U6534 ( .A(n5011), .B(SI_5_), .ZN(n4996) );
  XNOR2_X1 U6535 ( .A(n5010), .B(n4996), .ZN(n6541) );
  OR2_X1 U6536 ( .A1(n6541), .A2(n5071), .ZN(n4998) );
  OR2_X1 U6537 ( .A1(n7751), .A2(n6540), .ZN(n4997) );
  OAI211_X1 U6538 ( .C1(n5015), .C2(n9511), .A(n4998), .B(n4997), .ZN(n6961)
         );
  NAND2_X1 U6539 ( .A1(n5468), .A2(n6961), .ZN(n5467) );
  NAND2_X1 U6540 ( .A1(n6954), .A2(n5467), .ZN(n4999) );
  INV_X1 U6541 ( .A(n6961), .ZN(n9708) );
  NAND2_X1 U6542 ( .A1(n9653), .A2(n9708), .ZN(n7840) );
  NAND2_X1 U6543 ( .A1(n4967), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U6544 ( .A1(n7731), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U6545 ( .A1(n5002), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5062) );
  OAI21_X1 U6546 ( .B1(n5002), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5062), .ZN(
        n5003) );
  INV_X1 U6547 ( .A(n5003), .ZN(n9639) );
  NAND2_X1 U6548 ( .A1(n5340), .A2(n9639), .ZN(n5005) );
  NAND2_X1 U6549 ( .A1(n7732), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5004) );
  NAND4_X1 U6550 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n8911)
         );
  INV_X1 U6551 ( .A(n8911), .ZN(n6957) );
  INV_X1 U6552 ( .A(SI_5_), .ZN(n5008) );
  NAND2_X1 U6553 ( .A1(n5011), .A2(n5008), .ZN(n5009) );
  INV_X1 U6554 ( .A(n5011), .ZN(n5012) );
  NAND2_X1 U6555 ( .A1(n5012), .A2(SI_5_), .ZN(n5013) );
  INV_X1 U6556 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6545) );
  INV_X1 U6557 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6542) );
  MUX2_X1 U6558 ( .A(n6545), .B(n6542), .S(n7725), .Z(n5025) );
  XNOR2_X1 U6559 ( .A(n5024), .B(n5023), .ZN(n6544) );
  OR2_X1 U6560 ( .A1(n6544), .A2(n5071), .ZN(n5022) );
  INV_X1 U6561 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6562 ( .A1(n5017), .A2(n5016), .ZN(n5039) );
  NAND2_X1 U6563 ( .A1(n5039), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5019) );
  INV_X1 U6564 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U6565 ( .A1(n5019), .A2(n5018), .ZN(n5072) );
  OR2_X1 U6566 ( .A1(n5019), .A2(n5018), .ZN(n5020) );
  AOI22_X1 U6567 ( .A1(n5256), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6560), .B2(
        n6633), .ZN(n5021) );
  NAND2_X1 U6568 ( .A1(n5022), .A2(n5021), .ZN(n5781) );
  NAND2_X1 U6569 ( .A1(n6957), .A2(n5781), .ZN(n7768) );
  NAND2_X1 U6570 ( .A1(n7639), .A2(n7768), .ZN(n7008) );
  INV_X1 U6571 ( .A(n5025), .ZN(n5026) );
  INV_X1 U6572 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6551) );
  MUX2_X1 U6573 ( .A(n6554), .B(n6551), .S(n7725), .Z(n5027) );
  XNOR2_X1 U6574 ( .A(n5027), .B(SI_7_), .ZN(n5070) );
  INV_X1 U6575 ( .A(n5027), .ZN(n5028) );
  NAND2_X1 U6576 ( .A1(n5028), .A2(SI_7_), .ZN(n5029) );
  MUX2_X1 U6577 ( .A(n6559), .B(n6556), .S(n7725), .Z(n5031) );
  INV_X1 U6578 ( .A(SI_8_), .ZN(n5030) );
  NAND2_X1 U6579 ( .A1(n5031), .A2(n5030), .ZN(n5034) );
  INV_X1 U6580 ( .A(n5031), .ZN(n5032) );
  NAND2_X1 U6581 ( .A1(n5032), .A2(SI_8_), .ZN(n5033) );
  NAND2_X1 U6582 ( .A1(n5034), .A2(n5033), .ZN(n5050) );
  MUX2_X1 U6583 ( .A(n6567), .B(n6571), .S(n7725), .Z(n5036) );
  INV_X1 U6584 ( .A(SI_9_), .ZN(n5035) );
  NAND2_X1 U6585 ( .A1(n5036), .A2(n5035), .ZN(n5082) );
  INV_X1 U6586 ( .A(n5036), .ZN(n5037) );
  NAND2_X1 U6587 ( .A1(n5037), .A2(SI_9_), .ZN(n5038) );
  NAND2_X1 U6588 ( .A1(n6566), .A2(n5318), .ZN(n5042) );
  NAND2_X1 U6589 ( .A1(n5085), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5040) );
  XNOR2_X1 U6590 ( .A(n5040), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6846) );
  AOI22_X1 U6591 ( .A1(n5256), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6560), .B2(
        n6846), .ZN(n5041) );
  NAND2_X1 U6592 ( .A1(n7731), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6593 ( .A1(n4967), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6594 ( .A1(n5064), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6595 ( .A1(n5056), .A2(n5043), .ZN(n5044) );
  AND2_X1 U6596 ( .A1(n5092), .A2(n5044), .ZN(n7264) );
  NAND2_X1 U6597 ( .A1(n5340), .A2(n7264), .ZN(n5046) );
  NAND2_X1 U6598 ( .A1(n7732), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5045) );
  NAND4_X1 U6599 ( .A1(n5048), .A2(n5047), .A3(n5046), .A4(n5045), .ZN(n8909)
         );
  INV_X1 U6600 ( .A(n8909), .ZN(n9617) );
  XNOR2_X1 U6601 ( .A(n5049), .B(n5050), .ZN(n6555) );
  NAND2_X1 U6602 ( .A1(n6555), .A2(n5318), .ZN(n5054) );
  NAND2_X1 U6603 ( .A1(n5051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5052) );
  XNOR2_X1 U6604 ( .A(n5052), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6637) );
  AOI22_X1 U6605 ( .A1(n5256), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6560), .B2(
        n6637), .ZN(n5053) );
  NAND2_X1 U6606 ( .A1(n5054), .A2(n5053), .ZN(n7181) );
  NAND2_X1 U6607 ( .A1(n4967), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6608 ( .A1(n4966), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5059) );
  OR2_X1 U6609 ( .A1(n5064), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5055) );
  AND2_X1 U6610 ( .A1(n5056), .A2(n5055), .ZN(n9626) );
  NAND2_X1 U6611 ( .A1(n5340), .A2(n9626), .ZN(n5058) );
  NAND2_X1 U6612 ( .A1(n7732), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5057) );
  NAND4_X1 U6613 ( .A1(n5060), .A2(n5059), .A3(n5058), .A4(n5057), .ZN(n8910)
         );
  INV_X1 U6614 ( .A(n8910), .ZN(n7265) );
  OR2_X1 U6615 ( .A1(n7181), .A2(n7265), .ZN(n7644) );
  NAND2_X1 U6616 ( .A1(n7648), .A2(n7644), .ZN(n7653) );
  NAND2_X1 U6617 ( .A1(n7731), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6618 ( .A1(n4967), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5067) );
  AND2_X1 U6619 ( .A1(n5062), .A2(n5061), .ZN(n5063) );
  NOR2_X1 U6620 ( .A1(n5064), .A2(n5063), .ZN(n7042) );
  NAND2_X1 U6621 ( .A1(n5340), .A2(n7042), .ZN(n5066) );
  NAND2_X1 U6622 ( .A1(n7732), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5065) );
  NAND4_X1 U6623 ( .A1(n5068), .A2(n5067), .A3(n5066), .A4(n5065), .ZN(n9637)
         );
  XNOR2_X1 U6624 ( .A(n5069), .B(n5070), .ZN(n6553) );
  OR2_X1 U6625 ( .A1(n6553), .A2(n5071), .ZN(n5075) );
  NAND2_X1 U6626 ( .A1(n5072), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5073) );
  XNOR2_X1 U6627 ( .A(n5073), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6635) );
  AOI22_X1 U6628 ( .A1(n5256), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6560), .B2(
        n6635), .ZN(n5074) );
  NAND2_X1 U6629 ( .A1(n5075), .A2(n5074), .ZN(n7045) );
  NAND2_X1 U6630 ( .A1(n9714), .A2(n8911), .ZN(n7640) );
  NAND2_X1 U6631 ( .A1(n7643), .A2(n7640), .ZN(n5076) );
  NOR2_X1 U6632 ( .A1(n7653), .A2(n5076), .ZN(n7844) );
  NAND2_X1 U6633 ( .A1(n7008), .A2(n7844), .ZN(n5080) );
  INV_X1 U6634 ( .A(n7653), .ZN(n5077) );
  NAND2_X1 U6635 ( .A1(n7181), .A2(n7265), .ZN(n7646) );
  NAND2_X1 U6636 ( .A1(n7045), .A2(n9619), .ZN(n7009) );
  NAND2_X1 U6637 ( .A1(n5077), .A2(n4874), .ZN(n5079) );
  NAND2_X1 U6638 ( .A1(n5078), .A2(n9617), .ZN(n7652) );
  AND2_X1 U6639 ( .A1(n5079), .A2(n7652), .ZN(n7772) );
  NAND2_X1 U6640 ( .A1(n5081), .A2(n4289), .ZN(n5083) );
  INV_X1 U6641 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5084) );
  MUX2_X1 U6642 ( .A(n6580), .B(n5084), .S(n7725), .Z(n5100) );
  XNOR2_X1 U6643 ( .A(n5100), .B(SI_10_), .ZN(n5099) );
  XNOR2_X1 U6644 ( .A(n5104), .B(n5099), .ZN(n6568) );
  NAND2_X1 U6645 ( .A1(n6568), .A2(n5318), .ZN(n5090) );
  OAI21_X1 U6646 ( .B1(n5085), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5087) );
  INV_X1 U6647 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6648 ( .A1(n5087), .A2(n5086), .ZN(n5111) );
  OR2_X1 U6649 ( .A1(n5087), .A2(n5086), .ZN(n5088) );
  AOI22_X1 U6650 ( .A1(n5256), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6560), .B2(
        n9406), .ZN(n5089) );
  NAND2_X1 U6651 ( .A1(n7733), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6652 ( .A1(n7731), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6653 ( .A1(n5092), .A2(n5091), .ZN(n5093) );
  AND2_X1 U6654 ( .A1(n5116), .A2(n5093), .ZN(n7427) );
  NAND2_X1 U6655 ( .A1(n5340), .A2(n7427), .ZN(n5095) );
  NAND2_X1 U6656 ( .A1(n7732), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5094) );
  NAND4_X1 U6657 ( .A1(n5097), .A2(n5096), .A3(n5095), .A4(n5094), .ZN(n8908)
         );
  INV_X1 U6658 ( .A(n8908), .ZN(n5098) );
  OR2_X1 U6659 ( .A1(n5476), .A2(n5098), .ZN(n7845) );
  NAND2_X1 U6660 ( .A1(n5476), .A2(n5098), .ZN(n7655) );
  NAND2_X1 U6661 ( .A1(n7845), .A2(n7655), .ZN(n6997) );
  NAND2_X1 U6662 ( .A1(n7842), .A2(n7773), .ZN(n7078) );
  INV_X1 U6663 ( .A(n5099), .ZN(n5103) );
  INV_X1 U6664 ( .A(n5100), .ZN(n5101) );
  NAND2_X1 U6665 ( .A1(n5101), .A2(SI_10_), .ZN(n5102) );
  INV_X1 U6666 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5106) );
  INV_X1 U6667 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5105) );
  MUX2_X1 U6668 ( .A(n5106), .B(n5105), .S(n7725), .Z(n5108) );
  INV_X1 U6669 ( .A(SI_11_), .ZN(n5107) );
  INV_X1 U6670 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6671 ( .A1(n5109), .A2(SI_11_), .ZN(n5110) );
  NAND2_X1 U6672 ( .A1(n5124), .A2(n5110), .ZN(n5125) );
  NAND2_X1 U6673 ( .A1(n6583), .A2(n5318), .ZN(n5114) );
  NAND2_X1 U6674 ( .A1(n5111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5112) );
  AOI22_X1 U6675 ( .A1(n5256), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6560), .B2(
        n9531), .ZN(n5113) );
  NAND2_X1 U6676 ( .A1(n7731), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6677 ( .A1(n7733), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5120) );
  AND2_X1 U6678 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  NOR2_X1 U6679 ( .A1(n5132), .A2(n5117), .ZN(n7488) );
  NAND2_X1 U6680 ( .A1(n5340), .A2(n7488), .ZN(n5119) );
  NAND2_X1 U6681 ( .A1(n7732), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5118) );
  NAND4_X1 U6682 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n8907)
         );
  INV_X1 U6683 ( .A(n8907), .ZN(n7400) );
  NAND2_X1 U6684 ( .A1(n7086), .A2(n7400), .ZN(n7656) );
  NAND2_X1 U6685 ( .A1(n7078), .A2(n5122), .ZN(n5123) );
  NAND2_X1 U6686 ( .A1(n5123), .A2(n7848), .ZN(n7092) );
  MUX2_X1 U6687 ( .A(n5127), .B(n6605), .S(n7725), .Z(n5139) );
  XNOR2_X1 U6688 ( .A(n5139), .B(SI_12_), .ZN(n5138) );
  XNOR2_X1 U6689 ( .A(n5142), .B(n5138), .ZN(n6599) );
  NAND2_X1 U6690 ( .A1(n6599), .A2(n5318), .ZN(n5131) );
  OR2_X1 U6691 ( .A1(n5128), .A2(n9384), .ZN(n5129) );
  XNOR2_X1 U6692 ( .A(n5129), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8934) );
  AOI22_X1 U6693 ( .A1(n5256), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6560), .B2(
        n8934), .ZN(n5130) );
  NAND2_X1 U6694 ( .A1(n4967), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6695 ( .A1(n4966), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5136) );
  OR2_X1 U6696 ( .A1(n5132), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6697 ( .A1(n5132), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5148) );
  AND2_X1 U6698 ( .A1(n5133), .A2(n5148), .ZN(n7399) );
  NAND2_X1 U6699 ( .A1(n5340), .A2(n7399), .ZN(n5135) );
  NAND2_X1 U6700 ( .A1(n7732), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5134) );
  NAND4_X1 U6701 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), .ZN(n7474)
         );
  OR2_X1 U6702 ( .A1(n7100), .A2(n7489), .ZN(n7658) );
  NAND2_X1 U6703 ( .A1(n7100), .A2(n7489), .ZN(n7852) );
  NAND2_X1 U6704 ( .A1(n7658), .A2(n7852), .ZN(n7093) );
  INV_X1 U6705 ( .A(n7093), .ZN(n7775) );
  INV_X1 U6706 ( .A(n7658), .ZN(n7851) );
  AOI21_X1 U6707 ( .B1(n7092), .B2(n7775), .A(n7851), .ZN(n7191) );
  INV_X1 U6708 ( .A(n5139), .ZN(n5140) );
  MUX2_X1 U6709 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7725), .Z(n5157) );
  XNOR2_X1 U6710 ( .A(n5157), .B(SI_13_), .ZN(n5154) );
  XNOR2_X1 U6711 ( .A(n5156), .B(n5154), .ZN(n6607) );
  NAND2_X1 U6712 ( .A1(n6607), .A2(n5318), .ZN(n5146) );
  NAND2_X1 U6713 ( .A1(n5143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5144) );
  XNOR2_X1 U6714 ( .A(n5144), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9556) );
  AOI22_X1 U6715 ( .A1(n5256), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6560), .B2(
        n9556), .ZN(n5145) );
  NAND2_X1 U6716 ( .A1(n7733), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U6717 ( .A1(n7732), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6718 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  AND2_X1 U6719 ( .A1(n5171), .A2(n5149), .ZN(n7196) );
  NAND2_X1 U6720 ( .A1(n5340), .A2(n7196), .ZN(n5151) );
  NAND2_X1 U6721 ( .A1(n7731), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5150) );
  NAND4_X1 U6722 ( .A1(n5153), .A2(n5152), .A3(n5151), .A4(n5150), .ZN(n8906)
         );
  INV_X1 U6723 ( .A(n8906), .ZN(n8757) );
  OR2_X1 U6724 ( .A1(n7201), .A2(n8757), .ZN(n7666) );
  NAND2_X1 U6725 ( .A1(n7201), .A2(n8757), .ZN(n7662) );
  AND2_X2 U6726 ( .A1(n7191), .A2(n7777), .ZN(n7250) );
  INV_X1 U6727 ( .A(n5154), .ZN(n5155) );
  NAND2_X1 U6728 ( .A1(n5156), .A2(n5155), .ZN(n5159) );
  NAND2_X1 U6729 ( .A1(n5157), .A2(SI_13_), .ZN(n5158) );
  MUX2_X1 U6730 ( .A(n6655), .B(n5160), .S(n7725), .Z(n5162) );
  INV_X1 U6731 ( .A(SI_14_), .ZN(n5161) );
  INV_X1 U6732 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6733 ( .A1(n5163), .A2(SI_14_), .ZN(n5164) );
  NAND2_X1 U6734 ( .A1(n5179), .A2(n5164), .ZN(n5180) );
  NAND2_X1 U6735 ( .A1(n6651), .A2(n5318), .ZN(n5169) );
  NAND2_X1 U6736 ( .A1(n4348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6737 ( .A1(n5166), .A2(n5165), .ZN(n5182) );
  OR2_X1 U6738 ( .A1(n5166), .A2(n5165), .ZN(n5167) );
  AOI22_X1 U6739 ( .A1(n5256), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6560), .B2(
        n9568), .ZN(n5168) );
  NAND2_X1 U6740 ( .A1(n5169), .A2(n5168), .ZN(n5177) );
  NAND2_X1 U6741 ( .A1(n7733), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6742 ( .A1(n7731), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5175) );
  AND2_X1 U6743 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  NOR2_X1 U6744 ( .A1(n5187), .A2(n5172), .ZN(n8755) );
  NAND2_X1 U6745 ( .A1(n5340), .A2(n8755), .ZN(n5174) );
  NAND2_X1 U6746 ( .A1(n7732), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5173) );
  NAND4_X1 U6747 ( .A1(n5176), .A2(n5175), .A3(n5174), .A4(n5173), .ZN(n8905)
         );
  OR2_X1 U6748 ( .A1(n5177), .A2(n8892), .ZN(n7661) );
  NAND2_X1 U6749 ( .A1(n5177), .A2(n8892), .ZN(n7663) );
  INV_X1 U6750 ( .A(n7662), .ZN(n7856) );
  MUX2_X1 U6751 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7725), .Z(n5194) );
  NAND2_X1 U6752 ( .A1(n5182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5184) );
  XNOR2_X1 U6753 ( .A(n5184), .B(n5183), .ZN(n8937) );
  INV_X1 U6754 ( .A(n8937), .ZN(n9581) );
  AOI22_X1 U6755 ( .A1(n5256), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6560), .B2(
        n9581), .ZN(n5185) );
  NAND2_X1 U6756 ( .A1(n4966), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6757 ( .A1(n4967), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5191) );
  NOR2_X1 U6758 ( .A1(n5187), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5188) );
  NOR2_X1 U6759 ( .A1(n5205), .A2(n5188), .ZN(n8888) );
  NAND2_X1 U6760 ( .A1(n5340), .A2(n8888), .ZN(n5190) );
  NAND2_X1 U6761 ( .A1(n7732), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5189) );
  NAND4_X1 U6762 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n8904)
         );
  NAND2_X1 U6763 ( .A1(n5194), .A2(SI_15_), .ZN(n5195) );
  MUX2_X1 U6764 ( .A(n6774), .B(n9274), .S(n7746), .Z(n5199) );
  INV_X1 U6765 ( .A(SI_16_), .ZN(n5198) );
  NAND2_X1 U6766 ( .A1(n5199), .A2(n5198), .ZN(n5211) );
  INV_X1 U6767 ( .A(n5199), .ZN(n5200) );
  NAND2_X1 U6768 ( .A1(n5200), .A2(SI_16_), .ZN(n5201) );
  NAND2_X1 U6769 ( .A1(n5211), .A2(n5201), .ZN(n5212) );
  XNOR2_X1 U6770 ( .A(n5213), .B(n5212), .ZN(n6770) );
  NAND2_X1 U6771 ( .A1(n6770), .A2(n5318), .ZN(n5204) );
  NAND2_X1 U6772 ( .A1(n4350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5202) );
  XNOR2_X1 U6773 ( .A(n5202), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8955) );
  AOI22_X1 U6774 ( .A1(n5256), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6560), .B2(
        n8955), .ZN(n5203) );
  NAND2_X1 U6775 ( .A1(n7733), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6776 ( .A1(n7731), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5209) );
  OR2_X1 U6777 ( .A1(n5205), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5206) );
  AND2_X1 U6778 ( .A1(n5223), .A2(n5206), .ZN(n8808) );
  NAND2_X1 U6779 ( .A1(n5340), .A2(n8808), .ZN(n5208) );
  NAND2_X1 U6780 ( .A1(n7732), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5207) );
  NAND4_X1 U6781 ( .A1(n5210), .A2(n5209), .A3(n5208), .A4(n5207), .ZN(n8903)
         );
  INV_X1 U6782 ( .A(n8903), .ZN(n9143) );
  NAND2_X1 U6783 ( .A1(n9219), .A2(n9143), .ZN(n7671) );
  INV_X1 U6784 ( .A(n7671), .ZN(n9141) );
  INV_X1 U6785 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5214) );
  MUX2_X1 U6786 ( .A(n6775), .B(n5214), .S(n7725), .Z(n5216) );
  INV_X1 U6787 ( .A(SI_17_), .ZN(n5215) );
  INV_X1 U6788 ( .A(n5216), .ZN(n5217) );
  NAND2_X1 U6789 ( .A1(n5217), .A2(SI_17_), .ZN(n5218) );
  XNOR2_X1 U6790 ( .A(n5231), .B(n5230), .ZN(n6733) );
  NAND2_X1 U6791 ( .A1(n6733), .A2(n5318), .ZN(n5221) );
  XNOR2_X1 U6792 ( .A(n5234), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9593) );
  AOI22_X1 U6793 ( .A1(n5256), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6560), .B2(
        n9593), .ZN(n5220) );
  NAND2_X1 U6794 ( .A1(n7733), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6795 ( .A1(n7731), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5227) );
  INV_X1 U6796 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6797 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  AND2_X1 U6798 ( .A1(n5241), .A2(n5224), .ZN(n9135) );
  NAND2_X1 U6799 ( .A1(n5340), .A2(n9135), .ZN(n5226) );
  NAND2_X1 U6800 ( .A1(n7732), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5225) );
  NAND4_X1 U6801 ( .A1(n5228), .A2(n5227), .A3(n5226), .A4(n5225), .ZN(n9124)
         );
  INV_X1 U6802 ( .A(n9124), .ZN(n7374) );
  OR2_X1 U6803 ( .A1(n9213), .A2(n7374), .ZN(n7677) );
  NAND2_X1 U6804 ( .A1(n9213), .A2(n7374), .ZN(n7679) );
  NAND2_X1 U6805 ( .A1(n7677), .A2(n7679), .ZN(n9140) );
  INV_X1 U6806 ( .A(n7677), .ZN(n5229) );
  NOR2_X1 U6807 ( .A1(n9139), .A2(n5229), .ZN(n9123) );
  INV_X1 U6808 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5233) );
  MUX2_X1 U6809 ( .A(n6919), .B(n5233), .S(n7725), .Z(n5246) );
  XNOR2_X1 U6810 ( .A(n5246), .B(SI_18_), .ZN(n5245) );
  XNOR2_X1 U6811 ( .A(n5250), .B(n5245), .ZN(n6799) );
  NAND2_X1 U6812 ( .A1(n6799), .A2(n5318), .ZN(n5239) );
  NAND2_X1 U6813 ( .A1(n5234), .A2(n5406), .ZN(n5235) );
  OR2_X1 U6814 ( .A1(n5236), .A2(n5405), .ZN(n5237) );
  AND2_X1 U6815 ( .A1(n5255), .A2(n5237), .ZN(n9606) );
  AOI22_X1 U6816 ( .A1(n5256), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6560), .B2(
        n9606), .ZN(n5238) );
  INV_X1 U6817 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5240) );
  AND2_X1 U6818 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  OR2_X1 U6819 ( .A1(n5242), .A2(n5259), .ZN(n8865) );
  AOI22_X1 U6820 ( .A1(n7731), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n7733), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6821 ( .A1(n7732), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5243) );
  OAI211_X1 U6822 ( .C1(n8865), .C2(n5287), .A(n5244), .B(n5243), .ZN(n8902)
         );
  INV_X1 U6823 ( .A(n8902), .ZN(n9144) );
  OR2_X1 U6824 ( .A1(n9208), .A2(n9144), .ZN(n7681) );
  NAND2_X1 U6825 ( .A1(n9208), .A2(n9144), .ZN(n7680) );
  NAND2_X1 U6826 ( .A1(n9123), .A2(n9122), .ZN(n9121) );
  NAND2_X2 U6827 ( .A1(n9121), .A2(n7680), .ZN(n9110) );
  INV_X1 U6828 ( .A(n5245), .ZN(n5249) );
  INV_X1 U6829 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6830 ( .A1(n5247), .A2(SI_18_), .ZN(n5248) );
  MUX2_X1 U6831 ( .A(n7068), .B(n7926), .S(n7725), .Z(n5252) );
  INV_X1 U6832 ( .A(SI_19_), .ZN(n5251) );
  NAND2_X1 U6833 ( .A1(n5252), .A2(n5251), .ZN(n5263) );
  INV_X1 U6834 ( .A(n5252), .ZN(n5253) );
  NAND2_X1 U6835 ( .A1(n5253), .A2(SI_19_), .ZN(n5254) );
  NAND2_X1 U6836 ( .A1(n5263), .A2(n5254), .ZN(n5264) );
  XNOR2_X1 U6837 ( .A(n5265), .B(n5264), .ZN(n7066) );
  NAND2_X1 U6838 ( .A1(n7066), .A2(n5318), .ZN(n5258) );
  AOI22_X1 U6839 ( .A1(n5256), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9027), .B2(
        n6560), .ZN(n5257) );
  NAND2_X1 U6840 ( .A1(n5259), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5284) );
  OR2_X1 U6841 ( .A1(n5259), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U6842 ( .A1(n5284), .A2(n5260), .ZN(n9105) );
  AOI22_X1 U6843 ( .A1(n7731), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n7733), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6844 ( .A1(n7732), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5261) );
  OAI211_X1 U6845 ( .C1(n9105), .C2(n5287), .A(n5262), .B(n5261), .ZN(n9125)
         );
  INV_X1 U6846 ( .A(n9125), .ZN(n9089) );
  OR2_X1 U6847 ( .A1(n9204), .A2(n9089), .ZN(n7688) );
  NAND2_X1 U6848 ( .A1(n9204), .A2(n9089), .ZN(n7867) );
  INV_X1 U6849 ( .A(n7867), .ZN(n7683) );
  MUX2_X1 U6850 ( .A(n9349), .B(n9350), .S(n7746), .Z(n5267) );
  INV_X1 U6851 ( .A(SI_20_), .ZN(n5266) );
  NAND2_X1 U6852 ( .A1(n5267), .A2(n5266), .ZN(n5270) );
  INV_X1 U6853 ( .A(n5267), .ZN(n5268) );
  NAND2_X1 U6854 ( .A1(n5268), .A2(SI_20_), .ZN(n5269) );
  NAND2_X1 U6855 ( .A1(n5281), .A2(n5280), .ZN(n5271) );
  MUX2_X1 U6856 ( .A(n7161), .B(n7169), .S(n7725), .Z(n5294) );
  XNOR2_X1 U6857 ( .A(n5294), .B(SI_21_), .ZN(n5293) );
  XNOR2_X1 U6858 ( .A(n5298), .B(n5293), .ZN(n7160) );
  NAND2_X1 U6859 ( .A1(n7160), .A2(n5318), .ZN(n5273) );
  OR2_X1 U6860 ( .A1(n7751), .A2(n7169), .ZN(n5272) );
  INV_X1 U6861 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8845) );
  INV_X1 U6862 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U6863 ( .A1(n5286), .A2(n8789), .ZN(n5274) );
  INV_X1 U6864 ( .A(n5305), .ZN(n5306) );
  NAND2_X1 U6865 ( .A1(n5274), .A2(n5306), .ZN(n9078) );
  OR2_X1 U6866 ( .A1(n9078), .A2(n5287), .ZN(n5279) );
  INV_X1 U6867 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U6868 ( .A1(n4967), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6869 ( .A1(n7732), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5275) );
  OAI211_X1 U6870 ( .C1(n9229), .C2(n5000), .A(n5276), .B(n5275), .ZN(n5277)
         );
  INV_X1 U6871 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6872 ( .A1(n5279), .A2(n5278), .ZN(n9059) );
  INV_X1 U6873 ( .A(n9059), .ZN(n9090) );
  OR2_X1 U6874 ( .A1(n9194), .A2(n9090), .ZN(n7695) );
  XNOR2_X1 U6875 ( .A(n5281), .B(n5280), .ZN(n7133) );
  NAND2_X1 U6876 ( .A1(n7133), .A2(n5318), .ZN(n5283) );
  OR2_X1 U6877 ( .A1(n7751), .A2(n9350), .ZN(n5282) );
  NAND2_X1 U6878 ( .A1(n5284), .A2(n8845), .ZN(n5285) );
  NAND2_X1 U6879 ( .A1(n5286), .A2(n5285), .ZN(n9092) );
  OR2_X1 U6880 ( .A1(n9092), .A2(n5287), .ZN(n5292) );
  INV_X1 U6881 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U6882 ( .A1(n7732), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6883 ( .A1(n7733), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5288) );
  OAI211_X1 U6884 ( .C1(n5000), .C2(n9236), .A(n5289), .B(n5288), .ZN(n5290)
         );
  INV_X1 U6885 ( .A(n5290), .ZN(n5291) );
  NAND2_X1 U6886 ( .A1(n5292), .A2(n5291), .ZN(n8901) );
  INV_X1 U6887 ( .A(n8901), .ZN(n9112) );
  OR2_X1 U6888 ( .A1(n9199), .A2(n9112), .ZN(n7687) );
  NAND2_X1 U6889 ( .A1(n7695), .A2(n7687), .ZN(n7804) );
  AND2_X1 U6890 ( .A1(n9199), .A2(n9112), .ZN(n7690) );
  AND2_X1 U6891 ( .A1(n9194), .A2(n9090), .ZN(n7697) );
  AOI21_X1 U6892 ( .B1(n7690), .B2(n7695), .A(n7697), .ZN(n7807) );
  INV_X1 U6893 ( .A(n5293), .ZN(n5297) );
  INV_X1 U6894 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U6895 ( .A1(n5295), .A2(SI_21_), .ZN(n5296) );
  MUX2_X1 U6896 ( .A(n9297), .B(n7233), .S(n7725), .Z(n5300) );
  INV_X1 U6897 ( .A(SI_22_), .ZN(n5299) );
  NAND2_X1 U6898 ( .A1(n5300), .A2(n5299), .ZN(n5311) );
  INV_X1 U6899 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U6900 ( .A1(n5301), .A2(SI_22_), .ZN(n5302) );
  NAND2_X1 U6901 ( .A1(n5311), .A2(n5302), .ZN(n5312) );
  XNOR2_X1 U6902 ( .A(n5313), .B(n5312), .ZN(n7232) );
  NAND2_X1 U6903 ( .A1(n7232), .A2(n5318), .ZN(n5304) );
  OR2_X1 U6904 ( .A1(n7751), .A2(n7233), .ZN(n5303) );
  NAND2_X1 U6905 ( .A1(n7733), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6906 ( .A1(n7731), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5309) );
  INV_X1 U6907 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8857) );
  NAND2_X1 U6908 ( .A1(n5305), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5322) );
  AOI21_X1 U6909 ( .B1(n8857), .B2(n5306), .A(n5321), .ZN(n9056) );
  NAND2_X1 U6910 ( .A1(n5340), .A2(n9056), .ZN(n5308) );
  NAND2_X1 U6911 ( .A1(n7732), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5307) );
  NAND4_X1 U6912 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n9047)
         );
  XNOR2_X1 U6913 ( .A(n9188), .B(n9074), .ZN(n9062) );
  NOR2_X1 U6914 ( .A1(n9188), .A2(n9074), .ZN(n7700) );
  MUX2_X1 U6915 ( .A(n7300), .B(n7296), .S(n7746), .Z(n5315) );
  INV_X1 U6916 ( .A(SI_23_), .ZN(n5314) );
  NAND2_X1 U6917 ( .A1(n5315), .A2(n5314), .ZN(n5329) );
  INV_X1 U6918 ( .A(n5315), .ZN(n5316) );
  NAND2_X1 U6919 ( .A1(n5316), .A2(SI_23_), .ZN(n5317) );
  NAND2_X1 U6920 ( .A1(n7297), .A2(n5318), .ZN(n5320) );
  OR2_X1 U6921 ( .A1(n7751), .A2(n7296), .ZN(n5319) );
  NAND2_X1 U6922 ( .A1(n4967), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6923 ( .A1(n7731), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5325) );
  INV_X1 U6924 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8770) );
  AOI21_X1 U6925 ( .B1(n8770), .B2(n5322), .A(n5337), .ZN(n9042) );
  NAND2_X1 U6926 ( .A1(n5340), .A2(n9042), .ZN(n5324) );
  NAND2_X1 U6927 ( .A1(n7732), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5323) );
  NAND4_X1 U6928 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n9065)
         );
  INV_X1 U6929 ( .A(n9065), .ZN(n8827) );
  OR2_X1 U6930 ( .A1(n9183), .A2(n8827), .ZN(n7705) );
  NAND2_X1 U6931 ( .A1(n9183), .A2(n8827), .ZN(n7704) );
  NAND2_X1 U6932 ( .A1(n9045), .A2(n9046), .ZN(n9044) );
  NAND2_X1 U6933 ( .A1(n5330), .A2(n5329), .ZN(n5346) );
  MUX2_X1 U6934 ( .A(n7382), .B(n7392), .S(n7725), .Z(n5332) );
  INV_X1 U6935 ( .A(SI_24_), .ZN(n5331) );
  NAND2_X1 U6936 ( .A1(n5332), .A2(n5331), .ZN(n5347) );
  INV_X1 U6937 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U6938 ( .A1(n5333), .A2(SI_24_), .ZN(n5334) );
  XNOR2_X1 U6939 ( .A(n5346), .B(n5345), .ZN(n7381) );
  NAND2_X1 U6940 ( .A1(n7381), .A2(n5318), .ZN(n5336) );
  OR2_X1 U6941 ( .A1(n7751), .A2(n7392), .ZN(n5335) );
  NAND2_X1 U6942 ( .A1(n7733), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6943 ( .A1(n7732), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5343) );
  INV_X1 U6944 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8826) );
  INV_X1 U6945 ( .A(n5354), .ZN(n5338) );
  AOI21_X1 U6946 ( .B1(n8826), .B2(n5339), .A(n5338), .ZN(n9028) );
  NAND2_X1 U6947 ( .A1(n5340), .A2(n9028), .ZN(n5342) );
  NAND2_X1 U6948 ( .A1(n7731), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5341) );
  NAND4_X1 U6949 ( .A1(n5344), .A2(n5343), .A3(n5342), .A4(n5341), .ZN(n9048)
         );
  NAND2_X1 U6950 ( .A1(n9178), .A2(n8798), .ZN(n7809) );
  NAND2_X1 U6951 ( .A1(n7799), .A2(n7809), .ZN(n9033) );
  INV_X1 U6952 ( .A(n7799), .ZN(n7710) );
  INV_X1 U6953 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7447) );
  INV_X1 U6954 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7449) );
  MUX2_X1 U6955 ( .A(n7447), .B(n7449), .S(n7725), .Z(n5349) );
  INV_X1 U6956 ( .A(SI_25_), .ZN(n5348) );
  NAND2_X1 U6957 ( .A1(n5349), .A2(n5348), .ZN(n5362) );
  INV_X1 U6958 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6959 ( .A1(n5350), .A2(SI_25_), .ZN(n5351) );
  XNOR2_X1 U6960 ( .A(n5361), .B(n5360), .ZN(n7446) );
  NAND2_X1 U6961 ( .A1(n7446), .A2(n5318), .ZN(n5353) );
  OR2_X1 U6962 ( .A1(n7751), .A2(n7449), .ZN(n5352) );
  NAND2_X1 U6963 ( .A1(n7733), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6964 ( .A1(n7731), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5357) );
  INV_X1 U6965 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8797) );
  AOI21_X1 U6966 ( .B1(n8797), .B2(n5354), .A(n5369), .ZN(n9013) );
  NAND2_X1 U6967 ( .A1(n5340), .A2(n9013), .ZN(n5356) );
  NAND2_X1 U6968 ( .A1(n7732), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5355) );
  NAND4_X1 U6969 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n9036)
         );
  INV_X1 U6970 ( .A(n9036), .ZN(n5491) );
  NAND2_X1 U6971 ( .A1(n9173), .A2(n5491), .ZN(n7810) );
  NAND2_X1 U6972 ( .A1(n7803), .A2(n7810), .ZN(n9017) );
  INV_X1 U6973 ( .A(n7803), .ZN(n5359) );
  NOR2_X1 U6974 ( .A1(n9016), .A2(n5359), .ZN(n9004) );
  INV_X1 U6975 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7478) );
  MUX2_X1 U6976 ( .A(n7478), .B(n9228), .S(n7725), .Z(n5364) );
  INV_X1 U6977 ( .A(SI_26_), .ZN(n5363) );
  NAND2_X1 U6978 ( .A1(n5364), .A2(n5363), .ZN(n5377) );
  INV_X1 U6979 ( .A(n5364), .ZN(n5365) );
  NAND2_X1 U6980 ( .A1(n5365), .A2(SI_26_), .ZN(n5366) );
  XNOR2_X1 U6981 ( .A(n5376), .B(n5375), .ZN(n7477) );
  NAND2_X1 U6982 ( .A1(n7477), .A2(n5318), .ZN(n5368) );
  OR2_X1 U6983 ( .A1(n7751), .A2(n9228), .ZN(n5367) );
  NAND2_X1 U6984 ( .A1(n5369), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5385) );
  OAI21_X1 U6985 ( .B1(n5369), .B2(P1_REG3_REG_26__SCAN_IN), .A(n5385), .ZN(
        n5370) );
  INV_X1 U6986 ( .A(n5370), .ZN(n8999) );
  NAND2_X1 U6987 ( .A1(n5340), .A2(n8999), .ZN(n5374) );
  NAND2_X1 U6988 ( .A1(n7733), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6989 ( .A1(n7732), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6990 ( .A1(n7731), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U6991 ( .A(n9168), .B(n9020), .ZN(n9003) );
  INV_X1 U6992 ( .A(n9020), .ZN(n7637) );
  NAND2_X1 U6993 ( .A1(n9168), .A2(n7637), .ZN(n7870) );
  NAND2_X1 U6994 ( .A1(n5378), .A2(n5377), .ZN(n5391) );
  INV_X1 U6995 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7541) );
  INV_X1 U6996 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7925) );
  MUX2_X1 U6997 ( .A(n7541), .B(n7925), .S(n7746), .Z(n5380) );
  INV_X1 U6998 ( .A(SI_27_), .ZN(n5379) );
  NAND2_X1 U6999 ( .A1(n5380), .A2(n5379), .ZN(n5392) );
  INV_X1 U7000 ( .A(n5380), .ZN(n5381) );
  NAND2_X1 U7001 ( .A1(n5381), .A2(SI_27_), .ZN(n5382) );
  NAND2_X1 U7002 ( .A1(n7540), .A2(n5318), .ZN(n5384) );
  OR2_X1 U7003 ( .A1(n7751), .A2(n7925), .ZN(n5383) );
  NAND2_X1 U7004 ( .A1(n7733), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U7005 ( .A1(n7732), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5388) );
  INV_X1 U7006 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9277) );
  AOI21_X1 U7007 ( .B1(n9277), .B2(n5385), .A(n5398), .ZN(n8991) );
  NAND2_X1 U7008 ( .A1(n5340), .A2(n8991), .ZN(n5387) );
  NAND2_X1 U7009 ( .A1(n7731), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5386) );
  NAND4_X1 U7010 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(n9005)
         );
  INV_X1 U7011 ( .A(n9005), .ZN(n5493) );
  NAND2_X1 U7012 ( .A1(n9164), .A2(n5493), .ZN(n7635) );
  NAND2_X1 U7013 ( .A1(n7798), .A2(n7635), .ZN(n7762) );
  NAND2_X1 U7014 ( .A1(n5391), .A2(n5390), .ZN(n5393) );
  NAND2_X1 U7015 ( .A1(n5393), .A2(n5392), .ZN(n6407) );
  INV_X1 U7016 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7592) );
  INV_X1 U7017 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7614) );
  MUX2_X1 U7018 ( .A(n7592), .B(n7614), .S(n7725), .Z(n6409) );
  XNOR2_X1 U7019 ( .A(n6409), .B(SI_28_), .ZN(n6406) );
  NAND2_X1 U7020 ( .A1(n7591), .A2(n5318), .ZN(n5395) );
  OR2_X1 U7021 ( .A1(n7751), .A2(n7614), .ZN(n5394) );
  NAND2_X1 U7022 ( .A1(n7733), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U7023 ( .A1(n7731), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5402) );
  INV_X1 U7024 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5397) );
  INV_X1 U7025 ( .A(n5398), .ZN(n5396) );
  NAND2_X1 U7026 ( .A1(n5397), .A2(n5396), .ZN(n5399) );
  NAND2_X1 U7027 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n5398), .ZN(n5418) );
  NAND2_X1 U7028 ( .A1(n5340), .A2(n5964), .ZN(n5401) );
  NAND2_X1 U7029 ( .A1(n7732), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U7030 ( .A1(n9157), .A2(n6441), .ZN(n7636) );
  NAND2_X1 U7031 ( .A1(n7795), .A2(n7636), .ZN(n7761) );
  NAND2_X1 U7032 ( .A1(n5411), .A2(n5413), .ZN(n5409) );
  INV_X1 U7033 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U7034 ( .A1(n9027), .A2(n7898), .ZN(n7757) );
  INV_X1 U7035 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U7036 ( .A1(n5412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U7037 ( .A1(n5495), .A2(n7895), .ZN(n5494) );
  INV_X1 U7038 ( .A(n6452), .ZN(n5425) );
  NAND2_X1 U7039 ( .A1(n7898), .A2(n5495), .ZN(n7823) );
  OR2_X1 U7040 ( .A1(n7823), .A2(n5417), .ZN(n9618) );
  NAND2_X1 U7041 ( .A1(n7731), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U7042 ( .A1(n7733), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5421) );
  INV_X1 U7043 ( .A(n5418), .ZN(n7904) );
  NAND2_X1 U7044 ( .A1(n5340), .A2(n7904), .ZN(n5420) );
  NAND2_X1 U7045 ( .A1(n7732), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5419) );
  NAND4_X1 U7046 ( .A1(n5422), .A2(n5421), .A3(n5420), .A4(n5419), .ZN(n8900)
         );
  INV_X1 U7047 ( .A(n5417), .ZN(n9473) );
  AOI22_X1 U7048 ( .A1(n9651), .A2(n9005), .B1(n8900), .B2(n9652), .ZN(n5423)
         );
  NAND2_X1 U7049 ( .A1(n4322), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5427) );
  XNOR2_X1 U7050 ( .A(n5427), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5452) );
  INV_X1 U7051 ( .A(n5452), .ZN(n7451) );
  NAND2_X1 U7052 ( .A1(n7451), .A2(P1_B_REG_SCAN_IN), .ZN(n5431) );
  NAND2_X1 U7053 ( .A1(n5447), .A2(n5450), .ZN(n5428) );
  MUX2_X1 U7054 ( .A(n5431), .B(P1_B_REG_SCAN_IN), .S(n5455), .Z(n5433) );
  OR2_X1 U7055 ( .A1(n9379), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5434) );
  INV_X1 U7056 ( .A(n5455), .ZN(n7394) );
  INV_X1 U7057 ( .A(n5453), .ZN(n7480) );
  NAND2_X1 U7058 ( .A1(n7394), .A2(n7480), .ZN(n9382) );
  OR2_X1 U7059 ( .A1(n9379), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U7060 ( .A1(n7480), .A2(n7451), .ZN(n9381) );
  NOR4_X1 U7061 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5439) );
  NOR4_X1 U7062 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5438) );
  NOR4_X1 U7063 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5437) );
  NOR4_X1 U7064 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5436) );
  NAND4_X1 U7065 ( .A1(n5439), .A2(n5438), .A3(n5437), .A4(n5436), .ZN(n5445)
         );
  NOR2_X1 U7066 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5443) );
  NOR4_X1 U7067 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5442) );
  NOR4_X1 U7068 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5441) );
  NOR4_X1 U7069 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5440) );
  NAND4_X1 U7070 ( .A1(n5443), .A2(n5442), .A3(n5441), .A4(n5440), .ZN(n5444)
         );
  NOR2_X1 U7071 ( .A1(n5445), .A2(n5444), .ZN(n5446) );
  OR2_X1 U7072 ( .A1(n9379), .A2(n5446), .ZN(n5942) );
  NAND2_X1 U7073 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  NAND2_X1 U7074 ( .A1(n5449), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U7075 ( .A1(n6562), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6492) );
  INV_X1 U7076 ( .A(n7823), .ZN(n6561) );
  AND2_X1 U7077 ( .A1(n6561), .A2(n5943), .ZN(n5954) );
  NOR2_X1 U7078 ( .A1(n7896), .A2(n5954), .ZN(n5456) );
  NAND3_X1 U7079 ( .A1(n6473), .A2(n6470), .A3(n6471), .ZN(n5501) );
  INV_X1 U7080 ( .A(n7898), .ZN(n7235) );
  NAND2_X1 U7081 ( .A1(n5740), .A2(n6908), .ZN(n6904) );
  NAND2_X1 U7082 ( .A1(n6903), .A2(n6904), .ZN(n5458) );
  NAND2_X1 U7083 ( .A1(n6819), .A2(n9683), .ZN(n5457) );
  NAND2_X1 U7084 ( .A1(n5458), .A2(n5457), .ZN(n6821) );
  NAND2_X1 U7085 ( .A1(n6821), .A2(n7763), .ZN(n5460) );
  NAND2_X1 U7086 ( .A1(n7835), .A2(n9689), .ZN(n5459) );
  NAND2_X1 U7087 ( .A1(n5460), .A2(n5459), .ZN(n6811) );
  NAND2_X1 U7088 ( .A1(n6811), .A2(n7764), .ZN(n5463) );
  NAND2_X1 U7089 ( .A1(n6820), .A2(n9695), .ZN(n5462) );
  NAND2_X1 U7090 ( .A1(n5463), .A2(n5462), .ZN(n9662) );
  NAND2_X1 U7091 ( .A1(n5464), .A2(n7839), .ZN(n9663) );
  NAND2_X1 U7092 ( .A1(n9662), .A2(n9663), .ZN(n5466) );
  NAND2_X1 U7093 ( .A1(n6956), .A2(n9701), .ZN(n5465) );
  NAND2_X1 U7094 ( .A1(n5466), .A2(n5465), .ZN(n6958) );
  NAND2_X1 U7095 ( .A1(n5467), .A2(n7840), .ZN(n7769) );
  NAND2_X1 U7096 ( .A1(n6958), .A2(n7769), .ZN(n5470) );
  NAND2_X1 U7097 ( .A1(n5468), .A2(n9708), .ZN(n5469) );
  NAND2_X1 U7098 ( .A1(n5470), .A2(n5469), .ZN(n9642) );
  NAND2_X1 U7099 ( .A1(n7768), .A2(n7640), .ZN(n9643) );
  NAND2_X1 U7100 ( .A1(n6957), .A2(n9714), .ZN(n5471) );
  NAND2_X1 U7101 ( .A1(n7643), .A2(n7009), .ZN(n7645) );
  NAND2_X1 U7102 ( .A1(n7644), .A2(n7646), .ZN(n7010) );
  NAND2_X1 U7103 ( .A1(n9620), .A2(n7010), .ZN(n5473) );
  OR2_X1 U7104 ( .A1(n7181), .A2(n8910), .ZN(n5472) );
  NAND2_X1 U7105 ( .A1(n5473), .A2(n5472), .ZN(n7015) );
  NAND2_X1 U7106 ( .A1(n7648), .A2(n7652), .ZN(n7016) );
  NAND2_X1 U7107 ( .A1(n7015), .A2(n7016), .ZN(n5475) );
  OR2_X1 U7108 ( .A1(n5078), .A2(n8909), .ZN(n5474) );
  NOR2_X1 U7109 ( .A1(n5476), .A2(n8908), .ZN(n5477) );
  NOR2_X1 U7110 ( .A1(n5177), .A2(n8905), .ZN(n5479) );
  NAND2_X1 U7111 ( .A1(n9213), .A2(n9124), .ZN(n5480) );
  INV_X1 U7112 ( .A(n9213), .ZN(n9137) );
  NAND2_X1 U7113 ( .A1(n9120), .A2(n9144), .ZN(n5481) );
  NAND2_X1 U7114 ( .A1(n9116), .A2(n5481), .ZN(n5482) );
  INV_X1 U7115 ( .A(n9208), .ZN(n9120) );
  NAND2_X1 U7116 ( .A1(n5482), .A2(n4867), .ZN(n9099) );
  NAND2_X1 U7117 ( .A1(n9099), .A2(n5483), .ZN(n5484) );
  INV_X1 U7118 ( .A(n9199), .ZN(n9096) );
  INV_X1 U7119 ( .A(n9194), .ZN(n9082) );
  NAND2_X1 U7120 ( .A1(n5486), .A2(n4868), .ZN(n9053) );
  INV_X1 U7121 ( .A(n9188), .ZN(n9058) );
  NOR2_X1 U7122 ( .A1(n9058), .A2(n9074), .ZN(n5488) );
  OAI21_X1 U7123 ( .B1(n9053), .B2(n5488), .A(n5487), .ZN(n9040) );
  AOI21_X1 U7124 ( .B1(n8827), .B2(n4531), .A(n9040), .ZN(n5489) );
  AOI21_X1 U7125 ( .B1(n9065), .B2(n9183), .A(n5489), .ZN(n9024) );
  NAND2_X1 U7126 ( .A1(n9178), .A2(n9048), .ZN(n5490) );
  INV_X1 U7127 ( .A(n9173), .ZN(n9015) );
  NAND2_X1 U7128 ( .A1(n9015), .A2(n5491), .ZN(n5492) );
  INV_X1 U7129 ( .A(n9168), .ZN(n9001) );
  INV_X1 U7130 ( .A(n9164), .ZN(n8994) );
  XNOR2_X1 U7131 ( .A(n6444), .B(n7761), .ZN(n9161) );
  OR2_X1 U7132 ( .A1(n7898), .A2(n5494), .ZN(n7890) );
  NAND3_X1 U7133 ( .A1(n7890), .A2(n6802), .A3(n7928), .ZN(n5497) );
  NAND2_X1 U7134 ( .A1(n7898), .A2(n7928), .ZN(n5728) );
  INV_X1 U7135 ( .A(n5728), .ZN(n5496) );
  AND2_X1 U7136 ( .A1(n5496), .A2(n5498), .ZN(n6801) );
  INV_X1 U7137 ( .A(n5498), .ZN(n5727) );
  AND2_X1 U7138 ( .A1(n9622), .A2(n6905), .ZN(n5499) );
  INV_X1 U7139 ( .A(n7045), .ZN(n9723) );
  NAND2_X1 U7140 ( .A1(n9644), .A2(n9723), .ZN(n9630) );
  INV_X1 U7141 ( .A(n5476), .ZN(n9743) );
  INV_X1 U7142 ( .A(n7086), .ZN(n9749) );
  INV_X1 U7143 ( .A(n8895), .ZN(n7350) );
  INV_X1 U7144 ( .A(n9219), .ZN(n8814) );
  NAND2_X1 U7145 ( .A1(n9103), .A2(n9117), .ZN(n9100) );
  AOI21_X1 U7146 ( .B1(n9157), .B2(n8988), .A(n8967), .ZN(n9158) );
  NOR2_X1 U7147 ( .A1(n8982), .A2(n9769), .ZN(n7907) );
  INV_X1 U7148 ( .A(n9157), .ZN(n6442) );
  OR2_X1 U7149 ( .A1(n6802), .A2(n7146), .ZN(n5958) );
  OR2_X2 U7150 ( .A1(n9658), .A2(n5958), .ZN(n9660) );
  INV_X2 U7151 ( .A(n9104), .ZN(n9656) );
  AOI22_X1 U7152 ( .A1(n9673), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n5964), .B2(
        n9656), .ZN(n5502) );
  OAI21_X1 U7153 ( .B1(n6442), .B2(n9660), .A(n5502), .ZN(n5503) );
  AOI21_X1 U7154 ( .B1(n9158), .B2(n7907), .A(n5503), .ZN(n5504) );
  NOR3_X1 U7155 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n5513) );
  NOR2_X1 U7156 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5512) );
  NOR2_X1 U7157 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5511) );
  NAND2_X1 U7158 ( .A1(n5556), .A2(n5510), .ZN(n5551) );
  INV_X1 U7159 ( .A(n5551), .ZN(n5533) );
  NAND2_X1 U7160 ( .A1(n5531), .A2(n4274), .ZN(n5537) );
  INV_X1 U7161 ( .A(n5537), .ZN(n5515) );
  INV_X1 U7162 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5517) );
  INV_X1 U7163 ( .A(n5519), .ZN(n5518) );
  NAND2_X1 U7164 ( .A1(n5518), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7165 ( .A1(n5519), .A2(n9238), .ZN(n5520) );
  NAND2_X1 U7166 ( .A1(n5524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5522) );
  INV_X1 U7167 ( .A(n7448), .ZN(n5527) );
  NAND2_X1 U7168 ( .A1(n4321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5523) );
  MUX2_X1 U7169 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5523), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n5525) );
  NAND2_X1 U7170 ( .A1(n5525), .A2(n5524), .ZN(n7383) );
  INV_X1 U7171 ( .A(n7383), .ZN(n5526) );
  NAND2_X1 U7172 ( .A1(n5539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5529) );
  INV_X1 U7173 ( .A(n6595), .ZN(n5530) );
  NOR2_X1 U7174 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5532) );
  NAND2_X1 U7175 ( .A1(n6306), .A2(n6305), .ZN(n5535) );
  NAND2_X1 U7176 ( .A1(n5535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7177 ( .A1(n5537), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5538) );
  MUX2_X1 U7178 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5538), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5540) );
  NAND2_X1 U7179 ( .A1(n5540), .A2(n5539), .ZN(n8359) );
  NAND2_X1 U7180 ( .A1(n6747), .A2(n8278), .ZN(n5541) );
  NAND2_X1 U7181 ( .A1(n5541), .A2(n6746), .ZN(n5639) );
  NAND2_X1 U7182 ( .A1(n9238), .A2(n5545), .ZN(n5548) );
  NAND2_X1 U7183 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n5543) );
  NAND2_X1 U7184 ( .A1(n5543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5544) );
  OAI21_X1 U7185 ( .B1(n5545), .B2(P2_IR_REG_31__SCAN_IN), .A(n5544), .ZN(
        n5546) );
  OAI211_X2 U7186 ( .C1(n5549), .C2(n5548), .A(n5547), .B(n5546), .ZN(n5641)
         );
  NAND2_X1 U7187 ( .A1(n5639), .A2(n5989), .ZN(n5550) );
  NAND2_X1 U7188 ( .A1(n5550), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U7189 ( .A1(n5562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7190 ( .A1(n5551), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7191 ( .A1(n5557), .A2(n5552), .ZN(n5624) );
  OAI21_X1 U7192 ( .B1(n5624), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5553) );
  XNOR2_X1 U7193 ( .A(n5553), .B(P2_IR_REG_17__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7194 ( .A1(n5557), .A2(n5556), .ZN(n5554) );
  NAND2_X1 U7195 ( .A1(n5554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5555) );
  XNOR2_X1 U7196 ( .A(n5555), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U7197 ( .A(n5557), .B(n5556), .ZN(n6653) );
  INV_X1 U7198 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U7199 ( .A1(n5559), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5561) );
  MUX2_X1 U7200 ( .A(n5561), .B(P2_IR_REG_31__SCAN_IN), .S(n5560), .Z(n5563)
         );
  NAND2_X1 U7201 ( .A1(n5563), .A2(n5562), .ZN(n6649) );
  OR2_X1 U7202 ( .A1(n5564), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7203 ( .A1(n5569), .A2(n5565), .ZN(n5572) );
  OAI21_X1 U7204 ( .B1(n5572), .B2(P2_IR_REG_11__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U7205 ( .A(n5567), .B(n5566), .ZN(n6600) );
  NAND2_X1 U7206 ( .A1(n5572), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5568) );
  XNOR2_X1 U7207 ( .A(n5568), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7509) );
  NOR2_X1 U7208 ( .A1(n5569), .A2(n5974), .ZN(n5570) );
  MUX2_X1 U7209 ( .A(n5974), .B(n5570), .S(P2_IR_REG_10__SCAN_IN), .Z(n5571)
         );
  INV_X1 U7210 ( .A(n5571), .ZN(n5573) );
  NAND2_X1 U7211 ( .A1(n5573), .A2(n5572), .ZN(n6581) );
  NAND2_X1 U7212 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5574) );
  MUX2_X1 U7213 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5574), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5576) );
  INV_X1 U7214 ( .A(n5644), .ZN(n5575) );
  INV_X1 U7215 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9239) );
  AND2_X1 U7216 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n9239), .ZN(n5577) );
  NAND2_X1 U7217 ( .A1(n5644), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5578) );
  INV_X1 U7218 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9809) );
  INV_X1 U7219 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7031) );
  XNOR2_X1 U7220 ( .A(n4269), .B(n7031), .ZN(n6696) );
  NAND2_X1 U7221 ( .A1(n6695), .A2(n6696), .ZN(n6694) );
  NAND2_X1 U7222 ( .A1(n4269), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7223 ( .A1(n6694), .A2(n5581), .ZN(n5584) );
  NAND2_X1 U7224 ( .A1(n5582), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5583) );
  INV_X1 U7225 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9869) );
  INV_X1 U7226 ( .A(n5586), .ZN(n5590) );
  NAND2_X1 U7227 ( .A1(n5587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5588) );
  MUX2_X1 U7228 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5588), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5589) );
  NAND2_X1 U7229 ( .A1(n5590), .A2(n5589), .ZN(n9838) );
  INV_X1 U7230 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7129) );
  XNOR2_X1 U7231 ( .A(n9838), .B(n7129), .ZN(n9832) );
  NAND2_X1 U7232 ( .A1(n9838), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7233 ( .A1(n9837), .A2(n5591), .ZN(n5594) );
  OR2_X1 U7234 ( .A1(n5586), .A2(n5974), .ZN(n5593) );
  XNOR2_X1 U7235 ( .A(n5593), .B(n5592), .ZN(n6538) );
  INV_X1 U7236 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6708) );
  NOR2_X1 U7237 ( .A1(n5595), .A2(n5974), .ZN(n5596) );
  MUX2_X1 U7238 ( .A(n5974), .B(n5596), .S(P2_IR_REG_6__SCAN_IN), .Z(n5598) );
  INV_X1 U7239 ( .A(n5564), .ZN(n5597) );
  INV_X1 U7240 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6065) );
  XNOR2_X1 U7241 ( .A(n6543), .B(n6065), .ZN(n6788) );
  NAND2_X1 U7242 ( .A1(n5599), .A2(n6788), .ZN(n6786) );
  NAND2_X1 U7243 ( .A1(n6543), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7244 ( .A1(n5564), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5602) );
  XNOR2_X1 U7245 ( .A(n5602), .B(n5601), .ZN(n6552) );
  NAND2_X1 U7246 ( .A1(n6504), .A2(n5604), .ZN(n6522) );
  INV_X1 U7247 ( .A(n6522), .ZN(n5605) );
  INV_X1 U7248 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U7249 ( .A1(n6524), .A2(n6504), .ZN(n5609) );
  INV_X1 U7250 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7251 ( .A1(n5606), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5607) );
  XNOR2_X1 U7252 ( .A(n5607), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6093) );
  MUX2_X1 U7253 ( .A(n5608), .B(P2_REG2_REG_8__SCAN_IN), .S(n6093), .Z(n6503)
         );
  NAND2_X1 U7254 ( .A1(n5609), .A2(n6503), .ZN(n6507) );
  OR2_X1 U7255 ( .A1(n6093), .A2(n5608), .ZN(n5610) );
  NAND2_X1 U7256 ( .A1(n5611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5612) );
  XNOR2_X1 U7257 ( .A(n5612), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6094) );
  XNOR2_X1 U7258 ( .A(n5613), .B(n6094), .ZN(n7114) );
  NAND2_X1 U7259 ( .A1(n7114), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7116) );
  INV_X1 U7260 ( .A(n6094), .ZN(n7113) );
  NAND2_X1 U7261 ( .A1(n5613), .A2(n7113), .ZN(n5614) );
  NAND2_X1 U7262 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6581), .ZN(n5615) );
  OAI21_X1 U7263 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6581), .A(n5615), .ZN(
        n7220) );
  NOR2_X1 U7264 ( .A1(n7221), .A2(n7220), .ZN(n7219) );
  AOI21_X1 U7265 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6581), .A(n7219), .ZN(
        n5616) );
  NOR2_X1 U7266 ( .A1(n7509), .A2(n5616), .ZN(n5617) );
  INV_X1 U7267 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U7268 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6600), .ZN(n5618) );
  OAI21_X1 U7269 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6600), .A(n5618), .ZN(
        n7594) );
  INV_X1 U7270 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7560) );
  INV_X1 U7271 ( .A(n6649), .ZN(n7561) );
  NOR2_X1 U7272 ( .A1(n7561), .A2(n5619), .ZN(n5620) );
  NAND2_X1 U7273 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6653), .ZN(n5621) );
  OAI21_X1 U7274 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6653), .A(n5621), .ZN(
        n8396) );
  NOR2_X1 U7275 ( .A1(n8417), .A2(n5622), .ZN(n5623) );
  INV_X1 U7276 ( .A(n8417), .ZN(n6677) );
  INV_X1 U7277 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8416) );
  XNOR2_X1 U7278 ( .A(n5624), .B(P2_IR_REG_16__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U7279 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n6772), .ZN(n5625) );
  OAI21_X1 U7280 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n6772), .A(n5625), .ZN(
        n8434) );
  NOR2_X1 U7281 ( .A1(n5990), .A2(n5627), .ZN(n5628) );
  INV_X1 U7282 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8453) );
  XNOR2_X1 U7283 ( .A(n5627), .B(n5990), .ZN(n8452) );
  NOR2_X1 U7284 ( .A1(n8453), .A2(n8452), .ZN(n8451) );
  NAND2_X1 U7285 ( .A1(n5629), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5630) );
  XNOR2_X1 U7286 ( .A(n5630), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8484) );
  INV_X1 U7287 ( .A(n8484), .ZN(n8475) );
  NAND2_X1 U7288 ( .A1(n8475), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5631) );
  OAI21_X1 U7289 ( .B1(n8475), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5631), .ZN(
        n8480) );
  NOR2_X1 U7290 ( .A1(n8481), .A2(n8480), .ZN(n8479) );
  INV_X1 U7291 ( .A(n5631), .ZN(n5632) );
  NOR2_X1 U7292 ( .A1(n8479), .A2(n5632), .ZN(n5638) );
  INV_X1 U7293 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7294 ( .A1(n5633), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5635) );
  INV_X1 U7295 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5634) );
  MUX2_X1 U7296 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n5636), .S(n7067), .Z(n5715)
         );
  INV_X1 U7297 ( .A(n5715), .ZN(n5637) );
  XNOR2_X1 U7298 ( .A(n5638), .B(n5637), .ZN(n5643) );
  NAND2_X1 U7299 ( .A1(n5639), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5721) );
  NOR2_X1 U7300 ( .A1(n5721), .A2(n8370), .ZN(n9806) );
  INV_X2 U7301 ( .A(n5641), .ZN(n8371) );
  NAND2_X1 U7302 ( .A1(n9806), .A2(n8371), .ZN(n9822) );
  AND2_X1 U7303 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n9239), .ZN(n5645) );
  NAND2_X1 U7304 ( .A1(n5644), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5646) );
  OAI21_X1 U7305 ( .B1(n9818), .B2(n5645), .A(n5646), .ZN(n9814) );
  INV_X1 U7306 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9813) );
  XNOR2_X1 U7307 ( .A(n6532), .B(n9937), .ZN(n6693) );
  NAND2_X1 U7308 ( .A1(n6692), .A2(n6693), .ZN(n6691) );
  NAND2_X1 U7309 ( .A1(n4269), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7310 ( .A1(n6691), .A2(n5647), .ZN(n5648) );
  INV_X1 U7311 ( .A(n6546), .ZN(n6666) );
  XNOR2_X1 U7312 ( .A(n5648), .B(n6666), .ZN(n6661) );
  NAND2_X1 U7313 ( .A1(n6661), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7314 ( .A1(n5648), .A2(n6546), .ZN(n5649) );
  NAND2_X1 U7315 ( .A1(n5650), .A2(n5649), .ZN(n9849) );
  INV_X1 U7316 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6034) );
  XNOR2_X1 U7317 ( .A(n9838), .B(n6034), .ZN(n9850) );
  NAND2_X1 U7318 ( .A1(n9849), .A2(n9850), .ZN(n9848) );
  NAND2_X1 U7319 ( .A1(n9838), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5651) );
  INV_X1 U7320 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9941) );
  INV_X1 U7321 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5653) );
  XNOR2_X1 U7322 ( .A(n6543), .B(n5653), .ZN(n6780) );
  NAND2_X1 U7323 ( .A1(n5654), .A2(n6780), .ZN(n6785) );
  NAND2_X1 U7324 ( .A1(n6543), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7325 ( .A1(n6785), .A2(n5655), .ZN(n5656) );
  INV_X1 U7326 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9273) );
  MUX2_X1 U7327 ( .A(n9273), .B(P2_REG1_REG_8__SCAN_IN), .S(n6093), .Z(n6498)
         );
  NAND2_X1 U7328 ( .A1(n5657), .A2(n6498), .ZN(n6502) );
  OR2_X1 U7329 ( .A1(n6093), .A2(n9273), .ZN(n5658) );
  NAND2_X1 U7330 ( .A1(n6502), .A2(n5658), .ZN(n5659) );
  XNOR2_X1 U7331 ( .A(n5659), .B(n6094), .ZN(n7110) );
  NAND2_X1 U7332 ( .A1(n7110), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U7333 ( .A1(n5659), .A2(n7113), .ZN(n5660) );
  NAND2_X1 U7334 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6581), .ZN(n5661) );
  OAI21_X1 U7335 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6581), .A(n5661), .ZN(
        n7217) );
  AOI21_X1 U7336 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6581), .A(n7216), .ZN(
        n5662) );
  NOR2_X1 U7337 ( .A1(n7509), .A2(n5662), .ZN(n5663) );
  INV_X1 U7338 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9948) );
  XNOR2_X1 U7339 ( .A(n5662), .B(n7509), .ZN(n7496) );
  NOR2_X1 U7340 ( .A1(n9948), .A2(n7496), .ZN(n7495) );
  NAND2_X1 U7341 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6600), .ZN(n5664) );
  OAI21_X1 U7342 ( .B1(n6600), .B2(P2_REG1_REG_12__SCAN_IN), .A(n5664), .ZN(
        n7606) );
  NOR2_X1 U7343 ( .A1(n7561), .A2(n5665), .ZN(n5667) );
  INV_X1 U7344 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9459) );
  NOR2_X1 U7345 ( .A1(n9459), .A2(n7567), .ZN(n7566) );
  NOR2_X1 U7346 ( .A1(n5667), .A2(n7566), .ZN(n8407) );
  NAND2_X1 U7347 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6653), .ZN(n5668) );
  OAI21_X1 U7348 ( .B1(n6653), .B2(P2_REG1_REG_14__SCAN_IN), .A(n5668), .ZN(
        n8406) );
  NOR2_X1 U7349 ( .A1(n8407), .A2(n8406), .ZN(n8405) );
  NOR2_X1 U7350 ( .A1(n8417), .A2(n5669), .ZN(n5670) );
  INV_X1 U7351 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8424) );
  XNOR2_X1 U7352 ( .A(n6772), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8443) );
  NOR2_X1 U7353 ( .A1(n5990), .A2(n5671), .ZN(n5672) );
  INV_X1 U7354 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U7355 ( .A1(n8475), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5673) );
  OAI21_X1 U7356 ( .B1(n8475), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5673), .ZN(
        n8470) );
  INV_X1 U7357 ( .A(n5673), .ZN(n5674) );
  INV_X1 U7358 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n6210) );
  XNOR2_X1 U7359 ( .A(n7067), .B(n6210), .ZN(n5716) );
  XNOR2_X1 U7360 ( .A(n5675), .B(n5716), .ZN(n5725) );
  INV_X4 U7361 ( .A(n8371), .ZN(n7542) );
  NAND2_X1 U7362 ( .A1(n9806), .A2(n7542), .ZN(n8485) );
  MUX2_X1 U7363 ( .A(n8453), .B(n8458), .S(n7542), .Z(n5676) );
  NAND2_X1 U7364 ( .A1(n5676), .A2(n5990), .ZN(n5709) );
  INV_X1 U7365 ( .A(n5990), .ZN(n8463) );
  XNOR2_X1 U7366 ( .A(n5676), .B(n8463), .ZN(n8456) );
  MUX2_X1 U7367 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n7542), .Z(n5677) );
  OR2_X1 U7368 ( .A1(n6772), .A2(n5677), .ZN(n5708) );
  INV_X1 U7369 ( .A(n6772), .ZN(n8448) );
  XNOR2_X1 U7370 ( .A(n5677), .B(n8448), .ZN(n8437) );
  MUX2_X1 U7371 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n7542), .Z(n5707) );
  XNOR2_X1 U7372 ( .A(n5707), .B(n8417), .ZN(n8421) );
  MUX2_X1 U7373 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n7542), .Z(n5678) );
  OR2_X1 U7374 ( .A1(n5678), .A2(n6653), .ZN(n5706) );
  INV_X1 U7375 ( .A(n6653), .ZN(n8411) );
  XNOR2_X1 U7376 ( .A(n5678), .B(n8411), .ZN(n8399) );
  MUX2_X1 U7377 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n7542), .Z(n5704) );
  OR2_X1 U7378 ( .A1(n5704), .A2(n6649), .ZN(n5705) );
  MUX2_X1 U7379 ( .A(n7505), .B(n9948), .S(n7542), .Z(n5702) );
  INV_X1 U7380 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5679) );
  INV_X1 U7381 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9946) );
  MUX2_X1 U7382 ( .A(n5679), .B(n9946), .S(n7542), .Z(n5700) );
  INV_X1 U7383 ( .A(n6581), .ZN(n7225) );
  AND2_X1 U7384 ( .A1(n5700), .A2(n7225), .ZN(n5701) );
  INV_X1 U7385 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6102) );
  INV_X1 U7386 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6098) );
  MUX2_X1 U7387 ( .A(n6102), .B(n6098), .S(n7542), .Z(n5698) );
  MUX2_X1 U7388 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n7542), .Z(n5685) );
  MUX2_X1 U7389 ( .A(n9809), .B(n9813), .S(n5641), .Z(n5680) );
  XNOR2_X1 U7390 ( .A(n5680), .B(n9818), .ZN(n9825) );
  INV_X1 U7391 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6003) );
  MUX2_X1 U7392 ( .A(n6003), .B(n9935), .S(n7542), .Z(n9804) );
  NAND2_X1 U7393 ( .A1(n9804), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9826) );
  INV_X1 U7394 ( .A(n5680), .ZN(n5681) );
  AOI22_X1 U7395 ( .A1(n9825), .A2(n9826), .B1(n9818), .B2(n5681), .ZN(n6690)
         );
  MUX2_X1 U7396 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n7542), .Z(n5682) );
  XNOR2_X1 U7397 ( .A(n5682), .B(n4269), .ZN(n6689) );
  INV_X1 U7398 ( .A(n4269), .ZN(n6702) );
  INV_X1 U7399 ( .A(n5682), .ZN(n5683) );
  MUX2_X1 U7400 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n7542), .Z(n5684) );
  XNOR2_X1 U7401 ( .A(n5684), .B(n6546), .ZN(n6657) );
  XNOR2_X1 U7402 ( .A(n5685), .B(n9838), .ZN(n9846) );
  NOR2_X1 U7403 ( .A1(n9845), .A2(n9846), .ZN(n9843) );
  AOI21_X1 U7404 ( .B1(n5685), .B2(n9838), .A(n9843), .ZN(n6706) );
  MUX2_X1 U7405 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n7542), .Z(n5686) );
  XNOR2_X1 U7406 ( .A(n5686), .B(n6538), .ZN(n6705) );
  INV_X1 U7407 ( .A(n5686), .ZN(n5687) );
  MUX2_X1 U7408 ( .A(n6065), .B(n5653), .S(n7542), .Z(n5688) );
  INV_X1 U7409 ( .A(n6543), .ZN(n6796) );
  NAND2_X1 U7410 ( .A1(n5688), .A2(n6796), .ZN(n5689) );
  OAI21_X1 U7411 ( .B1(n5688), .B2(n6796), .A(n5689), .ZN(n6778) );
  NOR2_X1 U7412 ( .A1(n6779), .A2(n6778), .ZN(n6777) );
  INV_X1 U7413 ( .A(n5689), .ZN(n6515) );
  INV_X1 U7414 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6074) );
  MUX2_X1 U7415 ( .A(n6521), .B(n6074), .S(n7542), .Z(n5690) );
  NAND2_X1 U7416 ( .A1(n5690), .A2(n4747), .ZN(n6495) );
  INV_X1 U7417 ( .A(n5690), .ZN(n5691) );
  NAND2_X1 U7418 ( .A1(n5691), .A2(n6552), .ZN(n5692) );
  AND2_X1 U7419 ( .A1(n6495), .A2(n5692), .ZN(n6514) );
  MUX2_X1 U7420 ( .A(n5608), .B(n9273), .S(n7542), .Z(n5693) );
  NAND2_X1 U7421 ( .A1(n5693), .A2(n6093), .ZN(n5696) );
  INV_X1 U7422 ( .A(n5693), .ZN(n5694) );
  INV_X1 U7423 ( .A(n6093), .ZN(n6557) );
  NAND2_X1 U7424 ( .A1(n5694), .A2(n6557), .ZN(n5695) );
  NAND2_X1 U7425 ( .A1(n5696), .A2(n5695), .ZN(n6494) );
  INV_X1 U7426 ( .A(n5696), .ZN(n5697) );
  NOR2_X1 U7427 ( .A1(n6493), .A2(n5697), .ZN(n7108) );
  XNOR2_X1 U7428 ( .A(n5698), .B(n6094), .ZN(n7107) );
  NOR2_X1 U7429 ( .A1(n7108), .A2(n7107), .ZN(n7106) );
  INV_X1 U7430 ( .A(n5701), .ZN(n5699) );
  OAI21_X1 U7431 ( .B1(n7225), .B2(n5700), .A(n5699), .ZN(n7214) );
  NOR2_X1 U7432 ( .A1(n7215), .A2(n7214), .ZN(n7213) );
  NOR2_X1 U7433 ( .A1(n5701), .A2(n7213), .ZN(n7498) );
  XNOR2_X1 U7434 ( .A(n5702), .B(n7509), .ZN(n7499) );
  NOR2_X1 U7435 ( .A1(n7498), .A2(n7499), .ZN(n7497) );
  INV_X1 U7436 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7327) );
  INV_X1 U7437 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6143) );
  MUX2_X1 U7438 ( .A(n7327), .B(n6143), .S(n7542), .Z(n5703) );
  INV_X1 U7439 ( .A(n6600), .ZN(n7611) );
  NAND2_X1 U7440 ( .A1(n5703), .A2(n7611), .ZN(n7595) );
  NOR2_X1 U7441 ( .A1(n7611), .A2(n5703), .ZN(n7596) );
  XNOR2_X1 U7442 ( .A(n5704), .B(n7561), .ZN(n7564) );
  NAND2_X1 U7443 ( .A1(n7563), .A2(n7564), .ZN(n7562) );
  NAND2_X1 U7444 ( .A1(n5705), .A2(n7562), .ZN(n8398) );
  NAND2_X1 U7445 ( .A1(n8399), .A2(n8398), .ZN(n8397) );
  NAND2_X1 U7446 ( .A1(n5706), .A2(n8397), .ZN(n8420) );
  NAND2_X1 U7447 ( .A1(n8421), .A2(n8420), .ZN(n8419) );
  OAI21_X1 U7448 ( .B1(n5707), .B2(n6677), .A(n8419), .ZN(n8436) );
  NAND2_X1 U7449 ( .A1(n8437), .A2(n8436), .ZN(n8435) );
  NAND2_X1 U7450 ( .A1(n5708), .A2(n8435), .ZN(n8455) );
  NAND2_X1 U7451 ( .A1(n8456), .A2(n8455), .ZN(n8454) );
  NAND2_X1 U7452 ( .A1(n5709), .A2(n8454), .ZN(n5710) );
  INV_X1 U7453 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8611) );
  INV_X1 U7454 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8669) );
  MUX2_X1 U7455 ( .A(n8611), .B(n8669), .S(n7542), .Z(n5711) );
  NAND2_X1 U7456 ( .A1(n5710), .A2(n5711), .ZN(n8471) );
  NAND2_X1 U7457 ( .A1(n8471), .A2(n8475), .ZN(n5714) );
  INV_X1 U7458 ( .A(n5710), .ZN(n5713) );
  INV_X1 U7459 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7460 ( .A1(n5713), .A2(n5712), .ZN(n8472) );
  NAND2_X1 U7461 ( .A1(n5714), .A2(n8472), .ZN(n5718) );
  MUX2_X1 U7462 ( .A(n5716), .B(n5715), .S(n8371), .Z(n5717) );
  NAND2_X1 U7463 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8015) );
  INV_X1 U7464 ( .A(n6746), .ZN(n7298) );
  NOR2_X1 U7465 ( .A1(n6747), .A2(n7298), .ZN(n5719) );
  NAND2_X1 U7466 ( .A1(n9841), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5720) );
  MUX2_X1 U7467 ( .A(n8474), .B(n5721), .S(n8370), .Z(n5722) );
  NOR2_X2 U7468 ( .A1(n5722), .A2(n6204), .ZN(n9839) );
  OAI21_X1 U7469 ( .B1(n5725), .B2(n8485), .A(n5724), .ZN(n5726) );
  AND2_X1 U7470 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  NAND2_X1 U7471 ( .A1(n5732), .A2(n5908), .ZN(n5731) );
  NAND2_X1 U7472 ( .A1(n5732), .A2(n5885), .ZN(n5734) );
  NAND2_X1 U7473 ( .A1(n5939), .A2(n6907), .ZN(n5733) );
  NAND2_X1 U7474 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  NOR2_X1 U7475 ( .A1(n5737), .A2(n5745), .ZN(n6726) );
  NAND2_X1 U7476 ( .A1(n5746), .A2(n6908), .ZN(n5739) );
  NAND2_X1 U7477 ( .A1(n5912), .A2(n5740), .ZN(n5738) );
  AND2_X1 U7478 ( .A1(n5739), .A2(n5738), .ZN(n5744) );
  INV_X1 U7479 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U7480 ( .A1(n5744), .A2(n4861), .ZN(n6670) );
  NAND2_X1 U7481 ( .A1(n5740), .A2(n5885), .ZN(n5742) );
  NAND2_X1 U7482 ( .A1(n5742), .A2(n5741), .ZN(n6669) );
  AOI22_X1 U7483 ( .A1(n6670), .A2(n6669), .B1(n5744), .B2(n4377), .ZN(n6727)
         );
  NAND2_X1 U7484 ( .A1(n6726), .A2(n6727), .ZN(n6725) );
  INV_X1 U7485 ( .A(n5745), .ZN(n6718) );
  NAND2_X1 U7486 ( .A1(n6911), .A2(n5908), .ZN(n5748) );
  NAND2_X1 U7487 ( .A1(n5746), .A2(n7834), .ZN(n5747) );
  NAND2_X1 U7488 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  AND2_X1 U7489 ( .A1(n5939), .A2(n7834), .ZN(n5750) );
  AOI21_X1 U7490 ( .B1(n6911), .B2(n5885), .A(n5750), .ZN(n5751) );
  NAND2_X1 U7491 ( .A1(n5752), .A2(n4879), .ZN(n6717) );
  INV_X1 U7492 ( .A(n5752), .ZN(n5753) );
  NOR2_X1 U7493 ( .A1(n6720), .A2(n5753), .ZN(n6680) );
  AOI22_X1 U7494 ( .A1(n5754), .A2(n5885), .B1(n5939), .B2(n5755), .ZN(n5760)
         );
  NAND2_X1 U7495 ( .A1(n5754), .A2(n5912), .ZN(n5757) );
  NAND2_X1 U7496 ( .A1(n5746), .A2(n5755), .ZN(n5756) );
  NAND2_X1 U7497 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  XNOR2_X1 U7498 ( .A(n5758), .B(n5937), .ZN(n5759) );
  XOR2_X1 U7499 ( .A(n5760), .B(n5759), .Z(n6679) );
  NOR2_X1 U7500 ( .A1(n6680), .A2(n6679), .ZN(n6678) );
  INV_X1 U7501 ( .A(n5759), .ZN(n5761) );
  AOI22_X1 U7502 ( .A1(n8912), .A2(n5885), .B1(n5939), .B2(n5762), .ZN(n5764)
         );
  AOI22_X1 U7503 ( .A1(n8912), .A2(n5939), .B1(n5762), .B2(n5746), .ZN(n5763)
         );
  XNOR2_X1 U7504 ( .A(n5763), .B(n5937), .ZN(n5765) );
  XOR2_X1 U7505 ( .A(n5764), .B(n5765), .Z(n8834) );
  OR2_X1 U7506 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  NAND2_X1 U7507 ( .A1(n9653), .A2(n5908), .ZN(n5768) );
  NAND2_X1 U7508 ( .A1(n5746), .A2(n6961), .ZN(n5767) );
  NAND2_X1 U7509 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  XNOR2_X1 U7510 ( .A(n5769), .B(n5937), .ZN(n6736) );
  INV_X1 U7511 ( .A(n6736), .ZN(n5773) );
  NAND2_X1 U7512 ( .A1(n9653), .A2(n5885), .ZN(n5771) );
  NAND2_X1 U7513 ( .A1(n6961), .A2(n5908), .ZN(n5770) );
  NAND2_X1 U7514 ( .A1(n5771), .A2(n5770), .ZN(n5775) );
  INV_X1 U7515 ( .A(n5775), .ZN(n5772) );
  NAND2_X1 U7516 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  NAND2_X1 U7517 ( .A1(n6736), .A2(n5775), .ZN(n5776) );
  NAND2_X1 U7518 ( .A1(n5777), .A2(n5776), .ZN(n6947) );
  NAND2_X1 U7519 ( .A1(n8911), .A2(n5908), .ZN(n5779) );
  NAND2_X1 U7520 ( .A1(n5781), .A2(n5746), .ZN(n5778) );
  NAND2_X1 U7521 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  XNOR2_X1 U7522 ( .A(n5780), .B(n4377), .ZN(n5783) );
  AOI22_X1 U7523 ( .A1(n8911), .A2(n5885), .B1(n5781), .B2(n5912), .ZN(n5782)
         );
  NAND2_X1 U7524 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  OAI21_X1 U7525 ( .B1(n5783), .B2(n5782), .A(n5784), .ZN(n6948) );
  INV_X1 U7526 ( .A(n5784), .ZN(n5785) );
  NAND2_X1 U7527 ( .A1(n7045), .A2(n5746), .ZN(n5787) );
  NAND2_X1 U7528 ( .A1(n9637), .A2(n5908), .ZN(n5786) );
  NAND2_X1 U7529 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  XNOR2_X1 U7530 ( .A(n5788), .B(n4377), .ZN(n5790) );
  AOI22_X1 U7531 ( .A1(n7045), .A2(n5912), .B1(n5885), .B2(n9637), .ZN(n5789)
         );
  NAND2_X1 U7532 ( .A1(n5790), .A2(n5789), .ZN(n7069) );
  NAND2_X1 U7533 ( .A1(n7181), .A2(n5746), .ZN(n5793) );
  NAND2_X1 U7534 ( .A1(n8910), .A2(n5939), .ZN(n5792) );
  NAND2_X1 U7535 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  XNOR2_X1 U7536 ( .A(n5794), .B(n5937), .ZN(n5796) );
  AOI22_X1 U7537 ( .A1(n7181), .A2(n5912), .B1(n5885), .B2(n8910), .ZN(n7183)
         );
  NAND2_X1 U7538 ( .A1(n5078), .A2(n5746), .ZN(n5799) );
  NAND2_X1 U7539 ( .A1(n8909), .A2(n5912), .ZN(n5798) );
  NAND2_X1 U7540 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  XNOR2_X1 U7541 ( .A(n5800), .B(n5937), .ZN(n5801) );
  AOI22_X1 U7542 ( .A1(n5078), .A2(n5939), .B1(n5885), .B2(n8909), .ZN(n5802)
         );
  XNOR2_X1 U7543 ( .A(n5801), .B(n5802), .ZN(n7262) );
  INV_X1 U7544 ( .A(n5801), .ZN(n5803) );
  AOI22_X1 U7545 ( .A1(n7086), .A2(n5746), .B1(n5939), .B2(n8907), .ZN(n5804)
         );
  XNOR2_X1 U7546 ( .A(n5804), .B(n5937), .ZN(n7483) );
  AND2_X1 U7547 ( .A1(n8907), .A2(n5885), .ZN(n5805) );
  AOI21_X1 U7548 ( .B1(n7086), .B2(n5939), .A(n5805), .ZN(n7484) );
  NAND2_X1 U7549 ( .A1(n5476), .A2(n5746), .ZN(n5807) );
  NAND2_X1 U7550 ( .A1(n8908), .A2(n5912), .ZN(n5806) );
  NAND2_X1 U7551 ( .A1(n5807), .A2(n5806), .ZN(n5808) );
  XNOR2_X1 U7552 ( .A(n5808), .B(n5937), .ZN(n7482) );
  INV_X1 U7553 ( .A(n7482), .ZN(n7423) );
  NAND2_X1 U7554 ( .A1(n5476), .A2(n5912), .ZN(n5810) );
  NAND2_X1 U7555 ( .A1(n8908), .A2(n5885), .ZN(n5809) );
  NAND2_X1 U7556 ( .A1(n5810), .A2(n5809), .ZN(n5811) );
  INV_X1 U7557 ( .A(n5811), .ZN(n7425) );
  AOI22_X1 U7558 ( .A1(n7483), .A2(n7484), .B1(n7423), .B2(n7425), .ZN(n5815)
         );
  NAND2_X1 U7559 ( .A1(n7482), .A2(n5811), .ZN(n5812) );
  AOI21_X1 U7560 ( .B1(n7484), .B2(n5812), .A(n7483), .ZN(n5814) );
  NOR3_X1 U7561 ( .A1(n7484), .A2(n7423), .A3(n7425), .ZN(n5813) );
  AOI22_X1 U7562 ( .A1(n7100), .A2(n5746), .B1(n5939), .B2(n7474), .ZN(n5816)
         );
  XOR2_X1 U7563 ( .A(n5937), .B(n5816), .Z(n5819) );
  OAI22_X1 U7564 ( .A1(n9757), .A2(n5791), .B1(n7489), .B2(n5817), .ZN(n5818)
         );
  NOR2_X1 U7565 ( .A1(n5819), .A2(n5818), .ZN(n5820) );
  AOI21_X1 U7566 ( .B1(n5819), .B2(n5818), .A(n5820), .ZN(n7396) );
  NAND2_X1 U7567 ( .A1(n7201), .A2(n5746), .ZN(n5822) );
  NAND2_X1 U7568 ( .A1(n8906), .A2(n5908), .ZN(n5821) );
  NAND2_X1 U7569 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  XNOR2_X1 U7570 ( .A(n5823), .B(n5937), .ZN(n5826) );
  AOI22_X1 U7571 ( .A1(n7201), .A2(n5908), .B1(n5885), .B2(n8906), .ZN(n5824)
         );
  XNOR2_X1 U7572 ( .A(n5826), .B(n5824), .ZN(n7469) );
  NAND2_X1 U7573 ( .A1(n7468), .A2(n7469), .ZN(n7467) );
  INV_X1 U7574 ( .A(n5824), .ZN(n5825) );
  NAND2_X1 U7575 ( .A1(n7467), .A2(n5827), .ZN(n5830) );
  AOI22_X1 U7576 ( .A1(n5177), .A2(n5746), .B1(n5939), .B2(n8905), .ZN(n5828)
         );
  XNOR2_X1 U7577 ( .A(n5828), .B(n5937), .ZN(n5829) );
  OAI22_X1 U7578 ( .A1(n9768), .A2(n5791), .B1(n8892), .B2(n5817), .ZN(n8754)
         );
  AOI22_X1 U7579 ( .A1(n8895), .A2(n5746), .B1(n5939), .B2(n8904), .ZN(n5834)
         );
  XNOR2_X1 U7580 ( .A(n5834), .B(n5937), .ZN(n5835) );
  OAI22_X1 U7581 ( .A1(n7350), .A2(n5791), .B1(n8809), .B2(n5817), .ZN(n8886)
         );
  NAND2_X1 U7582 ( .A1(n8884), .A2(n5836), .ZN(n8804) );
  NAND2_X1 U7583 ( .A1(n9219), .A2(n5746), .ZN(n5838) );
  NAND2_X1 U7584 ( .A1(n8903), .A2(n5908), .ZN(n5837) );
  NAND2_X1 U7585 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  XNOR2_X1 U7586 ( .A(n5839), .B(n5937), .ZN(n5842) );
  AOI22_X1 U7587 ( .A1(n9219), .A2(n5912), .B1(n5885), .B2(n8903), .ZN(n5840)
         );
  XNOR2_X1 U7588 ( .A(n5842), .B(n5840), .ZN(n8806) );
  INV_X1 U7589 ( .A(n5840), .ZN(n5841) );
  NAND2_X1 U7590 ( .A1(n9213), .A2(n5746), .ZN(n5845) );
  NAND2_X1 U7591 ( .A1(n9124), .A2(n5912), .ZN(n5844) );
  NAND2_X1 U7592 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  XNOR2_X1 U7593 ( .A(n5846), .B(n5937), .ZN(n5850) );
  NAND2_X1 U7594 ( .A1(n9213), .A2(n5912), .ZN(n5848) );
  NAND2_X1 U7595 ( .A1(n9124), .A2(n5885), .ZN(n5847) );
  NAND2_X1 U7596 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  NAND2_X1 U7597 ( .A1(n5850), .A2(n5849), .ZN(n8815) );
  NAND2_X1 U7598 ( .A1(n9208), .A2(n5746), .ZN(n5852) );
  NAND2_X1 U7599 ( .A1(n8902), .A2(n5908), .ZN(n5851) );
  NAND2_X1 U7600 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  XNOR2_X1 U7601 ( .A(n5853), .B(n5937), .ZN(n8863) );
  NAND2_X1 U7602 ( .A1(n9208), .A2(n5939), .ZN(n5855) );
  NAND2_X1 U7603 ( .A1(n8902), .A2(n5885), .ZN(n5854) );
  NAND2_X1 U7604 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  INV_X1 U7605 ( .A(n8863), .ZN(n5857) );
  INV_X1 U7606 ( .A(n5856), .ZN(n8862) );
  NAND2_X1 U7607 ( .A1(n9204), .A2(n5746), .ZN(n5860) );
  NAND2_X1 U7608 ( .A1(n9125), .A2(n5908), .ZN(n5859) );
  NAND2_X1 U7609 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  XNOR2_X1 U7610 ( .A(n5861), .B(n4377), .ZN(n5867) );
  AND2_X1 U7611 ( .A1(n9125), .A2(n5885), .ZN(n5862) );
  AOI21_X1 U7612 ( .B1(n9204), .B2(n5939), .A(n5862), .ZN(n5866) );
  NOR2_X1 U7613 ( .A1(n5867), .A2(n5866), .ZN(n8777) );
  NAND2_X1 U7614 ( .A1(n9199), .A2(n5746), .ZN(n5864) );
  NAND2_X1 U7615 ( .A1(n8901), .A2(n5939), .ZN(n5863) );
  NAND2_X1 U7616 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  XNOR2_X1 U7617 ( .A(n5865), .B(n5937), .ZN(n5870) );
  AOI22_X1 U7618 ( .A1(n9199), .A2(n5912), .B1(n5885), .B2(n8901), .ZN(n5871)
         );
  XNOR2_X1 U7619 ( .A(n5870), .B(n5871), .ZN(n8843) );
  INV_X1 U7620 ( .A(n8843), .ZN(n5868) );
  NAND2_X1 U7621 ( .A1(n5867), .A2(n5866), .ZN(n8840) );
  OR2_X1 U7622 ( .A1(n5868), .A2(n8840), .ZN(n5869) );
  INV_X1 U7623 ( .A(n5870), .ZN(n5872) );
  NAND2_X1 U7624 ( .A1(n5872), .A2(n5871), .ZN(n8785) );
  NAND2_X1 U7625 ( .A1(n9194), .A2(n5746), .ZN(n5874) );
  NAND2_X1 U7626 ( .A1(n9059), .A2(n5908), .ZN(n5873) );
  NAND2_X1 U7627 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  XNOR2_X1 U7628 ( .A(n5875), .B(n5937), .ZN(n5890) );
  INV_X1 U7629 ( .A(n5890), .ZN(n5876) );
  AOI22_X1 U7630 ( .A1(n9194), .A2(n5912), .B1(n5885), .B2(n9059), .ZN(n5889)
         );
  NAND2_X1 U7631 ( .A1(n5876), .A2(n5889), .ZN(n5888) );
  NAND2_X1 U7632 ( .A1(n9188), .A2(n5908), .ZN(n5878) );
  NAND2_X1 U7633 ( .A1(n9047), .A2(n5885), .ZN(n5877) );
  NAND2_X1 U7634 ( .A1(n5878), .A2(n5877), .ZN(n8854) );
  NAND2_X1 U7635 ( .A1(n9188), .A2(n5746), .ZN(n5880) );
  NAND2_X1 U7636 ( .A1(n9047), .A2(n5908), .ZN(n5879) );
  NAND2_X1 U7637 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  XNOR2_X1 U7638 ( .A(n5881), .B(n5937), .ZN(n5895) );
  NAND2_X1 U7639 ( .A1(n9183), .A2(n5746), .ZN(n5883) );
  NAND2_X1 U7640 ( .A1(n9065), .A2(n5912), .ZN(n5882) );
  NAND2_X1 U7641 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  XNOR2_X1 U7642 ( .A(n5884), .B(n4377), .ZN(n8767) );
  NAND2_X1 U7643 ( .A1(n9183), .A2(n5908), .ZN(n5887) );
  NAND2_X1 U7644 ( .A1(n9065), .A2(n5885), .ZN(n5886) );
  NOR2_X1 U7645 ( .A1(n8767), .A2(n8766), .ZN(n8765) );
  AOI21_X1 U7646 ( .B1(n8854), .B2(n5895), .A(n8765), .ZN(n5892) );
  INV_X1 U7647 ( .A(n5888), .ZN(n5891) );
  XNOR2_X1 U7648 ( .A(n5890), .B(n5889), .ZN(n8787) );
  AND2_X1 U7649 ( .A1(n5892), .A2(n8761), .ZN(n5893) );
  NAND2_X1 U7650 ( .A1(n5894), .A2(n5893), .ZN(n5902) );
  INV_X1 U7651 ( .A(n8854), .ZN(n5896) );
  AOI21_X1 U7652 ( .B1(n8762), .B2(n5896), .A(n8766), .ZN(n5899) );
  INV_X1 U7653 ( .A(n8767), .ZN(n5898) );
  NAND3_X1 U7654 ( .A1(n8766), .A2(n5896), .A3(n8762), .ZN(n5897) );
  NAND2_X1 U7655 ( .A1(n5902), .A2(n5901), .ZN(n8822) );
  AOI22_X1 U7656 ( .A1(n9178), .A2(n5746), .B1(n5939), .B2(n9048), .ZN(n5903)
         );
  XOR2_X1 U7657 ( .A(n5937), .B(n5903), .Z(n5905) );
  OAI22_X1 U7658 ( .A1(n9030), .A2(n5791), .B1(n8798), .B2(n5817), .ZN(n5904)
         );
  NOR2_X1 U7659 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  AOI21_X1 U7660 ( .B1(n5905), .B2(n5904), .A(n5906), .ZN(n8824) );
  INV_X1 U7661 ( .A(n5906), .ZN(n5907) );
  NAND2_X1 U7662 ( .A1(n9173), .A2(n5746), .ZN(n5910) );
  NAND2_X1 U7663 ( .A1(n9036), .A2(n5908), .ZN(n5909) );
  NAND2_X1 U7664 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  XNOR2_X1 U7665 ( .A(n5911), .B(n5937), .ZN(n5919) );
  AOI22_X1 U7666 ( .A1(n9173), .A2(n5912), .B1(n5885), .B2(n9036), .ZN(n5917)
         );
  XNOR2_X1 U7667 ( .A(n5919), .B(n5917), .ZN(n8795) );
  NAND2_X1 U7668 ( .A1(n9168), .A2(n5746), .ZN(n5914) );
  NAND2_X1 U7669 ( .A1(n9020), .A2(n5908), .ZN(n5913) );
  NAND2_X1 U7670 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  XNOR2_X1 U7671 ( .A(n5915), .B(n4377), .ZN(n5928) );
  AND2_X1 U7672 ( .A1(n9020), .A2(n5885), .ZN(n5916) );
  AOI21_X1 U7673 ( .B1(n9168), .B2(n5912), .A(n5916), .ZN(n5929) );
  XNOR2_X1 U7674 ( .A(n5928), .B(n5929), .ZN(n8872) );
  INV_X1 U7675 ( .A(n5917), .ZN(n5918) );
  NOR2_X1 U7676 ( .A1(n5919), .A2(n5918), .ZN(n8873) );
  NOR2_X1 U7677 ( .A1(n8872), .A2(n8873), .ZN(n5920) );
  NAND2_X1 U7678 ( .A1(n9164), .A2(n5746), .ZN(n5922) );
  NAND2_X1 U7679 ( .A1(n9005), .A2(n5912), .ZN(n5921) );
  NAND2_X1 U7680 ( .A1(n5922), .A2(n5921), .ZN(n5923) );
  XNOR2_X1 U7681 ( .A(n5923), .B(n5937), .ZN(n5927) );
  NAND2_X1 U7682 ( .A1(n9164), .A2(n5908), .ZN(n5925) );
  NAND2_X1 U7683 ( .A1(n9005), .A2(n5885), .ZN(n5924) );
  NAND2_X1 U7684 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  NOR2_X1 U7685 ( .A1(n5927), .A2(n5926), .ZN(n5948) );
  AOI21_X1 U7686 ( .B1(n5927), .B2(n5926), .A(n5948), .ZN(n6477) );
  INV_X1 U7687 ( .A(n6477), .ZN(n5933) );
  INV_X1 U7688 ( .A(n5928), .ZN(n5931) );
  INV_X1 U7689 ( .A(n5929), .ZN(n5930) );
  NAND2_X1 U7690 ( .A1(n5931), .A2(n5930), .ZN(n6478) );
  INV_X1 U7691 ( .A(n6478), .ZN(n5932) );
  NOR2_X1 U7692 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  INV_X1 U7693 ( .A(n6480), .ZN(n5947) );
  NAND2_X1 U7694 ( .A1(n9157), .A2(n5912), .ZN(n5936) );
  NAND2_X1 U7695 ( .A1(n8985), .A2(n5885), .ZN(n5935) );
  NAND2_X1 U7696 ( .A1(n5936), .A2(n5935), .ZN(n5938) );
  XNOR2_X1 U7697 ( .A(n5938), .B(n5937), .ZN(n5941) );
  AOI22_X1 U7698 ( .A1(n9157), .A2(n5746), .B1(n5939), .B2(n8985), .ZN(n5940)
         );
  XNOR2_X1 U7699 ( .A(n5941), .B(n5940), .ZN(n5949) );
  INV_X1 U7700 ( .A(n5949), .ZN(n5946) );
  INV_X1 U7701 ( .A(n5948), .ZN(n5944) );
  NAND3_X1 U7702 ( .A1(n6486), .A2(n6470), .A3(n5942), .ZN(n5951) );
  INV_X1 U7703 ( .A(n5943), .ZN(n7886) );
  AND2_X1 U7704 ( .A1(n9767), .A2(n7823), .ZN(n5952) );
  NAND3_X1 U7705 ( .A1(n6480), .A2(n8876), .A3(n5949), .ZN(n5971) );
  NAND3_X1 U7706 ( .A1(n5949), .A2(n8876), .A3(n5948), .ZN(n5970) );
  INV_X1 U7707 ( .A(n5963), .ZN(n5950) );
  INV_X1 U7708 ( .A(n5951), .ZN(n5961) );
  INV_X1 U7709 ( .A(n5952), .ZN(n5953) );
  NOR2_X1 U7710 ( .A1(n5961), .A2(n5953), .ZN(n5957) );
  INV_X1 U7711 ( .A(n6562), .ZN(n5955) );
  NOR4_X1 U7712 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n5962)
         );
  INV_X1 U7713 ( .A(n5958), .ZN(n5959) );
  AOI22_X1 U7714 ( .A1(n9380), .A2(n6801), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5959), .ZN(n5960) );
  OAI22_X2 U7715 ( .A1(n5962), .A2(P1_U3086), .B1(n5961), .B2(n5960), .ZN(
        n8889) );
  AOI22_X1 U7716 ( .A1(n8889), .A2(n5964), .B1(n8887), .B2(n8900), .ZN(n5967)
         );
  AOI22_X1 U7717 ( .A1(n8878), .A2(n9005), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5966) );
  NAND2_X1 U7718 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  AOI21_X1 U7719 ( .B1(n9157), .B2(n8894), .A(n5968), .ZN(n5969) );
  NAND4_X1 U7720 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(
        P1_U3220) );
  NAND2_X1 U7721 ( .A1(n5976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5978) );
  AND2_X4 U7722 ( .A1(n5979), .A2(n5980), .ZN(n6183) );
  NAND2_X1 U7723 ( .A1(n6183), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7724 ( .A1(n4271), .A2(n8458), .ZN(n5987) );
  OR2_X1 U7725 ( .A1(n6077), .A2(n8453), .ZN(n5986) );
  NAND2_X1 U7726 ( .A1(n6049), .A2(n6048), .ZN(n6063) );
  NOR2_X2 U7727 ( .A1(n6144), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6154) );
  INV_X1 U7728 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7729 ( .A1(n6154), .A2(n6153), .ZN(n6163) );
  INV_X1 U7730 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6184) );
  INV_X1 U7731 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5983) );
  OR2_X1 U7732 ( .A1(n6187), .A2(n5983), .ZN(n5984) );
  AND2_X1 U7733 ( .A1(n6197), .A2(n5984), .ZN(n8619) );
  OR2_X1 U7734 ( .A1(n4268), .A2(n8619), .ZN(n5985) );
  INV_X1 U7735 ( .A(n8604), .ZN(n8382) );
  INV_X2 U7736 ( .A(n6082), .ZN(n6095) );
  NAND2_X1 U7737 ( .A1(n6733), .A2(n6095), .ZN(n5992) );
  NAND2_X4 U7738 ( .A1(n5989), .A2(n7725), .ZN(n8291) );
  INV_X2 U7739 ( .A(n8291), .ZN(n6205) );
  AOI22_X1 U7740 ( .A1(n6205), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6204), .B2(
        n5990), .ZN(n5991) );
  NAND2_X1 U7741 ( .A1(n5992), .A2(n5991), .ZN(n8067) );
  NAND2_X1 U7742 ( .A1(n6183), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5996) );
  OR2_X1 U7743 ( .A1(n6077), .A2(n9809), .ZN(n5995) );
  INV_X1 U7744 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5993) );
  OR2_X1 U7745 ( .A1(n8291), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6001) );
  OR2_X1 U7746 ( .A1(n6082), .A2(n5998), .ZN(n6000) );
  NAND2_X1 U7747 ( .A1(n6204), .A2(n9818), .ZN(n5999) );
  NAND2_X1 U7748 ( .A1(n6183), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6007) );
  INV_X1 U7749 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6002) );
  OR2_X1 U7750 ( .A1(n6101), .A2(n6002), .ZN(n6006) );
  OR2_X1 U7751 ( .A1(n4271), .A2(n9935), .ZN(n6005) );
  OR2_X1 U7752 ( .A1(n6077), .A2(n6003), .ZN(n6004) );
  NAND4_X1 U7753 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n8394)
         );
  NAND2_X1 U7754 ( .A1(n6008), .A2(SI_0_), .ZN(n6010) );
  INV_X1 U7755 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7756 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  AND2_X1 U7757 ( .A1(n6012), .A2(n6011), .ZN(n6530) );
  MUX2_X1 U7758 ( .A(P2_IR_REG_0__SCAN_IN), .B(n6530), .S(n5989), .Z(n9875) );
  NAND2_X1 U7759 ( .A1(n8394), .A2(n9875), .ZN(n6835) );
  NAND2_X1 U7760 ( .A1(n6834), .A2(n6835), .ZN(n6015) );
  NAND2_X1 U7761 ( .A1(n6929), .A2(n6013), .ZN(n6014) );
  NAND2_X1 U7762 ( .A1(n6015), .A2(n6014), .ZN(n7025) );
  INV_X1 U7763 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7764 ( .A1(n6077), .A2(n7031), .ZN(n6020) );
  INV_X1 U7765 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6018) );
  OR2_X1 U7766 ( .A1(n6101), .A2(n6018), .ZN(n6019) );
  OR2_X1 U7767 ( .A1(n6082), .A2(n6535), .ZN(n6023) );
  INV_X1 U7768 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6021) );
  OAI211_X1 U7769 ( .C1(n5989), .C2(n4269), .A(n6023), .B(n6022), .ZN(n6870)
         );
  NAND2_X1 U7770 ( .A1(n6881), .A2(n6870), .ZN(n8159) );
  NAND2_X1 U7771 ( .A1(n6922), .A2(n9879), .ZN(n8158) );
  NAND2_X1 U7772 ( .A1(n8159), .A2(n8158), .ZN(n8315) );
  NAND2_X1 U7773 ( .A1(n7025), .A2(n8315), .ZN(n6025) );
  NAND2_X1 U7774 ( .A1(n6881), .A2(n9879), .ZN(n6024) );
  NAND2_X1 U7775 ( .A1(n6183), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6030) );
  OR2_X1 U7776 ( .A1(n6101), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6029) );
  INV_X1 U7777 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6026) );
  OR2_X1 U7778 ( .A1(n4271), .A2(n6026), .ZN(n6028) );
  OR2_X1 U7779 ( .A1(n6077), .A2(n9869), .ZN(n6027) );
  OR2_X1 U7780 ( .A1(n6082), .A2(n6547), .ZN(n6032) );
  OR2_X1 U7781 ( .A1(n8291), .A2(n6548), .ZN(n6031) );
  OAI211_X1 U7782 ( .C1(n5989), .C2(n6546), .A(n6032), .B(n6031), .ZN(n6033)
         );
  NAND2_X1 U7783 ( .A1(n6183), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6039) );
  OR2_X1 U7784 ( .A1(n4271), .A2(n6034), .ZN(n6038) );
  AND2_X1 U7785 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6035) );
  NOR2_X1 U7786 ( .A1(n6049), .A2(n6035), .ZN(n6899) );
  OR2_X1 U7787 ( .A1(n6101), .A2(n6899), .ZN(n6037) );
  OR2_X1 U7788 ( .A1(n6077), .A2(n7129), .ZN(n6036) );
  OR2_X1 U7789 ( .A1(n6082), .A2(n6549), .ZN(n6042) );
  OR2_X1 U7790 ( .A1(n8291), .A2(n6550), .ZN(n6041) );
  OR2_X1 U7791 ( .A1(n5989), .A2(n9838), .ZN(n6040) );
  NAND2_X1 U7792 ( .A1(n8165), .A2(n9890), .ZN(n6057) );
  NAND2_X1 U7793 ( .A1(n6877), .A2(n8166), .ZN(n6043) );
  INV_X1 U7794 ( .A(n8316), .ZN(n6044) );
  NAND2_X1 U7795 ( .A1(n8393), .A2(n6033), .ZN(n7124) );
  AND2_X1 U7796 ( .A1(n6044), .A2(n7124), .ZN(n6055) );
  NAND2_X1 U7797 ( .A1(n7126), .A2(n6057), .ZN(n7151) );
  OR2_X1 U7798 ( .A1(n6082), .A2(n6541), .ZN(n6047) );
  OR2_X1 U7799 ( .A1(n8291), .A2(n6539), .ZN(n6046) );
  OR2_X1 U7800 ( .A1(n5989), .A2(n6538), .ZN(n6045) );
  NAND2_X1 U7801 ( .A1(n6183), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7802 ( .A1(n4271), .A2(n9941), .ZN(n6053) );
  OR2_X1 U7803 ( .A1(n6077), .A2(n6708), .ZN(n6052) );
  OR2_X1 U7804 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  AND2_X1 U7805 ( .A1(n6063), .A2(n6050), .ZN(n6939) );
  OR2_X1 U7806 ( .A1(n4268), .A2(n6939), .ZN(n6051) );
  OAI21_X1 U7807 ( .B1(n7151), .B2(n6942), .A(n7172), .ZN(n6061) );
  AND2_X1 U7808 ( .A1(n6055), .A2(n6942), .ZN(n6056) );
  NAND2_X1 U7809 ( .A1(n6056), .A2(n7125), .ZN(n6059) );
  INV_X1 U7810 ( .A(n6942), .ZN(n9894) );
  OR2_X1 U7811 ( .A1(n9894), .A2(n6057), .ZN(n6058) );
  AND2_X1 U7812 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  NAND2_X1 U7813 ( .A1(n6061), .A2(n6060), .ZN(n7171) );
  INV_X1 U7814 ( .A(n7171), .ZN(n6073) );
  NAND2_X1 U7815 ( .A1(n6420), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6069) );
  INV_X1 U7816 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6062) );
  OR2_X1 U7817 ( .A1(n6199), .A2(n6062), .ZN(n6068) );
  NAND2_X1 U7818 ( .A1(n6063), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6064) );
  AND2_X1 U7819 ( .A1(n6075), .A2(n6064), .ZN(n7175) );
  OR2_X1 U7820 ( .A1(n6101), .A2(n7175), .ZN(n6067) );
  OR2_X1 U7821 ( .A1(n6077), .A2(n6065), .ZN(n6066) );
  OR2_X1 U7822 ( .A1(n6082), .A2(n6544), .ZN(n6071) );
  OR2_X1 U7823 ( .A1(n8291), .A2(n6545), .ZN(n6070) );
  OAI211_X1 U7824 ( .C1(n5989), .C2(n6543), .A(n6071), .B(n6070), .ZN(n7177)
         );
  NAND2_X1 U7825 ( .A1(n7283), .A2(n7177), .ZN(n8178) );
  INV_X1 U7826 ( .A(n7177), .ZN(n9900) );
  NAND2_X1 U7827 ( .A1(n8391), .A2(n9900), .ZN(n8175) );
  NAND2_X1 U7828 ( .A1(n6183), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6081) );
  OR2_X1 U7829 ( .A1(n4271), .A2(n6074), .ZN(n6080) );
  AND2_X1 U7830 ( .A1(n6075), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6076) );
  NOR2_X1 U7831 ( .A1(n6087), .A2(n6076), .ZN(n7289) );
  OR2_X1 U7832 ( .A1(n6101), .A2(n7289), .ZN(n6079) );
  OR2_X1 U7833 ( .A1(n6077), .A2(n6521), .ZN(n6078) );
  OR2_X1 U7834 ( .A1(n6553), .A2(n6082), .ZN(n6084) );
  OR2_X1 U7835 ( .A1(n8291), .A2(n6554), .ZN(n6083) );
  OAI211_X1 U7836 ( .C1(n5989), .C2(n6552), .A(n6084), .B(n6083), .ZN(n6085)
         );
  NAND2_X1 U7837 ( .A1(n7919), .A2(n6085), .ZN(n8189) );
  INV_X1 U7838 ( .A(n7919), .ZN(n8390) );
  NAND2_X1 U7839 ( .A1(n8390), .A2(n9903), .ZN(n7307) );
  NAND2_X1 U7840 ( .A1(n8189), .A2(n7307), .ZN(n8323) );
  NAND2_X1 U7841 ( .A1(n6183), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6092) );
  NOR2_X1 U7842 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  OR2_X1 U7843 ( .A1(n6101), .A2(n4857), .ZN(n6090) );
  OR2_X1 U7844 ( .A1(n6077), .A2(n5608), .ZN(n6089) );
  AOI22_X1 U7845 ( .A1(n6205), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6204), .B2(
        n6093), .ZN(n6108) );
  NAND2_X1 U7846 ( .A1(n6555), .A2(n6095), .ZN(n6107) );
  AND2_X1 U7847 ( .A1(n6108), .A2(n6107), .ZN(n7310) );
  NAND2_X1 U7848 ( .A1(n7282), .A2(n7310), .ZN(n7358) );
  AOI22_X1 U7849 ( .A1(n6205), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6204), .B2(
        n6094), .ZN(n6097) );
  NAND2_X1 U7850 ( .A1(n6566), .A2(n6095), .ZN(n6096) );
  NAND2_X1 U7851 ( .A1(n6183), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6106) );
  OR2_X1 U7852 ( .A1(n4271), .A2(n6098), .ZN(n6105) );
  OR2_X1 U7853 ( .A1(n6099), .A2(n7111), .ZN(n6100) );
  AND2_X1 U7854 ( .A1(n6116), .A2(n6100), .ZN(n7365) );
  OR2_X1 U7855 ( .A1(n4268), .A2(n7365), .ZN(n6104) );
  OR2_X1 U7856 ( .A1(n6077), .A2(n6102), .ZN(n6103) );
  NAND2_X1 U7857 ( .A1(n9908), .A2(n7916), .ZN(n6110) );
  INV_X1 U7858 ( .A(n6124), .ZN(n6109) );
  NAND2_X1 U7859 ( .A1(n6108), .A2(n6107), .ZN(n7239) );
  NAND2_X1 U7860 ( .A1(n7282), .A2(n7239), .ZN(n8190) );
  INV_X1 U7861 ( .A(n7282), .ZN(n8389) );
  NAND2_X1 U7862 ( .A1(n8389), .A2(n7310), .ZN(n8182) );
  INV_X1 U7863 ( .A(n6110), .ZN(n6112) );
  INV_X1 U7864 ( .A(n9908), .ZN(n6111) );
  NAND2_X1 U7865 ( .A1(n6568), .A2(n6095), .ZN(n6115) );
  AOI22_X1 U7866 ( .A1(n6205), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6204), .B2(
        n7225), .ZN(n6114) );
  NAND2_X1 U7867 ( .A1(n6115), .A2(n6114), .ZN(n7411) );
  NAND2_X1 U7868 ( .A1(n6183), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6121) );
  OR2_X1 U7869 ( .A1(n4271), .A2(n9946), .ZN(n6120) );
  NAND2_X1 U7870 ( .A1(n6116), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6117) );
  AND2_X1 U7871 ( .A1(n6135), .A2(n6117), .ZN(n7415) );
  OR2_X1 U7872 ( .A1(n6101), .A2(n7415), .ZN(n6119) );
  OR2_X1 U7873 ( .A1(n6077), .A2(n5679), .ZN(n6118) );
  NAND4_X1 U7874 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), .ZN(n8388)
         );
  NAND2_X1 U7875 ( .A1(n7411), .A2(n8388), .ZN(n8202) );
  NAND2_X1 U7876 ( .A1(n8391), .A2(n7177), .ZN(n7272) );
  NOR2_X1 U7877 ( .A1(n7411), .A2(n8388), .ZN(n7331) );
  INV_X1 U7878 ( .A(n7331), .ZN(n6129) );
  NAND2_X1 U7879 ( .A1(n7919), .A2(n9903), .ZN(n7301) );
  AND2_X1 U7880 ( .A1(n7301), .A2(n6124), .ZN(n6125) );
  AND2_X1 U7881 ( .A1(n6129), .A2(n7336), .ZN(n6130) );
  INV_X1 U7882 ( .A(n8202), .ZN(n7332) );
  NAND2_X1 U7883 ( .A1(n6583), .A2(n6095), .ZN(n6134) );
  AOI22_X1 U7884 ( .A1(n6205), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6204), .B2(
        n7509), .ZN(n6133) );
  NAND2_X1 U7885 ( .A1(n6134), .A2(n6133), .ZN(n9920) );
  NAND2_X1 U7886 ( .A1(n6183), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7887 ( .A1(n4271), .A2(n9948), .ZN(n6139) );
  NAND2_X1 U7888 ( .A1(n6135), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6136) );
  AND2_X1 U7889 ( .A1(n6144), .A2(n6136), .ZN(n7461) );
  OR2_X1 U7890 ( .A1(n6101), .A2(n7461), .ZN(n6138) );
  OR2_X1 U7891 ( .A1(n6077), .A2(n7505), .ZN(n6137) );
  NAND4_X1 U7892 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n8387)
         );
  NAND2_X1 U7893 ( .A1(n6599), .A2(n6095), .ZN(n6142) );
  AOI22_X1 U7894 ( .A1(n6205), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6204), .B2(
        n7611), .ZN(n6141) );
  NAND2_X1 U7895 ( .A1(n6183), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6149) );
  OR2_X1 U7896 ( .A1(n4271), .A2(n6143), .ZN(n6148) );
  AND2_X1 U7897 ( .A1(n6144), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6145) );
  NOR2_X1 U7898 ( .A1(n6154), .A2(n6145), .ZN(n7519) );
  OR2_X1 U7899 ( .A1(n6101), .A2(n7519), .ZN(n6147) );
  OR2_X1 U7900 ( .A1(n6077), .A2(n7327), .ZN(n6146) );
  NAND4_X1 U7901 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n8386)
         );
  XNOR2_X1 U7902 ( .A(n9930), .B(n8386), .ZN(n8209) );
  NAND2_X1 U7903 ( .A1(n9930), .A2(n8386), .ZN(n6150) );
  NAND2_X1 U7904 ( .A1(n6607), .A2(n6095), .ZN(n6152) );
  AOI22_X1 U7905 ( .A1(n6205), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6204), .B2(
        n7561), .ZN(n6151) );
  NAND2_X1 U7906 ( .A1(n6152), .A2(n6151), .ZN(n7632) );
  NAND2_X1 U7907 ( .A1(n6183), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6159) );
  OR2_X1 U7908 ( .A1(n4271), .A2(n9459), .ZN(n6158) );
  OR2_X1 U7909 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  AND2_X1 U7910 ( .A1(n6155), .A2(n6163), .ZN(n7630) );
  OR2_X1 U7911 ( .A1(n4268), .A2(n7630), .ZN(n6157) );
  OR2_X1 U7912 ( .A1(n6077), .A2(n7560), .ZN(n6156) );
  NAND4_X1 U7913 ( .A1(n6159), .A2(n6158), .A3(n6157), .A4(n6156), .ZN(n8385)
         );
  OR2_X1 U7914 ( .A1(n7632), .A2(n8385), .ZN(n6160) );
  NAND2_X1 U7915 ( .A1(n7437), .A2(n6160), .ZN(n7433) );
  NAND2_X1 U7916 ( .A1(n7632), .A2(n8385), .ZN(n7434) );
  NAND2_X1 U7917 ( .A1(n7433), .A2(n7434), .ZN(n7524) );
  NAND2_X1 U7918 ( .A1(n6651), .A2(n6095), .ZN(n6162) );
  AOI22_X1 U7919 ( .A1(n6205), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6204), .B2(
        n8411), .ZN(n6161) );
  NAND2_X1 U7920 ( .A1(n6183), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6168) );
  INV_X1 U7921 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7528) );
  OR2_X1 U7922 ( .A1(n4271), .A2(n7528), .ZN(n6167) );
  INV_X1 U7923 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7535) );
  OR2_X1 U7924 ( .A1(n6077), .A2(n7535), .ZN(n6166) );
  NAND2_X1 U7925 ( .A1(n6163), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6164) );
  AND2_X1 U7926 ( .A1(n6173), .A2(n6164), .ZN(n7536) );
  OR2_X1 U7927 ( .A1(n6101), .A2(n7536), .ZN(n6165) );
  NAND4_X1 U7928 ( .A1(n6168), .A2(n6167), .A3(n6166), .A4(n6165), .ZN(n8384)
         );
  OR2_X1 U7929 ( .A1(n7990), .A2(n8384), .ZN(n6169) );
  NAND2_X1 U7930 ( .A1(n7990), .A2(n8384), .ZN(n6170) );
  NAND2_X1 U7931 ( .A1(n6675), .A2(n6095), .ZN(n6172) );
  AOI22_X1 U7932 ( .A1(n6205), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6204), .B2(
        n8417), .ZN(n6171) );
  NAND2_X1 U7933 ( .A1(n6183), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6178) );
  OR2_X1 U7934 ( .A1(n4271), .A2(n8424), .ZN(n6177) );
  AND2_X1 U7935 ( .A1(n6173), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6174) );
  NOR2_X1 U7936 ( .A1(n6185), .A2(n6174), .ZN(n7554) );
  OR2_X1 U7937 ( .A1(n6101), .A2(n7554), .ZN(n6176) );
  OR2_X1 U7938 ( .A1(n6077), .A2(n8416), .ZN(n6175) );
  NAND4_X1 U7939 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(n8383)
         );
  AND2_X1 U7940 ( .A1(n8225), .A2(n8383), .ZN(n7543) );
  INV_X1 U7941 ( .A(n7543), .ZN(n6179) );
  OR2_X1 U7942 ( .A1(n8225), .A2(n8383), .ZN(n7544) );
  NAND2_X1 U7943 ( .A1(n6180), .A2(n7544), .ZN(n7576) );
  INV_X1 U7944 ( .A(n7576), .ZN(n6194) );
  NAND2_X1 U7945 ( .A1(n6770), .A2(n6095), .ZN(n6182) );
  AOI22_X1 U7946 ( .A1(n6205), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6204), .B2(
        n8448), .ZN(n6181) );
  NAND2_X1 U7947 ( .A1(n6183), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6192) );
  INV_X1 U7948 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7583) );
  OR2_X1 U7949 ( .A1(n4271), .A2(n7583), .ZN(n6191) );
  NOR2_X1 U7950 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  OR2_X1 U7951 ( .A1(n6187), .A2(n6186), .ZN(n8063) );
  INV_X1 U7952 ( .A(n8063), .ZN(n6188) );
  OR2_X1 U7953 ( .A1(n4268), .A2(n6188), .ZN(n6190) );
  INV_X1 U7954 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7586) );
  OR2_X1 U7955 ( .A1(n6077), .A2(n7586), .ZN(n6189) );
  NAND2_X1 U7956 ( .A1(n8053), .A2(n8139), .ZN(n8230) );
  INV_X1 U7957 ( .A(n8335), .ZN(n6193) );
  NAND2_X1 U7958 ( .A1(n6194), .A2(n6193), .ZN(n8623) );
  NAND2_X1 U7959 ( .A1(n8053), .A2(n8626), .ZN(n8621) );
  OR2_X1 U7960 ( .A1(n8067), .A2(n8604), .ZN(n8236) );
  NAND2_X1 U7961 ( .A1(n8067), .A2(n8604), .ZN(n8234) );
  NAND2_X1 U7962 ( .A1(n6799), .A2(n6095), .ZN(n6196) );
  AOI22_X1 U7963 ( .A1(n6205), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6204), .B2(
        n8484), .ZN(n6195) );
  NAND2_X1 U7964 ( .A1(n6197), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7965 ( .A1(n6208), .A2(n6198), .ZN(n8609) );
  NAND2_X1 U7966 ( .A1(n6307), .A2(n8609), .ZN(n6203) );
  INV_X1 U7967 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8732) );
  OR2_X1 U7968 ( .A1(n6199), .A2(n8732), .ZN(n6202) );
  OR2_X1 U7969 ( .A1(n4271), .A2(n8669), .ZN(n6201) );
  OR2_X1 U7970 ( .A1(n6077), .A2(n8611), .ZN(n6200) );
  NAND4_X1 U7971 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(n8625)
         );
  INV_X1 U7972 ( .A(n8668), .ZN(n8123) );
  NAND2_X1 U7973 ( .A1(n7066), .A2(n6095), .ZN(n6207) );
  AOI22_X1 U7974 ( .A1(n6205), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8368), .B2(
        n6204), .ZN(n6206) );
  AND2_X1 U7975 ( .A1(n6208), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6209) );
  NOR2_X2 U7976 ( .A1(n6208), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6218) );
  OR2_X1 U7977 ( .A1(n6209), .A2(n6218), .ZN(n8014) );
  NAND2_X1 U7978 ( .A1(n6307), .A2(n8014), .ZN(n6214) );
  INV_X1 U7979 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9298) );
  OR2_X1 U7980 ( .A1(n6199), .A2(n9298), .ZN(n6213) );
  OR2_X1 U7981 ( .A1(n4271), .A2(n6210), .ZN(n6212) );
  OR2_X1 U7982 ( .A1(n6077), .A2(n5636), .ZN(n6211) );
  NAND2_X1 U7983 ( .A1(n8661), .A2(n8606), .ZN(n8243) );
  NAND2_X1 U7984 ( .A1(n8575), .A2(n8243), .ZN(n8313) );
  INV_X1 U7985 ( .A(n8606), .ZN(n8582) );
  NAND2_X1 U7986 ( .A1(n7133), .A2(n6095), .ZN(n6216) );
  OR2_X1 U7987 ( .A1(n8291), .A2(n9349), .ZN(n6215) );
  INV_X1 U7988 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8584) );
  INV_X1 U7989 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6217) );
  NOR2_X1 U7990 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  OR2_X1 U7991 ( .A1(n6227), .A2(n6219), .ZN(n8585) );
  NAND2_X1 U7992 ( .A1(n8585), .A2(n6307), .ZN(n6223) );
  NAND2_X1 U7993 ( .A1(n6183), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7994 ( .A1(n6420), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6220) );
  AND2_X1 U7995 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  OAI211_X1 U7996 ( .C1(n6077), .C2(n8584), .A(n6223), .B(n6222), .ZN(n8589)
         );
  NAND2_X1 U7997 ( .A1(n7955), .A2(n8589), .ZN(n8245) );
  INV_X1 U7998 ( .A(n8589), .ZN(n8042) );
  NAND2_X1 U7999 ( .A1(n8726), .A2(n8042), .ZN(n8244) );
  NAND2_X1 U8000 ( .A1(n8245), .A2(n8244), .ZN(n8579) );
  NAND2_X1 U8001 ( .A1(n8580), .A2(n8579), .ZN(n8578) );
  NAND2_X1 U8002 ( .A1(n7955), .A2(n8042), .ZN(n8563) );
  NAND2_X1 U8003 ( .A1(n7160), .A2(n6095), .ZN(n6225) );
  OR2_X1 U8004 ( .A1(n8291), .A2(n7161), .ZN(n6224) );
  INV_X1 U8005 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6226) );
  OR2_X1 U8006 ( .A1(n6227), .A2(n6226), .ZN(n6228) );
  NAND2_X1 U8007 ( .A1(n6234), .A2(n6228), .ZN(n8570) );
  NAND2_X1 U8008 ( .A1(n8570), .A2(n6307), .ZN(n6231) );
  AOI22_X1 U8009 ( .A1(n6183), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n6420), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U8010 ( .A1(n6419), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U8011 ( .A1(n8719), .A2(n7957), .ZN(n8249) );
  NOR2_X1 U8012 ( .A1(n8719), .A2(n8581), .ZN(n8552) );
  NAND2_X1 U8013 ( .A1(n7232), .A2(n6095), .ZN(n6233) );
  OR2_X1 U8014 ( .A1(n8291), .A2(n9297), .ZN(n6232) );
  NAND2_X1 U8015 ( .A1(n6234), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U8016 ( .A1(n6242), .A2(n6235), .ZN(n8558) );
  NAND2_X1 U8017 ( .A1(n8558), .A2(n6307), .ZN(n6238) );
  AOI22_X1 U8018 ( .A1(n6183), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n6420), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U8019 ( .A1(n6419), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U8020 ( .A1(n8713), .A2(n8542), .ZN(n8254) );
  NAND2_X1 U8021 ( .A1(n8253), .A2(n8254), .ZN(n8551) );
  NAND2_X1 U8022 ( .A1(n8554), .A2(n6239), .ZN(n8539) );
  NAND2_X1 U8023 ( .A1(n7297), .A2(n6095), .ZN(n6241) );
  OR2_X1 U8024 ( .A1(n8291), .A2(n7300), .ZN(n6240) );
  NAND2_X1 U8025 ( .A1(n6242), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U8026 ( .A1(n6253), .A2(n6243), .ZN(n8545) );
  NAND2_X1 U8027 ( .A1(n8545), .A2(n6307), .ZN(n6248) );
  INV_X1 U8028 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U8029 ( .A1(n6420), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U8030 ( .A1(n6419), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6244) );
  OAI211_X1 U8031 ( .C1(n9327), .C2(n6199), .A(n6245), .B(n6244), .ZN(n6246)
         );
  INV_X1 U8032 ( .A(n6246), .ZN(n6247) );
  NAND2_X1 U8033 ( .A1(n6248), .A2(n6247), .ZN(n8555) );
  NAND2_X1 U8034 ( .A1(n8546), .A2(n8555), .ZN(n6250) );
  NAND2_X1 U8035 ( .A1(n7381), .A2(n6095), .ZN(n6252) );
  OR2_X1 U8036 ( .A1(n8291), .A2(n7382), .ZN(n6251) );
  NOR2_X2 U8037 ( .A1(n6253), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6265) );
  INV_X1 U8038 ( .A(n6265), .ZN(n6255) );
  NAND2_X1 U8039 ( .A1(n6253), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U8040 ( .A1(n6255), .A2(n6254), .ZN(n8534) );
  NAND2_X1 U8041 ( .A1(n8534), .A2(n6307), .ZN(n6260) );
  INV_X1 U8042 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U8043 ( .A1(n6419), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U8044 ( .A1(n6420), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6256) );
  OAI211_X1 U8045 ( .C1(n6199), .C2(n8701), .A(n6257), .B(n6256), .ZN(n6258)
         );
  INV_X1 U8046 ( .A(n6258), .ZN(n6259) );
  NAND2_X1 U8047 ( .A1(n8528), .A2(n6261), .ZN(n6262) );
  INV_X1 U8048 ( .A(n8702), .ZN(n8646) );
  NAND2_X1 U8049 ( .A1(n7446), .A2(n6095), .ZN(n6264) );
  OR2_X1 U8050 ( .A1(n8291), .A2(n7447), .ZN(n6263) );
  NAND2_X1 U8051 ( .A1(n6265), .A2(n9230), .ZN(n6276) );
  OR2_X1 U8052 ( .A1(n6265), .A2(n9230), .ZN(n6266) );
  NAND2_X1 U8053 ( .A1(n6276), .A2(n6266), .ZN(n8522) );
  NAND2_X1 U8054 ( .A1(n8522), .A2(n6307), .ZN(n6271) );
  INV_X1 U8055 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U8056 ( .A1(n6420), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U8057 ( .A1(n6183), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6267) );
  OAI211_X1 U8058 ( .C1(n8521), .C2(n6077), .A(n6268), .B(n6267), .ZN(n6269)
         );
  INV_X1 U8059 ( .A(n6269), .ZN(n6270) );
  NOR2_X1 U8060 ( .A1(n7977), .A2(n8531), .ZN(n6273) );
  NAND2_X1 U8061 ( .A1(n7477), .A2(n6095), .ZN(n6275) );
  OR2_X1 U8062 ( .A1(n8291), .A2(n7478), .ZN(n6274) );
  NAND2_X1 U8063 ( .A1(n6276), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U8064 ( .A1(n6286), .A2(n6277), .ZN(n8511) );
  NAND2_X1 U8065 ( .A1(n8511), .A2(n6307), .ZN(n6282) );
  INV_X1 U8066 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U8067 ( .A1(n6419), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U8068 ( .A1(n6420), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6278) );
  OAI211_X1 U8069 ( .C1(n6199), .C2(n9325), .A(n6279), .B(n6278), .ZN(n6280)
         );
  INV_X1 U8070 ( .A(n6280), .ZN(n6281) );
  NAND2_X2 U8071 ( .A1(n6282), .A2(n6281), .ZN(n8518) );
  NOR2_X1 U8072 ( .A1(n8512), .A2(n8518), .ZN(n6283) );
  INV_X1 U8073 ( .A(n8512), .ZN(n8690) );
  NAND2_X1 U8074 ( .A1(n7540), .A2(n6095), .ZN(n6285) );
  OR2_X1 U8075 ( .A1(n8291), .A2(n7541), .ZN(n6284) );
  INV_X1 U8076 ( .A(n6297), .ZN(n6288) );
  NAND2_X1 U8077 ( .A1(n6286), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U8078 ( .A1(n6288), .A2(n6287), .ZN(n8501) );
  NAND2_X1 U8079 ( .A1(n8501), .A2(n6307), .ZN(n6293) );
  INV_X1 U8080 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U8081 ( .A1(n6420), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U8082 ( .A1(n6419), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6289) );
  OAI211_X1 U8083 ( .C1(n8684), .C2(n6199), .A(n6290), .B(n6289), .ZN(n6291)
         );
  INV_X1 U8084 ( .A(n6291), .ZN(n6292) );
  NOR2_X1 U8085 ( .A1(n8271), .A2(n8508), .ZN(n6294) );
  INV_X1 U8086 ( .A(n8508), .ZN(n8380) );
  NAND2_X1 U8087 ( .A1(n7591), .A2(n6095), .ZN(n6296) );
  OR2_X1 U8088 ( .A1(n8291), .A2(n7592), .ZN(n6295) );
  INV_X1 U8089 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8027) );
  NOR2_X1 U8090 ( .A1(n6297), .A2(n8027), .ZN(n6298) );
  NAND2_X1 U8091 ( .A1(n8028), .A2(n6307), .ZN(n6304) );
  INV_X1 U8092 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U8093 ( .A1(n6419), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U8094 ( .A1(n6420), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6299) );
  OAI211_X1 U8095 ( .C1(n6199), .C2(n6301), .A(n6300), .B(n6299), .ZN(n6302)
         );
  INV_X1 U8096 ( .A(n6302), .ZN(n6303) );
  NAND2_X2 U8097 ( .A1(n6304), .A2(n6303), .ZN(n8498) );
  XNOR2_X2 U8098 ( .A(n8286), .B(n8498), .ZN(n8308) );
  XNOR2_X1 U8099 ( .A(n6405), .B(n8308), .ZN(n6317) );
  INV_X1 U8100 ( .A(n8303), .ZN(n8360) );
  NAND2_X1 U8101 ( .A1(n6858), .A2(n8360), .ZN(n8355) );
  NAND2_X1 U8102 ( .A1(n8368), .A2(n8373), .ZN(n6377) );
  NAND2_X1 U8103 ( .A1(n8487), .A2(n6307), .ZN(n8300) );
  INV_X1 U8104 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U8105 ( .A1(n6420), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U8106 ( .A1(n6419), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6308) );
  OAI211_X1 U8107 ( .C1(n9247), .C2(n6199), .A(n6309), .B(n6308), .ZN(n6310)
         );
  INV_X1 U8108 ( .A(n6310), .ZN(n6311) );
  INV_X1 U8109 ( .A(n8370), .ZN(n6312) );
  NAND2_X1 U8110 ( .A1(n8371), .A2(n6312), .ZN(n6313) );
  NAND2_X1 U8111 ( .A1(n5989), .A2(n6313), .ZN(n6757) );
  NOR2_X1 U8112 ( .A1(n8030), .A2(n8607), .ZN(n6315) );
  INV_X1 U8113 ( .A(n6757), .ZN(n6871) );
  OAI21_X1 U8114 ( .B1(n6317), .B2(n9872), .A(n6316), .ZN(n6392) );
  NAND2_X1 U8115 ( .A1(n8303), .A2(n8368), .ZN(n6380) );
  NOR2_X1 U8116 ( .A1(n9913), .A2(n6380), .ZN(n6324) );
  XNOR2_X1 U8117 ( .A(n7383), .B(P2_B_REG_SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8118 ( .A1(n6318), .A2(n7448), .ZN(n6319) );
  INV_X1 U8119 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U8120 ( .A1(n6588), .A2(n6596), .ZN(n6321) );
  NAND2_X1 U8121 ( .A1(n6325), .A2(n7383), .ZN(n6593) );
  NAND2_X1 U8122 ( .A1(n6858), .A2(n8303), .ZN(n6859) );
  NAND2_X1 U8123 ( .A1(n6859), .A2(n8359), .ZN(n6322) );
  NAND2_X1 U8124 ( .A1(n6322), .A2(n7067), .ZN(n6368) );
  OR2_X1 U8125 ( .A1(n6368), .A2(n8303), .ZN(n6323) );
  AND2_X1 U8126 ( .A1(n6323), .A2(n8278), .ZN(n6390) );
  OAI21_X1 U8127 ( .B1(n6324), .B2(n6862), .A(n6390), .ZN(n6329) );
  INV_X1 U8128 ( .A(n6390), .ZN(n6327) );
  INV_X1 U8129 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U8130 ( .A1(n6588), .A2(n6592), .ZN(n6326) );
  NAND2_X1 U8131 ( .A1(n6325), .A2(n7448), .ZN(n6590) );
  NAND2_X1 U8132 ( .A1(n6326), .A2(n6590), .ZN(n6387) );
  NAND2_X1 U8133 ( .A1(n6327), .A2(n6387), .ZN(n6328) );
  INV_X1 U8134 ( .A(n6387), .ZN(n6330) );
  NAND2_X1 U8135 ( .A1(n6391), .A2(n6330), .ZN(n6375) );
  NOR2_X1 U8136 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .ZN(
        n6334) );
  NOR4_X1 U8137 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6333) );
  NOR4_X1 U8138 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6332) );
  NOR4_X1 U8139 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6331) );
  NAND4_X1 U8140 ( .A1(n6334), .A2(n6333), .A3(n6332), .A4(n6331), .ZN(n6340)
         );
  NOR4_X1 U8141 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6338) );
  NOR4_X1 U8142 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6337) );
  NOR4_X1 U8143 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6336) );
  NOR4_X1 U8144 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6335) );
  NAND4_X1 U8145 ( .A1(n6338), .A2(n6337), .A3(n6336), .A4(n6335), .ZN(n6339)
         );
  OAI21_X1 U8146 ( .B1(n6340), .B2(n6339), .A(n6588), .ZN(n6379) );
  OR2_X1 U8147 ( .A1(n8278), .A2(n6369), .ZN(n6748) );
  AND3_X1 U8148 ( .A1(n6752), .A2(n6379), .A3(n6748), .ZN(n6341) );
  MUX2_X1 U8149 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n6392), .S(n9952), .Z(n6343)
         );
  INV_X1 U8150 ( .A(n6343), .ZN(n6373) );
  INV_X1 U8151 ( .A(n8394), .ZN(n6923) );
  NAND2_X1 U8152 ( .A1(n6923), .A2(n9875), .ZN(n8151) );
  NAND2_X1 U8153 ( .A1(n6833), .A2(n8152), .ZN(n7023) );
  INV_X1 U8154 ( .A(n8315), .ZN(n6346) );
  NAND2_X1 U8155 ( .A1(n7023), .A2(n6346), .ZN(n6347) );
  NAND2_X1 U8156 ( .A1(n6347), .A2(n8159), .ZN(n9863) );
  XNOR2_X1 U8157 ( .A(n8393), .B(n6033), .ZN(n9862) );
  NAND2_X1 U8158 ( .A1(n9863), .A2(n9862), .ZN(n6348) );
  INV_X1 U8159 ( .A(n8393), .ZN(n6896) );
  NAND2_X1 U8160 ( .A1(n6348), .A2(n8164), .ZN(n7123) );
  NAND2_X1 U8161 ( .A1(n7123), .A2(n8316), .ZN(n6349) );
  NAND2_X1 U8162 ( .A1(n8165), .A2(n8166), .ZN(n8172) );
  NAND2_X1 U8163 ( .A1(n6349), .A2(n8172), .ZN(n7148) );
  NAND2_X1 U8164 ( .A1(n7172), .A2(n9894), .ZN(n8171) );
  INV_X1 U8165 ( .A(n7172), .ZN(n8392) );
  NAND2_X1 U8166 ( .A1(n8392), .A2(n6942), .ZN(n8176) );
  NAND2_X1 U8167 ( .A1(n7148), .A2(n8319), .ZN(n7147) );
  AND2_X1 U8168 ( .A1(n8171), .A2(n8178), .ZN(n7277) );
  INV_X1 U8169 ( .A(n8323), .ZN(n6350) );
  AND2_X1 U8170 ( .A1(n7277), .A2(n6350), .ZN(n6351) );
  NAND2_X1 U8171 ( .A1(n7147), .A2(n6351), .ZN(n7276) );
  AND2_X1 U8172 ( .A1(n7307), .A2(n8182), .ZN(n8188) );
  INV_X1 U8173 ( .A(n8178), .ZN(n6352) );
  OR2_X1 U8174 ( .A1(n6352), .A2(n8318), .ZN(n7278) );
  OR2_X1 U8175 ( .A1(n8323), .A2(n7278), .ZN(n7275) );
  AND2_X1 U8176 ( .A1(n8188), .A2(n7275), .ZN(n6353) );
  NAND2_X1 U8177 ( .A1(n7276), .A2(n6353), .ZN(n7353) );
  INV_X1 U8178 ( .A(n8322), .ZN(n7355) );
  AND2_X1 U8179 ( .A1(n8190), .A2(n7355), .ZN(n6354) );
  NAND2_X1 U8180 ( .A1(n7353), .A2(n6354), .ZN(n7354) );
  OR2_X1 U8181 ( .A1(n7411), .A2(n8197), .ZN(n6355) );
  AND2_X1 U8182 ( .A1(n6355), .A2(n8183), .ZN(n8187) );
  NAND2_X1 U8183 ( .A1(n7354), .A2(n8187), .ZN(n6356) );
  NAND2_X1 U8184 ( .A1(n7411), .A2(n8197), .ZN(n8191) );
  NAND2_X1 U8185 ( .A1(n6356), .A2(n8191), .ZN(n7210) );
  OR2_X1 U8186 ( .A1(n9920), .A2(n7516), .ZN(n8207) );
  NAND2_X1 U8187 ( .A1(n9920), .A2(n7516), .ZN(n8206) );
  INV_X1 U8188 ( .A(n8209), .ZN(n8330) );
  INV_X1 U8189 ( .A(n8386), .ZN(n8210) );
  OR2_X1 U8190 ( .A1(n9930), .A2(n8210), .ZN(n8212) );
  NAND2_X1 U8191 ( .A1(n7632), .A2(n7999), .ZN(n8214) );
  NAND2_X1 U8192 ( .A1(n7443), .A2(n8214), .ZN(n6357) );
  OR2_X1 U8193 ( .A1(n7632), .A2(n7999), .ZN(n8215) );
  NAND2_X1 U8194 ( .A1(n6357), .A2(n8215), .ZN(n7523) );
  INV_X1 U8195 ( .A(n8384), .ZN(n7939) );
  NAND2_X1 U8196 ( .A1(n7990), .A2(n7939), .ZN(n8218) );
  NAND2_X1 U8197 ( .A1(n7523), .A2(n8218), .ZN(n6358) );
  OR2_X1 U8198 ( .A1(n7990), .A2(n7939), .ZN(n8219) );
  INV_X1 U8199 ( .A(n8383), .ZN(n8224) );
  NAND2_X1 U8200 ( .A1(n8225), .A2(n8224), .ZN(n6359) );
  NAND2_X1 U8201 ( .A1(n7545), .A2(n6359), .ZN(n6361) );
  OR2_X1 U8202 ( .A1(n8225), .A2(n8224), .ZN(n6360) );
  NAND2_X1 U8203 ( .A1(n6361), .A2(n6360), .ZN(n7575) );
  NAND2_X1 U8204 ( .A1(n7575), .A2(n8230), .ZN(n6362) );
  NAND2_X1 U8205 ( .A1(n8668), .A2(n8074), .ZN(n8238) );
  NAND2_X1 U8206 ( .A1(n8593), .A2(n8238), .ZN(n8602) );
  OR2_X1 U8207 ( .A1(n8313), .A2(n8593), .ZN(n8573) );
  AND2_X1 U8208 ( .A1(n8245), .A2(n8575), .ZN(n8240) );
  AND2_X1 U8209 ( .A1(n8573), .A2(n8240), .ZN(n6363) );
  NAND2_X1 U8210 ( .A1(n6364), .A2(n8244), .ZN(n8561) );
  INV_X1 U8211 ( .A(n8561), .ZN(n6365) );
  NAND2_X1 U8212 ( .A1(n6365), .A2(n8249), .ZN(n6366) );
  NAND2_X1 U8213 ( .A1(n6366), .A2(n8246), .ZN(n8550) );
  NAND2_X1 U8214 ( .A1(n8702), .A2(n8541), .ZN(n8309) );
  NAND2_X1 U8215 ( .A1(n8546), .A2(n8532), .ZN(n8525) );
  AND2_X1 U8216 ( .A1(n8309), .A2(n8525), .ZN(n8259) );
  NAND2_X1 U8217 ( .A1(n8696), .A2(n8531), .ZN(n8266) );
  NOR2_X1 U8218 ( .A1(n8512), .A2(n7979), .ZN(n8265) );
  NAND2_X1 U8219 ( .A1(n8512), .A2(n7979), .ZN(n8147) );
  OR2_X1 U8220 ( .A1(n8685), .A2(n8508), .ZN(n8270) );
  XNOR2_X1 U8221 ( .A(n6416), .B(n8308), .ZN(n6400) );
  INV_X1 U8222 ( .A(n6368), .ZN(n6370) );
  INV_X1 U8223 ( .A(n6369), .ZN(n6860) );
  OAI22_X1 U8224 ( .A1(n6400), .A2(n8673), .B1(n4437), .B2(n8672), .ZN(n6371)
         );
  INV_X1 U8225 ( .A(n6371), .ZN(n6372) );
  NAND2_X1 U8226 ( .A1(n6373), .A2(n6372), .ZN(P2_U3487) );
  INV_X1 U8227 ( .A(n6379), .ZN(n6374) );
  OR2_X1 U8228 ( .A1(n6375), .A2(n6374), .ZN(n6745) );
  INV_X1 U8229 ( .A(n6752), .ZN(n6376) );
  OR3_X1 U8230 ( .A1(n6858), .A2(n6377), .A3(n8303), .ZN(n6763) );
  NAND2_X1 U8231 ( .A1(n6756), .A2(n6763), .ZN(n6378) );
  NAND2_X1 U8232 ( .A1(n6762), .A2(n6378), .ZN(n6382) );
  AND3_X1 U8233 ( .A1(n6862), .A2(n6387), .A3(n6379), .ZN(n6753) );
  NAND2_X1 U8234 ( .A1(n6753), .A2(n6752), .ZN(n6764) );
  NAND3_X1 U8235 ( .A1(n9913), .A2(n6763), .A3(n8278), .ZN(n6760) );
  INV_X1 U8236 ( .A(n6380), .ZN(n6393) );
  AND2_X1 U8237 ( .A1(n6760), .A2(n7441), .ZN(n6743) );
  MUX2_X1 U8238 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n6392), .S(n9932), .Z(n6383)
         );
  INV_X1 U8239 ( .A(n6383), .ZN(n6386) );
  INV_X1 U8240 ( .A(n9921), .ZN(n9926) );
  OAI22_X1 U8241 ( .A1(n6400), .A2(n8738), .B1(n4437), .B2(n8736), .ZN(n6384)
         );
  INV_X1 U8242 ( .A(n6384), .ZN(n6385) );
  NAND2_X1 U8243 ( .A1(n6386), .A2(n6385), .ZN(P2_U3455) );
  NAND2_X1 U8244 ( .A1(n6390), .A2(n6387), .ZN(n6388) );
  NAND2_X1 U8245 ( .A1(n6392), .A2(n8608), .ZN(n6403) );
  AND2_X1 U8246 ( .A1(n6393), .A2(n6858), .ZN(n7024) );
  INV_X1 U8247 ( .A(n7024), .ZN(n6394) );
  NAND2_X1 U8248 ( .A1(n7364), .A2(n6394), .ZN(n6395) );
  AOI22_X1 U8249 ( .A1(n8286), .A2(n9864), .B1(n9865), .B2(n8028), .ZN(n6398)
         );
  INV_X1 U8250 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U8251 ( .A1(n6403), .A2(n6402), .ZN(P2_U3205) );
  NOR2_X1 U8252 ( .A1(n8286), .A2(n8498), .ZN(n6404) );
  OAI22_X1 U8253 ( .A1(n6405), .A2(n6404), .B1(n4438), .B2(n4437), .ZN(n6415)
         );
  INV_X1 U8254 ( .A(SI_28_), .ZN(n6408) );
  NAND2_X1 U8255 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  INV_X1 U8256 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8752) );
  INV_X1 U8257 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9393) );
  MUX2_X1 U8258 ( .A(n8752), .B(n9393), .S(n7725), .Z(n7721) );
  NAND2_X1 U8259 ( .A1(n8750), .A2(n6095), .ZN(n6413) );
  OR2_X1 U8260 ( .A1(n8291), .A2(n8752), .ZN(n6412) );
  NAND2_X1 U8261 ( .A1(n6414), .A2(n8030), .ZN(n8284) );
  XNOR2_X1 U8262 ( .A(n6415), .B(n8277), .ZN(n6429) );
  NAND2_X1 U8263 ( .A1(n6416), .A2(n8308), .ZN(n6418) );
  OR2_X1 U8264 ( .A1(n8286), .A2(n4438), .ZN(n6417) );
  XNOR2_X2 U8265 ( .A(n8351), .B(n8277), .ZN(n6430) );
  INV_X1 U8266 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U8267 ( .A1(n6419), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U8268 ( .A1(n6420), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6421) );
  OAI211_X1 U8269 ( .C1(n6199), .C2(n6423), .A(n6422), .B(n6421), .ZN(n6424)
         );
  INV_X1 U8270 ( .A(n6424), .ZN(n6425) );
  NAND2_X1 U8271 ( .A1(n8300), .A2(n6425), .ZN(n8379) );
  AND2_X1 U8272 ( .A1(n5989), .A2(P2_B_REG_SCAN_IN), .ZN(n6426) );
  NOR2_X1 U8273 ( .A1(n8607), .A2(n6426), .ZN(n8488) );
  AOI22_X1 U8274 ( .A1(n8498), .A2(n9858), .B1(n8379), .B2(n8488), .ZN(n6427)
         );
  OAI21_X1 U8275 ( .B1(n6430), .B2(n7364), .A(n6427), .ZN(n6428) );
  INV_X1 U8276 ( .A(n6414), .ZN(n6437) );
  NOR2_X1 U8277 ( .A1(n6437), .A2(n8736), .ZN(n6434) );
  NAND2_X1 U8278 ( .A1(n6436), .A2(n9952), .ZN(n6440) );
  NOR2_X1 U8279 ( .A1(n6437), .A2(n8672), .ZN(n6438) );
  NAND2_X1 U8280 ( .A1(n6440), .A2(n6439), .ZN(P2_U3488) );
  NAND2_X1 U8281 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  NAND2_X1 U8282 ( .A1(n6444), .A2(n6443), .ZN(n6446) );
  NAND2_X1 U8283 ( .A1(n9157), .A2(n8985), .ZN(n6445) );
  NAND2_X1 U8284 ( .A1(n6446), .A2(n6445), .ZN(n6450) );
  NAND2_X1 U8285 ( .A1(n8750), .A2(n5318), .ZN(n6448) );
  OR2_X1 U8286 ( .A1(n7751), .A2(n9393), .ZN(n6447) );
  INV_X1 U8287 ( .A(n8900), .ZN(n6449) );
  NAND2_X1 U8288 ( .A1(n6465), .A2(n6449), .ZN(n7818) );
  INV_X1 U8289 ( .A(n7888), .ZN(n7753) );
  NAND2_X1 U8290 ( .A1(n7753), .A2(n7146), .ZN(n9680) );
  NAND2_X1 U8291 ( .A1(n7903), .A2(n9773), .ZN(n6468) );
  INV_X1 U8292 ( .A(n7795), .ZN(n6451) );
  NOR2_X1 U8293 ( .A1(n6452), .A2(n6451), .ZN(n6454) );
  XNOR2_X1 U8294 ( .A(n6454), .B(n6453), .ZN(n6464) );
  NAND2_X1 U8295 ( .A1(n8985), .A2(n9651), .ZN(n6462) );
  NAND2_X1 U8296 ( .A1(n4966), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8297 ( .A1(n4951), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U8298 ( .A1(n7733), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6455) );
  NAND3_X1 U8299 ( .A1(n6457), .A2(n6456), .A3(n6455), .ZN(n8899) );
  INV_X1 U8300 ( .A(P1_B_REG_SCAN_IN), .ZN(n6459) );
  NOR2_X1 U8301 ( .A1(n9474), .A2(n6459), .ZN(n6460) );
  NOR2_X1 U8302 ( .A1(n9616), .A2(n6460), .ZN(n8971) );
  NAND2_X1 U8303 ( .A1(n8899), .A2(n8971), .ZN(n6461) );
  XOR2_X1 U8304 ( .A(n8967), .B(n8968), .Z(n7908) );
  AOI22_X1 U8305 ( .A1(n7908), .A2(n9666), .B1(n9734), .B2(n6465), .ZN(n6466)
         );
  NAND2_X1 U8306 ( .A1(n6468), .A2(n6467), .ZN(n6488) );
  NOR2_X1 U8307 ( .A1(n6470), .A2(n6469), .ZN(n6472) );
  NAND2_X1 U8308 ( .A1(n6488), .A2(n9777), .ZN(n6476) );
  NAND2_X1 U8309 ( .A1(n6476), .A2(n6475), .ZN(P1_U3519) );
  AOI21_X1 U8310 ( .B1(n8875), .B2(n6478), .A(n6477), .ZN(n6479) );
  NAND2_X1 U8311 ( .A1(n9164), .A2(n8894), .ZN(n6484) );
  AOI22_X1 U8312 ( .A1(n8889), .A2(n8991), .B1(n8887), .B2(n8985), .ZN(n6482)
         );
  AOI22_X1 U8313 ( .A1(n8878), .A2(n9020), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6481) );
  AND2_X1 U8314 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  NAND3_X1 U8315 ( .A1(n6485), .A2(n6484), .A3(n6483), .ZN(P1_U3214) );
  NAND2_X1 U8316 ( .A1(n6488), .A2(n9803), .ZN(n6491) );
  INV_X1 U8317 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6489) );
  OR2_X1 U8318 ( .A1(n9803), .A2(n6489), .ZN(n6490) );
  NAND2_X1 U8319 ( .A1(n6491), .A2(n6490), .ZN(P1_U3551) );
  OR2_X2 U8320 ( .A1(n6492), .A2(n5730), .ZN(n8913) );
  INV_X1 U8321 ( .A(n6493), .ZN(n6497) );
  NAND3_X1 U8322 ( .A1(n6517), .A2(n6495), .A3(n6494), .ZN(n6496) );
  AOI21_X1 U8323 ( .B1(n6497), .B2(n6496), .A(n9844), .ZN(n6513) );
  INV_X1 U8324 ( .A(n6498), .ZN(n6500) );
  NAND3_X1 U8325 ( .A1(n6520), .A2(n6500), .A3(n6499), .ZN(n6501) );
  AOI21_X1 U8326 ( .B1(n6502), .B2(n6501), .A(n8485), .ZN(n6512) );
  INV_X1 U8327 ( .A(n6503), .ZN(n6505) );
  NAND3_X1 U8328 ( .A1(n6524), .A2(n6505), .A3(n6504), .ZN(n6506) );
  AOI21_X1 U8329 ( .B1(n6507), .B2(n6506), .A(n9822), .ZN(n6511) );
  INV_X1 U8330 ( .A(n9839), .ZN(n8473) );
  NAND2_X1 U8331 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n7917) );
  INV_X1 U8332 ( .A(n7917), .ZN(n6508) );
  AOI21_X1 U8333 ( .B1(n9841), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6508), .ZN(
        n6509) );
  OAI21_X1 U8334 ( .B1(n8473), .B2(n6557), .A(n6509), .ZN(n6510) );
  OR4_X1 U8335 ( .A1(n6513), .A2(n6512), .A3(n6511), .A4(n6510), .ZN(P2_U3190)
         );
  OR3_X1 U8336 ( .A1(n6777), .A2(n6515), .A3(n6514), .ZN(n6516) );
  AOI21_X1 U8337 ( .B1(n6517), .B2(n6516), .A(n9844), .ZN(n6529) );
  NAND2_X1 U8338 ( .A1(n6518), .A2(n6074), .ZN(n6519) );
  AOI21_X1 U8339 ( .B1(n6520), .B2(n6519), .A(n8485), .ZN(n6528) );
  NAND2_X1 U8340 ( .A1(n6522), .A2(n6521), .ZN(n6523) );
  AOI21_X1 U8341 ( .B1(n6524), .B2(n6523), .A(n9822), .ZN(n6527) );
  NAND2_X1 U8342 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7139) );
  NAND2_X1 U8343 ( .A1(n9841), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6525) );
  OAI211_X1 U8344 ( .C1(n8473), .C2(n6552), .A(n7139), .B(n6525), .ZN(n6526)
         );
  OR4_X1 U8345 ( .A1(n6529), .A2(n6528), .A3(n6527), .A4(n6526), .ZN(P2_U3189)
         );
  NAND2_X1 U8346 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9239), .ZN(n9348) );
  OAI21_X1 U8347 ( .B1(n6530), .B2(P2_STATE_REG_SCAN_IN), .A(n9348), .ZN(n6531) );
  INV_X1 U8348 ( .A(n6531), .ZN(P2_U3295) );
  AND2_X1 U8349 ( .A1(n7746), .A2(P2_U3151), .ZN(n6585) );
  INV_X2 U8350 ( .A(n6585), .ZN(n8751) );
  NOR2_X1 U8351 ( .A1(n7746), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8748) );
  OAI222_X1 U8352 ( .A1(n8751), .A2(n4911), .B1(n7936), .B2(n6536), .C1(
        P2_U3151), .C2(n9818), .ZN(P2_U3294) );
  OAI222_X1 U8353 ( .A1(n4269), .A2(P2_U3151), .B1(n7936), .B2(n6535), .C1(
        n8751), .C2(n6021), .ZN(P2_U3293) );
  AND2_X1 U8354 ( .A1(n7725), .A2(P1_U3086), .ZN(n7294) );
  NOR2_X1 U8355 ( .A1(n7725), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9386) );
  OAI222_X1 U8356 ( .A1(n9435), .A2(P1_U3086), .B1(n9395), .B2(n6547), .C1(
        n6533), .C2(n9392), .ZN(P1_U3352) );
  INV_X2 U8357 ( .A(n7294), .ZN(n9395) );
  OAI222_X1 U8358 ( .A1(n9471), .A2(P1_U3086), .B1(n9395), .B2(n6535), .C1(
        n6534), .C2(n9392), .ZN(P1_U3353) );
  OAI222_X1 U8359 ( .A1(n6619), .A2(P1_U3086), .B1(n9395), .B2(n6536), .C1(
        n4909), .C2(n9392), .ZN(P1_U3354) );
  OAI222_X1 U8360 ( .A1(n9496), .A2(P1_U3086), .B1(n9395), .B2(n6549), .C1(
        n6537), .C2(n9392), .ZN(P1_U3351) );
  OAI222_X1 U8361 ( .A1(n8751), .A2(n6539), .B1(n7936), .B2(n6541), .C1(
        P2_U3151), .C2(n6538), .ZN(P2_U3290) );
  OAI222_X1 U8362 ( .A1(n9511), .A2(P1_U3086), .B1(n9395), .B2(n6541), .C1(
        n6540), .C2(n9392), .ZN(P1_U3350) );
  INV_X1 U8363 ( .A(n6633), .ZN(n9526) );
  OAI222_X1 U8364 ( .A1(n9526), .A2(P1_U3086), .B1(n9395), .B2(n6544), .C1(
        n6542), .C2(n9392), .ZN(P1_U3349) );
  OAI222_X1 U8365 ( .A1(n8751), .A2(n6545), .B1(n7936), .B2(n6544), .C1(
        P2_U3151), .C2(n6543), .ZN(P2_U3289) );
  OAI222_X1 U8366 ( .A1(n8751), .A2(n6548), .B1(n7936), .B2(n6547), .C1(
        P2_U3151), .C2(n6546), .ZN(P2_U3292) );
  OAI222_X1 U8367 ( .A1(n8751), .A2(n6550), .B1(n7936), .B2(n6549), .C1(
        P2_U3151), .C2(n9838), .ZN(P2_U3291) );
  INV_X1 U8368 ( .A(n6635), .ZN(n9420) );
  OAI222_X1 U8369 ( .A1(n9392), .A2(n6551), .B1(n9395), .B2(n6553), .C1(n9420), 
        .C2(P1_U3086), .ZN(P1_U3348) );
  OAI222_X1 U8370 ( .A1(n8751), .A2(n6554), .B1(n7936), .B2(n6553), .C1(
        P2_U3151), .C2(n6552), .ZN(P2_U3288) );
  INV_X1 U8371 ( .A(n6637), .ZN(n9450) );
  INV_X1 U8372 ( .A(n6555), .ZN(n6558) );
  OAI222_X1 U8373 ( .A1(n9450), .A2(P1_U3086), .B1(n9395), .B2(n6558), .C1(
        n6556), .C2(n9392), .ZN(P1_U3347) );
  OAI222_X1 U8374 ( .A1(n8751), .A2(n6559), .B1(n7936), .B2(n6558), .C1(
        P2_U3151), .C2(n6557), .ZN(P2_U3287) );
  AOI21_X1 U8375 ( .B1(n6561), .B2(n6562), .A(n6560), .ZN(n6572) );
  INV_X1 U8376 ( .A(n6572), .ZN(n6563) );
  OR2_X1 U8377 ( .A1(n6562), .A2(P1_U3086), .ZN(n7901) );
  NAND2_X1 U8378 ( .A1(n7896), .A2(n7901), .ZN(n6573) );
  AND2_X1 U8379 ( .A1(n6563), .A2(n6573), .ZN(n9486) );
  NOR2_X1 U8380 ( .A1(n9486), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8381 ( .A1(n7474), .A2(P1_U3973), .ZN(n6564) );
  OAI21_X1 U8382 ( .B1(n5127), .B2(P1_U3973), .A(n6564), .ZN(P1_U3566) );
  NAND2_X1 U8383 ( .A1(n6911), .A2(P1_U3973), .ZN(n6565) );
  OAI21_X1 U8384 ( .B1(P1_U3973), .B2(n6021), .A(n6565), .ZN(P1_U3556) );
  INV_X1 U8385 ( .A(n6566), .ZN(n6570) );
  OAI222_X1 U8386 ( .A1(n7936), .A2(n6570), .B1(n7113), .B2(P2_U3151), .C1(
        n6567), .C2(n8751), .ZN(P2_U3286) );
  INV_X1 U8387 ( .A(n6568), .ZN(n6582) );
  AOI22_X1 U8388 ( .A1(n9406), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9386), .ZN(n6569) );
  OAI21_X1 U8389 ( .B1(n6582), .B2(n9395), .A(n6569), .ZN(P1_U3345) );
  INV_X1 U8390 ( .A(n6846), .ZN(n6645) );
  OAI222_X1 U8391 ( .A1(n9392), .A2(n6571), .B1(n9395), .B2(n6570), .C1(
        P1_U3086), .C2(n6645), .ZN(P1_U3346) );
  INV_X1 U8392 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U8393 ( .A1(n6573), .A2(n6572), .ZN(n6641) );
  INV_X1 U8394 ( .A(n6641), .ZN(n6577) );
  INV_X1 U8395 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6808) );
  OAI21_X1 U8396 ( .B1(n9474), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9473), .ZN(
        n9479) );
  AOI21_X1 U8397 ( .B1(n9474), .B2(n6574), .A(n9479), .ZN(n6575) );
  XNOR2_X1 U8398 ( .A(n6575), .B(n9480), .ZN(n6576) );
  AOI22_X1 U8399 ( .A1(n6577), .A2(n6576), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6578) );
  OAI21_X1 U8400 ( .B1(n9613), .B2(n6579), .A(n6578), .ZN(P1_U3243) );
  OAI222_X1 U8401 ( .A1(n7936), .A2(n6582), .B1(n6581), .B2(P2_U3151), .C1(
        n6580), .C2(n8751), .ZN(P2_U3285) );
  INV_X1 U8402 ( .A(n6583), .ZN(n6587) );
  AOI22_X1 U8403 ( .A1(n9531), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9386), .ZN(n6584) );
  OAI21_X1 U8404 ( .B1(n6587), .B2(n9395), .A(n6584), .ZN(P1_U3344) );
  AOI22_X1 U8405 ( .A1(n7509), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6585), .ZN(n6586) );
  OAI21_X1 U8406 ( .B1(n6587), .B2(n7936), .A(n6586), .ZN(P2_U3284) );
  INV_X1 U8407 ( .A(n6588), .ZN(n6589) );
  INV_X1 U8408 ( .A(n6590), .ZN(n6591) );
  AOI22_X1 U8409 ( .A1(n6597), .A2(n6592), .B1(n6595), .B2(n6591), .ZN(
        P2_U3377) );
  INV_X1 U8410 ( .A(n6593), .ZN(n6594) );
  AOI22_X1 U8411 ( .A1(n6597), .A2(n6596), .B1(n6595), .B2(n6594), .ZN(
        P2_U3376) );
  AND2_X1 U8412 ( .A1(n6597), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8413 ( .A1(n6597), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8414 ( .A1(n6597), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8415 ( .A1(n6597), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8416 ( .A1(n6597), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8417 ( .A1(n6597), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8418 ( .A1(n6597), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8419 ( .A1(n6597), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8420 ( .A1(n6597), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8421 ( .A1(n6597), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8422 ( .A1(n6597), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8423 ( .A1(n6597), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8424 ( .A1(n6597), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8425 ( .A1(n6597), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8426 ( .A1(n6597), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8427 ( .A1(n6597), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8428 ( .A1(n6597), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8429 ( .A1(n6597), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8430 ( .A1(n6597), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8431 ( .A1(n6597), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8432 ( .A1(n6597), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8433 ( .A1(n6597), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8434 ( .A1(n6597), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8435 ( .A1(n6597), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8436 ( .A1(n6597), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8437 ( .A1(n6597), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8438 ( .A1(n6597), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8439 ( .A1(n6597), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  INV_X1 U8440 ( .A(n6597), .ZN(n6598) );
  INV_X1 U8441 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9287) );
  NOR2_X1 U8442 ( .A1(n6598), .A2(n9287), .ZN(P2_U3244) );
  INV_X1 U8443 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9254) );
  NOR2_X1 U8444 ( .A1(n6598), .A2(n9254), .ZN(P2_U3242) );
  INV_X1 U8445 ( .A(n6599), .ZN(n6606) );
  OAI222_X1 U8446 ( .A1(n7936), .A2(n6606), .B1(n8751), .B2(n5127), .C1(
        P2_U3151), .C2(n6600), .ZN(P2_U3283) );
  INV_X1 U8447 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6604) );
  AND2_X1 U8448 ( .A1(n5740), .A2(n6671), .ZN(n7832) );
  NOR2_X1 U8449 ( .A1(n6910), .A2(n7832), .ZN(n7766) );
  INV_X1 U8450 ( .A(n7766), .ZN(n6601) );
  OAI21_X1 U8451 ( .B1(n9655), .B2(n9773), .A(n6601), .ZN(n6602) );
  NAND2_X1 U8452 ( .A1(n5732), .A2(n9652), .ZN(n6803) );
  OAI211_X1 U8453 ( .C1(n6802), .C2(n6671), .A(n6602), .B(n6803), .ZN(n9223)
         );
  NAND2_X1 U8454 ( .A1(n9223), .A2(n9777), .ZN(n6603) );
  OAI21_X1 U8455 ( .B1(n9777), .B2(n6604), .A(n6603), .ZN(P1_U3453) );
  INV_X1 U8456 ( .A(n8934), .ZN(n6854) );
  OAI222_X1 U8457 ( .A1(P1_U3086), .A2(n6854), .B1(n9395), .B2(n6606), .C1(
        n6605), .C2(n9392), .ZN(P1_U3343) );
  INV_X1 U8458 ( .A(n6607), .ZN(n6650) );
  AOI22_X1 U8459 ( .A1(n9556), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9386), .ZN(n6608) );
  OAI21_X1 U8460 ( .B1(n6650), .B2(n9395), .A(n6608), .ZN(P1_U3342) );
  INV_X1 U8461 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6609) );
  AOI22_X1 U8462 ( .A1(n6846), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6609), .B2(
        n6645), .ZN(n6617) );
  INV_X1 U8463 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9309) );
  MUX2_X1 U8464 ( .A(n9309), .B(P1_REG2_REG_1__SCAN_IN), .S(n6619), .Z(n8915)
         );
  NOR2_X1 U8465 ( .A1(n9480), .A2(n6808), .ZN(n9477) );
  NAND2_X1 U8466 ( .A1(n8915), .A2(n9477), .ZN(n8914) );
  NAND2_X1 U8467 ( .A1(n4916), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U8468 ( .A1(n8914), .A2(n6610), .ZN(n9464) );
  INV_X1 U8469 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9280) );
  XNOR2_X1 U8470 ( .A(n6618), .B(n9280), .ZN(n9465) );
  NAND2_X1 U8471 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6624), .ZN(n6611) );
  OAI21_X1 U8472 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6624), .A(n6611), .ZN(
        n9427) );
  NAND2_X1 U8473 ( .A1(n6627), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6612) );
  OAI21_X1 U8474 ( .B1(n6627), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6612), .ZN(
        n9488) );
  NOR2_X1 U8475 ( .A1(n4294), .A2(n9488), .ZN(n9487) );
  AOI21_X1 U8476 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6627), .A(n9487), .ZN(
        n9502) );
  NAND2_X1 U8477 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6630), .ZN(n6613) );
  OAI21_X1 U8478 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6630), .A(n6613), .ZN(
        n9503) );
  NAND2_X1 U8479 ( .A1(n6633), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6614) );
  OAI21_X1 U8480 ( .B1(n6633), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6614), .ZN(
        n9518) );
  INV_X1 U8481 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7043) );
  AOI22_X1 U8482 ( .A1(n6635), .A2(n7043), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9420), .ZN(n9411) );
  NOR2_X1 U8483 ( .A1(n9412), .A2(n9411), .ZN(n9410) );
  NAND2_X1 U8484 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6637), .ZN(n6615) );
  OAI21_X1 U8485 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6637), .A(n6615), .ZN(
        n9442) );
  OAI21_X1 U8486 ( .B1(n6617), .B2(n6616), .A(n6840), .ZN(n6647) );
  OR2_X1 U8487 ( .A1(n5417), .A2(n9474), .ZN(n9476) );
  INV_X1 U8488 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9792) );
  AOI22_X1 U8489 ( .A1(n6846), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n9792), .B2(
        n6645), .ZN(n6639) );
  INV_X1 U8490 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9778) );
  MUX2_X1 U8491 ( .A(n9778), .B(P1_REG1_REG_1__SCAN_IN), .S(n6619), .Z(n8918)
         );
  NAND2_X1 U8492 ( .A1(n8918), .A2(n8917), .ZN(n8916) );
  NAND2_X1 U8493 ( .A1(n4916), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U8494 ( .A1(n8916), .A2(n6620), .ZN(n9467) );
  NAND2_X1 U8495 ( .A1(n9468), .A2(n9467), .ZN(n9466) );
  AND2_X1 U8496 ( .A1(n9466), .A2(n6621), .ZN(n9431) );
  OR2_X1 U8497 ( .A1(n6624), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U8498 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6624), .ZN(n6622) );
  NAND2_X1 U8499 ( .A1(n6623), .A2(n6622), .ZN(n9430) );
  NOR2_X1 U8500 ( .A1(n9431), .A2(n9430), .ZN(n9429) );
  OR2_X1 U8501 ( .A1(n6627), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U8502 ( .A1(n6627), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U8503 ( .A1(n6626), .A2(n6625), .ZN(n9492) );
  NOR2_X1 U8504 ( .A1(n9491), .A2(n9492), .ZN(n9490) );
  AOI21_X1 U8505 ( .B1(n6627), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9490), .ZN(
        n9506) );
  OR2_X1 U8506 ( .A1(n6630), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U8507 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6630), .ZN(n6628) );
  NAND2_X1 U8508 ( .A1(n6629), .A2(n6628), .ZN(n9507) );
  OR2_X1 U8509 ( .A1(n6633), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U8510 ( .A1(n6633), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U8511 ( .A1(n6632), .A2(n6631), .ZN(n9522) );
  INV_X1 U8512 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6634) );
  MUX2_X1 U8513 ( .A(n6634), .B(P1_REG1_REG_7__SCAN_IN), .S(n6635), .Z(n9416)
         );
  NOR2_X1 U8514 ( .A1(n9415), .A2(n9416), .ZN(n9414) );
  AOI21_X1 U8515 ( .B1(n6635), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9414), .ZN(
        n9446) );
  INV_X1 U8516 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6636) );
  MUX2_X1 U8517 ( .A(n6636), .B(P1_REG1_REG_8__SCAN_IN), .S(n6637), .Z(n9445)
         );
  NOR2_X1 U8518 ( .A1(n9446), .A2(n9445), .ZN(n9444) );
  OAI21_X1 U8519 ( .B1(n6639), .B2(n6638), .A(n6845), .ZN(n6642) );
  INV_X1 U8520 ( .A(n9474), .ZN(n6640) );
  NAND2_X1 U8521 ( .A1(n6642), .A2(n9591), .ZN(n6644) );
  AND2_X1 U8522 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7268) );
  AOI21_X1 U8523 ( .B1(n9486), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7268), .ZN(
        n6643) );
  OAI211_X1 U8524 ( .C1(n9543), .C2(n6645), .A(n6644), .B(n6643), .ZN(n6646)
         );
  AOI21_X1 U8525 ( .B1(n6647), .B2(n9598), .A(n6646), .ZN(n6648) );
  INV_X1 U8526 ( .A(n6648), .ZN(P1_U3252) );
  INV_X1 U8527 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9285) );
  OAI222_X1 U8528 ( .A1(n8751), .A2(n9285), .B1(n7936), .B2(n6650), .C1(
        P2_U3151), .C2(n6649), .ZN(P2_U3282) );
  INV_X1 U8529 ( .A(n6651), .ZN(n6654) );
  AOI22_X1 U8530 ( .A1(n9568), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9386), .ZN(n6652) );
  OAI21_X1 U8531 ( .B1(n6654), .B2(n9395), .A(n6652), .ZN(P1_U3341) );
  OAI222_X1 U8532 ( .A1(n8751), .A2(n6655), .B1(n7936), .B2(n6654), .C1(
        P2_U3151), .C2(n6653), .ZN(P2_U3281) );
  XOR2_X1 U8533 ( .A(n6657), .B(n6656), .Z(n6668) );
  INV_X1 U8534 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U8535 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n6988) );
  OAI21_X1 U8536 ( .B1(n9831), .B2(n6658), .A(n6988), .ZN(n6665) );
  INV_X1 U8537 ( .A(n9835), .ZN(n6659) );
  AOI21_X1 U8538 ( .B1(n9869), .B2(n6660), .A(n6659), .ZN(n6663) );
  XNOR2_X1 U8539 ( .A(n6661), .B(n6026), .ZN(n6662) );
  OAI22_X1 U8540 ( .A1(n6663), .A2(n9822), .B1(n8485), .B2(n6662), .ZN(n6664)
         );
  AOI211_X1 U8541 ( .C1(n6666), .C2(n9839), .A(n6665), .B(n6664), .ZN(n6667)
         );
  OAI21_X1 U8542 ( .B1(n9844), .B2(n6668), .A(n6667), .ZN(P2_U3185) );
  NOR2_X1 U8543 ( .A1(n8889), .A2(P1_U3086), .ZN(n6732) );
  INV_X1 U8544 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6674) );
  XNOR2_X1 U8545 ( .A(n6670), .B(n6669), .ZN(n9475) );
  OAI22_X1 U8546 ( .A1(n8851), .A2(n6671), .B1(n8897), .B2(n9475), .ZN(n6672)
         );
  AOI21_X1 U8547 ( .B1(n8887), .B2(n5732), .A(n6672), .ZN(n6673) );
  OAI21_X1 U8548 ( .B1(n6732), .B2(n6674), .A(n6673), .ZN(P1_U3232) );
  INV_X1 U8549 ( .A(n6675), .ZN(n6688) );
  INV_X1 U8550 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6676) );
  OAI222_X1 U8551 ( .A1(n7936), .A2(n6688), .B1(n6677), .B2(P2_U3151), .C1(
        n6676), .C2(n8751), .ZN(P2_U3280) );
  AOI21_X1 U8552 ( .B1(n6680), .B2(n6679), .A(n6678), .ZN(n6686) );
  AOI22_X1 U8553 ( .A1(n8878), .A2(n6911), .B1(n8887), .B2(n8912), .ZN(n6685)
         );
  INV_X1 U8554 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6683) );
  NAND2_X1 U8555 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9437) );
  INV_X1 U8556 ( .A(n9437), .ZN(n6682) );
  NOR2_X1 U8557 ( .A1(n8851), .A2(n9695), .ZN(n6681) );
  AOI211_X1 U8558 ( .C1(n6683), .C2(n8889), .A(n6682), .B(n6681), .ZN(n6684)
         );
  OAI211_X1 U8559 ( .C1(n6686), .C2(n8897), .A(n6685), .B(n6684), .ZN(P1_U3218) );
  INV_X1 U8560 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U8561 ( .A1(P1_U3086), .A2(n8937), .B1(n9395), .B2(n6688), .C1(
        n6687), .C2(n9392), .ZN(P1_U3340) );
  XNOR2_X1 U8562 ( .A(n6690), .B(n6689), .ZN(n6704) );
  INV_X1 U8563 ( .A(n8485), .ZN(n9852) );
  OAI21_X1 U8564 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(n6698) );
  OAI21_X1 U8565 ( .B1(n6696), .B2(n6695), .A(n6694), .ZN(n6697) );
  AOI22_X1 U8566 ( .A1(n9852), .A2(n6698), .B1(n5642), .B2(n6697), .ZN(n6700)
         );
  NAND2_X1 U8567 ( .A1(n9841), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n6699) );
  OAI211_X1 U8568 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6018), .A(n6700), .B(n6699), .ZN(n6701) );
  AOI21_X1 U8569 ( .B1(n6702), .B2(n9839), .A(n6701), .ZN(n6703) );
  OAI21_X1 U8570 ( .B1(n9844), .B2(n6704), .A(n6703), .ZN(P2_U3184) );
  XNOR2_X1 U8571 ( .A(n6706), .B(n6705), .ZN(n6716) );
  INV_X1 U8572 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U8573 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n6940) );
  OAI21_X1 U8574 ( .B1(n9831), .B2(n9313), .A(n6940), .ZN(n6714) );
  AOI21_X1 U8575 ( .B1(n6708), .B2(n6707), .A(n4360), .ZN(n6712) );
  INV_X1 U8576 ( .A(n6783), .ZN(n6709) );
  AOI21_X1 U8577 ( .B1(n9941), .B2(n6710), .A(n6709), .ZN(n6711) );
  OAI22_X1 U8578 ( .A1(n6712), .A2(n9822), .B1(n8485), .B2(n6711), .ZN(n6713)
         );
  AOI211_X1 U8579 ( .C1(n4752), .C2(n9839), .A(n6714), .B(n6713), .ZN(n6715)
         );
  OAI21_X1 U8580 ( .B1(n6716), .B2(n9844), .A(n6715), .ZN(P2_U3187) );
  INV_X1 U8581 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6825) );
  AND3_X1 U8582 ( .A1(n6725), .A2(n6718), .A3(n6717), .ZN(n6719) );
  OAI21_X1 U8583 ( .B1(n6720), .B2(n6719), .A(n8876), .ZN(n6723) );
  OAI22_X1 U8584 ( .A1(n8867), .A2(n6820), .B1(n9689), .B2(n8851), .ZN(n6721)
         );
  AOI21_X1 U8585 ( .B1(n8878), .B2(n5732), .A(n6721), .ZN(n6722) );
  OAI211_X1 U8586 ( .C1(n6732), .C2(n6825), .A(n6723), .B(n6722), .ZN(P1_U3237) );
  INV_X1 U8587 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6731) );
  OAI22_X1 U8588 ( .A1(n8867), .A2(n7835), .B1(n9683), .B2(n8851), .ZN(n6724)
         );
  AOI21_X1 U8589 ( .B1(n8878), .B2(n5740), .A(n6724), .ZN(n6730) );
  OAI21_X1 U8590 ( .B1(n6727), .B2(n6726), .A(n6725), .ZN(n6728) );
  NAND2_X1 U8591 ( .A1(n6728), .A2(n8876), .ZN(n6729) );
  OAI211_X1 U8592 ( .C1(n6732), .C2(n6731), .A(n6730), .B(n6729), .ZN(P1_U3222) );
  INV_X1 U8593 ( .A(n6733), .ZN(n6776) );
  AOI22_X1 U8594 ( .A1(n9593), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9386), .ZN(n6734) );
  OAI21_X1 U8595 ( .B1(n6776), .B2(n9395), .A(n6734), .ZN(P1_U3338) );
  XNOR2_X1 U8596 ( .A(n6736), .B(n5772), .ZN(n6737) );
  XNOR2_X1 U8597 ( .A(n6735), .B(n6737), .ZN(n6742) );
  AOI22_X1 U8598 ( .A1(n8878), .A2(n8912), .B1(n8887), .B2(n8911), .ZN(n6741)
         );
  NAND2_X1 U8599 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9513) );
  INV_X1 U8600 ( .A(n9513), .ZN(n6739) );
  NOR2_X1 U8601 ( .A1(n8851), .A2(n9708), .ZN(n6738) );
  AOI211_X1 U8602 ( .C1(n6962), .C2(n8889), .A(n6739), .B(n6738), .ZN(n6740)
         );
  OAI211_X1 U8603 ( .C1(n6742), .C2(n8897), .A(n6741), .B(n6740), .ZN(P1_U3227) );
  INV_X1 U8604 ( .A(n6743), .ZN(n6744) );
  NAND2_X1 U8605 ( .A1(n6745), .A2(n6744), .ZN(n6751) );
  AND3_X1 U8606 ( .A1(n6748), .A2(n6747), .A3(n6746), .ZN(n6750) );
  OR2_X1 U8607 ( .A1(n6753), .A2(n6763), .ZN(n6749) );
  NAND3_X1 U8608 ( .A1(n6751), .A2(n6750), .A3(n6749), .ZN(n6755) );
  INV_X1 U8609 ( .A(n6756), .ZN(n6930) );
  NAND2_X1 U8610 ( .A1(n6752), .A2(n6930), .ZN(n8372) );
  NOR2_X1 U8611 ( .A1(n6753), .A2(n8372), .ZN(n6754) );
  AOI21_X2 U8612 ( .B1(n6755), .B2(P2_STATE_REG_SCAN_IN), .A(n6754), .ZN(n8075) );
  NOR2_X1 U8613 ( .A1(n8141), .A2(P2_U3151), .ZN(n6924) );
  NOR2_X1 U8614 ( .A1(n6764), .A2(n6756), .ZN(n6872) );
  NAND2_X1 U8615 ( .A1(n6872), .A2(n6757), .ZN(n8138) );
  NAND2_X1 U8616 ( .A1(n6762), .A2(n9931), .ZN(n6759) );
  INV_X1 U8617 ( .A(n9875), .ZN(n6767) );
  INV_X1 U8618 ( .A(n6760), .ZN(n6761) );
  NAND2_X1 U8619 ( .A1(n6762), .A2(n6761), .ZN(n6766) );
  OR2_X1 U8620 ( .A1(n6764), .A2(n6763), .ZN(n6765) );
  NAND2_X1 U8621 ( .A1(n8394), .A2(n6767), .ZN(n8149) );
  AND2_X1 U8622 ( .A1(n8151), .A2(n8149), .ZN(n9871) );
  OAI22_X1 U8623 ( .A1(n8145), .A2(n6767), .B1(n8132), .B2(n9871), .ZN(n6768)
         );
  AOI21_X1 U8624 ( .B1(n8092), .B2(n6758), .A(n6768), .ZN(n6769) );
  OAI21_X1 U8625 ( .B1(n6924), .B2(n6002), .A(n6769), .ZN(P2_U3172) );
  INV_X1 U8626 ( .A(n8955), .ZN(n6771) );
  INV_X1 U8627 ( .A(n6770), .ZN(n6773) );
  OAI222_X1 U8628 ( .A1(n6771), .A2(P1_U3086), .B1(n9395), .B2(n6773), .C1(
        n9274), .C2(n9392), .ZN(P1_U3339) );
  OAI222_X1 U8629 ( .A1(n8751), .A2(n6774), .B1(n7936), .B2(n6773), .C1(
        P2_U3151), .C2(n6772), .ZN(P2_U3279) );
  OAI222_X1 U8630 ( .A1(n7936), .A2(n6776), .B1(n8463), .B2(P2_U3151), .C1(
        n6775), .C2(n8751), .ZN(P2_U3278) );
  AOI21_X1 U8631 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(n6798) );
  INV_X1 U8632 ( .A(n6780), .ZN(n6782) );
  NAND3_X1 U8633 ( .A1(n6783), .A2(n6782), .A3(n6781), .ZN(n6784) );
  AOI21_X1 U8634 ( .B1(n6785), .B2(n6784), .A(n8485), .ZN(n6795) );
  INV_X1 U8635 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6793) );
  INV_X1 U8636 ( .A(n6786), .ZN(n6791) );
  INV_X1 U8637 ( .A(n6787), .ZN(n6789) );
  NOR3_X1 U8638 ( .A1(n4360), .A2(n6789), .A3(n6788), .ZN(n6790) );
  OAI21_X1 U8639 ( .B1(n6791), .B2(n6790), .A(n5642), .ZN(n6792) );
  NAND2_X1 U8640 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n7061) );
  OAI211_X1 U8641 ( .C1(n9831), .C2(n6793), .A(n6792), .B(n7061), .ZN(n6794)
         );
  AOI211_X1 U8642 ( .C1(n9839), .C2(n6796), .A(n6795), .B(n6794), .ZN(n6797)
         );
  OAI21_X1 U8643 ( .B1(n6798), .B2(n9844), .A(n6797), .ZN(P2_U3188) );
  INV_X1 U8644 ( .A(n6799), .ZN(n6918) );
  AOI22_X1 U8645 ( .A1(n9606), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9386), .ZN(n6800) );
  OAI21_X1 U8646 ( .B1(n6918), .B2(n9395), .A(n6800), .ZN(P1_U3337) );
  OAI21_X1 U8647 ( .B1(n7202), .B2(n7907), .A(n6908), .ZN(n6807) );
  INV_X1 U8648 ( .A(n6801), .ZN(n7897) );
  NAND2_X1 U8649 ( .A1(n7897), .A2(n6802), .ZN(n6804) );
  OAI21_X1 U8650 ( .B1(n7766), .B2(n6804), .A(n6803), .ZN(n6805) );
  AOI22_X1 U8651 ( .A1(n9113), .A2(n6805), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9656), .ZN(n6806) );
  OAI211_X1 U8652 ( .C1(n6808), .C2(n9113), .A(n6807), .B(n6806), .ZN(P1_U3293) );
  XNOR2_X1 U8653 ( .A(n7764), .B(n6809), .ZN(n6810) );
  OAI222_X1 U8654 ( .A1(n9616), .A2(n6956), .B1(n9618), .B2(n7835), .C1(n6810), 
        .C2(n9138), .ZN(n9696) );
  INV_X1 U8655 ( .A(n9696), .ZN(n6816) );
  XNOR2_X1 U8656 ( .A(n7764), .B(n6811), .ZN(n9698) );
  OAI211_X1 U8657 ( .C1(n6822), .C2(n9695), .A(n9666), .B(n9664), .ZN(n9694)
         );
  OAI22_X1 U8658 ( .A1(n8982), .A2(n9694), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9104), .ZN(n6812) );
  AOI21_X1 U8659 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n9658), .A(n6812), .ZN(
        n6813) );
  OAI21_X1 U8660 ( .B1(n9695), .B2(n9660), .A(n6813), .ZN(n6814) );
  AOI21_X1 U8661 ( .B1(n9670), .B2(n9698), .A(n6814), .ZN(n6815) );
  OAI21_X1 U8662 ( .B1(n6816), .B2(n9658), .A(n6815), .ZN(P1_U3290) );
  XNOR2_X1 U8663 ( .A(n7763), .B(n6817), .ZN(n6818) );
  OAI222_X1 U8664 ( .A1(n9616), .A2(n6820), .B1(n9618), .B2(n6819), .C1(n9138), 
        .C2(n6818), .ZN(n9690) );
  INV_X1 U8665 ( .A(n9690), .ZN(n6831) );
  XNOR2_X1 U8666 ( .A(n7763), .B(n6821), .ZN(n9692) );
  INV_X1 U8667 ( .A(n6822), .ZN(n6824) );
  AOI21_X1 U8668 ( .B1(n6906), .B2(n7834), .A(n9769), .ZN(n6823) );
  NAND2_X1 U8669 ( .A1(n6824), .A2(n6823), .ZN(n9688) );
  OAI22_X1 U8670 ( .A1(n8982), .A2(n9688), .B1(n6825), .B2(n9104), .ZN(n6826)
         );
  INV_X1 U8671 ( .A(n6826), .ZN(n6828) );
  NAND2_X1 U8672 ( .A1(n9658), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6827) );
  OAI211_X1 U8673 ( .C1(n9660), .C2(n9689), .A(n6828), .B(n6827), .ZN(n6829)
         );
  AOI21_X1 U8674 ( .B1(n9670), .B2(n9692), .A(n6829), .ZN(n6830) );
  OAI21_X1 U8675 ( .B1(n6831), .B2(n9673), .A(n6830), .ZN(P1_U3291) );
  NAND2_X1 U8676 ( .A1(n6834), .A2(n8151), .ZN(n6832) );
  NAND2_X1 U8677 ( .A1(n6833), .A2(n6832), .ZN(n7166) );
  NOR2_X1 U8678 ( .A1(n6013), .A2(n9913), .ZN(n6837) );
  XNOR2_X1 U8679 ( .A(n6345), .B(n6835), .ZN(n6836) );
  OAI222_X1 U8680 ( .A1(n8605), .A2(n6923), .B1(n8607), .B2(n6881), .C1(n9872), 
        .C2(n6836), .ZN(n7162) );
  AOI211_X1 U8681 ( .C1(n9921), .C2(n7166), .A(n6837), .B(n7162), .ZN(n9877)
         );
  NAND2_X1 U8682 ( .A1(n9950), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8683 ( .B1(n9877), .B2(n9950), .A(n6838), .ZN(P2_U3460) );
  INV_X1 U8684 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9255) );
  AOI22_X1 U8685 ( .A1(n8934), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9255), .B2(
        n6854), .ZN(n6843) );
  NAND2_X1 U8686 ( .A1(n9406), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6839) );
  OAI21_X1 U8687 ( .B1(n9406), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6839), .ZN(
        n9402) );
  OAI21_X1 U8688 ( .B1(n6846), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6840), .ZN(
        n9403) );
  NOR2_X1 U8689 ( .A1(n9402), .A2(n9403), .ZN(n9401) );
  NAND2_X1 U8690 ( .A1(n9531), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6841) );
  OAI21_X1 U8691 ( .B1(n9531), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6841), .ZN(
        n9534) );
  OAI21_X1 U8692 ( .B1(n6843), .B2(n6842), .A(n8933), .ZN(n6856) );
  INV_X1 U8693 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6844) );
  MUX2_X1 U8694 ( .A(n6844), .B(P1_REG1_REG_10__SCAN_IN), .S(n9406), .Z(n9399)
         );
  INV_X1 U8695 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6847) );
  MUX2_X1 U8696 ( .A(n6847), .B(P1_REG1_REG_11__SCAN_IN), .S(n9531), .Z(n9538)
         );
  NOR2_X1 U8697 ( .A1(n9537), .A2(n9538), .ZN(n9536) );
  INV_X1 U8698 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9796) );
  AOI22_X1 U8699 ( .A1(n8934), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9796), .B2(
        n6854), .ZN(n6848) );
  OAI21_X1 U8700 ( .B1(n6849), .B2(n6848), .A(n8924), .ZN(n6850) );
  NAND2_X1 U8701 ( .A1(n6850), .A2(n9591), .ZN(n6853) );
  INV_X1 U8702 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6851) );
  NOR2_X1 U8703 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6851), .ZN(n7403) );
  AOI21_X1 U8704 ( .B1(n9486), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7403), .ZN(
        n6852) );
  OAI211_X1 U8705 ( .C1(n9543), .C2(n6854), .A(n6853), .B(n6852), .ZN(n6855)
         );
  AOI21_X1 U8706 ( .B1(n6856), .B2(n9598), .A(n6855), .ZN(n6857) );
  INV_X1 U8707 ( .A(n6857), .ZN(P1_U3255) );
  OR2_X1 U8708 ( .A1(n6858), .A2(n8303), .ZN(n8314) );
  AND2_X1 U8709 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  OAI21_X2 U8710 ( .B1(n6862), .B2(n8314), .A(n6861), .ZN(n6869) );
  OR2_X1 U8711 ( .A1(n6869), .A2(n9875), .ZN(n6864) );
  NAND2_X1 U8712 ( .A1(n6864), .A2(n8151), .ZN(n6921) );
  XNOR2_X1 U8713 ( .A(n6865), .B(n6869), .ZN(n6866) );
  XNOR2_X1 U8714 ( .A(n6758), .B(n6866), .ZN(n6920) );
  NAND2_X1 U8715 ( .A1(n6921), .A2(n6920), .ZN(n6868) );
  NAND2_X1 U8716 ( .A1(n6866), .A2(n6929), .ZN(n6867) );
  NAND2_X1 U8717 ( .A1(n6868), .A2(n6867), .ZN(n6879) );
  XNOR2_X1 U8718 ( .A(n6880), .B(n6881), .ZN(n6878) );
  XOR2_X1 U8719 ( .A(n6879), .B(n6878), .Z(n6876) );
  NAND2_X1 U8720 ( .A1(n6872), .A2(n6871), .ZN(n8095) );
  OAI22_X1 U8721 ( .A1(n8145), .A2(n9879), .B1(n6929), .B2(n8095), .ZN(n6874)
         );
  NOR2_X1 U8722 ( .A1(n6924), .A2(n6018), .ZN(n6873) );
  AOI211_X1 U8723 ( .C1(n8092), .C2(n8393), .A(n6874), .B(n6873), .ZN(n6875)
         );
  OAI21_X1 U8724 ( .B1(n8132), .B2(n6876), .A(n6875), .ZN(P2_U3177) );
  XNOR2_X1 U8725 ( .A(n6869), .B(n9890), .ZN(n6935) );
  XNOR2_X1 U8726 ( .A(n6935), .B(n6877), .ZN(n6895) );
  NAND2_X1 U8727 ( .A1(n6879), .A2(n6878), .ZN(n6884) );
  INV_X1 U8728 ( .A(n6880), .ZN(n6882) );
  NAND2_X1 U8729 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  NAND2_X1 U8730 ( .A1(n6884), .A2(n6883), .ZN(n6991) );
  INV_X1 U8731 ( .A(n6991), .ZN(n6886) );
  XNOR2_X1 U8732 ( .A(n6869), .B(n6033), .ZN(n6887) );
  XNOR2_X1 U8733 ( .A(n6887), .B(n6896), .ZN(n6992) );
  NAND2_X1 U8734 ( .A1(n6886), .A2(n6885), .ZN(n6892) );
  INV_X1 U8735 ( .A(n6887), .ZN(n6888) );
  NAND2_X1 U8736 ( .A1(n6888), .A2(n8393), .ZN(n6889) );
  NAND2_X1 U8737 ( .A1(n6892), .A2(n6889), .ZN(n6894) );
  INV_X1 U8738 ( .A(n6895), .ZN(n6890) );
  AND2_X1 U8739 ( .A1(n6890), .A2(n6889), .ZN(n6891) );
  NAND2_X1 U8740 ( .A1(n6892), .A2(n6891), .ZN(n6938) );
  INV_X1 U8741 ( .A(n6938), .ZN(n6893) );
  AOI21_X1 U8742 ( .B1(n6895), .B2(n6894), .A(n6893), .ZN(n6902) );
  NAND2_X1 U8743 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9855) );
  INV_X1 U8744 ( .A(n9855), .ZN(n6898) );
  OAI22_X1 U8745 ( .A1(n7172), .A2(n8138), .B1(n8095), .B2(n6896), .ZN(n6897)
         );
  AOI211_X1 U8746 ( .C1(n8166), .C2(n8129), .A(n6898), .B(n6897), .ZN(n6901)
         );
  INV_X1 U8747 ( .A(n6899), .ZN(n7130) );
  NAND2_X1 U8748 ( .A1(n8141), .A2(n7130), .ZN(n6900) );
  OAI211_X1 U8749 ( .C1(n6902), .C2(n8132), .A(n6901), .B(n6900), .ZN(P2_U3170) );
  XNOR2_X1 U8750 ( .A(n6903), .B(n6904), .ZN(n9686) );
  NOR2_X1 U8751 ( .A1(n9673), .A2(n6905), .ZN(n9634) );
  AOI211_X1 U8752 ( .C1(n6908), .C2(n6907), .A(n9769), .B(n4516), .ZN(n9681)
         );
  AOI22_X1 U8753 ( .A1(n9669), .A2(n9681), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9656), .ZN(n6909) );
  OAI21_X1 U8754 ( .B1(n9683), .B2(n9660), .A(n6909), .ZN(n6916) );
  XNOR2_X1 U8755 ( .A(n6903), .B(n6910), .ZN(n6914) );
  INV_X1 U8756 ( .A(n9622), .ZN(n7084) );
  NAND2_X1 U8757 ( .A1(n9686), .A2(n7084), .ZN(n6913) );
  AOI22_X1 U8758 ( .A1(n9652), .A2(n6911), .B1(n5740), .B2(n9651), .ZN(n6912)
         );
  OAI211_X1 U8759 ( .C1(n6914), .C2(n9138), .A(n6913), .B(n6912), .ZN(n9684)
         );
  MUX2_X1 U8760 ( .A(n9684), .B(P1_REG2_REG_1__SCAN_IN), .S(n9658), .Z(n6915)
         );
  AOI211_X1 U8761 ( .C1(n9686), .C2(n9634), .A(n6916), .B(n6915), .ZN(n6917)
         );
  INV_X1 U8762 ( .A(n6917), .ZN(P1_U3292) );
  OAI222_X1 U8763 ( .A1(n8751), .A2(n6919), .B1(n8475), .B2(P2_U3151), .C1(
        n7936), .C2(n6918), .ZN(P2_U3277) );
  XOR2_X1 U8764 ( .A(n6921), .B(n6920), .Z(n6928) );
  OAI22_X1 U8765 ( .A1(n8145), .A2(n6013), .B1(n6923), .B2(n8095), .ZN(n6926)
         );
  NOR2_X1 U8766 ( .A1(n6924), .A2(n5993), .ZN(n6925) );
  AOI211_X1 U8767 ( .C1(n8092), .C2(n6922), .A(n6926), .B(n6925), .ZN(n6927)
         );
  OAI21_X1 U8768 ( .B1(n8132), .B2(n6928), .A(n6927), .ZN(P2_U3162) );
  NOR2_X1 U8769 ( .A1(n6929), .A2(n8607), .ZN(n9874) );
  NOR3_X1 U8770 ( .A1(n9871), .A2(n9931), .A3(n6930), .ZN(n6931) );
  AOI211_X1 U8771 ( .C1(n9865), .C2(P2_REG3_REG_0__SCAN_IN), .A(n9874), .B(
        n6931), .ZN(n6933) );
  AOI22_X1 U8772 ( .A1(n9870), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9864), .B2(
        n9875), .ZN(n6932) );
  OAI21_X1 U8773 ( .B1(n6933), .B2(n9870), .A(n6932), .ZN(P2_U3233) );
  NAND2_X1 U8774 ( .A1(n8474), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6934) );
  OAI21_X1 U8775 ( .B1(n8030), .B2(n8474), .A(n6934), .ZN(P2_U3520) );
  INV_X1 U8776 ( .A(n6935), .ZN(n6936) );
  NAND2_X1 U8777 ( .A1(n6936), .A2(n8165), .ZN(n6937) );
  NAND2_X1 U8778 ( .A1(n6938), .A2(n6937), .ZN(n7051) );
  INV_X2 U8779 ( .A(n6863), .ZN(n8024) );
  XNOR2_X1 U8780 ( .A(n8024), .B(n6942), .ZN(n7052) );
  XNOR2_X1 U8781 ( .A(n7052), .B(n7172), .ZN(n7050) );
  XOR2_X1 U8782 ( .A(n7051), .B(n7050), .Z(n6945) );
  INV_X1 U8783 ( .A(n6939), .ZN(n7156) );
  AOI22_X1 U8784 ( .A1(n8136), .A2(n6877), .B1(n8092), .B2(n8391), .ZN(n6941)
         );
  OAI211_X1 U8785 ( .C1(n6942), .C2(n8145), .A(n6941), .B(n6940), .ZN(n6943)
         );
  AOI21_X1 U8786 ( .B1(n7156), .B2(n8141), .A(n6943), .ZN(n6944) );
  OAI21_X1 U8787 ( .B1(n6945), .B2(n8132), .A(n6944), .ZN(P2_U3167) );
  AOI21_X1 U8788 ( .B1(n6948), .B2(n6947), .A(n6946), .ZN(n6953) );
  AOI22_X1 U8789 ( .A1(n8878), .A2(n9653), .B1(n8887), .B2(n9637), .ZN(n6952)
         );
  NAND2_X1 U8790 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9528) );
  INV_X1 U8791 ( .A(n9528), .ZN(n6950) );
  NOR2_X1 U8792 ( .A1(n8851), .A2(n9714), .ZN(n6949) );
  AOI211_X1 U8793 ( .C1(n9639), .C2(n8889), .A(n6950), .B(n6949), .ZN(n6951)
         );
  OAI211_X1 U8794 ( .C1(n6953), .C2(n8897), .A(n6952), .B(n6951), .ZN(P1_U3239) );
  XOR2_X1 U8795 ( .A(n6954), .B(n7769), .Z(n6955) );
  OAI222_X1 U8796 ( .A1(n9616), .A2(n6957), .B1(n9618), .B2(n6956), .C1(n9138), 
        .C2(n6955), .ZN(n9709) );
  INV_X1 U8797 ( .A(n9709), .ZN(n6967) );
  XNOR2_X1 U8798 ( .A(n6958), .B(n7769), .ZN(n9711) );
  INV_X1 U8799 ( .A(n9665), .ZN(n6960) );
  INV_X1 U8800 ( .A(n9646), .ZN(n6959) );
  OAI211_X1 U8801 ( .C1(n9708), .C2(n6960), .A(n6959), .B(n9666), .ZN(n9707)
         );
  NAND2_X1 U8802 ( .A1(n7202), .A2(n6961), .ZN(n6964) );
  AOI22_X1 U8803 ( .A1(n9673), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6962), .B2(
        n9656), .ZN(n6963) );
  OAI211_X1 U8804 ( .C1(n9707), .C2(n8982), .A(n6964), .B(n6963), .ZN(n6965)
         );
  AOI21_X1 U8805 ( .B1(n9711), .B2(n9670), .A(n6965), .ZN(n6966) );
  OAI21_X1 U8806 ( .B1(n6967), .B2(n9673), .A(n6966), .ZN(P1_U3288) );
  INV_X1 U8807 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9959) );
  INV_X1 U8808 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9597) );
  INV_X1 U8809 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9244) );
  AOI22_X1 U8810 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9597), .B2(n9244), .ZN(n9965) );
  NOR2_X1 U8811 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6968) );
  AOI21_X1 U8812 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6968), .ZN(n9968) );
  NOR2_X1 U8813 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6969) );
  AOI21_X1 U8814 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6969), .ZN(n9971) );
  NOR2_X1 U8815 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6970) );
  AOI21_X1 U8816 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6970), .ZN(n9974) );
  NOR2_X1 U8817 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6971) );
  AOI21_X1 U8818 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6971), .ZN(n9977) );
  NOR2_X1 U8819 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6972) );
  AOI21_X1 U8820 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6972), .ZN(n9980) );
  NOR2_X1 U8821 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6973) );
  AOI21_X1 U8822 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6973), .ZN(n9983) );
  NOR2_X1 U8823 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6974) );
  AOI21_X1 U8824 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6974), .ZN(n9986) );
  NOR2_X1 U8825 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n6975) );
  AOI21_X1 U8826 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n6975), .ZN(n9995) );
  NOR2_X1 U8827 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6976) );
  AOI21_X1 U8828 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6976), .ZN(n10001) );
  NOR2_X1 U8829 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6977) );
  AOI21_X1 U8830 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6977), .ZN(n9998) );
  NOR2_X1 U8831 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6978) );
  AOI21_X1 U8832 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6978), .ZN(n9989) );
  NOR2_X1 U8833 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6979) );
  AOI21_X1 U8834 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6979), .ZN(n9992) );
  AND2_X1 U8835 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6980) );
  NOR2_X1 U8836 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6980), .ZN(n9954) );
  INV_X1 U8837 ( .A(n9954), .ZN(n9955) );
  INV_X1 U8838 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9957) );
  NAND3_X1 U8839 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U8840 ( .A1(n9957), .A2(n9956), .ZN(n9953) );
  NAND2_X1 U8841 ( .A1(n9955), .A2(n9953), .ZN(n10004) );
  NAND2_X1 U8842 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6981) );
  OAI21_X1 U8843 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6981), .ZN(n10003) );
  NOR2_X1 U8844 ( .A1(n10004), .A2(n10003), .ZN(n10002) );
  AOI21_X1 U8845 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10002), .ZN(n10007) );
  NAND2_X1 U8846 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6982) );
  OAI21_X1 U8847 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6982), .ZN(n10006) );
  NOR2_X1 U8848 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  AOI21_X1 U8849 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10005), .ZN(n10010) );
  NOR2_X1 U8850 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6983) );
  AOI21_X1 U8851 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6983), .ZN(n10009) );
  NAND2_X1 U8852 ( .A1(n10010), .A2(n10009), .ZN(n10008) );
  OAI21_X1 U8853 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10008), .ZN(n9991) );
  NAND2_X1 U8854 ( .A1(n9992), .A2(n9991), .ZN(n9990) );
  OAI21_X1 U8855 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n9990), .ZN(n9988) );
  NAND2_X1 U8856 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  OAI21_X1 U8857 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n9987), .ZN(n9997) );
  NAND2_X1 U8858 ( .A1(n9998), .A2(n9997), .ZN(n9996) );
  OAI21_X1 U8859 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n9996), .ZN(n10000) );
  NAND2_X1 U8860 ( .A1(n10001), .A2(n10000), .ZN(n9999) );
  OAI21_X1 U8861 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n9999), .ZN(n9994) );
  NAND2_X1 U8862 ( .A1(n9995), .A2(n9994), .ZN(n9993) );
  OAI21_X1 U8863 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n9993), .ZN(n9985) );
  NAND2_X1 U8864 ( .A1(n9986), .A2(n9985), .ZN(n9984) );
  OAI21_X1 U8865 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9984), .ZN(n9982) );
  NAND2_X1 U8866 ( .A1(n9983), .A2(n9982), .ZN(n9981) );
  OAI21_X1 U8867 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9981), .ZN(n9979) );
  NAND2_X1 U8868 ( .A1(n9980), .A2(n9979), .ZN(n9978) );
  OAI21_X1 U8869 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9978), .ZN(n9976) );
  NAND2_X1 U8870 ( .A1(n9977), .A2(n9976), .ZN(n9975) );
  OAI21_X1 U8871 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9975), .ZN(n9973) );
  NAND2_X1 U8872 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  OAI21_X1 U8873 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9972), .ZN(n9970) );
  NAND2_X1 U8874 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  OAI21_X1 U8875 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9969), .ZN(n9967) );
  NAND2_X1 U8876 ( .A1(n9968), .A2(n9967), .ZN(n9966) );
  OAI21_X1 U8877 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9966), .ZN(n9964) );
  NAND2_X1 U8878 ( .A1(n9965), .A2(n9964), .ZN(n9963) );
  OAI21_X1 U8879 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9963), .ZN(n9960) );
  NOR2_X1 U8880 ( .A1(n9959), .A2(n9960), .ZN(n6984) );
  NAND2_X1 U8881 ( .A1(n9959), .A2(n9960), .ZN(n9958) );
  OAI21_X1 U8882 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6984), .A(n9958), .ZN(
        n6987) );
  XNOR2_X1 U8883 ( .A(n6985), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n6986) );
  XNOR2_X1 U8884 ( .A(n6987), .B(n6986), .ZN(ADD_1068_U4) );
  INV_X1 U8885 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9866) );
  INV_X1 U8886 ( .A(n6033), .ZN(n9884) );
  AOI22_X1 U8887 ( .A1(n8136), .A2(n6922), .B1(n8092), .B2(n6877), .ZN(n6989)
         );
  OAI211_X1 U8888 ( .C1(n9884), .C2(n8145), .A(n6989), .B(n6988), .ZN(n6994)
         );
  INV_X1 U8889 ( .A(n6892), .ZN(n6990) );
  AOI211_X1 U8890 ( .C1(n6992), .C2(n6991), .A(n8132), .B(n6990), .ZN(n6993)
         );
  AOI211_X1 U8891 ( .C1(n9866), .C2(n8141), .A(n6994), .B(n6993), .ZN(n6995)
         );
  INV_X1 U8892 ( .A(n6995), .ZN(P2_U3158) );
  XNOR2_X1 U8893 ( .A(n6996), .B(n6997), .ZN(n9746) );
  INV_X1 U8894 ( .A(n9746), .ZN(n7007) );
  OAI21_X1 U8895 ( .B1(n7773), .B2(n7842), .A(n7078), .ZN(n6998) );
  NAND2_X1 U8896 ( .A1(n6998), .A2(n9655), .ZN(n7000) );
  AOI22_X1 U8897 ( .A1(n9651), .A2(n8909), .B1(n8907), .B2(n9652), .ZN(n6999)
         );
  NAND2_X1 U8898 ( .A1(n7000), .A2(n6999), .ZN(n9745) );
  INV_X1 U8899 ( .A(n7085), .ZN(n7001) );
  OAI211_X1 U8900 ( .C1(n9743), .C2(n7002), .A(n7001), .B(n9666), .ZN(n9742)
         );
  AOI22_X1 U8901 ( .A1(n9673), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7427), .B2(
        n9656), .ZN(n7004) );
  NAND2_X1 U8902 ( .A1(n7202), .A2(n5476), .ZN(n7003) );
  OAI211_X1 U8903 ( .C1(n9742), .C2(n8982), .A(n7004), .B(n7003), .ZN(n7005)
         );
  AOI21_X1 U8904 ( .B1(n9745), .B2(n9113), .A(n7005), .ZN(n7006) );
  OAI21_X1 U8905 ( .B1(n7007), .B2(n9152), .A(n7006), .ZN(P1_U3283) );
  NAND2_X1 U8906 ( .A1(n7008), .A2(n7640), .ZN(n7035) );
  OR2_X1 U8907 ( .A1(n7035), .A2(n7645), .ZN(n7037) );
  NAND2_X1 U8908 ( .A1(n7037), .A2(n7009), .ZN(n9615) );
  INV_X1 U8909 ( .A(n7010), .ZN(n9621) );
  NAND2_X1 U8910 ( .A1(n9615), .A2(n9621), .ZN(n9614) );
  NAND2_X1 U8911 ( .A1(n9614), .A2(n7646), .ZN(n7012) );
  INV_X1 U8912 ( .A(n7016), .ZN(n7011) );
  XNOR2_X1 U8913 ( .A(n7012), .B(n7011), .ZN(n7014) );
  AND2_X1 U8914 ( .A1(n8910), .A2(n9651), .ZN(n7013) );
  AOI21_X1 U8915 ( .B1(n7014), .B2(n9655), .A(n7013), .ZN(n9740) );
  XNOR2_X1 U8916 ( .A(n7015), .B(n7016), .ZN(n9738) );
  XNOR2_X1 U8917 ( .A(n9631), .B(n4523), .ZN(n7018) );
  AND2_X1 U8918 ( .A1(n8908), .A2(n9652), .ZN(n7017) );
  AOI21_X1 U8919 ( .B1(n7018), .B2(n9666), .A(n7017), .ZN(n9736) );
  AOI22_X1 U8920 ( .A1(n9673), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7264), .B2(
        n9656), .ZN(n7020) );
  NAND2_X1 U8921 ( .A1(n7202), .A2(n5078), .ZN(n7019) );
  OAI211_X1 U8922 ( .C1(n9736), .C2(n8982), .A(n7020), .B(n7019), .ZN(n7021)
         );
  AOI21_X1 U8923 ( .B1(n9738), .B2(n9670), .A(n7021), .ZN(n7022) );
  OAI21_X1 U8924 ( .B1(n9740), .B2(n9673), .A(n7022), .ZN(P1_U3284) );
  XNOR2_X1 U8925 ( .A(n7023), .B(n6346), .ZN(n7026) );
  INV_X1 U8926 ( .A(n7026), .ZN(n9880) );
  NAND2_X1 U8927 ( .A1(n8608), .A2(n7024), .ZN(n7931) );
  XNOR2_X1 U8928 ( .A(n7025), .B(n6346), .ZN(n7029) );
  INV_X1 U8929 ( .A(n7364), .ZN(n7285) );
  NAND2_X1 U8930 ( .A1(n7026), .A2(n7285), .ZN(n7028) );
  AOI22_X1 U8931 ( .A1(n6758), .A2(n9858), .B1(n9859), .B2(n8393), .ZN(n7027)
         );
  OAI211_X1 U8932 ( .C1(n9872), .C2(n7029), .A(n7028), .B(n7027), .ZN(n9881)
         );
  OAI22_X1 U8933 ( .A1(n8618), .A2(n6018), .B1(n9879), .B2(n7441), .ZN(n7030)
         );
  NOR2_X1 U8934 ( .A1(n9881), .A2(n7030), .ZN(n7032) );
  MUX2_X1 U8935 ( .A(n7032), .B(n7031), .S(n9870), .Z(n7033) );
  OAI21_X1 U8936 ( .B1(n9880), .B2(n7931), .A(n7033), .ZN(P2_U3231) );
  XNOR2_X1 U8937 ( .A(n7034), .B(n7645), .ZN(n9720) );
  NAND2_X1 U8938 ( .A1(n9720), .A2(n7084), .ZN(n7041) );
  NAND2_X1 U8939 ( .A1(n7035), .A2(n7645), .ZN(n7036) );
  NAND2_X1 U8940 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  NAND2_X1 U8941 ( .A1(n7038), .A2(n9655), .ZN(n7040) );
  AOI22_X1 U8942 ( .A1(n9651), .A2(n8911), .B1(n8910), .B2(n9652), .ZN(n7039)
         );
  NAND3_X1 U8943 ( .A1(n7041), .A2(n7040), .A3(n7039), .ZN(n9725) );
  INV_X1 U8944 ( .A(n9725), .ZN(n7049) );
  OAI211_X1 U8945 ( .C1(n9644), .C2(n9723), .A(n9666), .B(n9630), .ZN(n9721)
         );
  INV_X1 U8946 ( .A(n7042), .ZN(n7072) );
  OAI22_X1 U8947 ( .A1(n9113), .A2(n7043), .B1(n7072), .B2(n9104), .ZN(n7044)
         );
  AOI21_X1 U8948 ( .B1(n7202), .B2(n7045), .A(n7044), .ZN(n7046) );
  OAI21_X1 U8949 ( .B1(n8982), .B2(n9721), .A(n7046), .ZN(n7047) );
  AOI21_X1 U8950 ( .B1(n9720), .B2(n9634), .A(n7047), .ZN(n7048) );
  OAI21_X1 U8951 ( .B1(n7049), .B2(n9658), .A(n7048), .ZN(P1_U3286) );
  NAND2_X1 U8952 ( .A1(n7051), .A2(n7050), .ZN(n7055) );
  INV_X1 U8953 ( .A(n7052), .ZN(n7053) );
  NAND2_X1 U8954 ( .A1(n7053), .A2(n7172), .ZN(n7054) );
  NAND2_X1 U8955 ( .A1(n7055), .A2(n7054), .ZN(n7056) );
  XNOR2_X1 U8956 ( .A(n8024), .B(n9900), .ZN(n7134) );
  XNOR2_X1 U8957 ( .A(n7134), .B(n8391), .ZN(n7057) );
  AOI21_X1 U8958 ( .B1(n7056), .B2(n7057), .A(n8132), .ZN(n7060) );
  INV_X1 U8959 ( .A(n7056), .ZN(n7059) );
  INV_X1 U8960 ( .A(n7057), .ZN(n7058) );
  NAND2_X1 U8961 ( .A1(n7060), .A2(n7136), .ZN(n7065) );
  INV_X1 U8962 ( .A(n7061), .ZN(n7063) );
  OAI22_X1 U8963 ( .A1(n8145), .A2(n9900), .B1(n7919), .B2(n8138), .ZN(n7062)
         );
  AOI211_X1 U8964 ( .C1(n8136), .C2(n8392), .A(n7063), .B(n7062), .ZN(n7064)
         );
  OAI211_X1 U8965 ( .C1(n7175), .C2(n8075), .A(n7065), .B(n7064), .ZN(P2_U3179) );
  INV_X1 U8966 ( .A(n7066), .ZN(n7927) );
  OAI222_X1 U8967 ( .A1(n8751), .A2(n7068), .B1(n7936), .B2(n7927), .C1(n7067), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  NAND2_X1 U8968 ( .A1(n4362), .A2(n7069), .ZN(n7070) );
  XNOR2_X1 U8969 ( .A(n4354), .B(n7070), .ZN(n7071) );
  NAND2_X1 U8970 ( .A1(n7071), .A2(n8876), .ZN(n7076) );
  NAND2_X1 U8971 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9422) );
  INV_X1 U8972 ( .A(n9422), .ZN(n7074) );
  OAI22_X1 U8973 ( .A1(n8846), .A2(n7072), .B1(n7265), .B2(n8867), .ZN(n7073)
         );
  AOI211_X1 U8974 ( .C1(n8878), .C2(n8911), .A(n7074), .B(n7073), .ZN(n7075)
         );
  OAI211_X1 U8975 ( .C1(n9723), .C2(n8851), .A(n7076), .B(n7075), .ZN(P1_U3213) );
  XNOR2_X1 U8976 ( .A(n7077), .B(n7776), .ZN(n9752) );
  NAND2_X1 U8977 ( .A1(n7078), .A2(n7655), .ZN(n7080) );
  INV_X1 U8978 ( .A(n7776), .ZN(n7079) );
  XNOR2_X1 U8979 ( .A(n7080), .B(n7079), .ZN(n7082) );
  AOI22_X1 U8980 ( .A1(n9651), .A2(n8908), .B1(n7474), .B2(n9652), .ZN(n7081)
         );
  OAI21_X1 U8981 ( .B1(n7082), .B2(n9138), .A(n7081), .ZN(n7083) );
  AOI21_X1 U8982 ( .B1(n9752), .B2(n7084), .A(n7083), .ZN(n9754) );
  OAI211_X1 U8983 ( .C1(n7085), .C2(n9749), .A(n9666), .B(n7097), .ZN(n9748)
         );
  AOI22_X1 U8984 ( .A1(n9673), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7488), .B2(
        n9656), .ZN(n7088) );
  NAND2_X1 U8985 ( .A1(n7086), .A2(n7202), .ZN(n7087) );
  OAI211_X1 U8986 ( .C1(n9748), .C2(n8982), .A(n7088), .B(n7087), .ZN(n7089)
         );
  AOI21_X1 U8987 ( .B1(n9752), .B2(n9634), .A(n7089), .ZN(n7090) );
  OAI21_X1 U8988 ( .B1(n9754), .B2(n9658), .A(n7090), .ZN(P1_U3282) );
  XNOR2_X1 U8989 ( .A(n7091), .B(n7093), .ZN(n9760) );
  INV_X1 U8990 ( .A(n9760), .ZN(n7105) );
  XNOR2_X1 U8991 ( .A(n7093), .B(n7092), .ZN(n7094) );
  NAND2_X1 U8992 ( .A1(n7094), .A2(n9655), .ZN(n7096) );
  AOI22_X1 U8993 ( .A1(n9651), .A2(n8907), .B1(n8906), .B2(n9652), .ZN(n7095)
         );
  NAND2_X1 U8994 ( .A1(n7096), .A2(n7095), .ZN(n9759) );
  INV_X1 U8995 ( .A(n7097), .ZN(n7099) );
  OAI211_X1 U8996 ( .C1(n7099), .C2(n9757), .A(n9666), .B(n7198), .ZN(n9756)
         );
  AOI22_X1 U8997 ( .A1(n9673), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7399), .B2(
        n9656), .ZN(n7102) );
  NAND2_X1 U8998 ( .A1(n7100), .A2(n7202), .ZN(n7101) );
  OAI211_X1 U8999 ( .C1(n9756), .C2(n8982), .A(n7102), .B(n7101), .ZN(n7103)
         );
  AOI21_X1 U9000 ( .B1(n9759), .B2(n9113), .A(n7103), .ZN(n7104) );
  OAI21_X1 U9001 ( .B1(n7105), .B2(n9152), .A(n7104), .ZN(P1_U3281) );
  AOI21_X1 U9002 ( .B1(n7108), .B2(n7107), .A(n7106), .ZN(n7122) );
  OAI21_X1 U9003 ( .B1(n7110), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7109), .ZN(
        n7120) );
  NOR2_X1 U9004 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7111), .ZN(n7241) );
  AOI21_X1 U9005 ( .B1(n9841), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7241), .ZN(
        n7112) );
  OAI21_X1 U9006 ( .B1(n8473), .B2(n7113), .A(n7112), .ZN(n7119) );
  INV_X1 U9007 ( .A(n7114), .ZN(n7115) );
  NAND2_X1 U9008 ( .A1(n7115), .A2(n6102), .ZN(n7117) );
  AOI21_X1 U9009 ( .B1(n7117), .B2(n7116), .A(n9822), .ZN(n7118) );
  AOI211_X1 U9010 ( .C1(n9852), .C2(n7120), .A(n7119), .B(n7118), .ZN(n7121)
         );
  OAI21_X1 U9011 ( .B1(n7122), .B2(n9844), .A(n7121), .ZN(P2_U3191) );
  XOR2_X1 U9012 ( .A(n7123), .B(n8316), .Z(n9888) );
  AND2_X1 U9013 ( .A1(n7125), .A2(n7124), .ZN(n7127) );
  OAI21_X1 U9014 ( .B1(n7127), .B2(n6044), .A(n7126), .ZN(n7128) );
  AOI222_X1 U9015 ( .A1(n9861), .A2(n7128), .B1(n8393), .B2(n9858), .C1(n8392), 
        .C2(n9859), .ZN(n9889) );
  MUX2_X1 U9016 ( .A(n7129), .B(n9889), .S(n8608), .Z(n7132) );
  AOI22_X1 U9017 ( .A1(n9864), .A2(n8166), .B1(n9865), .B2(n7130), .ZN(n7131)
         );
  OAI211_X1 U9018 ( .C1(n9888), .C2(n8615), .A(n7132), .B(n7131), .ZN(P2_U3229) );
  INV_X1 U9019 ( .A(n7133), .ZN(n7145) );
  OAI222_X1 U9020 ( .A1(n7936), .A2(n7145), .B1(P2_U3151), .B2(n8303), .C1(
        n9349), .C2(n8751), .ZN(P2_U3275) );
  NAND2_X1 U9021 ( .A1(n7134), .A2(n8391), .ZN(n7135) );
  XNOR2_X1 U9022 ( .A(n8024), .B(n9903), .ZN(n7236) );
  XNOR2_X1 U9023 ( .A(n7236), .B(n7919), .ZN(n7137) );
  OAI21_X1 U9024 ( .B1(n4359), .B2(n7137), .A(n7238), .ZN(n7138) );
  NAND2_X1 U9025 ( .A1(n7138), .A2(n8116), .ZN(n7144) );
  OR2_X1 U9026 ( .A1(n8095), .A2(n7283), .ZN(n7140) );
  OAI211_X1 U9027 ( .C1(n8138), .C2(n7282), .A(n7140), .B(n7139), .ZN(n7142)
         );
  NOR2_X1 U9028 ( .A1(n8075), .A2(n7289), .ZN(n7141) );
  NOR2_X1 U9029 ( .A1(n7142), .A2(n7141), .ZN(n7143) );
  OAI211_X1 U9030 ( .C1(n9903), .C2(n8145), .A(n7144), .B(n7143), .ZN(P2_U3153) );
  OAI222_X1 U9031 ( .A1(P1_U3086), .A2(n7146), .B1(n9395), .B2(n7145), .C1(
        n9350), .C2(n9392), .ZN(P1_U3335) );
  OR2_X1 U9032 ( .A1(n7148), .A2(n8319), .ZN(n7149) );
  NAND2_X1 U9033 ( .A1(n7147), .A2(n7149), .ZN(n9895) );
  INV_X1 U9034 ( .A(n9895), .ZN(n7159) );
  OAI22_X1 U9035 ( .A1(n8165), .A2(n8605), .B1(n7283), .B2(n8607), .ZN(n7150)
         );
  AOI21_X1 U9036 ( .B1(n9895), .B2(n7285), .A(n7150), .ZN(n7155) );
  INV_X1 U9037 ( .A(n8319), .ZN(n7152) );
  XNOR2_X1 U9038 ( .A(n7151), .B(n7152), .ZN(n7153) );
  NAND2_X1 U9039 ( .A1(n7153), .A2(n9861), .ZN(n7154) );
  AND2_X1 U9040 ( .A1(n7155), .A2(n7154), .ZN(n9897) );
  MUX2_X1 U9041 ( .A(n9897), .B(n6708), .S(n9870), .Z(n7158) );
  AOI22_X1 U9042 ( .A1(n9864), .A2(n9894), .B1(n9865), .B2(n7156), .ZN(n7157)
         );
  OAI211_X1 U9043 ( .C1(n7159), .C2(n7931), .A(n7158), .B(n7157), .ZN(P2_U3228) );
  INV_X1 U9044 ( .A(n7160), .ZN(n7170) );
  OAI222_X1 U9045 ( .A1(n7936), .A2(n7170), .B1(P2_U3151), .B2(n8361), .C1(
        n7161), .C2(n8751), .ZN(P2_U3274) );
  INV_X1 U9046 ( .A(n7162), .ZN(n7168) );
  OR2_X1 U9047 ( .A1(n8608), .A2(n9809), .ZN(n7164) );
  NAND2_X1 U9048 ( .A1(n9865), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7163) );
  OAI211_X1 U9049 ( .C1(n8620), .C2(n6013), .A(n7164), .B(n7163), .ZN(n7165)
         );
  AOI21_X1 U9050 ( .B1(n9867), .B2(n7166), .A(n7165), .ZN(n7167) );
  OAI21_X1 U9051 ( .B1(n7168), .B2(n9870), .A(n7167), .ZN(P2_U3232) );
  OAI222_X1 U9052 ( .A1(P1_U3086), .A2(n7837), .B1(n9395), .B2(n7170), .C1(
        n7169), .C2(n9392), .ZN(P1_U3334) );
  AOI21_X1 U9053 ( .B1(n7171), .B2(n8318), .A(n9872), .ZN(n7174) );
  OAI22_X1 U9054 ( .A1(n7172), .A2(n8605), .B1(n7919), .B2(n8607), .ZN(n7173)
         );
  AOI21_X1 U9055 ( .B1(n7174), .B2(n7273), .A(n7173), .ZN(n9899) );
  OAI22_X1 U9056 ( .A1(n8608), .A2(n6065), .B1(n7175), .B2(n8618), .ZN(n7176)
         );
  AOI21_X1 U9057 ( .B1(n9864), .B2(n7177), .A(n7176), .ZN(n7180) );
  NAND2_X1 U9058 ( .A1(n7147), .A2(n8171), .ZN(n7178) );
  XNOR2_X1 U9059 ( .A(n7178), .B(n8318), .ZN(n9902) );
  NAND2_X1 U9060 ( .A1(n9902), .A2(n9867), .ZN(n7179) );
  OAI211_X1 U9061 ( .C1(n9899), .C2(n9870), .A(n7180), .B(n7179), .ZN(P2_U3227) );
  INV_X1 U9062 ( .A(n7181), .ZN(n9728) );
  OAI21_X1 U9063 ( .B1(n7184), .B2(n7183), .A(n7182), .ZN(n7185) );
  NAND2_X1 U9064 ( .A1(n7185), .A2(n8876), .ZN(n7190) );
  NAND2_X1 U9065 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9452) );
  INV_X1 U9066 ( .A(n9452), .ZN(n7188) );
  INV_X1 U9067 ( .A(n9626), .ZN(n7186) );
  OAI22_X1 U9068 ( .A1(n8846), .A2(n7186), .B1(n9617), .B2(n8867), .ZN(n7187)
         );
  AOI211_X1 U9069 ( .C1(n8878), .C2(n9637), .A(n7188), .B(n7187), .ZN(n7189)
         );
  OAI211_X1 U9070 ( .C1(n9728), .C2(n8851), .A(n7190), .B(n7189), .ZN(P1_U3221) );
  NOR2_X1 U9071 ( .A1(n7191), .A2(n7777), .ZN(n7192) );
  OAI21_X1 U9072 ( .B1(n7192), .B2(n7250), .A(n9655), .ZN(n7194) );
  AOI22_X1 U9073 ( .A1(n9651), .A2(n7474), .B1(n8905), .B2(n9652), .ZN(n7193)
         );
  AND2_X1 U9074 ( .A1(n7194), .A2(n7193), .ZN(n9763) );
  XNOR2_X1 U9075 ( .A(n7195), .B(n7777), .ZN(n9765) );
  NAND2_X1 U9076 ( .A1(n9765), .A2(n9670), .ZN(n7204) );
  INV_X1 U9077 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7197) );
  INV_X1 U9078 ( .A(n7196), .ZN(n7471) );
  OAI22_X1 U9079 ( .A1(n9113), .A2(n7197), .B1(n7471), .B2(n9104), .ZN(n7200)
         );
  OAI211_X1 U9080 ( .C1(n7098), .C2(n5500), .A(n9666), .B(n7254), .ZN(n9762)
         );
  NOR2_X1 U9081 ( .A1(n9762), .A2(n8982), .ZN(n7199) );
  AOI211_X1 U9082 ( .C1(n7202), .C2(n7201), .A(n7200), .B(n7199), .ZN(n7203)
         );
  OAI211_X1 U9083 ( .C1(n9658), .C2(n9763), .A(n7204), .B(n7203), .ZN(P1_U3280) );
  XNOR2_X1 U9084 ( .A(n4282), .B(n8327), .ZN(n7208) );
  NAND2_X1 U9085 ( .A1(n8386), .A2(n9859), .ZN(n7206) );
  NAND2_X1 U9086 ( .A1(n8388), .A2(n9858), .ZN(n7205) );
  NAND2_X1 U9087 ( .A1(n7206), .A2(n7205), .ZN(n7207) );
  AOI21_X1 U9088 ( .B1(n7208), .B2(n9861), .A(n7207), .ZN(n9924) );
  OAI22_X1 U9089 ( .A1(n8608), .A2(n7505), .B1(n7461), .B2(n8618), .ZN(n7209)
         );
  AOI21_X1 U9090 ( .B1(n9864), .B2(n9920), .A(n7209), .ZN(n7212) );
  XNOR2_X1 U9091 ( .A(n7210), .B(n8327), .ZN(n9922) );
  NAND2_X1 U9092 ( .A1(n9922), .A2(n9867), .ZN(n7211) );
  OAI211_X1 U9093 ( .C1(n9924), .C2(n9870), .A(n7212), .B(n7211), .ZN(P2_U3222) );
  AOI21_X1 U9094 ( .B1(n7215), .B2(n7214), .A(n7213), .ZN(n7231) );
  AOI21_X1 U9095 ( .B1(n7218), .B2(n7217), .A(n7216), .ZN(n7228) );
  AOI21_X1 U9096 ( .B1(n7221), .B2(n7220), .A(n7219), .ZN(n7222) );
  OR2_X1 U9097 ( .A1(n7222), .A2(n9822), .ZN(n7227) );
  INV_X1 U9098 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9245) );
  AND2_X1 U9099 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7416) );
  INV_X1 U9100 ( .A(n7416), .ZN(n7223) );
  OAI21_X1 U9101 ( .B1(n9831), .B2(n9245), .A(n7223), .ZN(n7224) );
  AOI21_X1 U9102 ( .B1(n7225), .B2(n9839), .A(n7224), .ZN(n7226) );
  OAI211_X1 U9103 ( .C1(n7228), .C2(n8485), .A(n7227), .B(n7226), .ZN(n7229)
         );
  INV_X1 U9104 ( .A(n7229), .ZN(n7230) );
  OAI21_X1 U9105 ( .B1(n7231), .B2(n9844), .A(n7230), .ZN(P2_U3192) );
  INV_X1 U9106 ( .A(n7232), .ZN(n7234) );
  OAI222_X1 U9107 ( .A1(n8751), .A2(n9297), .B1(n7936), .B2(n7234), .C1(n8359), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9108 ( .A1(n7235), .A2(P1_U3086), .B1(n9395), .B2(n7234), .C1(
        n7233), .C2(n9392), .ZN(P1_U3333) );
  INV_X1 U9109 ( .A(n7236), .ZN(n7237) );
  XNOR2_X1 U9110 ( .A(n8024), .B(n7239), .ZN(n7912) );
  AND2_X1 U9111 ( .A1(n7912), .A2(n7282), .ZN(n7240) );
  XNOR2_X1 U9112 ( .A(n9908), .B(n8024), .ZN(n7408) );
  XNOR2_X1 U9113 ( .A(n7408), .B(n7916), .ZN(n7406) );
  XNOR2_X1 U9114 ( .A(n7407), .B(n7406), .ZN(n7248) );
  OR2_X1 U9115 ( .A1(n8095), .A2(n7282), .ZN(n7243) );
  INV_X1 U9116 ( .A(n7241), .ZN(n7242) );
  OAI211_X1 U9117 ( .C1(n8138), .C2(n8197), .A(n7243), .B(n7242), .ZN(n7245)
         );
  NOR2_X1 U9118 ( .A1(n8075), .A2(n7365), .ZN(n7244) );
  NOR2_X1 U9119 ( .A1(n7245), .A2(n7244), .ZN(n7247) );
  NAND2_X1 U9120 ( .A1(n8129), .A2(n6111), .ZN(n7246) );
  OAI211_X1 U9121 ( .C1(n7248), .C2(n8132), .A(n7247), .B(n7246), .ZN(P2_U3171) );
  XNOR2_X1 U9122 ( .A(n7249), .B(n7779), .ZN(n9774) );
  INV_X1 U9123 ( .A(n9774), .ZN(n7261) );
  OAI21_X1 U9124 ( .B1(n7250), .B2(n7856), .A(n7779), .ZN(n7251) );
  NAND3_X1 U9125 ( .A1(n4691), .A2(n9655), .A3(n7251), .ZN(n7253) );
  AOI22_X1 U9126 ( .A1(n9651), .A2(n8906), .B1(n8904), .B2(n9652), .ZN(n7252)
         );
  NAND2_X1 U9127 ( .A1(n7253), .A2(n7252), .ZN(n9772) );
  INV_X1 U9128 ( .A(n7254), .ZN(n7255) );
  OAI21_X1 U9129 ( .B1(n9768), .B2(n7255), .A(n4351), .ZN(n9770) );
  INV_X1 U9130 ( .A(n7907), .ZN(n7256) );
  NOR2_X1 U9131 ( .A1(n9770), .A2(n7256), .ZN(n7259) );
  AOI22_X1 U9132 ( .A1(n9673), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8755), .B2(
        n9656), .ZN(n7257) );
  OAI21_X1 U9133 ( .B1(n9768), .B2(n9660), .A(n7257), .ZN(n7258) );
  AOI211_X1 U9134 ( .C1(n9772), .C2(n9113), .A(n7259), .B(n7258), .ZN(n7260)
         );
  OAI21_X1 U9135 ( .B1(n7261), .B2(n9152), .A(n7260), .ZN(P1_U3279) );
  XOR2_X1 U9136 ( .A(n7263), .B(n7262), .Z(n7271) );
  INV_X1 U9137 ( .A(n7264), .ZN(n7266) );
  OAI22_X1 U9138 ( .A1(n8846), .A2(n7266), .B1(n7265), .B2(n8891), .ZN(n7267)
         );
  AOI211_X1 U9139 ( .C1(n8887), .C2(n8908), .A(n7268), .B(n7267), .ZN(n7270)
         );
  NAND2_X1 U9140 ( .A1(n8894), .A2(n5078), .ZN(n7269) );
  OAI211_X1 U9141 ( .C1(n7271), .C2(n8897), .A(n7270), .B(n7269), .ZN(P1_U3231) );
  NAND2_X1 U9142 ( .A1(n7335), .A2(n8323), .ZN(n7302) );
  OAI21_X1 U9143 ( .B1(n7335), .B2(n8323), .A(n7302), .ZN(n7274) );
  NAND2_X1 U9144 ( .A1(n7274), .A2(n9861), .ZN(n7287) );
  AND2_X1 U9145 ( .A1(n7276), .A2(n7275), .ZN(n7308) );
  NAND2_X1 U9146 ( .A1(n7147), .A2(n7277), .ZN(n7279) );
  AND2_X1 U9147 ( .A1(n7279), .A2(n7278), .ZN(n7280) );
  NAND2_X1 U9148 ( .A1(n7280), .A2(n8323), .ZN(n7281) );
  OAI22_X1 U9149 ( .A1(n7283), .A2(n8605), .B1(n7282), .B2(n8607), .ZN(n7284)
         );
  AOI21_X1 U9150 ( .B1(n9906), .B2(n7285), .A(n7284), .ZN(n7286) );
  NAND2_X1 U9151 ( .A1(n7287), .A2(n7286), .ZN(n9904) );
  MUX2_X1 U9152 ( .A(n9904), .B(P2_REG2_REG_7__SCAN_IN), .S(n9870), .Z(n7288)
         );
  INV_X1 U9153 ( .A(n7288), .ZN(n7293) );
  INV_X1 U9154 ( .A(n7931), .ZN(n7291) );
  OAI22_X1 U9155 ( .A1(n8620), .A2(n9903), .B1(n7289), .B2(n8618), .ZN(n7290)
         );
  AOI21_X1 U9156 ( .B1(n9906), .B2(n7291), .A(n7290), .ZN(n7292) );
  NAND2_X1 U9157 ( .A1(n7293), .A2(n7292), .ZN(P2_U3226) );
  NAND2_X1 U9158 ( .A1(n7297), .A2(n7294), .ZN(n7295) );
  OAI211_X1 U9159 ( .C1(n7296), .C2(n9392), .A(n7295), .B(n7901), .ZN(P1_U3332) );
  NAND2_X1 U9160 ( .A1(n7297), .A2(n8748), .ZN(n7299) );
  NAND2_X1 U9161 ( .A1(n7298), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8376) );
  OAI211_X1 U9162 ( .C1(n7300), .C2(n8751), .A(n7299), .B(n8376), .ZN(P2_U3272) );
  NAND2_X1 U9163 ( .A1(n7302), .A2(n7301), .ZN(n7357) );
  XNOR2_X1 U9164 ( .A(n7357), .B(n8321), .ZN(n7306) );
  NAND2_X1 U9165 ( .A1(n7303), .A2(n9859), .ZN(n7304) );
  OAI21_X1 U9166 ( .B1(n7919), .B2(n8605), .A(n7304), .ZN(n7305) );
  AOI21_X1 U9167 ( .B1(n7306), .B2(n9861), .A(n7305), .ZN(n7315) );
  MUX2_X1 U9168 ( .A(n5608), .B(n7315), .S(n8608), .Z(n7313) );
  NAND2_X1 U9169 ( .A1(n7308), .A2(n7307), .ZN(n7309) );
  XNOR2_X1 U9170 ( .A(n7309), .B(n8321), .ZN(n7314) );
  OAI22_X1 U9171 ( .A1(n8620), .A2(n7310), .B1(n4857), .B2(n8618), .ZN(n7311)
         );
  AOI21_X1 U9172 ( .B1(n7314), .B2(n9867), .A(n7311), .ZN(n7312) );
  NAND2_X1 U9173 ( .A1(n7313), .A2(n7312), .ZN(P2_U3225) );
  INV_X1 U9174 ( .A(n7314), .ZN(n7316) );
  OAI21_X1 U9175 ( .B1(n9926), .B2(n7316), .A(n7315), .ZN(n7321) );
  OAI22_X1 U9176 ( .A1(n8672), .A2(n7310), .B1(n9952), .B2(n9273), .ZN(n7317)
         );
  AOI21_X1 U9177 ( .B1(n7321), .B2(n9952), .A(n7317), .ZN(n7318) );
  INV_X1 U9178 ( .A(n7318), .ZN(P2_U3467) );
  INV_X1 U9179 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7319) );
  OAI22_X1 U9180 ( .A1(n7310), .A2(n8736), .B1(n9932), .B2(n7319), .ZN(n7320)
         );
  AOI21_X1 U9181 ( .B1(n7321), .B2(n9932), .A(n7320), .ZN(n7322) );
  INV_X1 U9182 ( .A(n7322), .ZN(P2_U3414) );
  OAI21_X1 U9183 ( .B1(n4339), .B2(n8209), .A(n7323), .ZN(n9927) );
  OAI211_X1 U9184 ( .C1(n4356), .C2(n8330), .A(n7324), .B(n9861), .ZN(n7326)
         );
  AOI22_X1 U9185 ( .A1(n9858), .A2(n8387), .B1(n8385), .B2(n9859), .ZN(n7325)
         );
  NAND2_X1 U9186 ( .A1(n7326), .A2(n7325), .ZN(n9928) );
  NAND2_X1 U9187 ( .A1(n9928), .A2(n8608), .ZN(n7330) );
  OAI22_X1 U9188 ( .A1(n8608), .A2(n7327), .B1(n7519), .B2(n8618), .ZN(n7328)
         );
  AOI21_X1 U9189 ( .B1(n9930), .B2(n9864), .A(n7328), .ZN(n7329) );
  OAI211_X1 U9190 ( .C1(n8615), .C2(n9927), .A(n7330), .B(n7329), .ZN(P2_U3221) );
  NAND2_X1 U9191 ( .A1(n7354), .A2(n8183), .ZN(n7333) );
  OR2_X1 U9192 ( .A1(n7332), .A2(n7331), .ZN(n8325) );
  XNOR2_X1 U9193 ( .A(n7333), .B(n8325), .ZN(n9916) );
  NAND2_X1 U9194 ( .A1(n7335), .A2(n7334), .ZN(n7337) );
  NAND2_X1 U9195 ( .A1(n7337), .A2(n7336), .ZN(n7338) );
  XOR2_X1 U9196 ( .A(n8325), .B(n7338), .Z(n7339) );
  NAND2_X1 U9197 ( .A1(n7339), .A2(n9861), .ZN(n7341) );
  AOI22_X1 U9198 ( .A1(n9858), .A2(n7303), .B1(n8387), .B2(n9859), .ZN(n7340)
         );
  OAI211_X1 U9199 ( .C1(n7364), .C2(n9916), .A(n7341), .B(n7340), .ZN(n9918)
         );
  NAND2_X1 U9200 ( .A1(n9918), .A2(n8608), .ZN(n7344) );
  OAI22_X1 U9201 ( .A1(n8608), .A2(n5679), .B1(n7415), .B2(n8618), .ZN(n7342)
         );
  AOI21_X1 U9202 ( .B1(n9864), .B2(n7411), .A(n7342), .ZN(n7343) );
  OAI211_X1 U9203 ( .C1(n9916), .C2(n7931), .A(n7344), .B(n7343), .ZN(P2_U3223) );
  XNOR2_X1 U9204 ( .A(n7345), .B(n4812), .ZN(n7387) );
  AOI21_X1 U9205 ( .B1(n4691), .B2(n7661), .A(n7781), .ZN(n7346) );
  NOR2_X1 U9206 ( .A1(n4338), .A2(n7346), .ZN(n7347) );
  OAI222_X1 U9207 ( .A1(n9618), .A2(n8892), .B1(n9616), .B2(n9143), .C1(n9138), 
        .C2(n7347), .ZN(n7384) );
  AOI211_X1 U9208 ( .C1(n8895), .C2(n4351), .A(n9769), .B(n7375), .ZN(n7385)
         );
  NAND2_X1 U9209 ( .A1(n7385), .A2(n9669), .ZN(n7349) );
  AOI22_X1 U9210 ( .A1(n9673), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8888), .B2(
        n9656), .ZN(n7348) );
  OAI211_X1 U9211 ( .C1(n7350), .C2(n9660), .A(n7349), .B(n7348), .ZN(n7351)
         );
  AOI21_X1 U9212 ( .B1(n7384), .B2(n9113), .A(n7351), .ZN(n7352) );
  OAI21_X1 U9213 ( .B1(n7387), .B2(n9152), .A(n7352), .ZN(P1_U3278) );
  AND2_X1 U9214 ( .A1(n7353), .A2(n8190), .ZN(n7356) );
  OAI21_X1 U9215 ( .B1(n7356), .B2(n7355), .A(n7354), .ZN(n9909) );
  NAND2_X1 U9216 ( .A1(n7357), .A2(n8321), .ZN(n7359) );
  NAND2_X1 U9217 ( .A1(n7359), .A2(n7358), .ZN(n7360) );
  XNOR2_X1 U9218 ( .A(n8322), .B(n7360), .ZN(n7361) );
  NAND2_X1 U9219 ( .A1(n7361), .A2(n9861), .ZN(n7363) );
  AOI22_X1 U9220 ( .A1(n8389), .A2(n9858), .B1(n9859), .B2(n8388), .ZN(n7362)
         );
  OAI211_X1 U9221 ( .C1(n7364), .C2(n9909), .A(n7363), .B(n7362), .ZN(n9911)
         );
  NAND2_X1 U9222 ( .A1(n9911), .A2(n8608), .ZN(n7368) );
  OAI22_X1 U9223 ( .A1(n8608), .A2(n6102), .B1(n7365), .B2(n8618), .ZN(n7366)
         );
  AOI21_X1 U9224 ( .B1(n9864), .B2(n6111), .A(n7366), .ZN(n7367) );
  OAI211_X1 U9225 ( .C1(n9909), .C2(n7931), .A(n7368), .B(n7367), .ZN(P2_U3224) );
  AOI21_X1 U9226 ( .B1(n7782), .B2(n7369), .A(n4343), .ZN(n7370) );
  INV_X1 U9227 ( .A(n7370), .ZN(n9221) );
  AOI21_X1 U9228 ( .B1(n7372), .B2(n7371), .A(n9142), .ZN(n7373) );
  OAI222_X1 U9229 ( .A1(n9616), .A2(n7374), .B1(n9618), .B2(n8809), .C1(n9138), 
        .C2(n7373), .ZN(n9217) );
  INV_X1 U9230 ( .A(n7375), .ZN(n7376) );
  AOI211_X1 U9231 ( .C1(n9219), .C2(n7376), .A(n9769), .B(n9132), .ZN(n9218)
         );
  NAND2_X1 U9232 ( .A1(n9218), .A2(n9669), .ZN(n7378) );
  AOI22_X1 U9233 ( .A1(n9673), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8808), .B2(
        n9656), .ZN(n7377) );
  OAI211_X1 U9234 ( .C1(n8814), .C2(n9660), .A(n7378), .B(n7377), .ZN(n7379)
         );
  AOI21_X1 U9235 ( .B1(n9217), .B2(n9113), .A(n7379), .ZN(n7380) );
  OAI21_X1 U9236 ( .B1(n9221), .B2(n9152), .A(n7380), .ZN(P1_U3277) );
  INV_X1 U9237 ( .A(n7381), .ZN(n7393) );
  OAI222_X1 U9238 ( .A1(n7936), .A2(n7393), .B1(P2_U3151), .B2(n7383), .C1(
        n7382), .C2(n8751), .ZN(P2_U3271) );
  INV_X1 U9239 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9574) );
  AOI211_X1 U9240 ( .C1(n9734), .C2(n8895), .A(n7385), .B(n7384), .ZN(n7386)
         );
  OAI21_X1 U9241 ( .B1(n9222), .B2(n7387), .A(n7386), .ZN(n7389) );
  NAND2_X1 U9242 ( .A1(n7389), .A2(n9803), .ZN(n7388) );
  OAI21_X1 U9243 ( .B1(n9803), .B2(n9574), .A(n7388), .ZN(P1_U3537) );
  INV_X1 U9244 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U9245 ( .A1(n7389), .A2(n9777), .ZN(n7390) );
  OAI21_X1 U9246 ( .B1(n9777), .B2(n7391), .A(n7390), .ZN(P1_U3498) );
  OAI222_X1 U9247 ( .A1(n7394), .A2(P1_U3086), .B1(n9395), .B2(n7393), .C1(
        n7392), .C2(n9392), .ZN(P1_U3331) );
  OAI21_X1 U9248 ( .B1(n7397), .B2(n7396), .A(n7395), .ZN(n7398) );
  NAND2_X1 U9249 ( .A1(n7398), .A2(n8876), .ZN(n7405) );
  INV_X1 U9250 ( .A(n7399), .ZN(n7401) );
  OAI22_X1 U9251 ( .A1(n8846), .A2(n7401), .B1(n7400), .B2(n8891), .ZN(n7402)
         );
  AOI211_X1 U9252 ( .C1(n8887), .C2(n8906), .A(n7403), .B(n7402), .ZN(n7404)
         );
  OAI211_X1 U9253 ( .C1(n9757), .C2(n8851), .A(n7405), .B(n7404), .ZN(P1_U3224) );
  INV_X1 U9254 ( .A(n7411), .ZN(n9914) );
  NAND2_X1 U9255 ( .A1(n7407), .A2(n7406), .ZN(n7410) );
  NAND2_X1 U9256 ( .A1(n7408), .A2(n7303), .ZN(n7409) );
  NAND2_X1 U9257 ( .A1(n7410), .A2(n7409), .ZN(n7452) );
  XNOR2_X1 U9258 ( .A(n7411), .B(n8024), .ZN(n7412) );
  OAI21_X1 U9259 ( .B1(n7413), .B2(n7412), .A(n7454), .ZN(n7414) );
  NAND2_X1 U9260 ( .A1(n7414), .A2(n8116), .ZN(n7421) );
  INV_X1 U9261 ( .A(n7415), .ZN(n7419) );
  AOI21_X1 U9262 ( .B1(n8136), .B2(n7303), .A(n7416), .ZN(n7417) );
  OAI21_X1 U9263 ( .B1(n7516), .B2(n8138), .A(n7417), .ZN(n7418) );
  AOI21_X1 U9264 ( .B1(n7419), .B2(n8141), .A(n7418), .ZN(n7420) );
  OAI211_X1 U9265 ( .C1(n9914), .C2(n8145), .A(n7421), .B(n7420), .ZN(P2_U3157) );
  XNOR2_X1 U9266 ( .A(n7422), .B(n7423), .ZN(n7424) );
  NAND2_X1 U9267 ( .A1(n7424), .A2(n7425), .ZN(n7481) );
  OAI21_X1 U9268 ( .B1(n7425), .B2(n7424), .A(n7481), .ZN(n7426) );
  NAND2_X1 U9269 ( .A1(n7426), .A2(n8876), .ZN(n7432) );
  NAND2_X1 U9270 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9407) );
  INV_X1 U9271 ( .A(n9407), .ZN(n7430) );
  INV_X1 U9272 ( .A(n7427), .ZN(n7428) );
  OAI22_X1 U9273 ( .A1(n8846), .A2(n7428), .B1(n9617), .B2(n8891), .ZN(n7429)
         );
  AOI211_X1 U9274 ( .C1(n8887), .C2(n8907), .A(n7430), .B(n7429), .ZN(n7431)
         );
  OAI211_X1 U9275 ( .C1(n9743), .C2(n8851), .A(n7432), .B(n7431), .ZN(P1_U3217) );
  INV_X1 U9276 ( .A(n8328), .ZN(n7438) );
  INV_X1 U9277 ( .A(n7433), .ZN(n7435) );
  NAND2_X1 U9278 ( .A1(n7435), .A2(n7434), .ZN(n7436) );
  OAI211_X1 U9279 ( .C1(n7438), .C2(n7437), .A(n7436), .B(n9861), .ZN(n7440)
         );
  AOI22_X1 U9280 ( .A1(n9858), .A2(n8386), .B1(n8384), .B2(n9859), .ZN(n7439)
         );
  NAND2_X1 U9281 ( .A1(n7440), .A2(n7439), .ZN(n9456) );
  INV_X1 U9282 ( .A(n7632), .ZN(n9455) );
  OAI22_X1 U9283 ( .A1(n9455), .A2(n7441), .B1(n7630), .B2(n8618), .ZN(n7442)
         );
  OAI21_X1 U9284 ( .B1(n9456), .B2(n7442), .A(n8608), .ZN(n7445) );
  XOR2_X1 U9285 ( .A(n8328), .B(n7443), .Z(n9458) );
  NAND2_X1 U9286 ( .A1(n9458), .A2(n9867), .ZN(n7444) );
  OAI211_X1 U9287 ( .C1(n7560), .C2(n8608), .A(n7445), .B(n7444), .ZN(P2_U3220) );
  INV_X1 U9288 ( .A(n7446), .ZN(n7450) );
  OAI222_X1 U9289 ( .A1(n7936), .A2(n7450), .B1(P2_U3151), .B2(n7448), .C1(
        n7447), .C2(n8751), .ZN(P2_U3270) );
  OAI222_X1 U9290 ( .A1(n7451), .A2(P1_U3086), .B1(n9395), .B2(n7450), .C1(
        n7449), .C2(n9392), .ZN(P1_U3330) );
  INV_X1 U9291 ( .A(n9920), .ZN(n7466) );
  OR2_X1 U9292 ( .A1(n7452), .A2(n8388), .ZN(n7453) );
  XNOR2_X1 U9293 ( .A(n9920), .B(n8024), .ZN(n7512) );
  XNOR2_X1 U9294 ( .A(n7512), .B(n7516), .ZN(n7456) );
  AOI21_X1 U9295 ( .B1(n7455), .B2(n7456), .A(n8132), .ZN(n7458) );
  INV_X1 U9296 ( .A(n7456), .ZN(n7457) );
  NAND2_X1 U9297 ( .A1(n7458), .A2(n7515), .ZN(n7465) );
  OR2_X1 U9298 ( .A1(n8138), .A2(n8210), .ZN(n7460) );
  INV_X1 U9299 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9276) );
  NOR2_X1 U9300 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9276), .ZN(n7500) );
  INV_X1 U9301 ( .A(n7500), .ZN(n7459) );
  OAI211_X1 U9302 ( .C1(n8095), .C2(n8197), .A(n7460), .B(n7459), .ZN(n7463)
         );
  NOR2_X1 U9303 ( .A1(n8075), .A2(n7461), .ZN(n7462) );
  NOR2_X1 U9304 ( .A1(n7463), .A2(n7462), .ZN(n7464) );
  OAI211_X1 U9305 ( .C1(n7466), .C2(n8145), .A(n7465), .B(n7464), .ZN(P2_U3176) );
  OAI21_X1 U9306 ( .B1(n7469), .B2(n7468), .A(n7467), .ZN(n7470) );
  NAND2_X1 U9307 ( .A1(n7470), .A2(n8876), .ZN(n7476) );
  NAND2_X1 U9308 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9557) );
  INV_X1 U9309 ( .A(n9557), .ZN(n7473) );
  OAI22_X1 U9310 ( .A1(n8846), .A2(n7471), .B1(n8892), .B2(n8867), .ZN(n7472)
         );
  AOI211_X1 U9311 ( .C1(n8878), .C2(n7474), .A(n7473), .B(n7472), .ZN(n7475)
         );
  OAI211_X1 U9312 ( .C1(n5500), .C2(n8851), .A(n7476), .B(n7475), .ZN(P1_U3234) );
  INV_X1 U9313 ( .A(n7477), .ZN(n7479) );
  OAI222_X1 U9314 ( .A1(n7936), .A2(n7479), .B1(P2_U3151), .B2(n6325), .C1(
        n7478), .C2(n8751), .ZN(P2_U3269) );
  OAI222_X1 U9315 ( .A1(n7480), .A2(P1_U3086), .B1(n9395), .B2(n7479), .C1(
        n9228), .C2(n9392), .ZN(P1_U3329) );
  OAI21_X1 U9316 ( .B1(n7422), .B2(n7482), .A(n7481), .ZN(n7486) );
  XOR2_X1 U9317 ( .A(n7484), .B(n7483), .Z(n7485) );
  XNOR2_X1 U9318 ( .A(n7486), .B(n7485), .ZN(n7487) );
  NAND2_X1 U9319 ( .A1(n7487), .A2(n8876), .ZN(n7494) );
  NAND2_X1 U9320 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9545) );
  INV_X1 U9321 ( .A(n9545), .ZN(n7492) );
  INV_X1 U9322 ( .A(n7488), .ZN(n7490) );
  OAI22_X1 U9323 ( .A1(n8846), .A2(n7490), .B1(n7489), .B2(n8867), .ZN(n7491)
         );
  AOI211_X1 U9324 ( .C1(n8878), .C2(n8908), .A(n7492), .B(n7491), .ZN(n7493)
         );
  OAI211_X1 U9325 ( .C1(n9749), .C2(n8851), .A(n7494), .B(n7493), .ZN(P1_U3236) );
  AOI21_X1 U9326 ( .B1(n9948), .B2(n7496), .A(n7495), .ZN(n7511) );
  AOI21_X1 U9327 ( .B1(n7499), .B2(n7498), .A(n7497), .ZN(n7502) );
  AOI21_X1 U9328 ( .B1(n9841), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7500), .ZN(
        n7501) );
  OAI21_X1 U9329 ( .B1(n7502), .B2(n9844), .A(n7501), .ZN(n7508) );
  AOI21_X1 U9330 ( .B1(n7505), .B2(n7504), .A(n7503), .ZN(n7506) );
  NOR2_X1 U9331 ( .A1(n7506), .A2(n9822), .ZN(n7507) );
  AOI211_X1 U9332 ( .C1(n9839), .C2(n7509), .A(n7508), .B(n7507), .ZN(n7510)
         );
  OAI21_X1 U9333 ( .B1(n7511), .B2(n8485), .A(n7510), .ZN(P2_U3193) );
  INV_X1 U9334 ( .A(n7512), .ZN(n7513) );
  NAND2_X1 U9335 ( .A1(n7513), .A2(n8387), .ZN(n7514) );
  NAND2_X1 U9336 ( .A1(n7515), .A2(n7514), .ZN(n7617) );
  XNOR2_X1 U9337 ( .A(n9930), .B(n8024), .ZN(n7618) );
  XNOR2_X1 U9338 ( .A(n7618), .B(n8386), .ZN(n7616) );
  XNOR2_X1 U9339 ( .A(n7617), .B(n7616), .ZN(n7522) );
  NAND2_X1 U9340 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .ZN(n7603) );
  OAI21_X1 U9341 ( .B1(n8095), .B2(n7516), .A(n7603), .ZN(n7517) );
  AOI21_X1 U9342 ( .B1(n8092), .B2(n8385), .A(n7517), .ZN(n7518) );
  OAI21_X1 U9343 ( .B1(n7519), .B2(n8075), .A(n7518), .ZN(n7520) );
  AOI21_X1 U9344 ( .B1(n9930), .B2(n8129), .A(n7520), .ZN(n7521) );
  OAI21_X1 U9345 ( .B1(n7522), .B2(n8132), .A(n7521), .ZN(P2_U3164) );
  NAND2_X1 U9346 ( .A1(n8219), .A2(n8218), .ZN(n8329) );
  XNOR2_X1 U9347 ( .A(n7523), .B(n8217), .ZN(n7539) );
  XNOR2_X1 U9348 ( .A(n7524), .B(n8217), .ZN(n7525) );
  NAND2_X1 U9349 ( .A1(n7525), .A2(n9861), .ZN(n7527) );
  AOI22_X1 U9350 ( .A1(n9858), .A2(n8385), .B1(n8383), .B2(n9859), .ZN(n7526)
         );
  MUX2_X1 U9351 ( .A(n7528), .B(n7534), .S(n9952), .Z(n7530) );
  NAND2_X1 U9352 ( .A1(n7990), .A2(n8658), .ZN(n7529) );
  OAI211_X1 U9353 ( .C1(n7539), .C2(n8673), .A(n7530), .B(n7529), .ZN(P2_U3473) );
  INV_X1 U9354 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7531) );
  MUX2_X1 U9355 ( .A(n7531), .B(n7534), .S(n9932), .Z(n7533) );
  NAND2_X1 U9356 ( .A1(n7990), .A2(n8725), .ZN(n7532) );
  OAI211_X1 U9357 ( .C1(n7539), .C2(n8738), .A(n7533), .B(n7532), .ZN(P2_U3432) );
  MUX2_X1 U9358 ( .A(n7535), .B(n7534), .S(n8608), .Z(n7538) );
  INV_X1 U9359 ( .A(n7536), .ZN(n8001) );
  AOI22_X1 U9360 ( .A1(n7990), .A2(n9864), .B1(n9865), .B2(n8001), .ZN(n7537)
         );
  OAI211_X1 U9361 ( .C1(n7539), .C2(n8615), .A(n7538), .B(n7537), .ZN(P2_U3219) );
  INV_X1 U9362 ( .A(n7540), .ZN(n7924) );
  OAI222_X1 U9363 ( .A1(n7936), .A2(n7924), .B1(n7542), .B2(P2_U3151), .C1(
        n7541), .C2(n8751), .ZN(P2_U3268) );
  XNOR2_X1 U9364 ( .A(n7545), .B(n8221), .ZN(n7557) );
  INV_X1 U9365 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7548) );
  XNOR2_X1 U9366 ( .A(n7546), .B(n8221), .ZN(n7547) );
  AOI222_X1 U9367 ( .A1(n9861), .A2(n7547), .B1(n8626), .B2(n9859), .C1(n8384), 
        .C2(n9858), .ZN(n7553) );
  MUX2_X1 U9368 ( .A(n7548), .B(n7553), .S(n9932), .Z(n7550) );
  NAND2_X1 U9369 ( .A1(n8225), .A2(n8725), .ZN(n7549) );
  OAI211_X1 U9370 ( .C1(n7557), .C2(n8738), .A(n7550), .B(n7549), .ZN(P2_U3435) );
  MUX2_X1 U9371 ( .A(n8424), .B(n7553), .S(n9952), .Z(n7552) );
  NAND2_X1 U9372 ( .A1(n8225), .A2(n8658), .ZN(n7551) );
  OAI211_X1 U9373 ( .C1(n8673), .C2(n7557), .A(n7552), .B(n7551), .ZN(P2_U3474) );
  MUX2_X1 U9374 ( .A(n8416), .B(n7553), .S(n8608), .Z(n7556) );
  INV_X1 U9375 ( .A(n7554), .ZN(n8142) );
  AOI22_X1 U9376 ( .A1(n8225), .A2(n9864), .B1(n9865), .B2(n8142), .ZN(n7555)
         );
  OAI211_X1 U9377 ( .C1(n7557), .C2(n8615), .A(n7556), .B(n7555), .ZN(P2_U3218) );
  AOI21_X1 U9378 ( .B1(n7560), .B2(n7559), .A(n7558), .ZN(n7574) );
  NAND2_X1 U9379 ( .A1(n9839), .A2(n7561), .ZN(n7572) );
  AND2_X1 U9380 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7628) );
  AOI21_X1 U9381 ( .B1(n9841), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7628), .ZN(
        n7571) );
  OAI21_X1 U9382 ( .B1(n7564), .B2(n7563), .A(n7562), .ZN(n7565) );
  NAND2_X1 U9383 ( .A1(n7565), .A2(n9827), .ZN(n7570) );
  AOI21_X1 U9384 ( .B1(n7567), .B2(n9459), .A(n7566), .ZN(n7568) );
  OR2_X1 U9385 ( .A1(n8485), .A2(n7568), .ZN(n7569) );
  OAI21_X1 U9386 ( .B1(n7574), .B2(n9822), .A(n7573), .ZN(P2_U3195) );
  XNOR2_X1 U9387 ( .A(n7575), .B(n8335), .ZN(n7590) );
  NAND2_X1 U9388 ( .A1(n7576), .A2(n8335), .ZN(n7577) );
  NAND3_X1 U9389 ( .A1(n8623), .A2(n9861), .A3(n7577), .ZN(n7579) );
  AOI22_X1 U9390 ( .A1(n8382), .A2(n9859), .B1(n9858), .B2(n8383), .ZN(n7578)
         );
  INV_X1 U9391 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7580) );
  MUX2_X1 U9392 ( .A(n7587), .B(n7580), .S(n9934), .Z(n7582) );
  NAND2_X1 U9393 ( .A1(n8053), .A2(n8725), .ZN(n7581) );
  OAI211_X1 U9394 ( .C1(n7590), .C2(n8738), .A(n7582), .B(n7581), .ZN(P2_U3438) );
  MUX2_X1 U9395 ( .A(n7583), .B(n7587), .S(n9952), .Z(n7585) );
  NAND2_X1 U9396 ( .A1(n8053), .A2(n8658), .ZN(n7584) );
  OAI211_X1 U9397 ( .C1(n7590), .C2(n8673), .A(n7585), .B(n7584), .ZN(P2_U3475) );
  MUX2_X1 U9398 ( .A(n7587), .B(n7586), .S(n9870), .Z(n7589) );
  AOI22_X1 U9399 ( .A1(n8053), .A2(n9864), .B1(n9865), .B2(n8063), .ZN(n7588)
         );
  OAI211_X1 U9400 ( .C1(n7590), .C2(n8615), .A(n7589), .B(n7588), .ZN(P2_U3217) );
  INV_X1 U9401 ( .A(n7591), .ZN(n7615) );
  OAI222_X1 U9402 ( .A1(n7936), .A2(n7615), .B1(n8370), .B2(P2_U3151), .C1(
        n7592), .C2(n8751), .ZN(P2_U3267) );
  AOI21_X1 U9403 ( .B1(n4357), .B2(n7594), .A(n7593), .ZN(n7613) );
  INV_X1 U9404 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7604) );
  INV_X1 U9405 ( .A(n7595), .ZN(n7597) );
  NOR2_X1 U9406 ( .A1(n7597), .A2(n7596), .ZN(n7599) );
  OAI21_X1 U9407 ( .B1(n7600), .B2(n7599), .A(n9827), .ZN(n7598) );
  AOI21_X1 U9408 ( .B1(n7600), .B2(n7599), .A(n7598), .ZN(n7601) );
  INV_X1 U9409 ( .A(n7601), .ZN(n7602) );
  OAI211_X1 U9410 ( .C1(n9831), .C2(n7604), .A(n7603), .B(n7602), .ZN(n7610)
         );
  AOI21_X1 U9411 ( .B1(n7607), .B2(n7606), .A(n7605), .ZN(n7608) );
  NOR2_X1 U9412 ( .A1(n7608), .A2(n8485), .ZN(n7609) );
  AOI211_X1 U9413 ( .C1(n9839), .C2(n7611), .A(n7610), .B(n7609), .ZN(n7612)
         );
  OAI21_X1 U9414 ( .B1(n7613), .B2(n9822), .A(n7612), .ZN(P2_U3194) );
  OAI222_X1 U9415 ( .A1(P1_U3086), .A2(n5417), .B1(n9395), .B2(n7615), .C1(
        n7614), .C2(n9392), .ZN(P1_U3327) );
  INV_X1 U9416 ( .A(n7618), .ZN(n7619) );
  NAND2_X1 U9417 ( .A1(n7619), .A2(n8386), .ZN(n7620) );
  XNOR2_X1 U9418 ( .A(n7632), .B(n8024), .ZN(n7621) );
  NAND2_X1 U9419 ( .A1(n7621), .A2(n7999), .ZN(n7991) );
  INV_X1 U9420 ( .A(n7621), .ZN(n7622) );
  NAND2_X1 U9421 ( .A1(n7622), .A2(n8385), .ZN(n7623) );
  NAND2_X1 U9422 ( .A1(n7991), .A2(n7623), .ZN(n7625) );
  INV_X1 U9423 ( .A(n7937), .ZN(n7994) );
  AOI21_X1 U9424 ( .B1(n7626), .B2(n7625), .A(n7994), .ZN(n7634) );
  NOR2_X1 U9425 ( .A1(n8095), .A2(n8210), .ZN(n7627) );
  AOI211_X1 U9426 ( .C1(n8092), .C2(n8384), .A(n7628), .B(n7627), .ZN(n7629)
         );
  OAI21_X1 U9427 ( .B1(n7630), .B2(n8075), .A(n7629), .ZN(n7631) );
  AOI21_X1 U9428 ( .B1(n7632), .B2(n8129), .A(n7631), .ZN(n7633) );
  OAI21_X1 U9429 ( .B1(n7634), .B2(n8132), .A(n7633), .ZN(P2_U3174) );
  NAND2_X1 U9430 ( .A1(n7636), .A2(n7635), .ZN(n7717) );
  INV_X1 U9431 ( .A(n7717), .ZN(n7814) );
  OR2_X1 U9432 ( .A1(n9168), .A2(n7637), .ZN(n7797) );
  OAI21_X1 U9433 ( .B1(n7797), .B2(n7888), .A(n7798), .ZN(n7714) );
  NAND3_X1 U9434 ( .A1(n9168), .A2(n7637), .A3(n7888), .ZN(n7638) );
  OAI211_X1 U9435 ( .C1(n7814), .C2(n7753), .A(n7795), .B(n7638), .ZN(n7713)
         );
  INV_X1 U9436 ( .A(n7640), .ZN(n7641) );
  INV_X1 U9437 ( .A(n7645), .ZN(n7642) );
  INV_X1 U9438 ( .A(n7655), .ZN(n7647) );
  AOI21_X1 U9439 ( .B1(n7654), .B2(n7648), .A(n7647), .ZN(n7650) );
  NAND2_X1 U9440 ( .A1(n7848), .A2(n7845), .ZN(n7649) );
  NAND2_X1 U9441 ( .A1(n7656), .A2(n7655), .ZN(n7849) );
  AOI21_X1 U9442 ( .B1(n7657), .B2(n7845), .A(n7849), .ZN(n7660) );
  NAND2_X1 U9443 ( .A1(n7658), .A2(n7848), .ZN(n7659) );
  NAND2_X1 U9444 ( .A1(n7661), .A2(n7666), .ZN(n7854) );
  AOI21_X1 U9445 ( .B1(n7667), .B2(n7662), .A(n7854), .ZN(n7664) );
  NAND3_X1 U9446 ( .A1(n7671), .A2(n7669), .A3(n7663), .ZN(n7831) );
  OAI21_X1 U9447 ( .B1(n7664), .B2(n7831), .A(n7858), .ZN(n7673) );
  OR2_X1 U9448 ( .A1(n8895), .A2(n7888), .ZN(n7668) );
  NAND2_X1 U9449 ( .A1(n7669), .A2(n7668), .ZN(n7674) );
  OAI21_X1 U9450 ( .B1(n7670), .B2(n7674), .A(n7858), .ZN(n7672) );
  INV_X1 U9451 ( .A(n7674), .ZN(n7675) );
  NOR3_X1 U9452 ( .A1(n9141), .A2(n8809), .A3(n7675), .ZN(n7676) );
  INV_X1 U9453 ( .A(n9140), .ZN(n9130) );
  INV_X1 U9454 ( .A(n7682), .ZN(n7678) );
  NAND2_X1 U9455 ( .A1(n7681), .A2(n7677), .ZN(n7860) );
  OAI211_X1 U9456 ( .C1(n7678), .C2(n7860), .A(n7867), .B(n7680), .ZN(n7686)
         );
  AND2_X1 U9457 ( .A1(n7680), .A2(n7679), .ZN(n7864) );
  NAND2_X1 U9458 ( .A1(n7688), .A2(n7681), .ZN(n7868) );
  INV_X1 U9459 ( .A(n7687), .ZN(n9070) );
  INV_X1 U9460 ( .A(n7688), .ZN(n7689) );
  OAI21_X1 U9461 ( .B1(n9070), .B2(n7689), .A(n7753), .ZN(n7693) );
  OR2_X1 U9462 ( .A1(n7697), .A2(n7690), .ZN(n7691) );
  MUX2_X1 U9463 ( .A(n7804), .B(n7691), .S(n7753), .Z(n7692) );
  INV_X1 U9464 ( .A(n7695), .ZN(n7696) );
  MUX2_X1 U9465 ( .A(n7697), .B(n7696), .S(n7753), .Z(n7698) );
  INV_X1 U9466 ( .A(n9062), .ZN(n7786) );
  INV_X1 U9467 ( .A(n7700), .ZN(n7701) );
  NAND2_X1 U9468 ( .A1(n7705), .A2(n7701), .ZN(n7702) );
  NAND2_X1 U9469 ( .A1(n7702), .A2(n7704), .ZN(n7800) );
  NAND2_X1 U9470 ( .A1(n9188), .A2(n9074), .ZN(n7703) );
  NAND2_X1 U9471 ( .A1(n7704), .A2(n7703), .ZN(n7806) );
  NAND2_X1 U9472 ( .A1(n7806), .A2(n7705), .ZN(n7706) );
  MUX2_X1 U9473 ( .A(n7800), .B(n7706), .S(n7888), .Z(n7707) );
  INV_X1 U9474 ( .A(n7809), .ZN(n7709) );
  MUX2_X1 U9475 ( .A(n7710), .B(n7709), .S(n7888), .Z(n7711) );
  NAND3_X1 U9476 ( .A1(n7870), .A2(n7753), .A3(n7810), .ZN(n7712) );
  NAND2_X1 U9477 ( .A1(n7715), .A2(n7810), .ZN(n7716) );
  NAND4_X1 U9478 ( .A1(n7716), .A2(n7797), .A3(n7803), .A4(n7888), .ZN(n7719)
         );
  OAI21_X1 U9479 ( .B1(n7717), .B2(n7798), .A(n7795), .ZN(n7718) );
  AOI22_X1 U9480 ( .A1(n7720), .A2(n7719), .B1(n7888), .B2(n7718), .ZN(n7737)
         );
  NAND2_X1 U9481 ( .A1(n7722), .A2(n7721), .ZN(n7723) );
  INV_X1 U9482 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8281) );
  INV_X1 U9483 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9390) );
  MUX2_X1 U9484 ( .A(n8281), .B(n9390), .S(n7725), .Z(n7727) );
  INV_X1 U9485 ( .A(SI_30_), .ZN(n7726) );
  NAND2_X1 U9486 ( .A1(n7727), .A2(n7726), .ZN(n7744) );
  INV_X1 U9487 ( .A(n7727), .ZN(n7728) );
  NAND2_X1 U9488 ( .A1(n7728), .A2(SI_30_), .ZN(n7729) );
  OR2_X1 U9489 ( .A1(n7751), .A2(n9390), .ZN(n7730) );
  INV_X1 U9490 ( .A(n8899), .ZN(n7739) );
  NOR2_X1 U9491 ( .A1(n8978), .A2(n7739), .ZN(n7880) );
  NAND2_X1 U9492 ( .A1(n7731), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U9493 ( .A1(n7732), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U9494 ( .A1(n7733), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7734) );
  NAND3_X1 U9495 ( .A1(n7736), .A2(n7735), .A3(n7734), .ZN(n8972) );
  INV_X1 U9496 ( .A(n7818), .ZN(n7877) );
  INV_X1 U9497 ( .A(n7796), .ZN(n7738) );
  MUX2_X1 U9498 ( .A(n7877), .B(n7738), .S(n7888), .Z(n7741) );
  NAND2_X1 U9499 ( .A1(n8978), .A2(n7739), .ZN(n7881) );
  INV_X1 U9500 ( .A(n8972), .ZN(n7756) );
  NAND2_X1 U9501 ( .A1(n8978), .A2(n7756), .ZN(n7740) );
  NAND2_X1 U9502 ( .A1(n7881), .A2(n7740), .ZN(n7821) );
  NAND2_X1 U9503 ( .A1(n7743), .A2(n7742), .ZN(n7745) );
  NAND2_X1 U9504 ( .A1(n7745), .A2(n7744), .ZN(n7749) );
  INV_X1 U9505 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8744) );
  INV_X1 U9506 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7750) );
  MUX2_X1 U9507 ( .A(n8744), .B(n7750), .S(n7746), .Z(n7747) );
  XNOR2_X1 U9508 ( .A(n7747), .B(SI_31_), .ZN(n7748) );
  NOR2_X1 U9509 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  AND2_X1 U9510 ( .A1(n9154), .A2(n8972), .ZN(n7891) );
  INV_X1 U9511 ( .A(n7820), .ZN(n7754) );
  INV_X1 U9512 ( .A(n9154), .ZN(n8969) );
  NAND2_X1 U9513 ( .A1(n8969), .A2(n7756), .ZN(n7887) );
  AOI21_X1 U9514 ( .B1(n7758), .B2(n7887), .A(n7757), .ZN(n7759) );
  AOI21_X1 U9515 ( .B1(n9027), .B2(n7837), .A(n7759), .ZN(n7828) );
  INV_X1 U9516 ( .A(n7880), .ZN(n7760) );
  AND2_X1 U9517 ( .A1(n7760), .A2(n7881), .ZN(n7794) );
  INV_X1 U9518 ( .A(n7761), .ZN(n7790) );
  XNOR2_X1 U9519 ( .A(n9194), .B(n9090), .ZN(n9071) );
  XNOR2_X1 U9520 ( .A(n9199), .B(n8901), .ZN(n9086) );
  NOR2_X1 U9521 ( .A1(n6903), .A2(n7763), .ZN(n7767) );
  INV_X1 U9522 ( .A(n7764), .ZN(n7765) );
  NAND4_X1 U9523 ( .A1(n7767), .A2(n7766), .A3(n7765), .A4(n7837), .ZN(n7770)
         );
  NOR4_X1 U9524 ( .A1(n7770), .A2(n4598), .A3(n7769), .A4(n9663), .ZN(n7771)
         );
  AND4_X1 U9525 ( .A1(n7773), .A2(n7844), .A3(n7772), .A4(n7771), .ZN(n7774)
         );
  NAND4_X1 U9526 ( .A1(n7777), .A2(n7776), .A3(n7775), .A4(n7774), .ZN(n7778)
         );
  NOR2_X1 U9527 ( .A1(n7779), .A2(n7778), .ZN(n7780) );
  NAND3_X1 U9528 ( .A1(n7782), .A2(n7781), .A3(n7780), .ZN(n7783) );
  NOR2_X1 U9529 ( .A1(n9140), .A2(n7783), .ZN(n7784) );
  NAND4_X1 U9530 ( .A1(n9086), .A2(n9109), .A3(n9122), .A4(n7784), .ZN(n7785)
         );
  NOR2_X1 U9531 ( .A1(n9071), .A2(n7785), .ZN(n7787) );
  NAND4_X1 U9532 ( .A1(n4617), .A2(n9046), .A3(n7787), .A4(n7786), .ZN(n7788)
         );
  NOR2_X1 U9533 ( .A1(n7788), .A2(n9017), .ZN(n7789) );
  NAND4_X1 U9534 ( .A1(n7790), .A2(n8984), .A3(n7789), .A4(n9003), .ZN(n7791)
         );
  NOR2_X1 U9535 ( .A1(n7792), .A2(n7791), .ZN(n7793) );
  AND4_X1 U9536 ( .A1(n4498), .A2(n7887), .A3(n7794), .A4(n7793), .ZN(n7827)
         );
  NAND2_X1 U9537 ( .A1(n7796), .A2(n7795), .ZN(n7829) );
  NAND2_X1 U9538 ( .A1(n7798), .A2(n7797), .ZN(n7875) );
  INV_X1 U9539 ( .A(n7875), .ZN(n7817) );
  NAND2_X1 U9540 ( .A1(n7800), .A2(n7799), .ZN(n7801) );
  NAND2_X1 U9541 ( .A1(n7801), .A2(n7809), .ZN(n7802) );
  AND2_X1 U9542 ( .A1(n7803), .A2(n7802), .ZN(n7813) );
  INV_X1 U9543 ( .A(n7813), .ZN(n7805) );
  OR2_X1 U9544 ( .A1(n7805), .A2(n7804), .ZN(n7830) );
  OAI21_X1 U9545 ( .B1(n9087), .B2(n7830), .A(n7870), .ZN(n7816) );
  INV_X1 U9546 ( .A(n7806), .ZN(n7808) );
  NAND3_X1 U9547 ( .A1(n7809), .A2(n7808), .A3(n7807), .ZN(n7812) );
  INV_X1 U9548 ( .A(n7810), .ZN(n7811) );
  AOI21_X1 U9549 ( .B1(n7813), .B2(n7812), .A(n7811), .ZN(n7815) );
  OAI21_X1 U9550 ( .B1(n7815), .B2(n7875), .A(n7814), .ZN(n7873) );
  AOI21_X1 U9551 ( .B1(n7817), .B2(n7816), .A(n7873), .ZN(n7819) );
  OAI21_X1 U9552 ( .B1(n7829), .B2(n7819), .A(n7818), .ZN(n7822) );
  OAI21_X1 U9553 ( .B1(n7822), .B2(n7821), .A(n7820), .ZN(n7824) );
  AOI211_X1 U9554 ( .C1(n4498), .C2(n7824), .A(n7823), .B(n4631), .ZN(n7825)
         );
  OAI21_X1 U9555 ( .B1(n7825), .B2(n7827), .A(n7928), .ZN(n7826) );
  OAI21_X1 U9556 ( .B1(n7828), .B2(n7827), .A(n7826), .ZN(n7894) );
  NOR2_X1 U9557 ( .A1(n7928), .A2(n7895), .ZN(n7885) );
  INV_X1 U9558 ( .A(n7829), .ZN(n7879) );
  INV_X1 U9559 ( .A(n7830), .ZN(n7872) );
  INV_X1 U9560 ( .A(n7831), .ZN(n7863) );
  INV_X1 U9561 ( .A(n7832), .ZN(n7833) );
  OAI21_X1 U9562 ( .B1(n7835), .B2(n7834), .A(n7833), .ZN(n7836) );
  AOI211_X1 U9563 ( .C1(n9683), .C2(n5732), .A(n7837), .B(n7836), .ZN(n7841)
         );
  AND4_X1 U9564 ( .A1(n7841), .A2(n7840), .A3(n7839), .A4(n7838), .ZN(n7843)
         );
  AOI21_X1 U9565 ( .B1(n7844), .B2(n7843), .A(n7842), .ZN(n7847) );
  INV_X1 U9566 ( .A(n7845), .ZN(n7846) );
  NOR2_X1 U9567 ( .A1(n7847), .A2(n7846), .ZN(n7850) );
  OAI21_X1 U9568 ( .B1(n7850), .B2(n7849), .A(n7848), .ZN(n7853) );
  AOI21_X1 U9569 ( .B1(n7853), .B2(n7852), .A(n7851), .ZN(n7857) );
  INV_X1 U9570 ( .A(n7854), .ZN(n7855) );
  OAI21_X1 U9571 ( .B1(n7857), .B2(n7856), .A(n7855), .ZN(n7862) );
  AOI21_X1 U9572 ( .B1(n7859), .B2(n7858), .A(n9141), .ZN(n7861) );
  AOI211_X1 U9573 ( .C1(n7863), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7866)
         );
  INV_X1 U9574 ( .A(n7864), .ZN(n7865) );
  NOR2_X1 U9575 ( .A1(n7866), .A2(n7865), .ZN(n7869) );
  OAI21_X1 U9576 ( .B1(n7869), .B2(n7868), .A(n7867), .ZN(n7871) );
  AOI21_X1 U9577 ( .B1(n7872), .B2(n7871), .A(n4704), .ZN(n7876) );
  INV_X1 U9578 ( .A(n7873), .ZN(n7874) );
  OAI21_X1 U9579 ( .B1(n7876), .B2(n7875), .A(n7874), .ZN(n7878) );
  AOI21_X1 U9580 ( .B1(n7879), .B2(n7878), .A(n7877), .ZN(n7882) );
  AOI21_X1 U9581 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7883) );
  AOI21_X1 U9582 ( .B1(n7883), .B2(n7887), .A(n7891), .ZN(n7884) );
  MUX2_X1 U9583 ( .A(n7886), .B(n7885), .S(n7884), .Z(n7893) );
  AOI211_X1 U9584 ( .C1(n7895), .C2(n7894), .A(n7893), .B(n7892), .ZN(n7902)
         );
  NOR3_X1 U9585 ( .A1(n7897), .A2(n7896), .A3(n9476), .ZN(n7900) );
  OAI21_X1 U9586 ( .B1(n7901), .B2(n7898), .A(P1_B_REG_SCAN_IN), .ZN(n7899) );
  OAI22_X1 U9587 ( .A1(n7902), .A2(n7901), .B1(n7900), .B2(n7899), .ZN(
        P1_U3242) );
  NAND2_X1 U9588 ( .A1(n7903), .A2(n9670), .ZN(n7910) );
  AOI22_X1 U9589 ( .A1(n9658), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n7904), .B2(
        n9656), .ZN(n7905) );
  OAI21_X1 U9590 ( .B1(n8968), .B2(n9660), .A(n7905), .ZN(n7906) );
  AOI21_X1 U9591 ( .B1(n7908), .B2(n7907), .A(n7906), .ZN(n7909) );
  OAI211_X1 U9592 ( .C1(n7911), .C2(n9658), .A(n7910), .B(n7909), .ZN(P1_U3356) );
  XNOR2_X1 U9593 ( .A(n8389), .B(n7912), .ZN(n7913) );
  XNOR2_X1 U9594 ( .A(n7914), .B(n7913), .ZN(n7915) );
  NAND2_X1 U9595 ( .A1(n7915), .A2(n8116), .ZN(n7923) );
  OR2_X1 U9596 ( .A1(n8138), .A2(n7916), .ZN(n7918) );
  OAI211_X1 U9597 ( .C1(n8095), .C2(n7919), .A(n7918), .B(n7917), .ZN(n7921)
         );
  NOR2_X1 U9598 ( .A1(n8075), .A2(n4857), .ZN(n7920) );
  NOR2_X1 U9599 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  OAI211_X1 U9600 ( .C1(n7310), .C2(n8145), .A(n7923), .B(n7922), .ZN(P2_U3161) );
  OAI222_X1 U9601 ( .A1(n9392), .A2(n7925), .B1(P1_U3086), .B2(n9474), .C1(
        n7924), .C2(n9395), .ZN(P1_U3328) );
  OAI222_X1 U9602 ( .A1(n7928), .A2(P1_U3086), .B1(n9395), .B2(n7927), .C1(
        n7926), .C2(n9392), .ZN(P1_U3336) );
  AOI22_X1 U9603 ( .A1(n8487), .A2(n9865), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9870), .ZN(n7930) );
  NAND2_X1 U9604 ( .A1(n6414), .A2(n9864), .ZN(n7929) );
  OAI211_X1 U9605 ( .C1(n6430), .C2(n7931), .A(n7930), .B(n7929), .ZN(n7932)
         );
  INV_X1 U9606 ( .A(n7932), .ZN(n7933) );
  OAI21_X1 U9607 ( .B1(n7934), .B2(n9870), .A(n7933), .ZN(P2_U3204) );
  INV_X1 U9608 ( .A(n8280), .ZN(n9391) );
  OAI222_X1 U9609 ( .A1(n7936), .A2(n9391), .B1(n5979), .B2(P2_U3151), .C1(
        n8281), .C2(n8751), .ZN(P2_U3265) );
  NAND2_X1 U9610 ( .A1(n7937), .A2(n7991), .ZN(n7938) );
  XNOR2_X1 U9611 ( .A(n7990), .B(n8024), .ZN(n7940) );
  XNOR2_X1 U9612 ( .A(n7940), .B(n8384), .ZN(n7992) );
  NAND2_X1 U9613 ( .A1(n7940), .A2(n7939), .ZN(n7941) );
  XNOR2_X1 U9614 ( .A(n8225), .B(n8024), .ZN(n7945) );
  XNOR2_X1 U9615 ( .A(n7945), .B(n8224), .ZN(n8133) );
  XNOR2_X1 U9616 ( .A(n8053), .B(n8024), .ZN(n7942) );
  NAND2_X1 U9617 ( .A1(n7942), .A2(n8139), .ZN(n8068) );
  INV_X1 U9618 ( .A(n7942), .ZN(n7943) );
  NAND2_X1 U9619 ( .A1(n7943), .A2(n8626), .ZN(n7944) );
  NAND2_X1 U9620 ( .A1(n8068), .A2(n7944), .ZN(n8057) );
  INV_X1 U9621 ( .A(n7945), .ZN(n7946) );
  AND2_X1 U9622 ( .A1(n7946), .A2(n8383), .ZN(n8056) );
  NOR2_X1 U9623 ( .A1(n8057), .A2(n8056), .ZN(n7947) );
  NAND2_X1 U9624 ( .A1(n8055), .A2(n7947), .ZN(n8054) );
  NAND2_X1 U9625 ( .A1(n8054), .A2(n8068), .ZN(n7951) );
  XNOR2_X1 U9626 ( .A(n8067), .B(n8024), .ZN(n7948) );
  NAND2_X1 U9627 ( .A1(n7948), .A2(n8604), .ZN(n8111) );
  INV_X1 U9628 ( .A(n7948), .ZN(n7949) );
  NAND2_X1 U9629 ( .A1(n7949), .A2(n8382), .ZN(n7950) );
  AND2_X1 U9630 ( .A1(n8111), .A2(n7950), .ZN(n8069) );
  NAND2_X1 U9631 ( .A1(n7951), .A2(n8069), .ZN(n8072) );
  NAND2_X1 U9632 ( .A1(n8072), .A2(n8111), .ZN(n7952) );
  XNOR2_X1 U9633 ( .A(n8668), .B(n8024), .ZN(n7953) );
  XNOR2_X1 U9634 ( .A(n7953), .B(n8625), .ZN(n8112) );
  NAND2_X1 U9635 ( .A1(n7952), .A2(n8112), .ZN(n8115) );
  NAND2_X1 U9636 ( .A1(n7953), .A2(n8074), .ZN(n7954) );
  XNOR2_X1 U9637 ( .A(n8661), .B(n8024), .ZN(n7958) );
  AND2_X1 U9638 ( .A1(n7958), .A2(n8606), .ZN(n8087) );
  XNOR2_X1 U9639 ( .A(n7955), .B(n8024), .ZN(n7960) );
  INV_X1 U9640 ( .A(n7960), .ZN(n7956) );
  AND2_X1 U9641 ( .A1(n7956), .A2(n8042), .ZN(n7963) );
  OR2_X1 U9642 ( .A1(n8087), .A2(n7963), .ZN(n8035) );
  XNOR2_X1 U9643 ( .A(n8719), .B(n8024), .ZN(n7964) );
  AND2_X1 U9644 ( .A1(n7964), .A2(n7957), .ZN(n7966) );
  OR2_X1 U9645 ( .A1(n8035), .A2(n7966), .ZN(n8099) );
  XNOR2_X1 U9646 ( .A(n8713), .B(n8024), .ZN(n7968) );
  XNOR2_X1 U9647 ( .A(n7968), .B(n8542), .ZN(n8102) );
  INV_X1 U9648 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U9649 ( .A1(n7959), .A2(n8582), .ZN(n8088) );
  XNOR2_X1 U9650 ( .A(n7960), .B(n8589), .ZN(n8091) );
  INV_X1 U9651 ( .A(n8091), .ZN(n7961) );
  AND2_X1 U9652 ( .A1(n8088), .A2(n7961), .ZN(n7962) );
  OR2_X1 U9653 ( .A1(n7963), .A2(n7962), .ZN(n8036) );
  XNOR2_X1 U9654 ( .A(n7964), .B(n8581), .ZN(n8039) );
  AND2_X1 U9655 ( .A1(n8036), .A2(n8039), .ZN(n7965) );
  OR2_X1 U9656 ( .A1(n7966), .A2(n7965), .ZN(n8100) );
  OR2_X1 U9657 ( .A1(n8102), .A2(n8100), .ZN(n7967) );
  INV_X1 U9658 ( .A(n7968), .ZN(n7969) );
  XNOR2_X1 U9659 ( .A(n8707), .B(n8024), .ZN(n7971) );
  XNOR2_X1 U9660 ( .A(n8702), .B(n8024), .ZN(n7975) );
  XNOR2_X1 U9661 ( .A(n7975), .B(n8519), .ZN(n8081) );
  XNOR2_X1 U9662 ( .A(n7977), .B(n8024), .ZN(n7978) );
  XNOR2_X1 U9663 ( .A(n7978), .B(n8381), .ZN(n8047) );
  XNOR2_X1 U9664 ( .A(n8512), .B(n8024), .ZN(n7980) );
  XNOR2_X1 U9665 ( .A(n7980), .B(n8518), .ZN(n8125) );
  XNOR2_X1 U9666 ( .A(n8271), .B(n6863), .ZN(n7982) );
  NOR2_X1 U9667 ( .A1(n7982), .A2(n8508), .ZN(n8021) );
  AOI21_X1 U9668 ( .B1(n8508), .B2(n7982), .A(n8021), .ZN(n7984) );
  OAI211_X1 U9669 ( .C1(n7983), .C2(n7984), .A(n8023), .B(n8116), .ZN(n7989)
         );
  INV_X1 U9670 ( .A(n8501), .ZN(n7986) );
  AOI22_X1 U9671 ( .A1(n8518), .A2(n8136), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7985) );
  OAI21_X1 U9672 ( .B1(n7986), .B2(n8075), .A(n7985), .ZN(n7987) );
  AOI21_X1 U9673 ( .B1(n8092), .B2(n8498), .A(n7987), .ZN(n7988) );
  OAI211_X1 U9674 ( .C1(n8271), .C2(n8145), .A(n7989), .B(n7988), .ZN(P2_U3154) );
  INV_X1 U9675 ( .A(n7990), .ZN(n8004) );
  INV_X1 U9676 ( .A(n7991), .ZN(n7993) );
  NOR3_X1 U9677 ( .A1(n7994), .A2(n7993), .A3(n7992), .ZN(n7997) );
  INV_X1 U9678 ( .A(n7995), .ZN(n7996) );
  OAI21_X1 U9679 ( .B1(n7997), .B2(n7996), .A(n8116), .ZN(n8003) );
  INV_X1 U9680 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9301) );
  NOR2_X1 U9681 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9301), .ZN(n8401) );
  AOI21_X1 U9682 ( .B1(n8092), .B2(n8383), .A(n8401), .ZN(n7998) );
  OAI21_X1 U9683 ( .B1(n7999), .B2(n8095), .A(n7998), .ZN(n8000) );
  AOI21_X1 U9684 ( .B1(n8001), .B2(n8141), .A(n8000), .ZN(n8002) );
  OAI211_X1 U9685 ( .C1(n8004), .C2(n8145), .A(n8003), .B(n8002), .ZN(P2_U3155) );
  XNOR2_X1 U9686 ( .A(n8005), .B(n8532), .ZN(n8010) );
  AOI22_X1 U9687 ( .A1(n8567), .A2(n8136), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8007) );
  NAND2_X1 U9688 ( .A1(n8141), .A2(n8545), .ZN(n8006) );
  OAI211_X1 U9689 ( .C1(n8541), .C2(n8138), .A(n8007), .B(n8006), .ZN(n8008)
         );
  AOI21_X1 U9690 ( .B1(n8546), .B2(n8129), .A(n8008), .ZN(n8009) );
  OAI21_X1 U9691 ( .B1(n8010), .B2(n8132), .A(n8009), .ZN(P2_U3156) );
  INV_X1 U9692 ( .A(n8087), .ZN(n8012) );
  NAND2_X1 U9693 ( .A1(n8012), .A2(n8088), .ZN(n8013) );
  XNOR2_X1 U9694 ( .A(n8011), .B(n8013), .ZN(n8020) );
  INV_X1 U9695 ( .A(n8014), .ZN(n8591) );
  OAI21_X1 U9696 ( .B1(n8095), .B2(n8074), .A(n8015), .ZN(n8016) );
  AOI21_X1 U9697 ( .B1(n8092), .B2(n8589), .A(n8016), .ZN(n8017) );
  OAI21_X1 U9698 ( .B1(n8591), .B2(n8075), .A(n8017), .ZN(n8018) );
  AOI21_X1 U9699 ( .B1(n8661), .B2(n8129), .A(n8018), .ZN(n8019) );
  OAI21_X1 U9700 ( .B1(n8020), .B2(n8132), .A(n8019), .ZN(P2_U3159) );
  INV_X1 U9701 ( .A(n8021), .ZN(n8022) );
  NAND2_X1 U9702 ( .A1(n8023), .A2(n8022), .ZN(n8026) );
  XNOR2_X1 U9703 ( .A(n8308), .B(n8024), .ZN(n8025) );
  XNOR2_X1 U9704 ( .A(n8026), .B(n8025), .ZN(n8034) );
  OAI22_X1 U9705 ( .A1(n8508), .A2(n8095), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8027), .ZN(n8032) );
  INV_X1 U9706 ( .A(n8028), .ZN(n8029) );
  OAI22_X1 U9707 ( .A1(n8030), .A2(n8138), .B1(n8029), .B2(n8075), .ZN(n8031)
         );
  AOI211_X1 U9708 ( .C1(n8286), .C2(n8129), .A(n8032), .B(n8031), .ZN(n8033)
         );
  OAI21_X1 U9709 ( .B1(n8034), .B2(n8132), .A(n8033), .ZN(P2_U3160) );
  OR2_X1 U9710 ( .A1(n8011), .A2(n8035), .ZN(n8037) );
  AND2_X1 U9711 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  XOR2_X1 U9712 ( .A(n8039), .B(n8038), .Z(n8045) );
  AOI22_X1 U9713 ( .A1(n8567), .A2(n8092), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8041) );
  NAND2_X1 U9714 ( .A1(n8141), .A2(n8570), .ZN(n8040) );
  OAI211_X1 U9715 ( .C1(n8042), .C2(n8095), .A(n8041), .B(n8040), .ZN(n8043)
         );
  AOI21_X1 U9716 ( .B1(n8719), .B2(n8129), .A(n8043), .ZN(n8044) );
  OAI21_X1 U9717 ( .B1(n8045), .B2(n8132), .A(n8044), .ZN(P2_U3163) );
  XOR2_X1 U9718 ( .A(n8047), .B(n8046), .Z(n8052) );
  AOI22_X1 U9719 ( .A1(n8518), .A2(n8092), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8049) );
  NAND2_X1 U9720 ( .A1(n8522), .A2(n8141), .ZN(n8048) );
  OAI211_X1 U9721 ( .C1(n8541), .C2(n8095), .A(n8049), .B(n8048), .ZN(n8050)
         );
  AOI21_X1 U9722 ( .B1(n8696), .B2(n8129), .A(n8050), .ZN(n8051) );
  OAI21_X1 U9723 ( .B1(n8052), .B2(n8132), .A(n8051), .ZN(P2_U3165) );
  INV_X1 U9724 ( .A(n8053), .ZN(n8066) );
  INV_X1 U9725 ( .A(n8054), .ZN(n8071) );
  INV_X1 U9726 ( .A(n8056), .ZN(n8059) );
  INV_X1 U9727 ( .A(n8057), .ZN(n8058) );
  AOI21_X1 U9728 ( .B1(n8055), .B2(n8059), .A(n8058), .ZN(n8060) );
  OAI21_X1 U9729 ( .B1(n8071), .B2(n8060), .A(n8116), .ZN(n8065) );
  NAND2_X1 U9730 ( .A1(n8136), .A2(n8383), .ZN(n8061) );
  NAND2_X1 U9731 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n8439) );
  OAI211_X1 U9732 ( .C1(n8604), .C2(n8138), .A(n8061), .B(n8439), .ZN(n8062)
         );
  AOI21_X1 U9733 ( .B1(n8063), .B2(n8141), .A(n8062), .ZN(n8064) );
  OAI211_X1 U9734 ( .C1(n8066), .C2(n8145), .A(n8065), .B(n8064), .ZN(P2_U3166) );
  INV_X1 U9735 ( .A(n8067), .ZN(n8737) );
  INV_X1 U9736 ( .A(n8068), .ZN(n8070) );
  NOR3_X1 U9737 ( .A1(n8071), .A2(n8070), .A3(n8069), .ZN(n8073) );
  INV_X1 U9738 ( .A(n8072), .ZN(n8114) );
  OAI21_X1 U9739 ( .B1(n8073), .B2(n8114), .A(n8116), .ZN(n8079) );
  NAND2_X1 U9740 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8461) );
  OAI21_X1 U9741 ( .B1(n8138), .B2(n8074), .A(n8461), .ZN(n8077) );
  NOR2_X1 U9742 ( .A1(n8075), .A2(n8619), .ZN(n8076) );
  AOI211_X1 U9743 ( .C1(n8136), .C2(n8626), .A(n8077), .B(n8076), .ZN(n8078)
         );
  OAI211_X1 U9744 ( .C1(n8737), .C2(n8145), .A(n8079), .B(n8078), .ZN(P2_U3168) );
  XOR2_X1 U9745 ( .A(n8081), .B(n8080), .Z(n8086) );
  AOI22_X1 U9746 ( .A1(n8381), .A2(n8092), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8083) );
  NAND2_X1 U9747 ( .A1(n8534), .A2(n8141), .ZN(n8082) );
  OAI211_X1 U9748 ( .C1(n8532), .C2(n8095), .A(n8083), .B(n8082), .ZN(n8084)
         );
  AOI21_X1 U9749 ( .B1(n8702), .B2(n8129), .A(n8084), .ZN(n8085) );
  OAI21_X1 U9750 ( .B1(n8086), .B2(n8132), .A(n8085), .ZN(P2_U3169) );
  OR2_X1 U9751 ( .A1(n8011), .A2(n8087), .ZN(n8089) );
  NAND2_X1 U9752 ( .A1(n8089), .A2(n8088), .ZN(n8090) );
  XOR2_X1 U9753 ( .A(n8091), .B(n8090), .Z(n8098) );
  AOI22_X1 U9754 ( .A1(n8092), .A2(n8581), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8094) );
  NAND2_X1 U9755 ( .A1(n8141), .A2(n8585), .ZN(n8093) );
  OAI211_X1 U9756 ( .C1(n8606), .C2(n8095), .A(n8094), .B(n8093), .ZN(n8096)
         );
  AOI21_X1 U9757 ( .B1(n8726), .B2(n8129), .A(n8096), .ZN(n8097) );
  OAI21_X1 U9758 ( .B1(n8098), .B2(n8132), .A(n8097), .ZN(P2_U3173) );
  INV_X1 U9759 ( .A(n8713), .ZN(n8110) );
  OR2_X1 U9760 ( .A1(n8011), .A2(n8099), .ZN(n8101) );
  AND2_X1 U9761 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  AOI21_X1 U9762 ( .B1(n8103), .B2(n8102), .A(n8132), .ZN(n8105) );
  NAND2_X1 U9763 ( .A1(n8105), .A2(n8104), .ZN(n8109) );
  AOI22_X1 U9764 ( .A1(n8136), .A2(n8581), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8106) );
  OAI21_X1 U9765 ( .B1(n8532), .B2(n8138), .A(n8106), .ZN(n8107) );
  AOI21_X1 U9766 ( .B1(n8558), .B2(n8141), .A(n8107), .ZN(n8108) );
  OAI211_X1 U9767 ( .C1(n8110), .C2(n8145), .A(n8109), .B(n8108), .ZN(P2_U3175) );
  INV_X1 U9768 ( .A(n8111), .ZN(n8113) );
  NOR3_X1 U9769 ( .A1(n8114), .A2(n8113), .A3(n8112), .ZN(n8118) );
  INV_X1 U9770 ( .A(n8115), .ZN(n8117) );
  OAI21_X1 U9771 ( .B1(n8118), .B2(n8117), .A(n8116), .ZN(n8122) );
  NAND2_X1 U9772 ( .A1(n8136), .A2(n8382), .ZN(n8119) );
  NAND2_X1 U9773 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8477) );
  OAI211_X1 U9774 ( .C1(n8606), .C2(n8138), .A(n8119), .B(n8477), .ZN(n8120)
         );
  AOI21_X1 U9775 ( .B1(n8609), .B2(n8141), .A(n8120), .ZN(n8121) );
  OAI211_X1 U9776 ( .C1(n8123), .C2(n8145), .A(n8122), .B(n8121), .ZN(P2_U3178) );
  XOR2_X1 U9777 ( .A(n8125), .B(n8124), .Z(n8131) );
  AOI22_X1 U9778 ( .A1(n8381), .A2(n8136), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8127) );
  NAND2_X1 U9779 ( .A1(n8511), .A2(n8141), .ZN(n8126) );
  OAI211_X1 U9780 ( .C1(n8508), .C2(n8138), .A(n8127), .B(n8126), .ZN(n8128)
         );
  AOI21_X1 U9781 ( .B1(n8512), .B2(n8129), .A(n8128), .ZN(n8130) );
  OAI21_X1 U9782 ( .B1(n8131), .B2(n8132), .A(n8130), .ZN(P2_U3180) );
  INV_X1 U9783 ( .A(n8225), .ZN(n8146) );
  AOI21_X1 U9784 ( .B1(n8134), .B2(n8133), .A(n8132), .ZN(n8135) );
  NAND2_X1 U9785 ( .A1(n8135), .A2(n8055), .ZN(n8144) );
  AND2_X1 U9786 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8418) );
  AOI21_X1 U9787 ( .B1(n8136), .B2(n8384), .A(n8418), .ZN(n8137) );
  OAI21_X1 U9788 ( .B1(n8139), .B2(n8138), .A(n8137), .ZN(n8140) );
  AOI21_X1 U9789 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8143) );
  OAI211_X1 U9790 ( .C1(n8146), .C2(n8145), .A(n8144), .B(n8143), .ZN(P2_U3181) );
  INV_X1 U9791 ( .A(n8147), .ZN(n8264) );
  MUX2_X1 U9792 ( .A(n8264), .B(n8265), .S(n8301), .Z(n8148) );
  NOR2_X1 U9793 ( .A1(n8497), .A2(n8148), .ZN(n8276) );
  AOI22_X1 U9794 ( .A1(n6345), .A2(n8149), .B1(n8278), .B2(n8152), .ZN(n8156)
         );
  INV_X1 U9795 ( .A(n8149), .ZN(n8150) );
  AOI211_X1 U9796 ( .C1(n8361), .C2(n8151), .A(n8301), .B(n8150), .ZN(n8155)
         );
  MUX2_X1 U9797 ( .A(n8153), .B(n8152), .S(n8301), .Z(n8154) );
  OAI211_X1 U9798 ( .C1(n8156), .C2(n8155), .A(n6346), .B(n8154), .ZN(n8157)
         );
  INV_X1 U9799 ( .A(n8157), .ZN(n8163) );
  NAND2_X1 U9800 ( .A1(n8393), .A2(n9884), .ZN(n8170) );
  NAND2_X1 U9801 ( .A1(n8170), .A2(n8158), .ZN(n8161) );
  NAND2_X1 U9802 ( .A1(n8159), .A2(n8164), .ZN(n8160) );
  NAND2_X1 U9803 ( .A1(n6877), .A2(n9890), .ZN(n8167) );
  OAI21_X1 U9804 ( .B1(n8169), .B2(n8168), .A(n8175), .ZN(n8181) );
  INV_X1 U9805 ( .A(n8170), .ZN(n8173) );
  OAI211_X1 U9806 ( .C1(n8174), .C2(n8173), .A(n8172), .B(n8171), .ZN(n8177)
         );
  NAND3_X1 U9807 ( .A1(n8177), .A2(n8176), .A3(n8175), .ZN(n8179) );
  NAND2_X1 U9808 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  MUX2_X1 U9809 ( .A(n8181), .B(n8180), .S(n8278), .Z(n8186) );
  NAND2_X1 U9810 ( .A1(n8192), .A2(n8190), .ZN(n8185) );
  NAND2_X1 U9811 ( .A1(n8183), .A2(n8182), .ZN(n8184) );
  MUX2_X1 U9812 ( .A(n8185), .B(n8184), .S(n8301), .Z(n8194) );
  OAI21_X1 U9813 ( .B1(n8194), .B2(n8188), .A(n8187), .ZN(n8196) );
  AND2_X1 U9814 ( .A1(n8190), .A2(n8189), .ZN(n8193) );
  OAI211_X1 U9815 ( .C1(n8194), .C2(n8193), .A(n8192), .B(n8191), .ZN(n8195)
         );
  MUX2_X1 U9816 ( .A(n8196), .B(n8195), .S(n8301), .Z(n8204) );
  INV_X1 U9817 ( .A(n8327), .ZN(n8201) );
  NAND2_X1 U9818 ( .A1(n8207), .A2(n8197), .ZN(n8199) );
  NAND2_X1 U9819 ( .A1(n8206), .A2(n9914), .ZN(n8198) );
  MUX2_X1 U9820 ( .A(n8199), .B(n8198), .S(n8278), .Z(n8200) );
  OAI21_X1 U9821 ( .B1(n8202), .B2(n8201), .A(n8200), .ZN(n8203) );
  MUX2_X1 U9822 ( .A(n8207), .B(n8206), .S(n8301), .Z(n8208) );
  NAND2_X1 U9823 ( .A1(n9930), .A2(n8210), .ZN(n8211) );
  MUX2_X1 U9824 ( .A(n8212), .B(n8211), .S(n8278), .Z(n8213) );
  MUX2_X1 U9825 ( .A(n8215), .B(n8214), .S(n8301), .Z(n8216) );
  MUX2_X1 U9826 ( .A(n8219), .B(n8218), .S(n8278), .Z(n8220) );
  NAND2_X1 U9827 ( .A1(n8223), .A2(n8222), .ZN(n8229) );
  NAND2_X1 U9828 ( .A1(n8383), .A2(n8278), .ZN(n8227) );
  NAND2_X1 U9829 ( .A1(n8224), .A2(n8301), .ZN(n8226) );
  MUX2_X1 U9830 ( .A(n8227), .B(n8226), .S(n8225), .Z(n8228) );
  NAND3_X1 U9831 ( .A1(n8229), .A2(n8335), .A3(n8228), .ZN(n8233) );
  MUX2_X1 U9832 ( .A(n8231), .B(n8230), .S(n8278), .Z(n8232) );
  NAND3_X1 U9833 ( .A1(n8233), .A2(n8622), .A3(n8232), .ZN(n8237) );
  NAND3_X1 U9834 ( .A1(n8237), .A2(n8238), .A3(n8234), .ZN(n8235) );
  NAND3_X1 U9835 ( .A1(n8237), .A2(n8236), .A3(n8593), .ZN(n8239) );
  INV_X1 U9836 ( .A(n8243), .ZN(n8241) );
  NAND3_X1 U9837 ( .A1(n8248), .A2(n8249), .A3(n8244), .ZN(n8242) );
  NAND2_X1 U9838 ( .A1(n8242), .A2(n8246), .ZN(n8252) );
  NAND2_X1 U9839 ( .A1(n8244), .A2(n8243), .ZN(n8247) );
  NAND2_X1 U9840 ( .A1(n8250), .A2(n8249), .ZN(n8251) );
  INV_X1 U9841 ( .A(n8551), .ZN(n8549) );
  INV_X1 U9842 ( .A(n8253), .ZN(n8256) );
  INV_X1 U9843 ( .A(n8254), .ZN(n8255) );
  MUX2_X1 U9844 ( .A(n8256), .B(n8255), .S(n8301), .Z(n8257) );
  AOI21_X1 U9845 ( .B1(n8258), .B2(n8549), .A(n8257), .ZN(n8260) );
  INV_X1 U9846 ( .A(n8525), .ZN(n8311) );
  OAI21_X1 U9847 ( .B1(n8260), .B2(n8312), .A(n8259), .ZN(n8261) );
  NAND2_X1 U9848 ( .A1(n8261), .A2(n8310), .ZN(n8262) );
  NAND2_X1 U9849 ( .A1(n8267), .A2(n8266), .ZN(n8517) );
  MUX2_X1 U9850 ( .A(n8267), .B(n8266), .S(n8301), .Z(n8268) );
  INV_X1 U9851 ( .A(n8270), .ZN(n8273) );
  NOR2_X1 U9852 ( .A1(n8271), .A2(n8380), .ZN(n8272) );
  MUX2_X1 U9853 ( .A(n8273), .B(n8272), .S(n8301), .Z(n8274) );
  MUX2_X1 U9854 ( .A(n8498), .B(n8286), .S(n8278), .Z(n8287) );
  INV_X1 U9855 ( .A(n8287), .ZN(n8279) );
  NAND2_X1 U9856 ( .A1(n8280), .A2(n6095), .ZN(n8283) );
  OR2_X1 U9857 ( .A1(n8291), .A2(n8281), .ZN(n8282) );
  INV_X1 U9858 ( .A(n8379), .ZN(n8285) );
  NAND2_X1 U9859 ( .A1(n8679), .A2(n8285), .ZN(n8307) );
  AND2_X1 U9860 ( .A1(n8288), .A2(n8287), .ZN(n8289) );
  NAND2_X1 U9861 ( .A1(n9383), .A2(n6095), .ZN(n8293) );
  OR2_X1 U9862 ( .A1(n8291), .A2(n8744), .ZN(n8292) );
  INV_X1 U9863 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U9864 ( .A1(n6183), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8296) );
  INV_X1 U9865 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8294) );
  OR2_X1 U9866 ( .A1(n6077), .A2(n8294), .ZN(n8295) );
  OAI211_X1 U9867 ( .C1(n4271), .C2(n8297), .A(n8296), .B(n8295), .ZN(n8298)
         );
  INV_X1 U9868 ( .A(n8298), .ZN(n8299) );
  NAND2_X1 U9869 ( .A1(n8305), .A2(n8490), .ZN(n8363) );
  NAND2_X1 U9870 ( .A1(n8307), .A2(n8301), .ZN(n8302) );
  NAND4_X1 U9871 ( .A1(n8363), .A2(n8303), .A3(n8354), .A4(n8302), .ZN(n8304)
         );
  OR2_X1 U9872 ( .A1(n8364), .A2(n8304), .ZN(n8367) );
  NOR2_X1 U9873 ( .A1(n8305), .A2(n8490), .ZN(n8352) );
  INV_X1 U9874 ( .A(n8352), .ZN(n8306) );
  NAND2_X1 U9875 ( .A1(n8306), .A2(n8363), .ZN(n8348) );
  INV_X1 U9876 ( .A(n8354), .ZN(n8347) );
  INV_X1 U9877 ( .A(n8307), .ZN(n8346) );
  INV_X1 U9878 ( .A(n8308), .ZN(n8343) );
  NOR2_X1 U9879 ( .A1(n8312), .A2(n8311), .ZN(n8538) );
  INV_X1 U9880 ( .A(n8313), .ZN(n8594) );
  INV_X1 U9881 ( .A(n8579), .ZN(n8576) );
  NOR2_X1 U9882 ( .A1(n8315), .A2(n8314), .ZN(n8317) );
  AND4_X1 U9883 ( .A1(n8317), .A2(n6345), .A3(n9871), .A4(n8316), .ZN(n8320)
         );
  NAND4_X1 U9884 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n9862), .ZN(n8324)
         );
  NOR4_X1 U9885 ( .A1(n8324), .A2(n8323), .A3(n8322), .A4(n8321), .ZN(n8326)
         );
  NAND4_X1 U9886 ( .A1(n8328), .A2(n8327), .A3(n8326), .A4(n8325), .ZN(n8331)
         );
  OR3_X1 U9887 ( .A1(n8331), .A2(n8330), .A3(n8329), .ZN(n8332) );
  NOR2_X1 U9888 ( .A1(n8333), .A2(n8332), .ZN(n8334) );
  NAND3_X1 U9889 ( .A1(n8622), .A2(n8335), .A3(n8334), .ZN(n8336) );
  NOR2_X1 U9890 ( .A1(n8602), .A2(n8336), .ZN(n8337) );
  NAND4_X1 U9891 ( .A1(n8564), .A2(n8594), .A3(n8576), .A4(n8337), .ZN(n8338)
         );
  NOR2_X1 U9892 ( .A1(n8551), .A2(n8338), .ZN(n8339) );
  NAND3_X1 U9893 ( .A1(n8529), .A2(n8538), .A3(n8339), .ZN(n8340) );
  OR3_X1 U9894 ( .A1(n8341), .A2(n8517), .A3(n8340), .ZN(n8342) );
  OR4_X1 U9895 ( .A1(n8344), .A2(n8343), .A3(n8342), .A4(n8497), .ZN(n8345) );
  NOR4_X1 U9896 ( .A1(n8348), .A2(n8347), .A3(n8346), .A4(n8345), .ZN(n8358)
         );
  INV_X1 U9897 ( .A(n8349), .ZN(n8350) );
  AOI21_X1 U9898 ( .B1(n8678), .B2(n8679), .A(n8352), .ZN(n8353) );
  INV_X1 U9899 ( .A(n8490), .ZN(n8378) );
  AOI21_X1 U9900 ( .B1(n8354), .B2(n8378), .A(n8678), .ZN(n8356) );
  NOR3_X1 U9901 ( .A1(n8361), .A2(n8360), .A3(n8359), .ZN(n8362) );
  NAND2_X1 U9902 ( .A1(n8364), .A2(n4875), .ZN(n8365) );
  NAND3_X1 U9903 ( .A1(n8367), .A2(n8366), .A3(n8365), .ZN(n8369) );
  XNOR2_X1 U9904 ( .A(n8369), .B(n8368), .ZN(n8377) );
  NOR3_X1 U9905 ( .A1(n8372), .A2(n8371), .A3(n8370), .ZN(n8375) );
  OAI21_X1 U9906 ( .B1(n8376), .B2(n8373), .A(P2_B_REG_SCAN_IN), .ZN(n8374) );
  OAI22_X1 U9907 ( .A1(n8377), .A2(n8376), .B1(n8375), .B2(n8374), .ZN(
        P2_U3296) );
  MUX2_X1 U9908 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8378), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9909 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8379), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9910 ( .A(n8498), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8474), .Z(
        P2_U3519) );
  MUX2_X1 U9911 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8380), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9912 ( .A(n8518), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8474), .Z(
        P2_U3517) );
  MUX2_X1 U9913 ( .A(n8381), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8474), .Z(
        P2_U3516) );
  MUX2_X1 U9914 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8519), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9915 ( .A(n8555), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8474), .Z(
        P2_U3514) );
  MUX2_X1 U9916 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8567), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9917 ( .A(n8581), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8474), .Z(
        P2_U3512) );
  MUX2_X1 U9918 ( .A(n8589), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8474), .Z(
        P2_U3511) );
  MUX2_X1 U9919 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8582), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9920 ( .A(n8625), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8474), .Z(
        P2_U3509) );
  MUX2_X1 U9921 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8382), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9922 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8626), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9923 ( .A(n8383), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8474), .Z(
        P2_U3506) );
  MUX2_X1 U9924 ( .A(n8384), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8474), .Z(
        P2_U3505) );
  MUX2_X1 U9925 ( .A(n8385), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8474), .Z(
        P2_U3504) );
  MUX2_X1 U9926 ( .A(n8386), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8474), .Z(
        P2_U3503) );
  MUX2_X1 U9927 ( .A(n8387), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8474), .Z(
        P2_U3502) );
  MUX2_X1 U9928 ( .A(n8388), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8474), .Z(
        P2_U3501) );
  MUX2_X1 U9929 ( .A(n7303), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8474), .Z(
        P2_U3500) );
  MUX2_X1 U9930 ( .A(n8389), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8474), .Z(
        P2_U3499) );
  MUX2_X1 U9931 ( .A(n8390), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8474), .Z(
        P2_U3498) );
  MUX2_X1 U9932 ( .A(n8391), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8474), .Z(
        P2_U3497) );
  MUX2_X1 U9933 ( .A(n8392), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8474), .Z(
        P2_U3496) );
  MUX2_X1 U9934 ( .A(n6877), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8474), .Z(
        P2_U3495) );
  MUX2_X1 U9935 ( .A(n8393), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8474), .Z(
        P2_U3494) );
  MUX2_X1 U9936 ( .A(n6922), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8474), .Z(
        P2_U3493) );
  MUX2_X1 U9937 ( .A(n6758), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8474), .Z(
        P2_U3492) );
  MUX2_X1 U9938 ( .A(n8394), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8474), .Z(
        P2_U3491) );
  AOI21_X1 U9939 ( .B1(n4342), .B2(n8396), .A(n8395), .ZN(n8413) );
  INV_X1 U9940 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8404) );
  OAI21_X1 U9941 ( .B1(n8399), .B2(n8398), .A(n8397), .ZN(n8400) );
  NAND2_X1 U9942 ( .A1(n8400), .A2(n9827), .ZN(n8403) );
  INV_X1 U9943 ( .A(n8401), .ZN(n8402) );
  OAI211_X1 U9944 ( .C1(n9831), .C2(n8404), .A(n8403), .B(n8402), .ZN(n8410)
         );
  AOI21_X1 U9945 ( .B1(n8407), .B2(n8406), .A(n8405), .ZN(n8408) );
  NOR2_X1 U9946 ( .A1(n8408), .A2(n8485), .ZN(n8409) );
  AOI211_X1 U9947 ( .C1(n9839), .C2(n8411), .A(n8410), .B(n8409), .ZN(n8412)
         );
  OAI21_X1 U9948 ( .B1(n8413), .B2(n9822), .A(n8412), .ZN(P2_U3196) );
  AOI21_X1 U9949 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8432) );
  NAND2_X1 U9950 ( .A1(n9839), .A2(n8417), .ZN(n8430) );
  AOI21_X1 U9951 ( .B1(n9841), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8418), .ZN(
        n8429) );
  OAI21_X1 U9952 ( .B1(n8421), .B2(n8420), .A(n8419), .ZN(n8422) );
  NAND2_X1 U9953 ( .A1(n8422), .A2(n9827), .ZN(n8428) );
  AOI21_X1 U9954 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n8426) );
  OR2_X1 U9955 ( .A1(n8485), .A2(n8426), .ZN(n8427) );
  OAI21_X1 U9956 ( .B1(n8432), .B2(n9822), .A(n8431), .ZN(P2_U3197) );
  AOI21_X1 U9957 ( .B1(n4340), .B2(n8434), .A(n8433), .ZN(n8450) );
  INV_X1 U9958 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8441) );
  OAI21_X1 U9959 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8438) );
  NAND2_X1 U9960 ( .A1(n8438), .A2(n9827), .ZN(n8440) );
  OAI211_X1 U9961 ( .C1(n9831), .C2(n8441), .A(n8440), .B(n8439), .ZN(n8447)
         );
  AOI21_X1 U9962 ( .B1(n8444), .B2(n8443), .A(n8442), .ZN(n8445) );
  NOR2_X1 U9963 ( .A1(n8445), .A2(n8485), .ZN(n8446) );
  AOI211_X1 U9964 ( .C1(n9839), .C2(n8448), .A(n8447), .B(n8446), .ZN(n8449)
         );
  OAI21_X1 U9965 ( .B1(n8450), .B2(n9822), .A(n8449), .ZN(P2_U3198) );
  AOI21_X1 U9966 ( .B1(n8453), .B2(n8452), .A(n8451), .ZN(n8468) );
  OAI21_X1 U9967 ( .B1(n8456), .B2(n8455), .A(n8454), .ZN(n8466) );
  AOI21_X1 U9968 ( .B1(n8459), .B2(n8458), .A(n8457), .ZN(n8462) );
  NAND2_X1 U9969 ( .A1(n9841), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8460) );
  OAI211_X1 U9970 ( .C1(n8485), .C2(n8462), .A(n8461), .B(n8460), .ZN(n8465)
         );
  NOR2_X1 U9971 ( .A1(n8473), .A2(n8463), .ZN(n8464) );
  AOI211_X1 U9972 ( .C1(n9827), .C2(n8466), .A(n8465), .B(n8464), .ZN(n8467)
         );
  OAI21_X1 U9973 ( .B1(n8468), .B2(n9822), .A(n8467), .ZN(P2_U3199) );
  AOI21_X1 U9974 ( .B1(n4304), .B2(n8470), .A(n8469), .ZN(n8486) );
  NAND2_X1 U9975 ( .A1(n8472), .A2(n8471), .ZN(n8476) );
  OAI21_X1 U9976 ( .B1(n8474), .B2(n8476), .A(n8473), .ZN(n8483) );
  INV_X1 U9977 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9961) );
  NAND3_X1 U9978 ( .A1(n8476), .A2(n9827), .A3(n8475), .ZN(n8478) );
  OAI211_X1 U9979 ( .C1(n9831), .C2(n9961), .A(n8478), .B(n8477), .ZN(n8482)
         );
  NAND2_X1 U9980 ( .A1(n8487), .A2(n9865), .ZN(n8491) );
  INV_X1 U9981 ( .A(n8488), .ZN(n8489) );
  AOI21_X1 U9982 ( .B1(n8491), .B2(n8676), .A(n9870), .ZN(n8493) );
  AOI21_X1 U9983 ( .B1(n9870), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8493), .ZN(
        n8492) );
  OAI21_X1 U9984 ( .B1(n8678), .B2(n8620), .A(n8492), .ZN(P2_U3202) );
  INV_X1 U9985 ( .A(n8679), .ZN(n8636) );
  AOI21_X1 U9986 ( .B1(n9870), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8493), .ZN(
        n8494) );
  OAI21_X1 U9987 ( .B1(n8636), .B2(n8620), .A(n8494), .ZN(P2_U3203) );
  XNOR2_X1 U9988 ( .A(n8495), .B(n8497), .ZN(n8688) );
  INV_X1 U9989 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8500) );
  XOR2_X1 U9990 ( .A(n8497), .B(n8496), .Z(n8499) );
  AOI222_X1 U9991 ( .A1(n9861), .A2(n8499), .B1(n8518), .B2(n9858), .C1(n8498), 
        .C2(n9859), .ZN(n8683) );
  MUX2_X1 U9992 ( .A(n8500), .B(n8683), .S(n8608), .Z(n8503) );
  AOI22_X1 U9993 ( .A1(n8685), .A2(n9864), .B1(n9865), .B2(n8501), .ZN(n8502)
         );
  OAI211_X1 U9994 ( .C1(n8688), .C2(n8615), .A(n8503), .B(n8502), .ZN(P2_U3206) );
  XNOR2_X1 U9995 ( .A(n8504), .B(n8505), .ZN(n8691) );
  INV_X1 U9996 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8510) );
  XNOR2_X1 U9997 ( .A(n8506), .B(n8505), .ZN(n8507) );
  OAI222_X1 U9998 ( .A1(n8607), .A2(n8508), .B1(n8605), .B2(n8531), .C1(n9872), 
        .C2(n8507), .ZN(n8689) );
  INV_X1 U9999 ( .A(n8689), .ZN(n8509) );
  MUX2_X1 U10000 ( .A(n8510), .B(n8509), .S(n8608), .Z(n8514) );
  AOI22_X1 U10001 ( .A1(n8512), .A2(n9864), .B1(n9865), .B2(n8511), .ZN(n8513)
         );
  OAI211_X1 U10002 ( .C1(n8691), .C2(n8615), .A(n8514), .B(n8513), .ZN(
        P2_U3207) );
  XOR2_X1 U10003 ( .A(n8517), .B(n8515), .Z(n8699) );
  XOR2_X1 U10004 ( .A(n8517), .B(n8516), .Z(n8520) );
  AOI222_X1 U10005 ( .A1(n9861), .A2(n8520), .B1(n8519), .B2(n9858), .C1(n8518), .C2(n9859), .ZN(n8694) );
  MUX2_X1 U10006 ( .A(n8521), .B(n8694), .S(n8608), .Z(n8524) );
  AOI22_X1 U10007 ( .A1(n8696), .A2(n9864), .B1(n9865), .B2(n8522), .ZN(n8523)
         );
  OAI211_X1 U10008 ( .C1(n8699), .C2(n8615), .A(n8524), .B(n8523), .ZN(
        P2_U3208) );
  NAND2_X1 U10009 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  XOR2_X1 U10010 ( .A(n8529), .B(n8527), .Z(n8705) );
  INV_X1 U10011 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8533) );
  XOR2_X1 U10012 ( .A(n8528), .B(n8529), .Z(n8530) );
  OAI222_X1 U10013 ( .A1(n8605), .A2(n8532), .B1(n8607), .B2(n8531), .C1(n9872), .C2(n8530), .ZN(n8645) );
  INV_X1 U10014 ( .A(n8645), .ZN(n8700) );
  MUX2_X1 U10015 ( .A(n8533), .B(n8700), .S(n8608), .Z(n8536) );
  AOI22_X1 U10016 ( .A1(n8702), .A2(n9864), .B1(n9865), .B2(n8534), .ZN(n8535)
         );
  OAI211_X1 U10017 ( .C1(n8705), .C2(n8615), .A(n8536), .B(n8535), .ZN(
        P2_U3209) );
  XNOR2_X1 U10018 ( .A(n8537), .B(n8538), .ZN(n8708) );
  INV_X1 U10019 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8544) );
  XNOR2_X1 U10020 ( .A(n8539), .B(n8538), .ZN(n8540) );
  OAI222_X1 U10021 ( .A1(n8605), .A2(n8542), .B1(n8607), .B2(n8541), .C1(n9872), .C2(n8540), .ZN(n8706) );
  INV_X1 U10022 ( .A(n8706), .ZN(n8543) );
  MUX2_X1 U10023 ( .A(n8544), .B(n8543), .S(n8608), .Z(n8548) );
  AOI22_X1 U10024 ( .A1(n8546), .A2(n9864), .B1(n9865), .B2(n8545), .ZN(n8547)
         );
  OAI211_X1 U10025 ( .C1(n8708), .C2(n8615), .A(n8548), .B(n8547), .ZN(
        P2_U3210) );
  XNOR2_X1 U10026 ( .A(n8550), .B(n8549), .ZN(n8716) );
  INV_X1 U10027 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8557) );
  OR3_X1 U10028 ( .A1(n8562), .A2(n8552), .A3(n8551), .ZN(n8553) );
  NAND2_X1 U10029 ( .A1(n8554), .A2(n8553), .ZN(n8556) );
  AOI222_X1 U10030 ( .A1(n9861), .A2(n8556), .B1(n8555), .B2(n9859), .C1(n8581), .C2(n9858), .ZN(n8711) );
  MUX2_X1 U10031 ( .A(n8557), .B(n8711), .S(n8608), .Z(n8560) );
  AOI22_X1 U10032 ( .A1(n8713), .A2(n9864), .B1(n9865), .B2(n8558), .ZN(n8559)
         );
  OAI211_X1 U10033 ( .C1(n8716), .C2(n8615), .A(n8560), .B(n8559), .ZN(
        P2_U3211) );
  XOR2_X1 U10034 ( .A(n8561), .B(n8564), .Z(n8722) );
  INV_X1 U10035 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8569) );
  INV_X1 U10036 ( .A(n8562), .ZN(n8566) );
  NAND3_X1 U10037 ( .A1(n8578), .A2(n8564), .A3(n8563), .ZN(n8565) );
  NAND2_X1 U10038 ( .A1(n8566), .A2(n8565), .ZN(n8568) );
  AOI222_X1 U10039 ( .A1(n9861), .A2(n8568), .B1(n8567), .B2(n9859), .C1(n8589), .C2(n9858), .ZN(n8717) );
  MUX2_X1 U10040 ( .A(n8569), .B(n8717), .S(n8608), .Z(n8572) );
  AOI22_X1 U10041 ( .A1(n8719), .A2(n9864), .B1(n9865), .B2(n8570), .ZN(n8571)
         );
  OAI211_X1 U10042 ( .C1(n8722), .C2(n8615), .A(n8572), .B(n8571), .ZN(
        P2_U3212) );
  NAND2_X1 U10043 ( .A1(n8662), .A2(n8575), .ZN(n8577) );
  XNOR2_X1 U10044 ( .A(n8577), .B(n8576), .ZN(n8729) );
  OAI21_X1 U10045 ( .B1(n8580), .B2(n8579), .A(n8578), .ZN(n8583) );
  AOI222_X1 U10046 ( .A1(n9861), .A2(n8583), .B1(n8582), .B2(n9858), .C1(n8581), .C2(n9859), .ZN(n8723) );
  MUX2_X1 U10047 ( .A(n8584), .B(n8723), .S(n8608), .Z(n8587) );
  AOI22_X1 U10048 ( .A1(n8726), .A2(n9864), .B1(n9865), .B2(n8585), .ZN(n8586)
         );
  OAI211_X1 U10049 ( .C1(n8729), .C2(n8615), .A(n8587), .B(n8586), .ZN(
        P2_U3213) );
  XNOR2_X1 U10050 ( .A(n8588), .B(n8594), .ZN(n8590) );
  AOI222_X1 U10051 ( .A1(n9861), .A2(n8590), .B1(n8589), .B2(n9859), .C1(n8625), .C2(n9858), .ZN(n8665) );
  OAI22_X1 U10052 ( .A1(n8608), .A2(n5636), .B1(n8591), .B2(n8618), .ZN(n8592)
         );
  AOI21_X1 U10053 ( .B1(n8661), .B2(n9864), .A(n8592), .ZN(n8597) );
  OR2_X1 U10054 ( .A1(n8598), .A2(n8602), .ZN(n8600) );
  NAND2_X1 U10055 ( .A1(n8600), .A2(n8593), .ZN(n8595) );
  NAND3_X1 U10056 ( .A1(n8663), .A2(n8662), .A3(n9867), .ZN(n8596) );
  OAI211_X1 U10057 ( .C1(n8665), .C2(n9870), .A(n8597), .B(n8596), .ZN(
        P2_U3214) );
  NAND2_X1 U10058 ( .A1(n8598), .A2(n8602), .ZN(n8599) );
  NAND2_X1 U10059 ( .A1(n8600), .A2(n8599), .ZN(n8734) );
  XOR2_X1 U10060 ( .A(n8602), .B(n8601), .Z(n8603) );
  OAI222_X1 U10061 ( .A1(n8607), .A2(n8606), .B1(n8605), .B2(n8604), .C1(n8603), .C2(n9872), .ZN(n8667) );
  NAND2_X1 U10062 ( .A1(n8667), .A2(n8608), .ZN(n8614) );
  INV_X1 U10063 ( .A(n8609), .ZN(n8610) );
  OAI22_X1 U10064 ( .A1(n8608), .A2(n8611), .B1(n8610), .B2(n8618), .ZN(n8612)
         );
  AOI21_X1 U10065 ( .B1(n8668), .B2(n9864), .A(n8612), .ZN(n8613) );
  OAI211_X1 U10066 ( .C1(n8734), .C2(n8615), .A(n8614), .B(n8613), .ZN(
        P2_U3215) );
  XNOR2_X1 U10067 ( .A(n8617), .B(n8616), .ZN(n8671) );
  OAI22_X1 U10068 ( .A1(n8737), .A2(n8620), .B1(n8619), .B2(n8618), .ZN(n8631)
         );
  NAND3_X1 U10069 ( .A1(n8623), .A2(n8622), .A3(n8621), .ZN(n8624) );
  NAND2_X1 U10070 ( .A1(n8624), .A2(n9861), .ZN(n8628) );
  AOI22_X1 U10071 ( .A1(n8626), .A2(n9858), .B1(n9859), .B2(n8625), .ZN(n8627)
         );
  OAI21_X1 U10072 ( .B1(n8629), .B2(n8628), .A(n8627), .ZN(n8735) );
  MUX2_X1 U10073 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8735), .S(n8608), .Z(n8630) );
  AOI211_X1 U10074 ( .C1(n9867), .C2(n8671), .A(n8631), .B(n8630), .ZN(n8632)
         );
  INV_X1 U10075 ( .A(n8632), .ZN(P2_U3216) );
  NOR2_X1 U10076 ( .A1(n8676), .A2(n9950), .ZN(n8634) );
  AOI21_X1 U10077 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9950), .A(n8634), .ZN(
        n8633) );
  OAI21_X1 U10078 ( .B1(n8678), .B2(n8672), .A(n8633), .ZN(P2_U3490) );
  AOI21_X1 U10079 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9950), .A(n8634), .ZN(
        n8635) );
  OAI21_X1 U10080 ( .B1(n8636), .B2(n8672), .A(n8635), .ZN(P2_U3489) );
  INV_X1 U10081 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8637) );
  MUX2_X1 U10082 ( .A(n8637), .B(n8683), .S(n9952), .Z(n8639) );
  NAND2_X1 U10083 ( .A1(n8685), .A2(n8658), .ZN(n8638) );
  OAI211_X1 U10084 ( .C1(n8688), .C2(n8673), .A(n8639), .B(n8638), .ZN(
        P2_U3486) );
  MUX2_X1 U10085 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8689), .S(n9952), .Z(n8641) );
  OAI22_X1 U10086 ( .A1(n8691), .A2(n8673), .B1(n8690), .B2(n8672), .ZN(n8640)
         );
  OR2_X1 U10087 ( .A1(n8641), .A2(n8640), .ZN(P2_U3485) );
  INV_X1 U10088 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8642) );
  MUX2_X1 U10089 ( .A(n8642), .B(n8694), .S(n9952), .Z(n8644) );
  NAND2_X1 U10090 ( .A1(n8696), .A2(n8658), .ZN(n8643) );
  OAI211_X1 U10091 ( .C1(n8699), .C2(n8673), .A(n8644), .B(n8643), .ZN(
        P2_U3484) );
  MUX2_X1 U10092 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8645), .S(n9952), .Z(n8648) );
  OAI22_X1 U10093 ( .A1(n8705), .A2(n8673), .B1(n8646), .B2(n8672), .ZN(n8647)
         );
  OR2_X1 U10094 ( .A1(n8648), .A2(n8647), .ZN(P2_U3483) );
  MUX2_X1 U10095 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8706), .S(n9952), .Z(n8650) );
  OAI22_X1 U10096 ( .A1(n8708), .A2(n8673), .B1(n8707), .B2(n8672), .ZN(n8649)
         );
  OR2_X1 U10097 ( .A1(n8650), .A2(n8649), .ZN(P2_U3482) );
  INV_X1 U10098 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8651) );
  MUX2_X1 U10099 ( .A(n8651), .B(n8711), .S(n9952), .Z(n8653) );
  NAND2_X1 U10100 ( .A1(n8713), .A2(n8658), .ZN(n8652) );
  OAI211_X1 U10101 ( .C1(n8716), .C2(n8673), .A(n8653), .B(n8652), .ZN(
        P2_U3481) );
  INV_X1 U10102 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8654) );
  MUX2_X1 U10103 ( .A(n8654), .B(n8717), .S(n9952), .Z(n8656) );
  NAND2_X1 U10104 ( .A1(n8719), .A2(n8658), .ZN(n8655) );
  OAI211_X1 U10105 ( .C1(n8673), .C2(n8722), .A(n8656), .B(n8655), .ZN(
        P2_U3480) );
  INV_X1 U10106 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8657) );
  MUX2_X1 U10107 ( .A(n8657), .B(n8723), .S(n9952), .Z(n8660) );
  NAND2_X1 U10108 ( .A1(n8726), .A2(n8658), .ZN(n8659) );
  OAI211_X1 U10109 ( .C1(n8729), .C2(n8673), .A(n8660), .B(n8659), .ZN(
        P2_U3479) );
  INV_X1 U10110 ( .A(n8661), .ZN(n8666) );
  NAND3_X1 U10111 ( .A1(n8663), .A2(n8662), .A3(n9921), .ZN(n8664) );
  OAI211_X1 U10112 ( .C1(n8666), .C2(n9913), .A(n8665), .B(n8664), .ZN(n8730)
         );
  MUX2_X1 U10113 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8730), .S(n9952), .Z(
        P2_U3478) );
  AOI21_X1 U10114 ( .B1(n9931), .B2(n8668), .A(n8667), .ZN(n8731) );
  MUX2_X1 U10115 ( .A(n8669), .B(n8731), .S(n9952), .Z(n8670) );
  OAI21_X1 U10116 ( .B1(n8673), .B2(n8734), .A(n8670), .ZN(P2_U3477) );
  MUX2_X1 U10117 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8735), .S(n9952), .Z(n8675) );
  INV_X1 U10118 ( .A(n8671), .ZN(n8739) );
  OAI22_X1 U10119 ( .A1(n8739), .A2(n8673), .B1(n8737), .B2(n8672), .ZN(n8674)
         );
  OR2_X1 U10120 ( .A1(n8675), .A2(n8674), .ZN(P2_U3476) );
  NOR2_X1 U10121 ( .A1(n8676), .A2(n9934), .ZN(n8680) );
  AOI21_X1 U10122 ( .B1(n9934), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8680), .ZN(
        n8677) );
  OAI21_X1 U10123 ( .B1(n8678), .B2(n8736), .A(n8677), .ZN(P2_U3458) );
  NAND2_X1 U10124 ( .A1(n8679), .A2(n8725), .ZN(n8682) );
  INV_X1 U10125 ( .A(n8680), .ZN(n8681) );
  OAI211_X1 U10126 ( .C1(n6423), .C2(n9932), .A(n8682), .B(n8681), .ZN(
        P2_U3457) );
  MUX2_X1 U10127 ( .A(n8684), .B(n8683), .S(n9932), .Z(n8687) );
  NAND2_X1 U10128 ( .A1(n8685), .A2(n8725), .ZN(n8686) );
  OAI211_X1 U10129 ( .C1(n8688), .C2(n8738), .A(n8687), .B(n8686), .ZN(
        P2_U3454) );
  MUX2_X1 U10130 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8689), .S(n9932), .Z(n8693) );
  OAI22_X1 U10131 ( .A1(n8691), .A2(n8738), .B1(n8690), .B2(n8736), .ZN(n8692)
         );
  OR2_X1 U10132 ( .A1(n8693), .A2(n8692), .ZN(P2_U3453) );
  INV_X1 U10133 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8695) );
  MUX2_X1 U10134 ( .A(n8695), .B(n8694), .S(n9932), .Z(n8698) );
  NAND2_X1 U10135 ( .A1(n8696), .A2(n8725), .ZN(n8697) );
  OAI211_X1 U10136 ( .C1(n8699), .C2(n8738), .A(n8698), .B(n8697), .ZN(
        P2_U3452) );
  MUX2_X1 U10137 ( .A(n8701), .B(n8700), .S(n9932), .Z(n8704) );
  NAND2_X1 U10138 ( .A1(n8702), .A2(n8725), .ZN(n8703) );
  OAI211_X1 U10139 ( .C1(n8705), .C2(n8738), .A(n8704), .B(n8703), .ZN(
        P2_U3451) );
  MUX2_X1 U10140 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8706), .S(n9932), .Z(n8710) );
  OAI22_X1 U10141 ( .A1(n8708), .A2(n8738), .B1(n8707), .B2(n8736), .ZN(n8709)
         );
  OR2_X1 U10142 ( .A1(n8710), .A2(n8709), .ZN(P2_U3450) );
  INV_X1 U10143 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8712) );
  MUX2_X1 U10144 ( .A(n8712), .B(n8711), .S(n9932), .Z(n8715) );
  NAND2_X1 U10145 ( .A1(n8713), .A2(n8725), .ZN(n8714) );
  OAI211_X1 U10146 ( .C1(n8716), .C2(n8738), .A(n8715), .B(n8714), .ZN(
        P2_U3449) );
  INV_X1 U10147 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8718) );
  MUX2_X1 U10148 ( .A(n8718), .B(n8717), .S(n9932), .Z(n8721) );
  NAND2_X1 U10149 ( .A1(n8719), .A2(n8725), .ZN(n8720) );
  OAI211_X1 U10150 ( .C1(n8722), .C2(n8738), .A(n8721), .B(n8720), .ZN(
        P2_U3448) );
  INV_X1 U10151 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8724) );
  MUX2_X1 U10152 ( .A(n8724), .B(n8723), .S(n9932), .Z(n8728) );
  NAND2_X1 U10153 ( .A1(n8726), .A2(n8725), .ZN(n8727) );
  OAI211_X1 U10154 ( .C1(n8729), .C2(n8738), .A(n8728), .B(n8727), .ZN(
        P2_U3447) );
  MUX2_X1 U10155 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8730), .S(n9932), .Z(
        P2_U3446) );
  MUX2_X1 U10156 ( .A(n8732), .B(n8731), .S(n9932), .Z(n8733) );
  OAI21_X1 U10157 ( .B1(n8734), .B2(n8738), .A(n8733), .ZN(P2_U3444) );
  MUX2_X1 U10158 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8735), .S(n9932), .Z(n8741) );
  OAI22_X1 U10159 ( .A1(n8739), .A2(n8738), .B1(n8737), .B2(n8736), .ZN(n8740)
         );
  OR2_X1 U10160 ( .A1(n8741), .A2(n8740), .ZN(P2_U3441) );
  INV_X1 U10161 ( .A(n8742), .ZN(n8746) );
  NAND3_X1 U10162 ( .A1(n8743), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8745) );
  OAI22_X1 U10163 ( .A1(n8746), .A2(n8745), .B1(n8744), .B2(n8751), .ZN(n8747)
         );
  AOI21_X1 U10164 ( .B1(n9383), .B2(n8748), .A(n8747), .ZN(n8749) );
  INV_X1 U10165 ( .A(n8749), .ZN(P2_U3264) );
  INV_X1 U10166 ( .A(n8750), .ZN(n9394) );
  OAI222_X1 U10167 ( .A1(n7936), .A2(n9394), .B1(n5980), .B2(P2_U3151), .C1(
        n8752), .C2(n8751), .ZN(P2_U3266) );
  AOI21_X1 U10168 ( .B1(n8754), .B2(n8753), .A(n4344), .ZN(n8760) );
  AOI22_X1 U10169 ( .A1(n8889), .A2(n8755), .B1(n8887), .B2(n8904), .ZN(n8756)
         );
  NAND2_X1 U10170 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9569) );
  OAI211_X1 U10171 ( .C1(n8757), .C2(n8891), .A(n8756), .B(n9569), .ZN(n8758)
         );
  AOI21_X1 U10172 ( .B1(n5177), .B2(n8894), .A(n8758), .ZN(n8759) );
  OAI21_X1 U10173 ( .B1(n8760), .B2(n8897), .A(n8759), .ZN(P1_U3215) );
  AOI21_X1 U10174 ( .B1(n8767), .B2(n8766), .A(n8765), .ZN(n8768) );
  XNOR2_X1 U10175 ( .A(n8769), .B(n8768), .ZN(n8775) );
  OAI22_X1 U10176 ( .A1(n8867), .A2(n8798), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8770), .ZN(n8773) );
  INV_X1 U10177 ( .A(n9042), .ZN(n8771) );
  OAI22_X1 U10178 ( .A1(n8846), .A2(n8771), .B1(n9074), .B2(n8891), .ZN(n8772)
         );
  AOI211_X1 U10179 ( .C1(n9183), .C2(n8894), .A(n8773), .B(n8772), .ZN(n8774)
         );
  OAI21_X1 U10180 ( .B1(n8775), .B2(n8897), .A(n8774), .ZN(P1_U3216) );
  OR2_X1 U10181 ( .A1(n8776), .A2(n8777), .ZN(n8841) );
  INV_X1 U10182 ( .A(n8840), .ZN(n8779) );
  OAI21_X1 U10183 ( .B1(n8777), .B2(n8779), .A(n8776), .ZN(n8778) );
  OAI21_X1 U10184 ( .B1(n8841), .B2(n8779), .A(n8778), .ZN(n8780) );
  NAND2_X1 U10185 ( .A1(n8780), .A2(n8876), .ZN(n8783) );
  AND2_X1 U10186 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8964) );
  OAI22_X1 U10187 ( .A1(n8846), .A2(n9105), .B1(n9144), .B2(n8891), .ZN(n8781)
         );
  AOI211_X1 U10188 ( .C1(n8887), .C2(n8901), .A(n8964), .B(n8781), .ZN(n8782)
         );
  OAI211_X1 U10189 ( .C1(n9103), .C2(n8851), .A(n8783), .B(n8782), .ZN(
        P1_U3219) );
  NAND2_X1 U10190 ( .A1(n8784), .A2(n8785), .ZN(n8786) );
  XOR2_X1 U10191 ( .A(n8787), .B(n8786), .Z(n8793) );
  NAND2_X1 U10192 ( .A1(n8887), .A2(n9047), .ZN(n8788) );
  OAI21_X1 U10193 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n8789), .A(n8788), .ZN(
        n8791) );
  OAI22_X1 U10194 ( .A1(n8846), .A2(n9078), .B1(n9112), .B2(n8891), .ZN(n8790)
         );
  AOI211_X1 U10195 ( .C1(n9194), .C2(n8894), .A(n8791), .B(n8790), .ZN(n8792)
         );
  OAI21_X1 U10196 ( .B1(n8793), .B2(n8897), .A(n8792), .ZN(P1_U3223) );
  OAI21_X1 U10197 ( .B1(n8795), .B2(n8794), .A(n8871), .ZN(n8796) );
  NAND2_X1 U10198 ( .A1(n8796), .A2(n8876), .ZN(n8803) );
  NOR2_X1 U10199 ( .A1(n8797), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8801) );
  INV_X1 U10200 ( .A(n9013), .ZN(n8799) );
  OAI22_X1 U10201 ( .A1(n8846), .A2(n8799), .B1(n8798), .B2(n8891), .ZN(n8800)
         );
  AOI211_X1 U10202 ( .C1(n8887), .C2(n9020), .A(n8801), .B(n8800), .ZN(n8802)
         );
  OAI211_X1 U10203 ( .C1(n9015), .C2(n8851), .A(n8803), .B(n8802), .ZN(
        P1_U3225) );
  OAI21_X1 U10204 ( .B1(n8806), .B2(n8804), .A(n8805), .ZN(n8807) );
  NAND2_X1 U10205 ( .A1(n8807), .A2(n8876), .ZN(n8813) );
  AND2_X1 U10206 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8943) );
  INV_X1 U10207 ( .A(n8808), .ZN(n8810) );
  OAI22_X1 U10208 ( .A1(n8846), .A2(n8810), .B1(n8809), .B2(n8891), .ZN(n8811)
         );
  AOI211_X1 U10209 ( .C1(n8887), .C2(n9124), .A(n8943), .B(n8811), .ZN(n8812)
         );
  OAI211_X1 U10210 ( .C1(n8814), .C2(n8851), .A(n8813), .B(n8812), .ZN(
        P1_U3226) );
  NAND2_X1 U10211 ( .A1(n4355), .A2(n8815), .ZN(n8816) );
  XNOR2_X1 U10212 ( .A(n8817), .B(n8816), .ZN(n8821) );
  AOI22_X1 U10213 ( .A1(n8889), .A2(n9135), .B1(n8878), .B2(n8903), .ZN(n8818)
         );
  NAND2_X1 U10214 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9595) );
  OAI211_X1 U10215 ( .C1(n9144), .C2(n8867), .A(n8818), .B(n9595), .ZN(n8819)
         );
  AOI21_X1 U10216 ( .B1(n9213), .B2(n8894), .A(n8819), .ZN(n8820) );
  OAI21_X1 U10217 ( .B1(n8821), .B2(n8897), .A(n8820), .ZN(P1_U3228) );
  OAI21_X1 U10218 ( .B1(n8824), .B2(n8822), .A(n8823), .ZN(n8825) );
  NAND2_X1 U10219 ( .A1(n8825), .A2(n8876), .ZN(n8832) );
  NOR2_X1 U10220 ( .A1(n8826), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8830) );
  INV_X1 U10221 ( .A(n9028), .ZN(n8828) );
  OAI22_X1 U10222 ( .A1(n8846), .A2(n8828), .B1(n8827), .B2(n8891), .ZN(n8829)
         );
  AOI211_X1 U10223 ( .C1(n8887), .C2(n9036), .A(n8830), .B(n8829), .ZN(n8831)
         );
  OAI211_X1 U10224 ( .C1(n9030), .C2(n8851), .A(n8832), .B(n8831), .ZN(
        P1_U3229) );
  OAI211_X1 U10225 ( .C1(n8835), .C2(n8834), .A(n8833), .B(n8876), .ZN(n8839)
         );
  AOI22_X1 U10226 ( .A1(n8878), .A2(n5754), .B1(n8887), .B2(n9653), .ZN(n8838)
         );
  AND2_X1 U10227 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9485) );
  NOR2_X1 U10228 ( .A1(n8851), .A2(n9701), .ZN(n8836) );
  AOI211_X1 U10229 ( .C1(n9657), .C2(n8889), .A(n9485), .B(n8836), .ZN(n8837)
         );
  NAND3_X1 U10230 ( .A1(n8839), .A2(n8838), .A3(n8837), .ZN(P1_U3230) );
  NAND2_X1 U10231 ( .A1(n8841), .A2(n8840), .ZN(n8842) );
  OAI21_X1 U10232 ( .B1(n8843), .B2(n8842), .A(n8784), .ZN(n8844) );
  NAND2_X1 U10233 ( .A1(n8844), .A2(n8876), .ZN(n8850) );
  NOR2_X1 U10234 ( .A1(n8845), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8848) );
  OAI22_X1 U10235 ( .A1(n8846), .A2(n9092), .B1(n9089), .B2(n8891), .ZN(n8847)
         );
  AOI211_X1 U10236 ( .C1(n8887), .C2(n9059), .A(n8848), .B(n8847), .ZN(n8849)
         );
  OAI211_X1 U10237 ( .C1(n9096), .C2(n8851), .A(n8850), .B(n8849), .ZN(
        P1_U3233) );
  AOI21_X1 U10238 ( .B1(n8852), .B2(n8854), .A(n8853), .ZN(n8860) );
  AOI22_X1 U10239 ( .A1(n8889), .A2(n9056), .B1(n8878), .B2(n9059), .ZN(n8856)
         );
  NAND2_X1 U10240 ( .A1(n8887), .A2(n9065), .ZN(n8855) );
  OAI211_X1 U10241 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n8857), .A(n8856), .B(
        n8855), .ZN(n8858) );
  AOI21_X1 U10242 ( .B1(n9188), .B2(n8894), .A(n8858), .ZN(n8859) );
  OAI21_X1 U10243 ( .B1(n8860), .B2(n8897), .A(n8859), .ZN(P1_U3235) );
  XNOR2_X1 U10244 ( .A(n8863), .B(n8862), .ZN(n8864) );
  XNOR2_X1 U10245 ( .A(n8861), .B(n8864), .ZN(n8870) );
  INV_X1 U10246 ( .A(n8865), .ZN(n9118) );
  AOI22_X1 U10247 ( .A1(n8889), .A2(n9118), .B1(n8878), .B2(n9124), .ZN(n8866)
         );
  NAND2_X1 U10248 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9611) );
  OAI211_X1 U10249 ( .C1(n9089), .C2(n8867), .A(n8866), .B(n9611), .ZN(n8868)
         );
  AOI21_X1 U10250 ( .B1(n9208), .B2(n8894), .A(n8868), .ZN(n8869) );
  OAI21_X1 U10251 ( .B1(n8870), .B2(n8897), .A(n8869), .ZN(P1_U3238) );
  INV_X1 U10252 ( .A(n8871), .ZN(n8874) );
  NAND3_X1 U10253 ( .A1(n8877), .A2(n8876), .A3(n8875), .ZN(n8882) );
  AOI22_X1 U10254 ( .A1(n8887), .A2(n9005), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8881) );
  AOI22_X1 U10255 ( .A1(n8889), .A2(n8999), .B1(n8878), .B2(n9036), .ZN(n8880)
         );
  NAND2_X1 U10256 ( .A1(n9168), .A2(n8894), .ZN(n8879) );
  NAND4_X1 U10257 ( .A1(n8882), .A2(n8881), .A3(n8880), .A4(n8879), .ZN(
        P1_U3240) );
  INV_X1 U10258 ( .A(n8884), .ZN(n8885) );
  AOI21_X1 U10259 ( .B1(n8883), .B2(n8886), .A(n8885), .ZN(n8898) );
  AOI22_X1 U10260 ( .A1(n8889), .A2(n8888), .B1(n8887), .B2(n8903), .ZN(n8890)
         );
  NAND2_X1 U10261 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9582) );
  OAI211_X1 U10262 ( .C1(n8892), .C2(n8891), .A(n8890), .B(n9582), .ZN(n8893)
         );
  AOI21_X1 U10263 ( .B1(n8895), .B2(n8894), .A(n8893), .ZN(n8896) );
  OAI21_X1 U10264 ( .B1(n8898), .B2(n8897), .A(n8896), .ZN(P1_U3241) );
  MUX2_X1 U10265 ( .A(n8972), .B(P1_DATAO_REG_31__SCAN_IN), .S(n8913), .Z(
        P1_U3585) );
  MUX2_X1 U10266 ( .A(n8899), .B(P1_DATAO_REG_30__SCAN_IN), .S(n8913), .Z(
        P1_U3584) );
  MUX2_X1 U10267 ( .A(n8900), .B(P1_DATAO_REG_29__SCAN_IN), .S(n8913), .Z(
        P1_U3583) );
  MUX2_X1 U10268 ( .A(n8985), .B(P1_DATAO_REG_28__SCAN_IN), .S(n8913), .Z(
        P1_U3582) );
  MUX2_X1 U10269 ( .A(n9005), .B(P1_DATAO_REG_27__SCAN_IN), .S(n8913), .Z(
        P1_U3581) );
  MUX2_X1 U10270 ( .A(n9020), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8913), .Z(
        P1_U3580) );
  MUX2_X1 U10271 ( .A(n9036), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8913), .Z(
        P1_U3579) );
  MUX2_X1 U10272 ( .A(n9048), .B(P1_DATAO_REG_24__SCAN_IN), .S(n8913), .Z(
        P1_U3578) );
  MUX2_X1 U10273 ( .A(n9065), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8913), .Z(
        P1_U3577) );
  MUX2_X1 U10274 ( .A(n9047), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8913), .Z(
        P1_U3576) );
  MUX2_X1 U10275 ( .A(n9059), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8913), .Z(
        P1_U3575) );
  MUX2_X1 U10276 ( .A(n8901), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8913), .Z(
        P1_U3574) );
  MUX2_X1 U10277 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9125), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10278 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n8902), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10279 ( .A(n9124), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8913), .Z(
        P1_U3571) );
  MUX2_X1 U10280 ( .A(n8903), .B(P1_DATAO_REG_16__SCAN_IN), .S(n8913), .Z(
        P1_U3570) );
  MUX2_X1 U10281 ( .A(n8904), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8913), .Z(
        P1_U3569) );
  MUX2_X1 U10282 ( .A(n8905), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8913), .Z(
        P1_U3568) );
  MUX2_X1 U10283 ( .A(n8906), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8913), .Z(
        P1_U3567) );
  MUX2_X1 U10284 ( .A(n8907), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8913), .Z(
        P1_U3565) );
  MUX2_X1 U10285 ( .A(n8908), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8913), .Z(
        P1_U3564) );
  MUX2_X1 U10286 ( .A(n8909), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8913), .Z(
        P1_U3563) );
  MUX2_X1 U10287 ( .A(n8910), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8913), .Z(
        P1_U3562) );
  MUX2_X1 U10288 ( .A(n9637), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8913), .Z(
        P1_U3561) );
  MUX2_X1 U10289 ( .A(n8911), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8913), .Z(
        P1_U3560) );
  MUX2_X1 U10290 ( .A(n9653), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8913), .Z(
        P1_U3559) );
  MUX2_X1 U10291 ( .A(n8912), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8913), .Z(
        P1_U3558) );
  MUX2_X1 U10292 ( .A(n5754), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8913), .Z(
        P1_U3557) );
  MUX2_X1 U10293 ( .A(n5732), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8913), .Z(
        P1_U3555) );
  MUX2_X1 U10294 ( .A(n5740), .B(P1_DATAO_REG_0__SCAN_IN), .S(n8913), .Z(
        P1_U3554) );
  OAI211_X1 U10295 ( .C1(n8915), .C2(n9477), .A(n9598), .B(n8914), .ZN(n8922)
         );
  OAI211_X1 U10296 ( .C1(n8918), .C2(n8917), .A(n9591), .B(n8916), .ZN(n8921)
         );
  AOI22_X1 U10297 ( .A1(n9486), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n8920) );
  INV_X1 U10298 ( .A(n9543), .ZN(n9605) );
  NAND2_X1 U10299 ( .A1(n9605), .A2(n4916), .ZN(n8919) );
  NAND4_X1 U10300 ( .A1(n8922), .A2(n8921), .A3(n8920), .A4(n8919), .ZN(
        P1_U3244) );
  NAND2_X1 U10301 ( .A1(n8955), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8923) );
  OAI21_X1 U10302 ( .B1(n8955), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8923), .ZN(
        n8932) );
  INV_X1 U10303 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9798) );
  NOR2_X1 U10304 ( .A1(n9556), .A2(n9798), .ZN(n8925) );
  AOI21_X1 U10305 ( .B1(n9556), .B2(n9798), .A(n8925), .ZN(n9550) );
  INV_X1 U10306 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9801) );
  NOR2_X1 U10307 ( .A1(n9568), .A2(n9801), .ZN(n8926) );
  AOI21_X1 U10308 ( .B1(n9568), .B2(n9801), .A(n8926), .ZN(n9562) );
  NOR2_X1 U10309 ( .A1(n9561), .A2(n9562), .ZN(n9560) );
  NOR2_X1 U10310 ( .A1(n8927), .A2(n8937), .ZN(n8928) );
  XNOR2_X1 U10311 ( .A(n8937), .B(n8927), .ZN(n9573) );
  NOR2_X1 U10312 ( .A1(n9574), .A2(n9573), .ZN(n9572) );
  NOR2_X1 U10313 ( .A1(n8928), .A2(n9572), .ZN(n8929) );
  INV_X1 U10314 ( .A(n8954), .ZN(n8930) );
  AOI21_X1 U10315 ( .B1(n8932), .B2(n8931), .A(n8930), .ZN(n8946) );
  OAI21_X1 U10316 ( .B1(n8934), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8933), .ZN(
        n9553) );
  XNOR2_X1 U10317 ( .A(n9556), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n9552) );
  NOR2_X1 U10318 ( .A1(n9553), .A2(n9552), .ZN(n9551) );
  NAND2_X1 U10319 ( .A1(n9568), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8935) );
  OAI21_X1 U10320 ( .B1(n9568), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8935), .ZN(
        n9564) );
  NOR2_X1 U10321 ( .A1(n8936), .A2(n8937), .ZN(n8938) );
  INV_X1 U10322 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9577) );
  NOR2_X1 U10323 ( .A1(n9577), .A2(n9578), .ZN(n9576) );
  NOR2_X1 U10324 ( .A1(n8938), .A2(n9576), .ZN(n8941) );
  XNOR2_X1 U10325 ( .A(n8955), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n8940) );
  INV_X1 U10326 ( .A(n8948), .ZN(n8939) );
  AOI211_X1 U10327 ( .C1(n8941), .C2(n8940), .A(n8939), .B(n9575), .ZN(n8942)
         );
  AOI211_X1 U10328 ( .C1(n9486), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n8943), .B(
        n8942), .ZN(n8945) );
  NAND2_X1 U10329 ( .A1(n9605), .A2(n8955), .ZN(n8944) );
  OAI211_X1 U10330 ( .C1(n8946), .C2(n9602), .A(n8945), .B(n8944), .ZN(
        P1_U3259) );
  NAND2_X1 U10331 ( .A1(n8955), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8947) );
  INV_X1 U10332 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8949) );
  XNOR2_X1 U10333 ( .A(n9593), .B(n8949), .ZN(n9587) );
  OR2_X1 U10334 ( .A1(n9593), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8950) );
  OR2_X1 U10335 ( .A1(n9606), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U10336 ( .A1(n9606), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8952) );
  AND2_X1 U10337 ( .A1(n8951), .A2(n8952), .ZN(n9600) );
  NAND2_X1 U10338 ( .A1(n9599), .A2(n8952), .ZN(n8953) );
  INV_X1 U10339 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9106) );
  XNOR2_X1 U10340 ( .A(n8953), .B(n9106), .ZN(n8961) );
  INV_X1 U10341 ( .A(n8961), .ZN(n8959) );
  NOR2_X1 U10342 ( .A1(n9593), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8956) );
  AOI21_X1 U10343 ( .B1(n9593), .B2(P1_REG1_REG_17__SCAN_IN), .A(n8956), .ZN(
        n9590) );
  OAI21_X1 U10344 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9593), .A(n9588), .ZN(
        n9604) );
  NAND2_X1 U10345 ( .A1(n9606), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8957) );
  OAI21_X1 U10346 ( .B1(n9606), .B2(P1_REG1_REG_18__SCAN_IN), .A(n8957), .ZN(
        n9603) );
  AOI21_X1 U10347 ( .B1(n8959), .B2(n9598), .A(n8958), .ZN(n8963) );
  AOI22_X1 U10348 ( .A1(n8961), .A2(n9598), .B1(n9591), .B2(n8960), .ZN(n8962)
         );
  MUX2_X1 U10349 ( .A(n8963), .B(n8962), .S(n7928), .Z(n8966) );
  INV_X1 U10350 ( .A(n8964), .ZN(n8965) );
  OAI211_X1 U10351 ( .C1(n6985), .C2(n9613), .A(n8966), .B(n8965), .ZN(
        P1_U3262) );
  XNOR2_X1 U10352 ( .A(n8969), .B(n8975), .ZN(n8970) );
  NAND2_X1 U10353 ( .A1(n8970), .A2(n9666), .ZN(n9153) );
  NAND2_X1 U10354 ( .A1(n8972), .A2(n8971), .ZN(n9155) );
  NOR2_X1 U10355 ( .A1(n9658), .A2(n9155), .ZN(n8980) );
  NOR2_X1 U10356 ( .A1(n9154), .A2(n9660), .ZN(n8973) );
  AOI211_X1 U10357 ( .C1(n9658), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8980), .B(
        n8973), .ZN(n8974) );
  OAI21_X1 U10358 ( .B1(n9153), .B2(n8982), .A(n8974), .ZN(P1_U3263) );
  AOI211_X1 U10359 ( .C1(n8978), .C2(n8976), .A(n8975), .B(n9769), .ZN(n8977)
         );
  INV_X1 U10360 ( .A(n8977), .ZN(n9156) );
  NOR2_X1 U10361 ( .A1(n4524), .A2(n9660), .ZN(n8979) );
  AOI211_X1 U10362 ( .C1(n9658), .C2(P1_REG2_REG_30__SCAN_IN), .A(n8980), .B(
        n8979), .ZN(n8981) );
  OAI21_X1 U10363 ( .B1(n9156), .B2(n8982), .A(n8981), .ZN(P1_U3264) );
  XNOR2_X1 U10364 ( .A(n8983), .B(n8984), .ZN(n9166) );
  OAI21_X1 U10365 ( .B1(n4303), .B2(n8984), .A(n9655), .ZN(n8987) );
  AOI22_X1 U10366 ( .A1(n9651), .A2(n9020), .B1(n8985), .B2(n9652), .ZN(n8986)
         );
  OAI21_X1 U10367 ( .B1(n8987), .B2(n4318), .A(n8986), .ZN(n9162) );
  INV_X1 U10368 ( .A(n8998), .ZN(n8990) );
  INV_X1 U10369 ( .A(n8988), .ZN(n8989) );
  AOI211_X1 U10370 ( .C1(n9164), .C2(n8990), .A(n9769), .B(n8989), .ZN(n9163)
         );
  NAND2_X1 U10371 ( .A1(n9163), .A2(n9669), .ZN(n8993) );
  AOI22_X1 U10372 ( .A1(n9658), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n8991), .B2(
        n9656), .ZN(n8992) );
  OAI211_X1 U10373 ( .C1(n8994), .C2(n9660), .A(n8993), .B(n8992), .ZN(n8995)
         );
  AOI21_X1 U10374 ( .B1(n9162), .B2(n9113), .A(n8995), .ZN(n8996) );
  OAI21_X1 U10375 ( .B1(n9166), .B2(n9152), .A(n8996), .ZN(P1_U3266) );
  XNOR2_X1 U10376 ( .A(n8997), .B(n9003), .ZN(n9171) );
  AOI211_X1 U10377 ( .C1(n9168), .C2(n9011), .A(n9769), .B(n8998), .ZN(n9167)
         );
  AOI22_X1 U10378 ( .A1(n9673), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9656), .B2(
        n8999), .ZN(n9000) );
  OAI21_X1 U10379 ( .B1(n9001), .B2(n9660), .A(n9000), .ZN(n9008) );
  OAI21_X1 U10380 ( .B1(n9004), .B2(n9003), .A(n9002), .ZN(n9006) );
  AOI222_X1 U10381 ( .A1(n9655), .A2(n9006), .B1(n9005), .B2(n9652), .C1(n9036), .C2(n9651), .ZN(n9170) );
  NOR2_X1 U10382 ( .A1(n9170), .A2(n9673), .ZN(n9007) );
  AOI211_X1 U10383 ( .C1(n9167), .C2(n9669), .A(n9008), .B(n9007), .ZN(n9009)
         );
  OAI21_X1 U10384 ( .B1(n9171), .B2(n9152), .A(n9009), .ZN(P1_U3267) );
  XNOR2_X1 U10385 ( .A(n9010), .B(n9017), .ZN(n9176) );
  INV_X1 U10386 ( .A(n9011), .ZN(n9012) );
  AOI211_X1 U10387 ( .C1(n9173), .C2(n9025), .A(n9769), .B(n9012), .ZN(n9172)
         );
  AOI22_X1 U10388 ( .A1(n9658), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9013), .B2(
        n9656), .ZN(n9014) );
  OAI21_X1 U10389 ( .B1(n9015), .B2(n9660), .A(n9014), .ZN(n9022) );
  AND2_X1 U10390 ( .A1(n9048), .A2(n9651), .ZN(n9019) );
  AOI211_X1 U10391 ( .C1(n4306), .C2(n9017), .A(n9138), .B(n9016), .ZN(n9018)
         );
  AOI211_X1 U10392 ( .C1(n9652), .C2(n9020), .A(n9019), .B(n9018), .ZN(n9175)
         );
  NOR2_X1 U10393 ( .A1(n9175), .A2(n9658), .ZN(n9021) );
  AOI211_X1 U10394 ( .C1(n9172), .C2(n9669), .A(n9022), .B(n9021), .ZN(n9023)
         );
  OAI21_X1 U10395 ( .B1(n9176), .B2(n9152), .A(n9023), .ZN(P1_U3268) );
  XNOR2_X1 U10396 ( .A(n9024), .B(n4617), .ZN(n9181) );
  INV_X1 U10397 ( .A(n9025), .ZN(n9026) );
  AOI211_X1 U10398 ( .C1(n9178), .C2(n4533), .A(n9769), .B(n9026), .ZN(n9177)
         );
  NOR2_X1 U10399 ( .A1(n9673), .A2(n9027), .ZN(n9150) );
  AOI22_X1 U10400 ( .A1(n9658), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9028), .B2(
        n9656), .ZN(n9029) );
  OAI21_X1 U10401 ( .B1(n9030), .B2(n9660), .A(n9029), .ZN(n9038) );
  AND2_X1 U10402 ( .A1(n9065), .A2(n9651), .ZN(n9035) );
  AOI211_X1 U10403 ( .C1(n9033), .C2(n9032), .A(n9138), .B(n9031), .ZN(n9034)
         );
  AOI211_X1 U10404 ( .C1(n9652), .C2(n9036), .A(n9035), .B(n9034), .ZN(n9180)
         );
  NOR2_X1 U10405 ( .A1(n9180), .A2(n9658), .ZN(n9037) );
  AOI211_X1 U10406 ( .C1(n9177), .C2(n9150), .A(n9038), .B(n9037), .ZN(n9039)
         );
  OAI21_X1 U10407 ( .B1(n9152), .B2(n9181), .A(n9039), .ZN(P1_U3269) );
  XNOR2_X1 U10408 ( .A(n9040), .B(n9046), .ZN(n9186) );
  AOI211_X1 U10409 ( .C1(n9183), .C2(n9054), .A(n9769), .B(n9041), .ZN(n9182)
         );
  AOI22_X1 U10410 ( .A1(n9658), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9042), .B2(
        n9656), .ZN(n9043) );
  OAI21_X1 U10411 ( .B1(n4531), .B2(n9660), .A(n9043), .ZN(n9051) );
  OAI21_X1 U10412 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9049) );
  AOI222_X1 U10413 ( .A1(n9655), .A2(n9049), .B1(n9048), .B2(n9652), .C1(n9047), .C2(n9651), .ZN(n9185) );
  NOR2_X1 U10414 ( .A1(n9185), .A2(n9658), .ZN(n9050) );
  AOI211_X1 U10415 ( .C1(n9182), .C2(n9669), .A(n9051), .B(n9050), .ZN(n9052)
         );
  OAI21_X1 U10416 ( .B1(n9186), .B2(n9152), .A(n9052), .ZN(P1_U3270) );
  XNOR2_X1 U10417 ( .A(n9053), .B(n9062), .ZN(n9191) );
  INV_X1 U10418 ( .A(n9054), .ZN(n9055) );
  AOI211_X1 U10419 ( .C1(n9188), .C2(n9075), .A(n9769), .B(n9055), .ZN(n9187)
         );
  AOI22_X1 U10420 ( .A1(n9658), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9056), .B2(
        n9656), .ZN(n9057) );
  OAI21_X1 U10421 ( .B1(n9058), .B2(n9660), .A(n9057), .ZN(n9067) );
  AND2_X1 U10422 ( .A1(n9059), .A2(n9651), .ZN(n9064) );
  AOI211_X1 U10423 ( .C1(n9062), .C2(n9061), .A(n9138), .B(n9060), .ZN(n9063)
         );
  AOI211_X1 U10424 ( .C1(n9652), .C2(n9065), .A(n9064), .B(n9063), .ZN(n9190)
         );
  NOR2_X1 U10425 ( .A1(n9190), .A2(n9673), .ZN(n9066) );
  AOI211_X1 U10426 ( .C1(n9187), .C2(n9669), .A(n9067), .B(n9066), .ZN(n9068)
         );
  OAI21_X1 U10427 ( .B1(n9191), .B2(n9152), .A(n9068), .ZN(P1_U3271) );
  XNOR2_X1 U10428 ( .A(n9069), .B(n9071), .ZN(n9196) );
  AOI21_X1 U10429 ( .B1(n9087), .B2(n9086), .A(n9070), .ZN(n9072) );
  XNOR2_X1 U10430 ( .A(n9072), .B(n9071), .ZN(n9073) );
  OAI222_X1 U10431 ( .A1(n9616), .A2(n9074), .B1(n9618), .B2(n9112), .C1(n9073), .C2(n9138), .ZN(n9192) );
  INV_X1 U10432 ( .A(n9091), .ZN(n9077) );
  INV_X1 U10433 ( .A(n9075), .ZN(n9076) );
  AOI211_X1 U10434 ( .C1(n9194), .C2(n9077), .A(n9769), .B(n9076), .ZN(n9193)
         );
  NAND2_X1 U10435 ( .A1(n9193), .A2(n9150), .ZN(n9081) );
  INV_X1 U10436 ( .A(n9078), .ZN(n9079) );
  AOI22_X1 U10437 ( .A1(n9658), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9079), .B2(
        n9656), .ZN(n9080) );
  OAI211_X1 U10438 ( .C1(n9082), .C2(n9660), .A(n9081), .B(n9080), .ZN(n9083)
         );
  AOI21_X1 U10439 ( .B1(n9192), .B2(n9113), .A(n9083), .ZN(n9084) );
  OAI21_X1 U10440 ( .B1(n9196), .B2(n9152), .A(n9084), .ZN(P1_U3272) );
  XOR2_X1 U10441 ( .A(n9086), .B(n9085), .Z(n9201) );
  XNOR2_X1 U10442 ( .A(n9087), .B(n9086), .ZN(n9088) );
  OAI222_X1 U10443 ( .A1(n9616), .A2(n9090), .B1(n9618), .B2(n9089), .C1(n9138), .C2(n9088), .ZN(n9197) );
  AOI211_X1 U10444 ( .C1(n9199), .C2(n9100), .A(n9769), .B(n9091), .ZN(n9198)
         );
  NAND2_X1 U10445 ( .A1(n9198), .A2(n9669), .ZN(n9095) );
  INV_X1 U10446 ( .A(n9092), .ZN(n9093) );
  AOI22_X1 U10447 ( .A1(n9658), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9093), .B2(
        n9656), .ZN(n9094) );
  OAI211_X1 U10448 ( .C1(n9096), .C2(n9660), .A(n9095), .B(n9094), .ZN(n9097)
         );
  AOI21_X1 U10449 ( .B1(n9197), .B2(n9113), .A(n9097), .ZN(n9098) );
  OAI21_X1 U10450 ( .B1(n9201), .B2(n9152), .A(n9098), .ZN(P1_U3273) );
  XOR2_X1 U10451 ( .A(n9099), .B(n9109), .Z(n9206) );
  INV_X1 U10452 ( .A(n9117), .ZN(n9102) );
  INV_X1 U10453 ( .A(n9100), .ZN(n9101) );
  AOI211_X1 U10454 ( .C1(n9204), .C2(n9102), .A(n9769), .B(n9101), .ZN(n9203)
         );
  NOR2_X1 U10455 ( .A1(n9103), .A2(n9660), .ZN(n9108) );
  OAI22_X1 U10456 ( .A1(n9113), .A2(n9106), .B1(n9105), .B2(n9104), .ZN(n9107)
         );
  AOI211_X1 U10457 ( .C1(n9203), .C2(n9669), .A(n9108), .B(n9107), .ZN(n9115)
         );
  XOR2_X1 U10458 ( .A(n9110), .B(n9109), .Z(n9111) );
  OAI222_X1 U10459 ( .A1(n9616), .A2(n9112), .B1(n9618), .B2(n9144), .C1(n9111), .C2(n9138), .ZN(n9202) );
  NAND2_X1 U10460 ( .A1(n9202), .A2(n9113), .ZN(n9114) );
  OAI211_X1 U10461 ( .C1(n9206), .C2(n9152), .A(n9115), .B(n9114), .ZN(
        P1_U3274) );
  XOR2_X1 U10462 ( .A(n9116), .B(n9122), .Z(n9211) );
  AOI211_X1 U10463 ( .C1(n9208), .C2(n9133), .A(n9769), .B(n9117), .ZN(n9207)
         );
  AOI22_X1 U10464 ( .A1(n9658), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9118), .B2(
        n9656), .ZN(n9119) );
  OAI21_X1 U10465 ( .B1(n9120), .B2(n9660), .A(n9119), .ZN(n9128) );
  OAI21_X1 U10466 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(n9126) );
  AOI222_X1 U10467 ( .A1(n9655), .A2(n9126), .B1(n9125), .B2(n9652), .C1(n9124), .C2(n9651), .ZN(n9210) );
  NOR2_X1 U10468 ( .A1(n9210), .A2(n9673), .ZN(n9127) );
  AOI211_X1 U10469 ( .C1(n9207), .C2(n9669), .A(n9128), .B(n9127), .ZN(n9129)
         );
  OAI21_X1 U10470 ( .B1(n9211), .B2(n9152), .A(n9129), .ZN(P1_U3275) );
  XNOR2_X1 U10471 ( .A(n9131), .B(n9130), .ZN(n9216) );
  INV_X1 U10472 ( .A(n9132), .ZN(n9134) );
  AOI211_X1 U10473 ( .C1(n9213), .C2(n9134), .A(n9769), .B(n4534), .ZN(n9212)
         );
  AOI22_X1 U10474 ( .A1(n9673), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9135), .B2(
        n9656), .ZN(n9136) );
  OAI21_X1 U10475 ( .B1(n9137), .B2(n9660), .A(n9136), .ZN(n9149) );
  NOR2_X1 U10476 ( .A1(n9139), .A2(n9138), .ZN(n9147) );
  OAI21_X1 U10477 ( .B1(n9142), .B2(n9141), .A(n9140), .ZN(n9146) );
  OAI22_X1 U10478 ( .A1(n9144), .A2(n9616), .B1(n9143), .B2(n9618), .ZN(n9145)
         );
  AOI21_X1 U10479 ( .B1(n9147), .B2(n9146), .A(n9145), .ZN(n9215) );
  NOR2_X1 U10480 ( .A1(n9215), .A2(n9673), .ZN(n9148) );
  AOI211_X1 U10481 ( .C1(n9212), .C2(n9150), .A(n9149), .B(n9148), .ZN(n9151)
         );
  OAI21_X1 U10482 ( .B1(n9152), .B2(n9216), .A(n9151), .ZN(P1_U3276) );
  OAI211_X1 U10483 ( .C1(n9154), .C2(n9767), .A(n9153), .B(n9155), .ZN(n9224)
         );
  MUX2_X1 U10484 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9224), .S(n9803), .Z(
        P1_U3553) );
  OAI211_X1 U10485 ( .C1(n4524), .C2(n9767), .A(n9156), .B(n9155), .ZN(n9225)
         );
  MUX2_X1 U10486 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9225), .S(n9803), .Z(
        P1_U3552) );
  AOI22_X1 U10487 ( .A1(n9158), .A2(n9666), .B1(n9734), .B2(n9157), .ZN(n9159)
         );
  OAI211_X1 U10488 ( .C1(n9161), .C2(n9222), .A(n9160), .B(n9159), .ZN(n9366)
         );
  MUX2_X1 U10489 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9366), .S(n9803), .Z(
        P1_U3550) );
  AOI211_X1 U10490 ( .C1(n9734), .C2(n9164), .A(n9163), .B(n9162), .ZN(n9165)
         );
  OAI21_X1 U10491 ( .B1(n9166), .B2(n9222), .A(n9165), .ZN(n9367) );
  MUX2_X1 U10492 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9367), .S(n9803), .Z(
        P1_U3549) );
  AOI21_X1 U10493 ( .B1(n9734), .B2(n9168), .A(n9167), .ZN(n9169) );
  OAI211_X1 U10494 ( .C1(n9171), .C2(n9222), .A(n9170), .B(n9169), .ZN(n9368)
         );
  MUX2_X1 U10495 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9368), .S(n9803), .Z(
        P1_U3548) );
  AOI21_X1 U10496 ( .B1(n9734), .B2(n9173), .A(n9172), .ZN(n9174) );
  OAI211_X1 U10497 ( .C1(n9176), .C2(n9222), .A(n9175), .B(n9174), .ZN(n9369)
         );
  MUX2_X1 U10498 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9369), .S(n9803), .Z(
        P1_U3547) );
  AOI21_X1 U10499 ( .B1(n9734), .B2(n9178), .A(n9177), .ZN(n9179) );
  OAI211_X1 U10500 ( .C1(n9181), .C2(n9222), .A(n9180), .B(n9179), .ZN(n9370)
         );
  MUX2_X1 U10501 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9370), .S(n9803), .Z(
        P1_U3546) );
  AOI21_X1 U10502 ( .B1(n9734), .B2(n9183), .A(n9182), .ZN(n9184) );
  OAI211_X1 U10503 ( .C1(n9186), .C2(n9222), .A(n9185), .B(n9184), .ZN(n9371)
         );
  MUX2_X1 U10504 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9371), .S(n9803), .Z(
        P1_U3545) );
  AOI21_X1 U10505 ( .B1(n9734), .B2(n9188), .A(n9187), .ZN(n9189) );
  OAI211_X1 U10506 ( .C1(n9191), .C2(n9222), .A(n9190), .B(n9189), .ZN(n9372)
         );
  MUX2_X1 U10507 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9372), .S(n9803), .Z(
        P1_U3544) );
  AOI211_X1 U10508 ( .C1(n9734), .C2(n9194), .A(n9193), .B(n9192), .ZN(n9195)
         );
  OAI21_X1 U10509 ( .B1(n9196), .B2(n9222), .A(n9195), .ZN(n9373) );
  MUX2_X1 U10510 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9373), .S(n9803), .Z(
        P1_U3543) );
  AOI211_X1 U10511 ( .C1(n9734), .C2(n9199), .A(n9198), .B(n9197), .ZN(n9200)
         );
  OAI21_X1 U10512 ( .B1(n9222), .B2(n9201), .A(n9200), .ZN(n9374) );
  MUX2_X1 U10513 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9374), .S(n9803), .Z(
        P1_U3542) );
  AOI211_X1 U10514 ( .C1(n9734), .C2(n9204), .A(n9203), .B(n9202), .ZN(n9205)
         );
  OAI21_X1 U10515 ( .B1(n9222), .B2(n9206), .A(n9205), .ZN(n9375) );
  MUX2_X1 U10516 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9375), .S(n9803), .Z(
        P1_U3541) );
  AOI21_X1 U10517 ( .B1(n9734), .B2(n9208), .A(n9207), .ZN(n9209) );
  OAI211_X1 U10518 ( .C1(n9211), .C2(n9222), .A(n9210), .B(n9209), .ZN(n9376)
         );
  MUX2_X1 U10519 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9376), .S(n9803), .Z(
        P1_U3540) );
  AOI21_X1 U10520 ( .B1(n9734), .B2(n9213), .A(n9212), .ZN(n9214) );
  OAI211_X1 U10521 ( .C1(n9216), .C2(n9222), .A(n9215), .B(n9214), .ZN(n9377)
         );
  MUX2_X1 U10522 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9377), .S(n9803), .Z(
        P1_U3539) );
  AOI211_X1 U10523 ( .C1(n9734), .C2(n9219), .A(n9218), .B(n9217), .ZN(n9220)
         );
  OAI21_X1 U10524 ( .B1(n9222), .B2(n9221), .A(n9220), .ZN(n9378) );
  MUX2_X1 U10525 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9378), .S(n9803), .Z(
        P1_U3538) );
  MUX2_X1 U10526 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9223), .S(n9803), .Z(
        P1_U3522) );
  MUX2_X1 U10527 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9224), .S(n9777), .Z(
        P1_U3521) );
  AOI22_X1 U10528 ( .A1(n6474), .A2(keyinput19), .B1(n5222), .B2(keyinput60), 
        .ZN(n9226) );
  OAI221_X1 U10529 ( .B1(n6474), .B2(keyinput19), .C1(n5222), .C2(keyinput60), 
        .A(n9226), .ZN(n9234) );
  AOI22_X1 U10530 ( .A1(n9229), .A2(keyinput49), .B1(n9228), .B2(keyinput39), 
        .ZN(n9227) );
  OAI221_X1 U10531 ( .B1(n9229), .B2(keyinput49), .C1(n9228), .C2(keyinput39), 
        .A(n9227), .ZN(n9233) );
  INV_X1 U10532 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9230) );
  XNOR2_X1 U10533 ( .A(keyinput16), .B(n9230), .ZN(n9232) );
  INV_X1 U10534 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9336) );
  XNOR2_X1 U10535 ( .A(keyinput17), .B(n9336), .ZN(n9231) );
  OR4_X1 U10536 ( .A1(n9234), .A2(n9233), .A3(n9232), .A4(n9231), .ZN(n9242)
         );
  AOI22_X1 U10537 ( .A1(n9792), .A2(keyinput62), .B1(n9236), .B2(keyinput47), 
        .ZN(n9235) );
  OAI221_X1 U10538 ( .B1(n9792), .B2(keyinput62), .C1(n9236), .C2(keyinput47), 
        .A(n9235), .ZN(n9241) );
  AOI22_X1 U10539 ( .A1(n9239), .A2(keyinput11), .B1(keyinput30), .B2(n9238), 
        .ZN(n9237) );
  OAI221_X1 U10540 ( .B1(n9239), .B2(keyinput11), .C1(n9238), .C2(keyinput30), 
        .A(n9237), .ZN(n9240) );
  NOR3_X1 U10541 ( .A1(n9242), .A2(n9241), .A3(n9240), .ZN(n9294) );
  AOI22_X1 U10542 ( .A1(n9245), .A2(keyinput63), .B1(keyinput22), .B2(n9244), 
        .ZN(n9243) );
  OAI221_X1 U10543 ( .B1(n9245), .B2(keyinput63), .C1(n9244), .C2(keyinput22), 
        .A(n9243), .ZN(n9252) );
  AOI22_X1 U10544 ( .A1(n5061), .A2(keyinput12), .B1(keyinput18), .B2(n9247), 
        .ZN(n9246) );
  OAI221_X1 U10545 ( .B1(n5061), .B2(keyinput12), .C1(n9247), .C2(keyinput18), 
        .A(n9246), .ZN(n9251) );
  INV_X1 U10546 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9249) );
  AOI22_X1 U10547 ( .A1(n9249), .A2(keyinput44), .B1(keyinput41), .B2(n9390), 
        .ZN(n9248) );
  OAI221_X1 U10548 ( .B1(n9249), .B2(keyinput44), .C1(n9390), .C2(keyinput41), 
        .A(n9248), .ZN(n9250) );
  NOR3_X1 U10549 ( .A1(n9252), .A2(n9251), .A3(n9250), .ZN(n9293) );
  AOI22_X1 U10550 ( .A1(n9254), .A2(keyinput28), .B1(n9349), .B2(keyinput37), 
        .ZN(n9253) );
  OAI221_X1 U10551 ( .B1(n9254), .B2(keyinput28), .C1(n9349), .C2(keyinput37), 
        .A(n9253), .ZN(n9271) );
  XOR2_X1 U10552 ( .A(n6003), .B(keyinput24), .Z(n9259) );
  XOR2_X1 U10553 ( .A(n9255), .B(keyinput20), .Z(n9258) );
  XNOR2_X1 U10554 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput57), .ZN(n9257) );
  XNOR2_X1 U10555 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput58), .ZN(n9256) );
  NAND4_X1 U10556 ( .A1(n9259), .A2(n9258), .A3(n9257), .A4(n9256), .ZN(n9270)
         );
  XNOR2_X1 U10557 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput2), .ZN(n9263) );
  XNOR2_X1 U10558 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput40), .ZN(n9262) );
  XNOR2_X1 U10559 ( .A(P1_REG3_REG_0__SCAN_IN), .B(keyinput59), .ZN(n9261) );
  XNOR2_X1 U10560 ( .A(SI_0_), .B(keyinput34), .ZN(n9260) );
  NAND4_X1 U10561 ( .A1(n9263), .A2(n9262), .A3(n9261), .A4(n9260), .ZN(n9269)
         );
  XNOR2_X1 U10562 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput10), .ZN(n9267) );
  XNOR2_X1 U10563 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput25), .ZN(n9266) );
  XNOR2_X1 U10564 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput50), .ZN(n9265) );
  XNOR2_X1 U10565 ( .A(SI_2_), .B(keyinput3), .ZN(n9264) );
  NAND4_X1 U10566 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(n9268)
         );
  NOR4_X1 U10567 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n9292)
         );
  AOI22_X1 U10568 ( .A1(n9274), .A2(keyinput21), .B1(keyinput27), .B2(n9273), 
        .ZN(n9272) );
  OAI221_X1 U10569 ( .B1(n9274), .B2(keyinput21), .C1(n9273), .C2(keyinput27), 
        .A(n9272), .ZN(n9283) );
  AOI22_X1 U10570 ( .A1(n9277), .A2(keyinput48), .B1(keyinput29), .B2(n9276), 
        .ZN(n9275) );
  OAI221_X1 U10571 ( .B1(n9277), .B2(keyinput48), .C1(n9276), .C2(keyinput29), 
        .A(n9275), .ZN(n9282) );
  INV_X1 U10572 ( .A(SI_12_), .ZN(n9279) );
  AOI22_X1 U10573 ( .A1(n9280), .A2(keyinput36), .B1(n9279), .B2(keyinput33), 
        .ZN(n9278) );
  OAI221_X1 U10574 ( .B1(n9280), .B2(keyinput36), .C1(n9279), .C2(keyinput33), 
        .A(n9278), .ZN(n9281) );
  OR3_X1 U10575 ( .A1(n9283), .A2(n9282), .A3(n9281), .ZN(n9290) );
  INV_X1 U10576 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9741) );
  AOI22_X1 U10577 ( .A1(n9285), .A2(keyinput53), .B1(keyinput32), .B2(n9741), 
        .ZN(n9284) );
  OAI221_X1 U10578 ( .B1(n9285), .B2(keyinput53), .C1(n9741), .C2(keyinput32), 
        .A(n9284), .ZN(n9289) );
  INV_X1 U10579 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U10580 ( .A1(n9677), .A2(keyinput4), .B1(keyinput38), .B2(n9287), 
        .ZN(n9286) );
  OAI221_X1 U10581 ( .B1(n9677), .B2(keyinput4), .C1(n9287), .C2(keyinput38), 
        .A(n9286), .ZN(n9288) );
  NOR3_X1 U10582 ( .A1(n9290), .A2(n9289), .A3(n9288), .ZN(n9291) );
  AND4_X1 U10583 ( .A1(n9294), .A2(n9293), .A3(n9292), .A4(n9291), .ZN(n9335)
         );
  INV_X1 U10584 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9676) );
  AOI22_X1 U10585 ( .A1(n5993), .A2(keyinput23), .B1(n9676), .B2(keyinput52), 
        .ZN(n9295) );
  OAI221_X1 U10586 ( .B1(n5993), .B2(keyinput23), .C1(n9676), .C2(keyinput52), 
        .A(n9295), .ZN(n9307) );
  AOI22_X1 U10587 ( .A1(n9298), .A2(keyinput15), .B1(n9297), .B2(keyinput31), 
        .ZN(n9296) );
  OAI221_X1 U10588 ( .B1(n9298), .B2(keyinput15), .C1(n9297), .C2(keyinput31), 
        .A(n9296), .ZN(n9306) );
  AOI22_X1 U10589 ( .A1(n9301), .A2(keyinput55), .B1(n9300), .B2(keyinput26), 
        .ZN(n9299) );
  OAI221_X1 U10590 ( .B1(n9301), .B2(keyinput55), .C1(n9300), .C2(keyinput26), 
        .A(n9299), .ZN(n9305) );
  INV_X1 U10591 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9303) );
  AOI22_X1 U10592 ( .A1(n8521), .A2(keyinput13), .B1(n9303), .B2(keyinput14), 
        .ZN(n9302) );
  OAI221_X1 U10593 ( .B1(n8521), .B2(keyinput13), .C1(n9303), .C2(keyinput14), 
        .A(n9302), .ZN(n9304) );
  NOR4_X1 U10594 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), .ZN(n9334)
         );
  INV_X1 U10595 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U10596 ( .A1(n9309), .A2(keyinput43), .B1(n9674), .B2(keyinput7), 
        .ZN(n9308) );
  OAI221_X1 U10597 ( .B1(n9309), .B2(keyinput43), .C1(n9674), .C2(keyinput7), 
        .A(n9308), .ZN(n9318) );
  INV_X1 U10598 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9311) );
  AOI22_X1 U10599 ( .A1(n8510), .A2(keyinput54), .B1(n9311), .B2(keyinput56), 
        .ZN(n9310) );
  OAI221_X1 U10600 ( .B1(n8510), .B2(keyinput54), .C1(n9311), .C2(keyinput56), 
        .A(n9310), .ZN(n9317) );
  INV_X1 U10601 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9693) );
  AOI22_X1 U10602 ( .A1(n9693), .A2(keyinput0), .B1(keyinput9), .B2(n9313), 
        .ZN(n9312) );
  OAI221_X1 U10603 ( .B1(n9693), .B2(keyinput0), .C1(n9313), .C2(keyinput9), 
        .A(n9312), .ZN(n9316) );
  INV_X1 U10604 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9675) );
  AOI22_X1 U10605 ( .A1(P2_U3151), .A2(keyinput1), .B1(n9675), .B2(keyinput42), 
        .ZN(n9314) );
  OAI221_X1 U10606 ( .B1(P2_U3151), .B2(keyinput1), .C1(n9675), .C2(keyinput42), .A(n9314), .ZN(n9315) );
  NOR4_X1 U10607 ( .A1(n9318), .A2(n9317), .A3(n9316), .A4(n9315), .ZN(n9333)
         );
  INV_X1 U10608 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9320) );
  AOI22_X1 U10609 ( .A1(n9350), .A2(keyinput6), .B1(keyinput35), .B2(n9320), 
        .ZN(n9319) );
  OAI221_X1 U10610 ( .B1(n9350), .B2(keyinput6), .C1(n9320), .C2(keyinput35), 
        .A(n9319), .ZN(n9331) );
  INV_X1 U10611 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9747) );
  INV_X1 U10612 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9322) );
  AOI22_X1 U10613 ( .A1(n9747), .A2(keyinput45), .B1(n9322), .B2(keyinput8), 
        .ZN(n9321) );
  OAI221_X1 U10614 ( .B1(n9747), .B2(keyinput45), .C1(n9322), .C2(keyinput8), 
        .A(n9321), .ZN(n9330) );
  INV_X1 U10615 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9324) );
  AOI22_X1 U10616 ( .A1(n9325), .A2(keyinput51), .B1(keyinput5), .B2(n9324), 
        .ZN(n9323) );
  OAI221_X1 U10617 ( .B1(n9325), .B2(keyinput51), .C1(n9324), .C2(keyinput5), 
        .A(n9323), .ZN(n9329) );
  INV_X1 U10618 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9733) );
  AOI22_X1 U10619 ( .A1(n9733), .A2(keyinput61), .B1(keyinput46), .B2(n9327), 
        .ZN(n9326) );
  OAI221_X1 U10620 ( .B1(n9733), .B2(keyinput61), .C1(n9327), .C2(keyinput46), 
        .A(n9326), .ZN(n9328) );
  NOR4_X1 U10621 ( .A1(n9331), .A2(n9330), .A3(n9329), .A4(n9328), .ZN(n9332)
         );
  NAND4_X1 U10622 ( .A1(n9335), .A2(n9334), .A3(n9333), .A4(n9332), .ZN(n9363)
         );
  NAND4_X1 U10623 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .A3(P2_REG3_REG_14__SCAN_IN), .A4(P2_REG2_REG_25__SCAN_IN), .ZN(n9346)
         );
  NAND4_X1 U10624 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(P2_REG0_REG_26__SCAN_IN), 
        .A3(P2_ADDR_REG_10__SCAN_IN), .A4(P2_ADDR_REG_17__SCAN_IN), .ZN(n9345)
         );
  NOR3_X1 U10625 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(P2_REG0_REG_19__SCAN_IN), 
        .A3(n9336), .ZN(n9338) );
  NOR3_X1 U10626 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .A3(P2_REG3_REG_11__SCAN_IN), .ZN(n9337) );
  NAND4_X1 U10627 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), 
        .A3(n9338), .A4(n9337), .ZN(n9344) );
  NOR4_X1 U10628 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG0_REG_23__SCAN_IN), .A4(P2_REG2_REG_0__SCAN_IN), .ZN(n9342)
         );
  NOR4_X1 U10629 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(P2_REG1_REG_8__SCAN_IN), 
        .A3(P2_REG1_REG_1__SCAN_IN), .A4(P2_REG3_REG_1__SCAN_IN), .ZN(n9341)
         );
  NOR4_X1 U10630 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG1_REG_20__SCAN_IN), 
        .A3(P1_REG0_REG_10__SCAN_IN), .A4(P1_REG0_REG_2__SCAN_IN), .ZN(n9340)
         );
  NOR4_X1 U10631 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(P1_REG1_REG_9__SCAN_IN), 
        .A3(P1_REG2_REG_2__SCAN_IN), .A4(P1_REG2_REG_1__SCAN_IN), .ZN(n9339)
         );
  NAND4_X1 U10632 ( .A1(n9342), .A2(n9341), .A3(n9340), .A4(n9339), .ZN(n9343)
         );
  NOR4_X1 U10633 ( .A1(n9346), .A2(n9345), .A3(n9344), .A4(n9343), .ZN(n9361)
         );
  NAND4_X1 U10634 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P2_DATAO_REG_26__SCAN_IN), 
        .A3(P1_D_REG_11__SCAN_IN), .A4(n9674), .ZN(n9347) );
  NOR4_X1 U10635 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .A3(n9348), .A4(n9347), .ZN(n9360) );
  NOR4_X1 U10636 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .A3(P1_D_REG_0__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9359) );
  NOR3_X1 U10637 ( .A1(SI_15_), .A2(P1_DATAO_REG_13__SCAN_IN), .A3(SI_2_), 
        .ZN(n9352) );
  NOR4_X1 U10638 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(P2_DATAO_REG_16__SCAN_IN), .A3(n9350), .A4(n9349), .ZN(n9351) );
  AND3_X1 U10639 ( .A1(SI_0_), .A2(n9352), .A3(n9351), .ZN(n9353) );
  NAND3_X1 U10640 ( .A1(n9353), .A2(SI_12_), .A3(P2_REG2_REG_26__SCAN_IN), 
        .ZN(n9357) );
  NAND4_X1 U10641 ( .A1(n9390), .A2(P2_REG2_REG_2__SCAN_IN), .A3(
        P1_REG0_REG_25__SCAN_IN), .A4(P1_REG3_REG_17__SCAN_IN), .ZN(n9356) );
  NAND4_X1 U10642 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(P1_REG0_REG_18__SCAN_IN), 
        .A3(P1_REG0_REG_8__SCAN_IN), .A4(P2_DATAO_REG_1__SCAN_IN), .ZN(n9355)
         );
  NAND2_X1 U10643 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(P1_REG0_REG_9__SCAN_IN), 
        .ZN(n9354) );
  NOR4_X1 U10644 ( .A1(n9357), .A2(n9356), .A3(n9355), .A4(n9354), .ZN(n9358)
         );
  NAND4_X1 U10645 ( .A1(n9361), .A2(n9360), .A3(n9359), .A4(n9358), .ZN(n9362)
         );
  XNOR2_X1 U10646 ( .A(n9363), .B(n9362), .ZN(n9364) );
  XNOR2_X1 U10647 ( .A(n9365), .B(n9364), .ZN(P1_U3520) );
  MUX2_X1 U10648 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9366), .S(n9777), .Z(
        P1_U3518) );
  MUX2_X1 U10649 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9367), .S(n9777), .Z(
        P1_U3517) );
  MUX2_X1 U10650 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9368), .S(n9777), .Z(
        P1_U3516) );
  MUX2_X1 U10651 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9369), .S(n9777), .Z(
        P1_U3515) );
  MUX2_X1 U10652 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9370), .S(n9777), .Z(
        P1_U3514) );
  MUX2_X1 U10653 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9371), .S(n9777), .Z(
        P1_U3513) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9372), .S(n9777), .Z(
        P1_U3512) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9373), .S(n9777), .Z(
        P1_U3511) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9374), .S(n9777), .Z(
        P1_U3510) );
  MUX2_X1 U10657 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9375), .S(n9777), .Z(
        P1_U3509) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9376), .S(n9777), .Z(
        P1_U3507) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9377), .S(n9777), .Z(
        P1_U3504) );
  MUX2_X1 U10660 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9378), .S(n9777), .Z(
        P1_U3501) );
  MUX2_X1 U10661 ( .A(P1_D_REG_1__SCAN_IN), .B(n9381), .S(n9678), .Z(P1_U3440)
         );
  MUX2_X1 U10662 ( .A(P1_D_REG_0__SCAN_IN), .B(n9382), .S(n9678), .Z(P1_U3439)
         );
  INV_X1 U10663 ( .A(n9383), .ZN(n9388) );
  NOR4_X1 U10664 ( .A1(n4896), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9384), .ZN(n9385) );
  AOI21_X1 U10665 ( .B1(n9386), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9385), .ZN(
        n9387) );
  OAI21_X1 U10666 ( .B1(n9388), .B2(n9395), .A(n9387), .ZN(P1_U3324) );
  OAI222_X1 U10667 ( .A1(P1_U3086), .A2(n9389), .B1(n9395), .B2(n9391), .C1(
        n9390), .C2(n9392), .ZN(P1_U3325) );
  OAI222_X1 U10668 ( .A1(P1_U3086), .A2(n9396), .B1(n9395), .B2(n9394), .C1(
        n9393), .C2(n9392), .ZN(P1_U3326) );
  INV_X1 U10669 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9409) );
  AOI211_X1 U10670 ( .C1(n9400), .C2(n9399), .A(n9398), .B(n9602), .ZN(n9405)
         );
  AOI211_X1 U10671 ( .C1(n9403), .C2(n9402), .A(n9401), .B(n9575), .ZN(n9404)
         );
  AOI211_X1 U10672 ( .C1(n9605), .C2(n9406), .A(n9405), .B(n9404), .ZN(n9408)
         );
  OAI211_X1 U10673 ( .C1(n9613), .C2(n9409), .A(n9408), .B(n9407), .ZN(
        P1_U3253) );
  INV_X1 U10674 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9424) );
  AOI21_X1 U10675 ( .B1(n9412), .B2(n9411), .A(n9410), .ZN(n9413) );
  NAND2_X1 U10676 ( .A1(n9598), .A2(n9413), .ZN(n9419) );
  AOI21_X1 U10677 ( .B1(n9416), .B2(n9415), .A(n9414), .ZN(n9417) );
  NAND2_X1 U10678 ( .A1(n9591), .A2(n9417), .ZN(n9418) );
  OAI211_X1 U10679 ( .C1(n9543), .C2(n9420), .A(n9419), .B(n9418), .ZN(n9421)
         );
  INV_X1 U10680 ( .A(n9421), .ZN(n9423) );
  OAI211_X1 U10681 ( .C1(n9613), .C2(n9424), .A(n9423), .B(n9422), .ZN(
        P1_U3250) );
  INV_X1 U10682 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9439) );
  AOI21_X1 U10683 ( .B1(n9427), .B2(n9426), .A(n9425), .ZN(n9428) );
  NAND2_X1 U10684 ( .A1(n9598), .A2(n9428), .ZN(n9434) );
  AOI21_X1 U10685 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n9432) );
  NAND2_X1 U10686 ( .A1(n9591), .A2(n9432), .ZN(n9433) );
  OAI211_X1 U10687 ( .C1(n9543), .C2(n9435), .A(n9434), .B(n9433), .ZN(n9436)
         );
  INV_X1 U10688 ( .A(n9436), .ZN(n9438) );
  OAI211_X1 U10689 ( .C1(n9439), .C2(n9613), .A(n9438), .B(n9437), .ZN(
        P1_U3246) );
  INV_X1 U10690 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9454) );
  AOI21_X1 U10691 ( .B1(n9442), .B2(n9441), .A(n9440), .ZN(n9443) );
  NAND2_X1 U10692 ( .A1(n9598), .A2(n9443), .ZN(n9449) );
  AOI21_X1 U10693 ( .B1(n9446), .B2(n9445), .A(n9444), .ZN(n9447) );
  NAND2_X1 U10694 ( .A1(n9591), .A2(n9447), .ZN(n9448) );
  OAI211_X1 U10695 ( .C1(n9543), .C2(n9450), .A(n9449), .B(n9448), .ZN(n9451)
         );
  INV_X1 U10696 ( .A(n9451), .ZN(n9453) );
  OAI211_X1 U10697 ( .C1(n9613), .C2(n9454), .A(n9453), .B(n9452), .ZN(
        P1_U3251) );
  NOR2_X1 U10698 ( .A1(n9455), .A2(n9913), .ZN(n9457) );
  AOI211_X1 U10699 ( .C1(n9921), .C2(n9458), .A(n9457), .B(n9456), .ZN(n9460)
         );
  AOI22_X1 U10700 ( .A1(n9952), .A2(n9460), .B1(n9459), .B2(n9950), .ZN(
        P2_U3472) );
  INV_X1 U10701 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9461) );
  AOI22_X1 U10702 ( .A1(n9934), .A2(n9461), .B1(n9460), .B2(n9932), .ZN(
        P2_U3429) );
  XNOR2_X1 U10703 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10704 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U10705 ( .A1(n9486), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9484) );
  INV_X1 U10706 ( .A(n9462), .ZN(n9463) );
  OAI211_X1 U10707 ( .C1(n9465), .C2(n9464), .A(n9598), .B(n9463), .ZN(n9470)
         );
  OAI211_X1 U10708 ( .C1(n9468), .C2(n9467), .A(n9591), .B(n9466), .ZN(n9469)
         );
  OAI211_X1 U10709 ( .C1(n9543), .C2(n9471), .A(n9470), .B(n9469), .ZN(n9472)
         );
  INV_X1 U10710 ( .A(n9472), .ZN(n9483) );
  NAND3_X1 U10711 ( .A1(n9475), .A2(n9474), .A3(n9473), .ZN(n9482) );
  INV_X1 U10712 ( .A(n9476), .ZN(n9478) );
  AOI22_X1 U10713 ( .A1(n9480), .A2(n9479), .B1(n9478), .B2(n9477), .ZN(n9481)
         );
  NAND3_X1 U10714 ( .A1(n9482), .A2(P1_U3973), .A3(n9481), .ZN(n9498) );
  NAND3_X1 U10715 ( .A1(n9484), .A2(n9483), .A3(n9498), .ZN(P1_U3245) );
  AOI21_X1 U10716 ( .B1(n9486), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9485), .ZN(
        n9500) );
  AOI21_X1 U10717 ( .B1(n9488), .B2(n4294), .A(n9487), .ZN(n9489) );
  NAND2_X1 U10718 ( .A1(n9598), .A2(n9489), .ZN(n9495) );
  AOI21_X1 U10719 ( .B1(n9492), .B2(n9491), .A(n9490), .ZN(n9493) );
  NAND2_X1 U10720 ( .A1(n9591), .A2(n9493), .ZN(n9494) );
  OAI211_X1 U10721 ( .C1(n9543), .C2(n9496), .A(n9495), .B(n9494), .ZN(n9497)
         );
  INV_X1 U10722 ( .A(n9497), .ZN(n9499) );
  NAND3_X1 U10723 ( .A1(n9500), .A2(n9499), .A3(n9498), .ZN(P1_U3247) );
  INV_X1 U10724 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9515) );
  AOI21_X1 U10725 ( .B1(n9503), .B2(n9502), .A(n9501), .ZN(n9504) );
  NAND2_X1 U10726 ( .A1(n9598), .A2(n9504), .ZN(n9510) );
  AOI21_X1 U10727 ( .B1(n9507), .B2(n9506), .A(n9505), .ZN(n9508) );
  NAND2_X1 U10728 ( .A1(n9591), .A2(n9508), .ZN(n9509) );
  OAI211_X1 U10729 ( .C1(n9543), .C2(n9511), .A(n9510), .B(n9509), .ZN(n9512)
         );
  INV_X1 U10730 ( .A(n9512), .ZN(n9514) );
  OAI211_X1 U10731 ( .C1(n9613), .C2(n9515), .A(n9514), .B(n9513), .ZN(
        P1_U3248) );
  INV_X1 U10732 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9530) );
  AOI21_X1 U10733 ( .B1(n9518), .B2(n9517), .A(n9516), .ZN(n9519) );
  NAND2_X1 U10734 ( .A1(n9598), .A2(n9519), .ZN(n9525) );
  AOI21_X1 U10735 ( .B1(n9522), .B2(n9521), .A(n9520), .ZN(n9523) );
  NAND2_X1 U10736 ( .A1(n9591), .A2(n9523), .ZN(n9524) );
  OAI211_X1 U10737 ( .C1(n9543), .C2(n9526), .A(n9525), .B(n9524), .ZN(n9527)
         );
  INV_X1 U10738 ( .A(n9527), .ZN(n9529) );
  OAI211_X1 U10739 ( .C1(n9613), .C2(n9530), .A(n9529), .B(n9528), .ZN(
        P1_U3249) );
  INV_X1 U10740 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9547) );
  INV_X1 U10741 ( .A(n9531), .ZN(n9542) );
  AOI21_X1 U10742 ( .B1(n9534), .B2(n9533), .A(n9532), .ZN(n9535) );
  NAND2_X1 U10743 ( .A1(n9598), .A2(n9535), .ZN(n9541) );
  AOI21_X1 U10744 ( .B1(n9538), .B2(n9537), .A(n9536), .ZN(n9539) );
  NAND2_X1 U10745 ( .A1(n9591), .A2(n9539), .ZN(n9540) );
  OAI211_X1 U10746 ( .C1(n9543), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9544)
         );
  INV_X1 U10747 ( .A(n9544), .ZN(n9546) );
  OAI211_X1 U10748 ( .C1(n9613), .C2(n9547), .A(n9546), .B(n9545), .ZN(
        P1_U3254) );
  INV_X1 U10749 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9559) );
  AOI211_X1 U10750 ( .C1(n9550), .C2(n9549), .A(n9602), .B(n9548), .ZN(n9555)
         );
  AOI211_X1 U10751 ( .C1(n9553), .C2(n9552), .A(n9575), .B(n9551), .ZN(n9554)
         );
  AOI211_X1 U10752 ( .C1(n9605), .C2(n9556), .A(n9555), .B(n9554), .ZN(n9558)
         );
  OAI211_X1 U10753 ( .C1(n9613), .C2(n9559), .A(n9558), .B(n9557), .ZN(
        P1_U3256) );
  INV_X1 U10754 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9571) );
  AOI211_X1 U10755 ( .C1(n9562), .C2(n9561), .A(n9602), .B(n9560), .ZN(n9567)
         );
  AOI211_X1 U10756 ( .C1(n9565), .C2(n9564), .A(n9563), .B(n9575), .ZN(n9566)
         );
  AOI211_X1 U10757 ( .C1(n9605), .C2(n9568), .A(n9567), .B(n9566), .ZN(n9570)
         );
  OAI211_X1 U10758 ( .C1(n9613), .C2(n9571), .A(n9570), .B(n9569), .ZN(
        P1_U3257) );
  INV_X1 U10759 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9584) );
  AOI211_X1 U10760 ( .C1(n9574), .C2(n9573), .A(n9572), .B(n9602), .ZN(n9580)
         );
  AOI211_X1 U10761 ( .C1(n9578), .C2(n9577), .A(n9576), .B(n9575), .ZN(n9579)
         );
  AOI211_X1 U10762 ( .C1(n9605), .C2(n9581), .A(n9580), .B(n9579), .ZN(n9583)
         );
  OAI211_X1 U10763 ( .C1(n9613), .C2(n9584), .A(n9583), .B(n9582), .ZN(
        P1_U3258) );
  OAI21_X1 U10764 ( .B1(n9587), .B2(n9586), .A(n9585), .ZN(n9594) );
  OAI21_X1 U10765 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9592) );
  AOI222_X1 U10766 ( .A1(n9594), .A2(n9598), .B1(n9593), .B2(n9605), .C1(n9592), .C2(n9591), .ZN(n9596) );
  OAI211_X1 U10767 ( .C1(n9613), .C2(n9597), .A(n9596), .B(n9595), .ZN(
        P1_U3260) );
  OAI211_X1 U10768 ( .C1(n9601), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9610)
         );
  AOI21_X1 U10769 ( .B1(n9604), .B2(n9603), .A(n9602), .ZN(n9608) );
  AOI22_X1 U10770 ( .A1(n9608), .A2(n9607), .B1(n9606), .B2(n9605), .ZN(n9609)
         );
  AND2_X1 U10771 ( .A1(n9610), .A2(n9609), .ZN(n9612) );
  OAI211_X1 U10772 ( .C1(n9613), .C2(n9959), .A(n9612), .B(n9611), .ZN(
        P1_U3261) );
  OAI21_X1 U10773 ( .B1(n9621), .B2(n9615), .A(n9614), .ZN(n9625) );
  OAI22_X1 U10774 ( .A1(n9619), .A2(n9618), .B1(n9617), .B2(n9616), .ZN(n9624)
         );
  XNOR2_X1 U10775 ( .A(n9620), .B(n9621), .ZN(n9629) );
  NOR2_X1 U10776 ( .A1(n9629), .A2(n9622), .ZN(n9623) );
  AOI211_X1 U10777 ( .C1(n9655), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9729)
         );
  AOI22_X1 U10778 ( .A1(n9658), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9626), .B2(
        n9656), .ZN(n9627) );
  OAI21_X1 U10779 ( .B1(n9660), .B2(n9728), .A(n9627), .ZN(n9628) );
  INV_X1 U10780 ( .A(n9628), .ZN(n9636) );
  INV_X1 U10781 ( .A(n9629), .ZN(n9732) );
  INV_X1 U10782 ( .A(n9630), .ZN(n9632) );
  OAI211_X1 U10783 ( .C1(n9632), .C2(n9728), .A(n9666), .B(n9631), .ZN(n9727)
         );
  INV_X1 U10784 ( .A(n9727), .ZN(n9633) );
  AOI22_X1 U10785 ( .A1(n9732), .A2(n9634), .B1(n9669), .B2(n9633), .ZN(n9635)
         );
  OAI211_X1 U10786 ( .C1(n9673), .C2(n9729), .A(n9636), .B(n9635), .ZN(
        P1_U3285) );
  XNOR2_X1 U10787 ( .A(n7639), .B(n9643), .ZN(n9638) );
  AOI222_X1 U10788 ( .A1(n9655), .A2(n9638), .B1(n9637), .B2(n9652), .C1(n9653), .C2(n9651), .ZN(n9715) );
  AOI22_X1 U10789 ( .A1(n9658), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9639), .B2(
        n9656), .ZN(n9640) );
  OAI21_X1 U10790 ( .B1(n9660), .B2(n9714), .A(n9640), .ZN(n9641) );
  INV_X1 U10791 ( .A(n9641), .ZN(n9649) );
  XNOR2_X1 U10792 ( .A(n9642), .B(n9643), .ZN(n9718) );
  INV_X1 U10793 ( .A(n9644), .ZN(n9645) );
  OAI211_X1 U10794 ( .C1(n9714), .C2(n9646), .A(n9645), .B(n9666), .ZN(n9713)
         );
  INV_X1 U10795 ( .A(n9713), .ZN(n9647) );
  AOI22_X1 U10796 ( .A1(n9718), .A2(n9670), .B1(n9669), .B2(n9647), .ZN(n9648)
         );
  OAI211_X1 U10797 ( .C1(n9658), .C2(n9715), .A(n9649), .B(n9648), .ZN(
        P1_U3287) );
  XNOR2_X1 U10798 ( .A(n9650), .B(n9663), .ZN(n9654) );
  AOI222_X1 U10799 ( .A1(n9655), .A2(n9654), .B1(n9653), .B2(n9652), .C1(n5754), .C2(n9651), .ZN(n9702) );
  AOI22_X1 U10800 ( .A1(n9658), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9657), .B2(
        n9656), .ZN(n9659) );
  OAI21_X1 U10801 ( .B1(n9660), .B2(n9701), .A(n9659), .ZN(n9661) );
  INV_X1 U10802 ( .A(n9661), .ZN(n9672) );
  XNOR2_X1 U10803 ( .A(n9663), .B(n9662), .ZN(n9705) );
  INV_X1 U10804 ( .A(n9664), .ZN(n9667) );
  OAI211_X1 U10805 ( .C1(n9667), .C2(n9701), .A(n9666), .B(n9665), .ZN(n9700)
         );
  INV_X1 U10806 ( .A(n9700), .ZN(n9668) );
  AOI22_X1 U10807 ( .A1(n9705), .A2(n9670), .B1(n9669), .B2(n9668), .ZN(n9671)
         );
  OAI211_X1 U10808 ( .C1(n9673), .C2(n9702), .A(n9672), .B(n9671), .ZN(
        P1_U3289) );
  AND2_X1 U10809 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9679), .ZN(P1_U3294) );
  AND2_X1 U10810 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9679), .ZN(P1_U3295) );
  AND2_X1 U10811 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9679), .ZN(P1_U3296) );
  AND2_X1 U10812 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9679), .ZN(P1_U3297) );
  AND2_X1 U10813 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9679), .ZN(P1_U3298) );
  AND2_X1 U10814 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9679), .ZN(P1_U3299) );
  AND2_X1 U10815 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9679), .ZN(P1_U3300) );
  AND2_X1 U10816 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9679), .ZN(P1_U3301) );
  AND2_X1 U10817 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9679), .ZN(P1_U3302) );
  AND2_X1 U10818 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9679), .ZN(P1_U3303) );
  AND2_X1 U10819 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9679), .ZN(P1_U3304) );
  AND2_X1 U10820 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9679), .ZN(P1_U3305) );
  NOR2_X1 U10821 ( .A1(n9678), .A2(n9674), .ZN(P1_U3306) );
  AND2_X1 U10822 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9679), .ZN(P1_U3307) );
  AND2_X1 U10823 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9679), .ZN(P1_U3308) );
  AND2_X1 U10824 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9679), .ZN(P1_U3309) );
  AND2_X1 U10825 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9679), .ZN(P1_U3310) );
  AND2_X1 U10826 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9679), .ZN(P1_U3311) );
  AND2_X1 U10827 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9679), .ZN(P1_U3312) );
  AND2_X1 U10828 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9679), .ZN(P1_U3313) );
  NOR2_X1 U10829 ( .A1(n9678), .A2(n9675), .ZN(P1_U3314) );
  AND2_X1 U10830 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9679), .ZN(P1_U3315) );
  AND2_X1 U10831 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9679), .ZN(P1_U3316) );
  AND2_X1 U10832 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9679), .ZN(P1_U3317) );
  AND2_X1 U10833 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9679), .ZN(P1_U3318) );
  NOR2_X1 U10834 ( .A1(n9678), .A2(n9676), .ZN(P1_U3319) );
  AND2_X1 U10835 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9679), .ZN(P1_U3320) );
  AND2_X1 U10836 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9679), .ZN(P1_U3321) );
  NOR2_X1 U10837 ( .A1(n9678), .A2(n9677), .ZN(P1_U3322) );
  AND2_X1 U10838 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9679), .ZN(P1_U3323) );
  INV_X1 U10839 ( .A(n9680), .ZN(n9751) );
  INV_X1 U10840 ( .A(n9681), .ZN(n9682) );
  OAI21_X1 U10841 ( .B1(n9683), .B2(n9767), .A(n9682), .ZN(n9685) );
  AOI211_X1 U10842 ( .C1(n9751), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9779)
         );
  INV_X1 U10843 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9687) );
  AOI22_X1 U10844 ( .A1(n9777), .A2(n9779), .B1(n9687), .B2(n9775), .ZN(
        P1_U3456) );
  OAI21_X1 U10845 ( .B1(n9689), .B2(n9767), .A(n9688), .ZN(n9691) );
  AOI211_X1 U10846 ( .C1(n9692), .C2(n9773), .A(n9691), .B(n9690), .ZN(n9781)
         );
  AOI22_X1 U10847 ( .A1(n9777), .A2(n9781), .B1(n9693), .B2(n9775), .ZN(
        P1_U3459) );
  OAI21_X1 U10848 ( .B1(n9695), .B2(n9767), .A(n9694), .ZN(n9697) );
  AOI211_X1 U10849 ( .C1(n9773), .C2(n9698), .A(n9697), .B(n9696), .ZN(n9783)
         );
  INV_X1 U10850 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U10851 ( .A1(n9777), .A2(n9783), .B1(n9699), .B2(n9775), .ZN(
        P1_U3462) );
  OAI21_X1 U10852 ( .B1(n9701), .B2(n9767), .A(n9700), .ZN(n9704) );
  INV_X1 U10853 ( .A(n9702), .ZN(n9703) );
  AOI211_X1 U10854 ( .C1(n9773), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9785)
         );
  INV_X1 U10855 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9706) );
  AOI22_X1 U10856 ( .A1(n9777), .A2(n9785), .B1(n9706), .B2(n9775), .ZN(
        P1_U3465) );
  OAI21_X1 U10857 ( .B1(n9708), .B2(n9767), .A(n9707), .ZN(n9710) );
  AOI211_X1 U10858 ( .C1(n9773), .C2(n9711), .A(n9710), .B(n9709), .ZN(n9787)
         );
  INV_X1 U10859 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9712) );
  AOI22_X1 U10860 ( .A1(n9777), .A2(n9787), .B1(n9712), .B2(n9775), .ZN(
        P1_U3468) );
  OAI21_X1 U10861 ( .B1(n9714), .B2(n9767), .A(n9713), .ZN(n9717) );
  INV_X1 U10862 ( .A(n9715), .ZN(n9716) );
  AOI211_X1 U10863 ( .C1(n9773), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9789)
         );
  INV_X1 U10864 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9719) );
  AOI22_X1 U10865 ( .A1(n9777), .A2(n9789), .B1(n9719), .B2(n9775), .ZN(
        P1_U3471) );
  NAND2_X1 U10866 ( .A1(n9720), .A2(n9751), .ZN(n9722) );
  OAI211_X1 U10867 ( .C1(n9723), .C2(n9767), .A(n9722), .B(n9721), .ZN(n9724)
         );
  NOR2_X1 U10868 ( .A1(n9725), .A2(n9724), .ZN(n9790) );
  INV_X1 U10869 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9726) );
  AOI22_X1 U10870 ( .A1(n9777), .A2(n9790), .B1(n9726), .B2(n9775), .ZN(
        P1_U3474) );
  OAI21_X1 U10871 ( .B1(n9728), .B2(n9767), .A(n9727), .ZN(n9731) );
  INV_X1 U10872 ( .A(n9729), .ZN(n9730) );
  AOI211_X1 U10873 ( .C1(n9751), .C2(n9732), .A(n9731), .B(n9730), .ZN(n9791)
         );
  AOI22_X1 U10874 ( .A1(n9777), .A2(n9791), .B1(n9733), .B2(n9775), .ZN(
        P1_U3477) );
  NAND2_X1 U10875 ( .A1(n5078), .A2(n9734), .ZN(n9735) );
  NAND2_X1 U10876 ( .A1(n9736), .A2(n9735), .ZN(n9737) );
  AOI21_X1 U10877 ( .B1(n9738), .B2(n9773), .A(n9737), .ZN(n9739) );
  AND2_X1 U10878 ( .A1(n9740), .A2(n9739), .ZN(n9793) );
  AOI22_X1 U10879 ( .A1(n9777), .A2(n9793), .B1(n9741), .B2(n9775), .ZN(
        P1_U3480) );
  OAI21_X1 U10880 ( .B1(n9743), .B2(n9767), .A(n9742), .ZN(n9744) );
  AOI211_X1 U10881 ( .C1(n9746), .C2(n9773), .A(n9745), .B(n9744), .ZN(n9794)
         );
  AOI22_X1 U10882 ( .A1(n9777), .A2(n9794), .B1(n9747), .B2(n9775), .ZN(
        P1_U3483) );
  OAI21_X1 U10883 ( .B1(n9749), .B2(n9767), .A(n9748), .ZN(n9750) );
  AOI21_X1 U10884 ( .B1(n9752), .B2(n9751), .A(n9750), .ZN(n9753) );
  AND2_X1 U10885 ( .A1(n9754), .A2(n9753), .ZN(n9795) );
  INV_X1 U10886 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9755) );
  AOI22_X1 U10887 ( .A1(n9777), .A2(n9795), .B1(n9755), .B2(n9775), .ZN(
        P1_U3486) );
  OAI21_X1 U10888 ( .B1(n9757), .B2(n9767), .A(n9756), .ZN(n9758) );
  AOI211_X1 U10889 ( .C1(n9760), .C2(n9773), .A(n9759), .B(n9758), .ZN(n9797)
         );
  INV_X1 U10890 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9761) );
  AOI22_X1 U10891 ( .A1(n9777), .A2(n9797), .B1(n9761), .B2(n9775), .ZN(
        P1_U3489) );
  OAI211_X1 U10892 ( .C1(n5500), .C2(n9767), .A(n9763), .B(n9762), .ZN(n9764)
         );
  AOI21_X1 U10893 ( .B1(n9765), .B2(n9773), .A(n9764), .ZN(n9799) );
  INV_X1 U10894 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9766) );
  AOI22_X1 U10895 ( .A1(n9777), .A2(n9799), .B1(n9766), .B2(n9775), .ZN(
        P1_U3492) );
  OAI22_X1 U10896 ( .A1(n9770), .A2(n9769), .B1(n9768), .B2(n9767), .ZN(n9771)
         );
  AOI211_X1 U10897 ( .C1(n9774), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9802)
         );
  INV_X1 U10898 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9776) );
  AOI22_X1 U10899 ( .A1(n9777), .A2(n9802), .B1(n9776), .B2(n9775), .ZN(
        P1_U3495) );
  AOI22_X1 U10900 ( .A1(n9803), .A2(n9779), .B1(n9778), .B2(n9800), .ZN(
        P1_U3523) );
  INV_X1 U10901 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U10902 ( .A1(n9803), .A2(n9781), .B1(n9780), .B2(n9800), .ZN(
        P1_U3524) );
  INV_X1 U10903 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9782) );
  AOI22_X1 U10904 ( .A1(n9803), .A2(n9783), .B1(n9782), .B2(n9800), .ZN(
        P1_U3525) );
  INV_X1 U10905 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U10906 ( .A1(n9803), .A2(n9785), .B1(n9784), .B2(n9800), .ZN(
        P1_U3526) );
  INV_X1 U10907 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9786) );
  AOI22_X1 U10908 ( .A1(n9803), .A2(n9787), .B1(n9786), .B2(n9800), .ZN(
        P1_U3527) );
  INV_X1 U10909 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9788) );
  AOI22_X1 U10910 ( .A1(n9803), .A2(n9789), .B1(n9788), .B2(n9800), .ZN(
        P1_U3528) );
  AOI22_X1 U10911 ( .A1(n9803), .A2(n9790), .B1(n6634), .B2(n9800), .ZN(
        P1_U3529) );
  AOI22_X1 U10912 ( .A1(n9803), .A2(n9791), .B1(n6636), .B2(n9800), .ZN(
        P1_U3530) );
  AOI22_X1 U10913 ( .A1(n9803), .A2(n9793), .B1(n9792), .B2(n9800), .ZN(
        P1_U3531) );
  AOI22_X1 U10914 ( .A1(n9803), .A2(n9794), .B1(n6844), .B2(n9800), .ZN(
        P1_U3532) );
  AOI22_X1 U10915 ( .A1(n9803), .A2(n9795), .B1(n6847), .B2(n9800), .ZN(
        P1_U3533) );
  AOI22_X1 U10916 ( .A1(n9803), .A2(n9797), .B1(n9796), .B2(n9800), .ZN(
        P1_U3534) );
  AOI22_X1 U10917 ( .A1(n9803), .A2(n9799), .B1(n9798), .B2(n9800), .ZN(
        P1_U3535) );
  AOI22_X1 U10918 ( .A1(n9803), .A2(n9802), .B1(n9801), .B2(n9800), .ZN(
        P1_U3536) );
  AOI22_X1 U10919 ( .A1(n9839), .A2(P2_IR_REG_0__SCAN_IN), .B1(n9841), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n9808) );
  OAI21_X1 U10920 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9804), .A(n9826), .ZN(
        n9805) );
  OAI21_X1 U10921 ( .B1(n9806), .B2(n9827), .A(n9805), .ZN(n9807) );
  OAI211_X1 U10922 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6002), .A(n9808), .B(
        n9807), .ZN(P2_U3182) );
  NAND2_X1 U10923 ( .A1(n9810), .A2(n9809), .ZN(n9811) );
  AND2_X1 U10924 ( .A1(n9812), .A2(n9811), .ZN(n9823) );
  NAND2_X1 U10925 ( .A1(n9814), .A2(n9813), .ZN(n9815) );
  NAND2_X1 U10926 ( .A1(n9816), .A2(n9815), .ZN(n9817) );
  AOI22_X1 U10927 ( .A1(n9852), .A2(n9817), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n9821) );
  INV_X1 U10928 ( .A(n9818), .ZN(n9819) );
  NAND2_X1 U10929 ( .A1(n9839), .A2(n9819), .ZN(n9820) );
  OAI211_X1 U10930 ( .C1(n9823), .C2(n9822), .A(n9821), .B(n9820), .ZN(n9824)
         );
  INV_X1 U10931 ( .A(n9824), .ZN(n9830) );
  XOR2_X1 U10932 ( .A(n9826), .B(n9825), .Z(n9828) );
  NAND2_X1 U10933 ( .A1(n9828), .A2(n9827), .ZN(n9829) );
  OAI211_X1 U10934 ( .C1(n9957), .C2(n9831), .A(n9830), .B(n9829), .ZN(
        P2_U3183) );
  INV_X1 U10935 ( .A(n9832), .ZN(n9834) );
  NAND3_X1 U10936 ( .A1(n9835), .A2(n9834), .A3(n9833), .ZN(n9836) );
  NAND2_X1 U10937 ( .A1(n9837), .A2(n9836), .ZN(n9842) );
  INV_X1 U10938 ( .A(n9838), .ZN(n9840) );
  AOI222_X1 U10939 ( .A1(n9842), .A2(n5642), .B1(n9841), .B2(
        P2_ADDR_REG_4__SCAN_IN), .C1(n9840), .C2(n9839), .ZN(n9856) );
  AOI211_X1 U10940 ( .C1(n9846), .C2(n9845), .A(n9844), .B(n9843), .ZN(n9847)
         );
  INV_X1 U10941 ( .A(n9847), .ZN(n9854) );
  OAI21_X1 U10942 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9851) );
  NAND2_X1 U10943 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  NAND4_X1 U10944 ( .A1(n9856), .A2(n9855), .A3(n9854), .A4(n9853), .ZN(
        P2_U3186) );
  XOR2_X1 U10945 ( .A(n9857), .B(n9862), .Z(n9860) );
  AOI222_X1 U10946 ( .A1(n9861), .A2(n9860), .B1(n6877), .B2(n9859), .C1(n6922), .C2(n9858), .ZN(n9883) );
  XNOR2_X1 U10947 ( .A(n9863), .B(n9862), .ZN(n9886) );
  AOI222_X1 U10948 ( .A1(n9886), .A2(n9867), .B1(n9866), .B2(n9865), .C1(n6033), .C2(n9864), .ZN(n9868) );
  OAI221_X1 U10949 ( .B1(n9870), .B2(n9883), .C1(n8608), .C2(n9869), .A(n9868), 
        .ZN(P2_U3230) );
  INV_X1 U10950 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9876) );
  AOI21_X1 U10951 ( .B1(n9872), .B2(n9926), .A(n9871), .ZN(n9873) );
  AOI211_X1 U10952 ( .C1(n9875), .C2(n9931), .A(n9874), .B(n9873), .ZN(n9936)
         );
  AOI22_X1 U10953 ( .A1(n9934), .A2(n9876), .B1(n9936), .B2(n9932), .ZN(
        P2_U3390) );
  INV_X1 U10954 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9878) );
  AOI22_X1 U10955 ( .A1(n9934), .A2(n9878), .B1(n9877), .B2(n9932), .ZN(
        P2_U3393) );
  OAI22_X1 U10956 ( .A1(n9880), .A2(n9915), .B1(n9879), .B2(n9913), .ZN(n9882)
         );
  NOR2_X1 U10957 ( .A1(n9882), .A2(n9881), .ZN(n9938) );
  AOI22_X1 U10958 ( .A1(n9934), .A2(n6016), .B1(n9938), .B2(n9932), .ZN(
        P2_U3396) );
  INV_X1 U10959 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9887) );
  OAI21_X1 U10960 ( .B1(n9884), .B2(n9913), .A(n9883), .ZN(n9885) );
  AOI21_X1 U10961 ( .B1(n9921), .B2(n9886), .A(n9885), .ZN(n9939) );
  AOI22_X1 U10962 ( .A1(n9934), .A2(n9887), .B1(n9939), .B2(n9932), .ZN(
        P2_U3399) );
  INV_X1 U10963 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9893) );
  INV_X1 U10964 ( .A(n9888), .ZN(n9892) );
  OAI21_X1 U10965 ( .B1(n9890), .B2(n9913), .A(n9889), .ZN(n9891) );
  AOI21_X1 U10966 ( .B1(n9921), .B2(n9892), .A(n9891), .ZN(n9940) );
  AOI22_X1 U10967 ( .A1(n9934), .A2(n9893), .B1(n9940), .B2(n9932), .ZN(
        P2_U3402) );
  INV_X1 U10968 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U10969 ( .A1(n9895), .A2(n6431), .B1(n9931), .B2(n9894), .ZN(n9896)
         );
  AND2_X1 U10970 ( .A1(n9897), .A2(n9896), .ZN(n9942) );
  AOI22_X1 U10971 ( .A1(n9934), .A2(n9898), .B1(n9942), .B2(n9932), .ZN(
        P2_U3405) );
  OAI21_X1 U10972 ( .B1(n9900), .B2(n9913), .A(n9899), .ZN(n9901) );
  AOI21_X1 U10973 ( .B1(n9902), .B2(n9921), .A(n9901), .ZN(n9943) );
  AOI22_X1 U10974 ( .A1(n9934), .A2(n6062), .B1(n9943), .B2(n9932), .ZN(
        P2_U3408) );
  INV_X1 U10975 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U10976 ( .A1(n9903), .A2(n9913), .ZN(n9905) );
  AOI211_X1 U10977 ( .C1(n9906), .C2(n6431), .A(n9905), .B(n9904), .ZN(n9944)
         );
  AOI22_X1 U10978 ( .A1(n9934), .A2(n9907), .B1(n9944), .B2(n9932), .ZN(
        P2_U3411) );
  INV_X1 U10979 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9912) );
  OAI22_X1 U10980 ( .A1(n9909), .A2(n9915), .B1(n9908), .B2(n9913), .ZN(n9910)
         );
  NOR2_X1 U10981 ( .A1(n9911), .A2(n9910), .ZN(n9945) );
  AOI22_X1 U10982 ( .A1(n9934), .A2(n9912), .B1(n9945), .B2(n9932), .ZN(
        P2_U3417) );
  INV_X1 U10983 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9919) );
  OAI22_X1 U10984 ( .A1(n9916), .A2(n9915), .B1(n9914), .B2(n9913), .ZN(n9917)
         );
  NOR2_X1 U10985 ( .A1(n9918), .A2(n9917), .ZN(n9947) );
  AOI22_X1 U10986 ( .A1(n9934), .A2(n9919), .B1(n9947), .B2(n9932), .ZN(
        P2_U3420) );
  INV_X1 U10987 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U10988 ( .A1(n9922), .A2(n9921), .B1(n9931), .B2(n9920), .ZN(n9923)
         );
  AND2_X1 U10989 ( .A1(n9924), .A2(n9923), .ZN(n9949) );
  AOI22_X1 U10990 ( .A1(n9934), .A2(n9925), .B1(n9949), .B2(n9932), .ZN(
        P2_U3423) );
  INV_X1 U10991 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U10992 ( .A1(n9927), .A2(n9926), .ZN(n9929) );
  AOI211_X1 U10993 ( .C1(n9931), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9951)
         );
  AOI22_X1 U10994 ( .A1(n9934), .A2(n9933), .B1(n9951), .B2(n9932), .ZN(
        P2_U3426) );
  INV_X1 U10995 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U10996 ( .A1(n9952), .A2(n9936), .B1(n9935), .B2(n9950), .ZN(
        P2_U3459) );
  INV_X1 U10997 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U10998 ( .A1(n9952), .A2(n9938), .B1(n9937), .B2(n9950), .ZN(
        P2_U3461) );
  AOI22_X1 U10999 ( .A1(n9952), .A2(n9939), .B1(n6026), .B2(n9950), .ZN(
        P2_U3462) );
  AOI22_X1 U11000 ( .A1(n9952), .A2(n9940), .B1(n6034), .B2(n9950), .ZN(
        P2_U3463) );
  AOI22_X1 U11001 ( .A1(n9952), .A2(n9942), .B1(n9941), .B2(n9950), .ZN(
        P2_U3464) );
  AOI22_X1 U11002 ( .A1(n9952), .A2(n9943), .B1(n5653), .B2(n9950), .ZN(
        P2_U3465) );
  AOI22_X1 U11003 ( .A1(n9952), .A2(n9944), .B1(n6074), .B2(n9950), .ZN(
        P2_U3466) );
  AOI22_X1 U11004 ( .A1(n9952), .A2(n9945), .B1(n6098), .B2(n9950), .ZN(
        P2_U3468) );
  AOI22_X1 U11005 ( .A1(n9952), .A2(n9947), .B1(n9946), .B2(n9950), .ZN(
        P2_U3469) );
  AOI22_X1 U11006 ( .A1(n9952), .A2(n9949), .B1(n9948), .B2(n9950), .ZN(
        P2_U3470) );
  AOI22_X1 U11007 ( .A1(n9952), .A2(n9951), .B1(n6143), .B2(n9950), .ZN(
        P2_U3471) );
  OAI222_X1 U11008 ( .A1(n9957), .A2(n9956), .B1(n9957), .B2(n9955), .C1(n9954), .C2(n9953), .ZN(ADD_1068_U5) );
  XOR2_X1 U11009 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11010 ( .B1(n9960), .B2(n9959), .A(n9958), .ZN(n9962) );
  XOR2_X1 U11011 ( .A(n9962), .B(n9961), .Z(ADD_1068_U55) );
  OAI21_X1 U11012 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(ADD_1068_U56) );
  OAI21_X1 U11013 ( .B1(n9968), .B2(n9967), .A(n9966), .ZN(ADD_1068_U57) );
  OAI21_X1 U11014 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(ADD_1068_U58) );
  OAI21_X1 U11015 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(ADD_1068_U59) );
  OAI21_X1 U11016 ( .B1(n9977), .B2(n9976), .A(n9975), .ZN(ADD_1068_U60) );
  OAI21_X1 U11017 ( .B1(n9980), .B2(n9979), .A(n9978), .ZN(ADD_1068_U61) );
  OAI21_X1 U11018 ( .B1(n9983), .B2(n9982), .A(n9981), .ZN(ADD_1068_U62) );
  OAI21_X1 U11019 ( .B1(n9986), .B2(n9985), .A(n9984), .ZN(ADD_1068_U63) );
  OAI21_X1 U11020 ( .B1(n9989), .B2(n9988), .A(n9987), .ZN(ADD_1068_U50) );
  OAI21_X1 U11021 ( .B1(n9992), .B2(n9991), .A(n9990), .ZN(ADD_1068_U51) );
  OAI21_X1 U11022 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(ADD_1068_U47) );
  OAI21_X1 U11023 ( .B1(n9998), .B2(n9997), .A(n9996), .ZN(ADD_1068_U49) );
  OAI21_X1 U11024 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(ADD_1068_U48) );
  AOI21_X1 U11025 ( .B1(n10004), .B2(n10003), .A(n10002), .ZN(ADD_1068_U54) );
  AOI21_X1 U11026 ( .B1(n10007), .B2(n10006), .A(n10005), .ZN(ADD_1068_U53) );
  OAI21_X1 U11027 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(ADD_1068_U52) );
  CLKBUF_X3 U4779 ( .A(n4951), .Z(n7732) );
  CLKBUF_X1 U4794 ( .A(n4927), .Z(n5015) );
  INV_X1 U4819 ( .A(n5979), .ZN(n5982) );
  INV_X1 U4821 ( .A(n6865), .ZN(n6013) );
  CLKBUF_X1 U4891 ( .A(n4967), .Z(n7733) );
  CLKBUF_X1 U4899 ( .A(n6532), .Z(n4269) );
endmodule

