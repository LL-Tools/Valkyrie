

module b14_C_gen_AntiSAT_k_256_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071;

  NAND2_X2 U2468 ( .A1(n2358), .A2(n2278), .ZN(n2513) );
  INV_X1 U2469 ( .A(n3569), .ZN(n3557) );
  NAND2_X1 U2470 ( .A1(n3257), .A2(n3256), .ZN(n2406) );
  BUF_X1 U2471 ( .A(n3009), .Z(n3561) );
  NAND2_X1 U2472 ( .A1(n3108), .A2(n2397), .ZN(n2399) );
  CLKBUF_X2 U2473 ( .A(n2516), .Z(n2631) );
  NAND2_X1 U2474 ( .A1(n2460), .A2(IR_REG_31__SCAN_IN), .ZN(n2461) );
  AND4_X1 U2475 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n3199)
         );
  NAND3_X1 U2476 ( .A1(n2804), .A2(n2853), .A3(n4446), .ZN(n3012) );
  XNOR2_X2 U2477 ( .A(n2461), .B(IR_REG_29__SCAN_IN), .ZN(n2469) );
  OAI21_X1 U2478 ( .B1(n3700), .B2(n2425), .A(n2422), .ZN(n3640) );
  INV_X2 U2479 ( .A(n3184), .ZN(n2291) );
  AND2_X1 U2480 ( .A1(n3607), .A2(n3541), .ZN(n3611) );
  NAND2_X1 U2481 ( .A1(n4478), .A2(n4474), .ZN(n3617) );
  NAND2_X1 U2482 ( .A1(n4475), .A2(n4473), .ZN(n4478) );
  AOI21_X1 U2483 ( .B1(n3595), .B2(n3597), .A(n2440), .ZN(n3721) );
  INV_X1 U2484 ( .A(n2502), .ZN(n3282) );
  NAND2_X1 U2485 ( .A1(n2497), .A2(n2239), .ZN(n2502) );
  NAND4_X1 U2486 ( .A1(n2509), .A2(n2508), .A3(n2507), .A4(n2506), .ZN(n3900)
         );
  NAND4_X1 U2487 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .ZN(n3901)
         );
  INV_X2 U2488 ( .A(n2476), .ZN(n2717) );
  INV_X2 U2489 ( .A(n3552), .ZN(n3570) );
  NAND2_X1 U2490 ( .A1(n2276), .A2(n3012), .ZN(n3099) );
  AND2_X1 U2491 ( .A1(n2826), .A2(n3832), .ZN(n4664) );
  NAND2_X2 U2492 ( .A1(n3012), .A2(n3046), .ZN(n3569) );
  BUF_X2 U2493 ( .A(n2463), .Z(n4445) );
  XNOR2_X1 U2494 ( .A(n2459), .B(IR_REG_30__SCAN_IN), .ZN(n2463) );
  XNOR2_X1 U2495 ( .A(n2799), .B(IR_REG_24__SCAN_IN), .ZN(n4446) );
  XNOR2_X1 U2496 ( .A(n2801), .B(IR_REG_26__SCAN_IN), .ZN(n2804) );
  INV_X1 U2497 ( .A(n2807), .ZN(n3874) );
  NAND2_X1 U2498 ( .A1(n2856), .A2(IR_REG_31__SCAN_IN), .ZN(n2459) );
  NOR2_X1 U2499 ( .A1(n2312), .A2(IR_REG_28__SCAN_IN), .ZN(n2311) );
  AND3_X1 U2500 ( .A1(n2393), .A2(n2392), .A3(n2390), .ZN(n4455) );
  AND2_X1 U2501 ( .A1(n2484), .A2(n2498), .ZN(n2511) );
  INV_X1 U2502 ( .A(IR_REG_13__SCAN_IN), .ZN(n4793) );
  NOR2_X1 U2503 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2454)
         );
  INV_X1 U2504 ( .A(IR_REG_3__SCAN_IN), .ZN(n2498) );
  INV_X1 U2505 ( .A(IR_REG_4__SCAN_IN), .ZN(n2510) );
  NOR2_X1 U2506 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2447)
         );
  NOR2_X1 U2507 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2448)
         );
  NOR2_X1 U2508 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2449)
         );
  NOR2_X1 U2509 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2450)
         );
  AND2_X2 U2510 ( .A1(n2453), .A2(n2511), .ZN(n2381) );
  XNOR2_X1 U2511 ( .A(n2970), .B(n3552), .ZN(n2985) );
  INV_X1 U2512 ( .A(n3046), .ZN(n2276) );
  NAND2_X1 U2513 ( .A1(n3832), .A2(n3874), .ZN(n3046) );
  AOI21_X1 U2514 ( .B1(n2329), .B2(n2328), .A(n2327), .ZN(n4014) );
  NOR2_X1 U2515 ( .A1(n2226), .A2(n2231), .ZN(n2328) );
  OAI21_X1 U2516 ( .B1(n2227), .B2(n2231), .A(n2261), .ZN(n2327) );
  OAI21_X1 U2517 ( .B1(n2835), .B2(n3825), .A(n2834), .ZN(n2836) );
  OR2_X1 U2518 ( .A1(n2838), .A2(n2744), .ZN(n2438) );
  NAND2_X1 U2519 ( .A1(n2345), .A2(n2258), .ZN(n2342) );
  AND2_X1 U2520 ( .A1(n4274), .A2(n3580), .ZN(n3868) );
  NOR2_X1 U2521 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2456)
         );
  NAND2_X1 U2522 ( .A1(n2246), .A2(n2456), .ZN(n2285) );
  AND2_X1 U2523 ( .A1(n2408), .A2(n2455), .ZN(n2380) );
  NOR2_X1 U2524 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2455)
         );
  INV_X1 U2525 ( .A(IR_REG_22__SCAN_IN), .ZN(n2733) );
  NOR2_X1 U2526 ( .A1(n2409), .A2(IR_REG_18__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U2527 ( .A1(n2454), .A2(n2410), .ZN(n2409) );
  INV_X1 U2528 ( .A(n2428), .ZN(n2423) );
  AOI21_X1 U2529 ( .B1(n2432), .B2(n2431), .A(n2429), .ZN(n2428) );
  AND2_X1 U2530 ( .A1(n3549), .A2(n3548), .ZN(n2429) );
  OAI22_X1 U2531 ( .A1(n3282), .A2(n3572), .B1(n3569), .B2(n3101), .ZN(n3100)
         );
  NAND2_X1 U2532 ( .A1(n3103), .A2(n3102), .ZN(n3108) );
  NAND2_X1 U2533 ( .A1(n2433), .A2(n2967), .ZN(n2970) );
  OAI22_X1 U2534 ( .A1(n3572), .A2(n3085), .B1(n3184), .B2(n2984), .ZN(n2275)
         );
  NAND2_X1 U2535 ( .A1(n4510), .A2(n4511), .ZN(n4509) );
  XNOR2_X1 U2536 ( .A(n3942), .B(n2319), .ZN(n4522) );
  NAND2_X1 U2537 ( .A1(n4531), .A2(n4532), .ZN(n4530) );
  XNOR2_X1 U2538 ( .A(n3945), .B(n2320), .ZN(n4543) );
  AOI21_X1 U2539 ( .B1(n2332), .B2(n2334), .A(n2248), .ZN(n2331) );
  INV_X1 U2540 ( .A(n2335), .ZN(n2332) );
  INV_X1 U2541 ( .A(n2334), .ZN(n2333) );
  NOR2_X1 U2542 ( .A1(n2373), .A2(n2559), .ZN(n2372) );
  INV_X1 U2543 ( .A(n2374), .ZN(n2373) );
  OR2_X1 U2544 ( .A1(n2845), .A2(n3839), .ZN(n4264) );
  OR2_X1 U2545 ( .A1(n4018), .A2(n3580), .ZN(n2845) );
  NAND2_X1 U2546 ( .A1(n4040), .A2(n4019), .ZN(n4018) );
  XNOR2_X1 U2547 ( .A(n2739), .B(n2738), .ZN(n3832) );
  INV_X1 U2548 ( .A(IR_REG_20__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U2549 ( .A1(n4006), .A2(n2260), .ZN(n2352) );
  NAND2_X1 U2550 ( .A1(n3839), .A2(n4366), .ZN(n2301) );
  NAND2_X1 U2551 ( .A1(n2300), .A2(n4699), .ZN(n2299) );
  NAND2_X1 U2552 ( .A1(n4001), .A2(n4676), .ZN(n2300) );
  AND2_X1 U2553 ( .A1(n3731), .A2(n4064), .ZN(n3863) );
  INV_X1 U2554 ( .A(n3237), .ZN(n3235) );
  NAND2_X1 U2555 ( .A1(n3690), .A2(n3691), .ZN(n2418) );
  AOI21_X1 U2556 ( .B1(n2416), .B2(n2418), .A(n2415), .ZN(n2414) );
  INV_X1 U2557 ( .A(n3597), .ZN(n2415) );
  INV_X1 U2558 ( .A(n2419), .ZN(n2416) );
  INV_X1 U2559 ( .A(n2418), .ZN(n2417) );
  INV_X1 U2560 ( .A(n3596), .ZN(n2413) );
  INV_X1 U2561 ( .A(n2463), .ZN(n2466) );
  NOR2_X1 U2562 ( .A1(n2296), .A2(n3766), .ZN(n2295) );
  NAND2_X1 U2563 ( .A1(n4065), .A2(n3863), .ZN(n2297) );
  OR2_X1 U2564 ( .A1(n4307), .A2(n4116), .ZN(n4090) );
  INV_X1 U2565 ( .A(n2238), .ZN(n2357) );
  INV_X1 U2566 ( .A(n2356), .ZN(n2355) );
  OAI21_X1 U2567 ( .B1(n4190), .B2(n2357), .A(n2662), .ZN(n2356) );
  NAND2_X1 U2568 ( .A1(n4472), .A2(n2661), .ZN(n2662) );
  OR2_X1 U2569 ( .A1(n4199), .A2(n4083), .ZN(n4162) );
  INV_X1 U2570 ( .A(n4246), .ZN(n3333) );
  NOR2_X1 U2571 ( .A1(n2379), .A2(n2547), .ZN(n2378) );
  INV_X1 U2572 ( .A(n2534), .ZN(n2379) );
  OAI21_X1 U2573 ( .B1(n2365), .B2(n2364), .A(n2360), .ZN(n3069) );
  NAND2_X1 U2574 ( .A1(n2242), .A2(n2485), .ZN(n2364) );
  AOI21_X1 U2575 ( .B1(n2242), .B2(n2362), .A(n2361), .ZN(n2360) );
  INV_X1 U2576 ( .A(n3086), .ZN(n2933) );
  OR2_X1 U2577 ( .A1(n4175), .A2(n4143), .ZN(n4127) );
  NAND2_X1 U2578 ( .A1(n5042), .A2(n2437), .ZN(n2436) );
  INV_X1 U2579 ( .A(IR_REG_25__SCAN_IN), .ZN(n2437) );
  NOR2_X1 U2580 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2317)
         );
  INV_X1 U2581 ( .A(n3294), .ZN(n2274) );
  AOI21_X1 U2582 ( .B1(n2241), .B2(n3294), .A(n2273), .ZN(n2272) );
  INV_X1 U2583 ( .A(n3347), .ZN(n2273) );
  XNOR2_X1 U2584 ( .A(n3008), .B(n3570), .ZN(n3104) );
  AND2_X1 U2585 ( .A1(n2969), .A2(n3046), .ZN(n3552) );
  AND2_X1 U2586 ( .A1(n3608), .A2(n3609), .ZN(n3541) );
  NAND2_X1 U2587 ( .A1(n3672), .A2(n3546), .ZN(n2430) );
  INV_X1 U2588 ( .A(n3701), .ZN(n2424) );
  NAND2_X1 U2589 ( .A1(n3545), .A2(n3546), .ZN(n2432) );
  INV_X1 U2590 ( .A(n3611), .ZN(n2277) );
  NAND2_X1 U2591 ( .A1(n2474), .A2(n2457), .ZN(n2358) );
  NAND2_X1 U2592 ( .A1(n2438), .A2(IR_REG_27__SCAN_IN), .ZN(n2278) );
  INV_X1 U2593 ( .A(n3148), .ZN(n2395) );
  NOR2_X1 U2594 ( .A1(n3149), .A2(n2398), .ZN(n2397) );
  INV_X1 U2595 ( .A(n3107), .ZN(n2398) );
  NAND2_X1 U2596 ( .A1(n2505), .A2(REG3_REG_5__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U2597 ( .A1(n2894), .A2(n2893), .ZN(n2896) );
  XNOR2_X1 U2598 ( .A(n3939), .B(n2314), .ZN(n4501) );
  NAND2_X1 U2599 ( .A1(n4509), .A2(n3967), .ZN(n3968) );
  NAND2_X1 U2600 ( .A1(n4512), .A2(n3941), .ZN(n3942) );
  NAND2_X1 U2601 ( .A1(n4522), .A2(REG2_REG_10__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U2602 ( .A1(n4533), .A2(n3944), .ZN(n3945) );
  NAND2_X1 U2603 ( .A1(n4543), .A2(REG2_REG_12__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U2604 ( .A1(n4530), .A2(n2256), .ZN(n3970) );
  NAND2_X1 U2605 ( .A1(n4590), .A2(n2264), .ZN(n2325) );
  AND2_X1 U2606 ( .A1(n2715), .A2(n2708), .ZN(n4043) );
  NOR2_X1 U2607 ( .A1(n2698), .A2(n2336), .ZN(n2335) );
  INV_X1 U2608 ( .A(n2691), .ZN(n2336) );
  NAND2_X1 U2609 ( .A1(n2251), .A2(n2338), .ZN(n2334) );
  AND3_X1 U2610 ( .A1(n2697), .A2(n2696), .A3(n2695), .ZN(n4097) );
  OAI21_X1 U2611 ( .B1(n2671), .B2(n2439), .A(n2670), .ZN(n4124) );
  INV_X1 U2612 ( .A(n3754), .ZN(n2670) );
  INV_X1 U2613 ( .A(n4307), .ZN(n4135) );
  NAND2_X1 U2614 ( .A1(n4183), .A2(n4190), .ZN(n4182) );
  OR2_X1 U2615 ( .A1(n4337), .A2(n4460), .ZN(n2630) );
  OAI21_X1 U2616 ( .B1(n3451), .B2(n2619), .A(n2618), .ZN(n4226) );
  OR2_X1 U2617 ( .A1(n2579), .A2(n5047), .ZN(n2591) );
  OR2_X1 U2618 ( .A1(n3333), .A2(n2763), .ZN(n2345) );
  NOR2_X1 U2619 ( .A1(n2589), .A2(n2344), .ZN(n2343) );
  INV_X1 U2620 ( .A(n2577), .ZN(n2344) );
  NAND2_X1 U2621 ( .A1(n2570), .A2(REG3_REG_11__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U2622 ( .A1(n2368), .A2(n2366), .ZN(n3332) );
  INV_X1 U2623 ( .A(n2367), .ZN(n2366) );
  NAND2_X1 U2624 ( .A1(n2535), .A2(n2229), .ZN(n2368) );
  OAI21_X1 U2625 ( .B1(n2372), .B2(n2370), .A(n2569), .ZN(n2367) );
  NAND2_X1 U2626 ( .A1(n2376), .A2(n2375), .ZN(n2374) );
  NOR2_X1 U2627 ( .A1(n2514), .A2(n2907), .ZN(n2525) );
  OAI21_X1 U2628 ( .B1(n3118), .B2(n3117), .A(n3795), .ZN(n3134) );
  AND2_X1 U2629 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2505) );
  NAND2_X1 U2630 ( .A1(n3012), .A2(n4641), .ZN(n3040) );
  AND2_X1 U2631 ( .A1(n4054), .A2(n4042), .ZN(n4040) );
  MUX2_X1 U2632 ( .A(n3960), .B(DATAI_9_), .S(n2513), .Z(n3306) );
  INV_X1 U2633 ( .A(n2285), .ZN(n2283) );
  AND3_X1 U2634 ( .A1(n2381), .A2(n2380), .A3(n2246), .ZN(n2797) );
  NAND2_X1 U2635 ( .A1(n2381), .A2(n2408), .ZN(n2659) );
  INV_X1 U2636 ( .A(IR_REG_31__SCAN_IN), .ZN(n2796) );
  AND2_X1 U2637 ( .A1(n2468), .A2(n2467), .ZN(n2472) );
  NAND2_X1 U2638 ( .A1(n2990), .A2(n2989), .ZN(n3005) );
  INV_X1 U2639 ( .A(n2993), .ZN(n2989) );
  OAI211_X1 U2640 ( .C1(n4100), .C2(n2486), .A(n2690), .B(n2689), .ZN(n4289)
         );
  INV_X1 U2641 ( .A(n4172), .ZN(n4334) );
  NAND4_X1 U2642 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n4368)
         );
  NAND4_X1 U2643 ( .A1(n2555), .A2(n2554), .A3(n2553), .A4(n2552), .ZN(n3896)
         );
  INV_X1 U2644 ( .A(n3321), .ZN(n3898) );
  XNOR2_X1 U2645 ( .A(n3970), .B(n2320), .ZN(n4548) );
  NAND2_X1 U2646 ( .A1(n4559), .A2(n4560), .ZN(n4558) );
  AND2_X1 U2647 ( .A1(n2880), .A2(n2881), .ZN(n4604) );
  INV_X1 U2648 ( .A(n2324), .ZN(n2323) );
  AOI21_X1 U2649 ( .B1(n2325), .B2(n4602), .A(n4600), .ZN(n2324) );
  NOR2_X1 U2650 ( .A1(n2325), .A2(n4602), .ZN(n4601) );
  OR2_X1 U2651 ( .A1(n4596), .A2(n2386), .ZN(n4605) );
  INV_X1 U2652 ( .A(n4252), .ZN(n4623) );
  INV_X1 U2653 ( .A(n2352), .ZN(n2350) );
  XNOR2_X1 U2654 ( .A(n2351), .B(n3763), .ZN(n4001) );
  OAI21_X1 U2655 ( .B1(n2833), .B2(n2832), .A(n2257), .ZN(n2351) );
  INV_X1 U2656 ( .A(n2347), .ZN(n2346) );
  OAI21_X1 U2657 ( .B1(n2352), .B2(n2348), .A(n2236), .ZN(n2347) );
  NAND2_X1 U2658 ( .A1(n4687), .A2(n4341), .ZN(n2348) );
  OAI21_X1 U2659 ( .B1(n2846), .B2(n4003), .A(n4264), .ZN(n4008) );
  NOR2_X1 U2660 ( .A1(n2754), .A2(n2363), .ZN(n2362) );
  INV_X1 U2661 ( .A(n2485), .ZN(n2363) );
  INV_X1 U2662 ( .A(IR_REG_16__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U2663 ( .A1(n2421), .A2(n2420), .ZN(n2419) );
  NAND2_X1 U2664 ( .A1(n3477), .A2(n3476), .ZN(n2268) );
  NAND2_X1 U2665 ( .A1(n2389), .A2(n2388), .ZN(n2955) );
  NAND2_X1 U2666 ( .A1(n4452), .A2(REG1_REG_5__SCAN_IN), .ZN(n2388) );
  INV_X1 U2667 ( .A(n2910), .ZN(n2389) );
  INV_X1 U2668 ( .A(n2863), .ZN(n2823) );
  OAI21_X1 U2669 ( .B1(n2295), .B2(n2294), .A(n2293), .ZN(n2292) );
  INV_X1 U2670 ( .A(n3861), .ZN(n2294) );
  AND2_X1 U2671 ( .A1(n2763), .A2(n3370), .ZN(n2282) );
  AND2_X1 U2672 ( .A1(n2289), .A2(n3235), .ZN(n2288) );
  AND2_X1 U2673 ( .A1(n3101), .A2(n3154), .ZN(n2290) );
  INV_X1 U2674 ( .A(IR_REG_19__SCAN_IN), .ZN(n2735) );
  OR2_X1 U2675 ( .A1(n2567), .A2(IR_REG_9__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U2676 ( .A1(n2270), .A2(n2418), .ZN(n3595) );
  NAND2_X1 U2677 ( .A1(n2269), .A2(n2267), .ZN(n2270) );
  AND2_X1 U2678 ( .A1(n2419), .A2(n2268), .ZN(n2267) );
  NAND2_X1 U2679 ( .A1(n3478), .A2(n3476), .ZN(n2269) );
  AND4_X1 U2680 ( .A1(n2928), .A2(n2927), .A3(n2926), .A4(n2925), .ZN(n2978)
         );
  INV_X1 U2681 ( .A(n3261), .ZN(n2405) );
  OR2_X1 U2682 ( .A1(n2663), .A2(n4822), .ZN(n2673) );
  NAND2_X1 U2683 ( .A1(n2407), .A2(n2247), .ZN(n3368) );
  INV_X1 U2684 ( .A(n4042), .ZN(n3713) );
  AOI21_X1 U2685 ( .B1(n2414), .B2(n2417), .A(n2413), .ZN(n2412) );
  OR2_X1 U2686 ( .A1(n2486), .A2(n2475), .ZN(n2928) );
  XNOR2_X1 U2687 ( .A(n2879), .B(n3065), .ZN(n3059) );
  NAND2_X1 U2688 ( .A1(n3059), .A2(REG1_REG_4__SCAN_IN), .ZN(n3062) );
  OAI21_X1 U2689 ( .B1(n3058), .B2(n2895), .A(n2897), .ZN(n2898) );
  XNOR2_X1 U2690 ( .A(n2955), .B(n4451), .ZN(n2912) );
  NAND2_X1 U2691 ( .A1(n2315), .A2(n2259), .ZN(n3939) );
  INV_X1 U2692 ( .A(n3937), .ZN(n2315) );
  NAND2_X1 U2693 ( .A1(n4501), .A2(REG2_REG_8__SCAN_IN), .ZN(n4500) );
  NAND2_X1 U2694 ( .A1(n4505), .A2(n3966), .ZN(n4510) );
  NAND2_X1 U2695 ( .A1(n4526), .A2(n3969), .ZN(n4531) );
  NAND2_X1 U2696 ( .A1(n4558), .A2(n3972), .ZN(n3974) );
  NAND2_X1 U2697 ( .A1(n4607), .A2(n2387), .ZN(n2386) );
  INV_X1 U2698 ( .A(n3982), .ZN(n2387) );
  INV_X1 U2699 ( .A(n2386), .ZN(n2385) );
  NAND2_X1 U2700 ( .A1(n2297), .A2(n2295), .ZN(n4032) );
  NAND2_X1 U2701 ( .A1(n2297), .A2(n3765), .ZN(n4048) );
  NAND2_X1 U2702 ( .A1(n2687), .A2(REG3_REG_23__SCAN_IN), .ZN(n2692) );
  INV_X1 U2703 ( .A(n4099), .ZN(n4094) );
  NOR2_X1 U2704 ( .A1(n2673), .A2(n2672), .ZN(n2683) );
  AOI21_X1 U2705 ( .B1(n2355), .B2(n2357), .A(n2230), .ZN(n2354) );
  OR2_X1 U2706 ( .A1(n4162), .A2(n4085), .ZN(n4153) );
  NAND2_X1 U2707 ( .A1(n2653), .A2(REG3_REG_19__SCAN_IN), .ZN(n2663) );
  AND4_X1 U2708 ( .A1(n2650), .A2(n2649), .A3(n2648), .A4(n2647), .ZN(n4172)
         );
  AND2_X1 U2709 ( .A1(n2645), .A2(REG3_REG_18__SCAN_IN), .ZN(n2653) );
  OR2_X1 U2710 ( .A1(n2620), .A2(n5041), .ZN(n2633) );
  NAND2_X1 U2711 ( .A1(n2610), .A2(REG3_REG_15__SCAN_IN), .ZN(n2620) );
  INV_X1 U2712 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4957) );
  OAI21_X1 U2713 ( .B1(n2578), .B2(n2342), .A(n2340), .ZN(n3380) );
  INV_X1 U2714 ( .A(n2341), .ZN(n2340) );
  OAI21_X1 U2715 ( .B1(n2343), .B2(n2342), .A(n2600), .ZN(n2341) );
  AOI21_X1 U2716 ( .B1(n2305), .B2(n2304), .A(n2303), .ZN(n2302) );
  INV_X1 U2717 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4847) );
  OAI21_X1 U2718 ( .B1(n3208), .B2(n2760), .A(n3786), .ZN(n3320) );
  NAND2_X1 U2719 ( .A1(n2309), .A2(n3782), .ZN(n3208) );
  NAND2_X1 U2720 ( .A1(n3134), .A2(n3794), .ZN(n2309) );
  OR2_X1 U2721 ( .A1(n3070), .A2(n2756), .ZN(n2757) );
  INV_X1 U2722 ( .A(n3110), .ZN(n3101) );
  NAND2_X1 U2723 ( .A1(n2308), .A2(n3771), .ZN(n3024) );
  NAND2_X1 U2724 ( .A1(n3181), .A2(n3180), .ZN(n2308) );
  NOR2_X1 U2725 ( .A1(n4264), .A2(n4267), .ZN(n4263) );
  AOI21_X1 U2726 ( .B1(n4014), .B2(n2723), .A(n2722), .ZN(n2833) );
  NOR2_X1 U2727 ( .A1(n3868), .A2(n3825), .ZN(n2832) );
  AND2_X1 U2728 ( .A1(n2732), .A2(n2731), .ZN(n4274) );
  AND2_X1 U2729 ( .A1(n4128), .A2(n2235), .ZN(n4054) );
  NAND2_X1 U2730 ( .A1(n4128), .A2(n2234), .ZN(n4070) );
  NAND2_X1 U2731 ( .A1(n2513), .A2(DATAI_23_), .ZN(n4099) );
  NAND2_X1 U2732 ( .A1(n4128), .A2(n2233), .ZN(n4098) );
  AND2_X1 U2733 ( .A1(n4128), .A2(n4116), .ZN(n4114) );
  NOR2_X1 U2734 ( .A1(n4127), .A2(n4306), .ZN(n4128) );
  INV_X1 U2735 ( .A(n4133), .ZN(n4306) );
  INV_X1 U2736 ( .A(n4316), .ZN(n4143) );
  NOR2_X1 U2737 ( .A1(n4203), .A2(n4483), .ZN(n4185) );
  NAND2_X1 U2738 ( .A1(n4185), .A2(n4173), .ZN(n4175) );
  NAND2_X1 U2739 ( .A1(n2287), .A2(n4211), .ZN(n4203) );
  AND4_X1 U2740 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(n4337)
         );
  INV_X1 U2741 ( .A(n4347), .ZN(n3456) );
  AND2_X1 U2742 ( .A1(n3391), .A2(n2281), .ZN(n3452) );
  AND2_X1 U2743 ( .A1(n2232), .A2(n3484), .ZN(n2281) );
  NAND2_X1 U2744 ( .A1(n3452), .A2(n3456), .ZN(n4229) );
  AND4_X1 U2745 ( .A1(n2606), .A2(n2605), .A3(n2604), .A4(n2603), .ZN(n4351)
         );
  NAND2_X1 U2746 ( .A1(n3391), .A2(n2282), .ZN(n4249) );
  NAND2_X1 U2747 ( .A1(n3391), .A2(n3370), .ZN(n3410) );
  AND4_X1 U2748 ( .A1(n2575), .A2(n2574), .A3(n2573), .A4(n2572), .ZN(n4372)
         );
  AND2_X1 U2749 ( .A1(n3393), .A2(n3396), .ZN(n3391) );
  NOR2_X1 U2750 ( .A1(n3317), .A2(n3306), .ZN(n3393) );
  OR2_X1 U2751 ( .A1(n3206), .A2(n3274), .ZN(n3317) );
  AND3_X1 U2752 ( .A1(n3076), .A2(n2290), .A3(n2289), .ZN(n3205) );
  AND4_X1 U2753 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n3321)
         );
  NAND2_X1 U2754 ( .A1(n3076), .A2(n2290), .ZN(n3136) );
  NAND2_X1 U2755 ( .A1(n3076), .A2(n3101), .ZN(n3123) );
  NOR2_X1 U2756 ( .A1(n3177), .A2(n3182), .ZN(n3176) );
  AND2_X1 U2757 ( .A1(n3176), .A2(n3194), .ZN(n3076) );
  INV_X1 U2758 ( .A(n4320), .ZN(n4371) );
  INV_X1 U2759 ( .A(n4664), .ZN(n4679) );
  AND3_X1 U2760 ( .A1(n2820), .A2(n2819), .A3(n2918), .ZN(n2828) );
  NAND2_X1 U2761 ( .A1(n2434), .A2(n2246), .ZN(n2312) );
  NOR2_X1 U2762 ( .A1(n2436), .A2(n2435), .ZN(n2434) );
  NAND2_X1 U2763 ( .A1(n2456), .A2(n2457), .ZN(n2435) );
  NAND2_X1 U2764 ( .A1(n2286), .A2(IR_REG_31__SCAN_IN), .ZN(n2838) );
  NOR2_X1 U2765 ( .A1(n2285), .A2(n2436), .ZN(n2284) );
  XNOR2_X1 U2766 ( .A(n2734), .B(n2733), .ZN(n2943) );
  XNOR2_X1 U2767 ( .A(n2741), .B(n2313), .ZN(n2807) );
  NOR2_X1 U2768 ( .A1(n2617), .A2(n2409), .ZN(n2651) );
  NOR2_X1 U2769 ( .A1(n2598), .A2(IR_REG_5__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U2770 ( .A1(n2249), .A2(IR_REG_1__SCAN_IN), .ZN(n2318) );
  NOR2_X1 U2771 ( .A1(n2317), .A2(n2482), .ZN(n2316) );
  NAND2_X1 U2772 ( .A1(n2402), .A2(n3709), .ZN(n3589) );
  NAND2_X1 U2773 ( .A1(n2407), .A2(n3352), .ZN(n3355) );
  NAND2_X1 U2774 ( .A1(n2402), .A2(n2400), .ZN(n2404) );
  NOR2_X1 U2775 ( .A1(n3588), .A2(n2401), .ZN(n2400) );
  INV_X1 U2776 ( .A(n3709), .ZN(n2401) );
  NAND2_X1 U2777 ( .A1(n2406), .A2(n3261), .ZN(n3292) );
  INV_X1 U2778 ( .A(n3085), .ZN(n3088) );
  INV_X1 U2779 ( .A(n2426), .ZN(n2425) );
  AOI21_X1 U2780 ( .B1(n2424), .B2(n2426), .A(n2423), .ZN(n2422) );
  AND2_X1 U2781 ( .A1(n3541), .A2(n2430), .ZN(n2426) );
  INV_X1 U2782 ( .A(n4228), .ZN(n4460) );
  NAND2_X1 U2783 ( .A1(n2399), .A2(n3148), .ZN(n3652) );
  OAI21_X1 U2784 ( .B1(n3611), .B2(n3549), .A(n3548), .ZN(n3671) );
  NAND2_X1 U2785 ( .A1(n2277), .A2(n2427), .ZN(n3670) );
  INV_X1 U2786 ( .A(n2432), .ZN(n2427) );
  NAND2_X1 U2787 ( .A1(n3108), .A2(n3107), .ZN(n3150) );
  OAI21_X1 U2788 ( .B1(n2271), .B2(n2241), .A(n3294), .ZN(n3348) );
  INV_X1 U2789 ( .A(n2406), .ZN(n2271) );
  INV_X1 U2790 ( .A(DATAI_0_), .ZN(n2279) );
  NAND2_X1 U2791 ( .A1(n3518), .A2(n3517), .ZN(n3519) );
  INV_X1 U2792 ( .A(n3515), .ZN(n3518) );
  NAND2_X1 U2793 ( .A1(n2266), .A2(n3476), .ZN(n3693) );
  OR2_X1 U2794 ( .A1(n3478), .A2(n3477), .ZN(n2266) );
  AND2_X1 U2795 ( .A1(n2681), .A2(n2680), .ZN(n4318) );
  NAND2_X1 U2796 ( .A1(n2986), .A2(n2275), .ZN(n2987) );
  INV_X1 U2797 ( .A(n4458), .ZN(n4481) );
  AOI21_X1 U2798 ( .B1(n3651), .B2(n2395), .A(n2245), .ZN(n2394) );
  INV_X1 U2799 ( .A(n3651), .ZN(n2396) );
  AOI21_X1 U2800 ( .B1(n3640), .B2(n3637), .A(n3636), .ZN(n3710) );
  AND2_X1 U2801 ( .A1(n3016), .A2(n3015), .ZN(n4488) );
  NAND2_X1 U2802 ( .A1(n2714), .A2(n2713), .ZN(n4271) );
  NAND2_X1 U2803 ( .A1(n2704), .A2(n2703), .ZN(n4037) );
  INV_X1 U2804 ( .A(n4097), .ZN(n3892) );
  OR2_X1 U2805 ( .A1(n3757), .A2(n4118), .ZN(n2685) );
  INV_X1 U2806 ( .A(n4318), .ZN(n4145) );
  NAND4_X1 U2807 ( .A1(n2669), .A2(n2668), .A3(n2667), .A4(n2666), .ZN(n4169)
         );
  INV_X1 U2808 ( .A(n4337), .ZN(n4348) );
  NAND4_X1 U2809 ( .A1(n2616), .A2(n2615), .A3(n2614), .A4(n2613), .ZN(n4217)
         );
  NAND4_X1 U2810 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n4246)
         );
  INV_X1 U2811 ( .A(n4372), .ZN(n3894) );
  NAND4_X1 U2812 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n3895)
         );
  NAND4_X1 U2813 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n3899)
         );
  NAND2_X1 U2814 ( .A1(n3908), .A2(n3909), .ZN(n3907) );
  NAND2_X1 U2815 ( .A1(n3920), .A2(n3921), .ZN(n3919) );
  NAND2_X1 U2816 ( .A1(n3918), .A2(n3917), .ZN(n3916) );
  XNOR2_X1 U2817 ( .A(n2896), .B(n4453), .ZN(n3058) );
  AND2_X1 U2818 ( .A1(n3062), .A2(n2382), .ZN(n2884) );
  NAND2_X1 U2819 ( .A1(n2879), .A2(n4453), .ZN(n2382) );
  NOR2_X1 U2820 ( .A1(n2961), .A2(n2960), .ZN(n3937) );
  XNOR2_X1 U2821 ( .A(n3968), .B(n2319), .ZN(n4527) );
  NAND2_X1 U2822 ( .A1(n4521), .A2(n3943), .ZN(n4534) );
  AND2_X1 U2823 ( .A1(n4496), .A2(n3884), .ZN(n4552) );
  NAND2_X1 U2824 ( .A1(n4542), .A2(n3946), .ZN(n4554) );
  NAND2_X1 U2825 ( .A1(n4547), .A2(n3971), .ZN(n4559) );
  XNOR2_X1 U2826 ( .A(n3974), .B(n4648), .ZN(n4568) );
  AOI21_X1 U2827 ( .B1(n4604), .B2(ADDR_REG_18__SCAN_IN), .A(n4603), .ZN(n2322) );
  AOI21_X1 U2828 ( .B1(n4594), .B2(n2385), .A(n2265), .ZN(n2384) );
  OAI21_X1 U2829 ( .B1(n4081), .B2(n2226), .A(n2227), .ZN(n4030) );
  NAND2_X1 U2830 ( .A1(n2330), .A2(n2334), .ZN(n4053) );
  NAND2_X1 U2831 ( .A1(n4081), .A2(n2335), .ZN(n2330) );
  NAND2_X1 U2832 ( .A1(n4081), .A2(n2691), .ZN(n2337) );
  NAND2_X1 U2833 ( .A1(n2513), .A2(DATAI_21_), .ZN(n4133) );
  NAND2_X1 U2834 ( .A1(n4182), .A2(n2238), .ZN(n4160) );
  NAND2_X1 U2835 ( .A1(n2339), .A2(n2345), .ZN(n4247) );
  NAND2_X1 U2836 ( .A1(n2578), .A2(n2343), .ZN(n2339) );
  NAND2_X1 U2837 ( .A1(n2371), .A2(n2558), .ZN(n3394) );
  NAND2_X1 U2838 ( .A1(n2377), .A2(n2372), .ZN(n2371) );
  NAND2_X1 U2839 ( .A1(n2377), .A2(n2374), .ZN(n3247) );
  NAND2_X1 U2840 ( .A1(n2535), .A2(n2534), .ZN(n3319) );
  INV_X1 U2841 ( .A(n4227), .ZN(n4259) );
  NAND2_X1 U2842 ( .A1(n4256), .A2(n3084), .ZN(n4252) );
  OAI21_X1 U2843 ( .B1(n2825), .B2(n3472), .A(n2845), .ZN(n3466) );
  AND2_X2 U2844 ( .A1(n2828), .A2(n3044), .ZN(n4687) );
  NAND2_X1 U2845 ( .A1(n2237), .A2(IR_REG_31__SCAN_IN), .ZN(n2801) );
  AND2_X1 U2846 ( .A1(n3011), .A2(STATE_REG_SCAN_IN), .ZN(n4641) );
  INV_X1 U2847 ( .A(n2943), .ZN(n4447) );
  XNOR2_X1 U2848 ( .A(n2736), .B(IR_REG_19__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U2849 ( .A1(n2796), .A2(n2391), .ZN(n2390) );
  INV_X1 U2850 ( .A(n2484), .ZN(n2393) );
  NAND2_X1 U2851 ( .A1(n2483), .A2(IR_REG_2__SCAN_IN), .ZN(n2392) );
  INV_X1 U2852 ( .A(n2321), .ZN(n4609) );
  OAI21_X1 U2853 ( .B1(n4601), .B2(n2323), .A(n2322), .ZN(n2321) );
  OR2_X1 U2854 ( .A1(n4008), .A2(n4377), .ZN(n2847) );
  OAI21_X1 U2855 ( .B1(n2352), .B2(n2299), .A(n2298), .ZN(n2848) );
  NAND2_X1 U2856 ( .A1(n4696), .A2(n2844), .ZN(n2298) );
  OAI21_X1 U2857 ( .B1(n2349), .B2(n4001), .A(n2346), .ZN(n2850) );
  NAND2_X1 U2858 ( .A1(n2350), .A2(n4687), .ZN(n2349) );
  OR2_X1 U2859 ( .A1(n2333), .A2(n2240), .ZN(n2226) );
  CLKBUF_X3 U2860 ( .A(n3099), .Z(n3572) );
  OR2_X1 U2861 ( .A1(n2331), .A2(n2240), .ZN(n2227) );
  INV_X1 U2862 ( .A(n3897), .ZN(n2375) );
  NAND2_X1 U2863 ( .A1(n2250), .A2(n2558), .ZN(n2370) );
  INV_X1 U2864 ( .A(n3765), .ZN(n2296) );
  NOR2_X1 U2865 ( .A1(n3127), .A2(n2524), .ZN(n2228) );
  AND2_X1 U2866 ( .A1(n2378), .A2(n2369), .ZN(n2229) );
  AND2_X1 U2867 ( .A1(n4151), .A2(n4173), .ZN(n2230) );
  AND2_X1 U2868 ( .A1(n4271), .A2(n3713), .ZN(n2231) );
  INV_X1 U2869 ( .A(n3787), .ZN(n2304) );
  AND2_X1 U2870 ( .A1(n2282), .A2(n4250), .ZN(n2232) );
  AND2_X1 U2871 ( .A1(n4099), .A2(n4116), .ZN(n2233) );
  AND2_X1 U2872 ( .A1(n2233), .A2(n4074), .ZN(n2234) );
  XNOR2_X1 U2873 ( .A(n2985), .B(n2275), .ZN(n2974) );
  NAND2_X1 U2874 ( .A1(n2381), .A2(n2454), .ZN(n2640) );
  AND2_X1 U2875 ( .A1(n2234), .A2(n4056), .ZN(n2235) );
  OR2_X1 U2876 ( .A1(n3033), .A2(n3832), .ZN(n4315) );
  INV_X1 U2877 ( .A(n4315), .ZN(n4366) );
  OR2_X1 U2878 ( .A1(n4687), .A2(REG0_REG_29__SCAN_IN), .ZN(n2236) );
  OR2_X1 U2879 ( .A1(n2793), .A2(IR_REG_25__SCAN_IN), .ZN(n2237) );
  AND2_X1 U2880 ( .A1(n2326), .A2(n4960), .ZN(n2484) );
  OR2_X1 U2881 ( .A1(n4334), .A2(n4483), .ZN(n2238) );
  AND3_X1 U2882 ( .A1(n2496), .A2(n2495), .A3(n2494), .ZN(n2239) );
  NOR2_X1 U2883 ( .A1(n4292), .A2(n4056), .ZN(n2240) );
  OR2_X1 U2884 ( .A1(n3293), .A2(n2405), .ZN(n2241) );
  OR2_X1 U2885 ( .A1(n3901), .A2(n3026), .ZN(n2242) );
  NAND2_X1 U2886 ( .A1(n4289), .A2(n4094), .ZN(n2243) );
  OR2_X1 U2887 ( .A1(n2740), .A2(IR_REG_21__SCAN_IN), .ZN(n2244) );
  OAI21_X1 U2888 ( .B1(n3660), .B2(n3661), .A(n3662), .ZN(n4475) );
  AND2_X1 U2890 ( .A1(n3158), .A2(n3157), .ZN(n2245) );
  NAND2_X1 U2891 ( .A1(n2381), .A2(n2380), .ZN(n2740) );
  AND2_X1 U2892 ( .A1(n2733), .A2(n2313), .ZN(n2246) );
  AND3_X1 U2893 ( .A1(n2473), .A2(n2472), .A3(n2471), .ZN(n3184) );
  INV_X1 U2894 ( .A(n2698), .ZN(n2338) );
  AND2_X1 U2895 ( .A1(n3353), .A2(n3352), .ZN(n2247) );
  NOR2_X1 U2896 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2482)
         );
  INV_X1 U2897 ( .A(n2370), .ZN(n2369) );
  AND2_X1 U2898 ( .A1(n4292), .A2(n4056), .ZN(n2248) );
  INV_X1 U2899 ( .A(IR_REG_28__SCAN_IN), .ZN(n2744) );
  AND2_X1 U2900 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2249)
         );
  NAND2_X1 U2901 ( .A1(n3895), .A2(n3358), .ZN(n2250) );
  NAND2_X1 U2902 ( .A1(n2699), .A2(n2243), .ZN(n2251) );
  INV_X1 U2903 ( .A(IR_REG_26__SCAN_IN), .ZN(n5042) );
  OR2_X1 U2904 ( .A1(n3899), .A2(n3166), .ZN(n2252) );
  AND2_X1 U2905 ( .A1(n2337), .A2(n2243), .ZN(n2253) );
  AND2_X1 U2906 ( .A1(n3861), .A2(n3863), .ZN(n2254) );
  NOR2_X1 U2907 ( .A1(n4596), .A2(n3982), .ZN(n2255) );
  INV_X1 U2908 ( .A(n3964), .ZN(n2314) );
  INV_X1 U2909 ( .A(n3166), .ZN(n2289) );
  INV_X1 U2910 ( .A(n4151), .ZN(n4472) );
  INV_X1 U2911 ( .A(n3274), .ZN(n2376) );
  AOI21_X1 U2912 ( .B1(n3504), .B2(n3505), .A(n3503), .ZN(n3660) );
  INV_X1 U2913 ( .A(IR_REG_21__SCAN_IN), .ZN(n2313) );
  INV_X1 U2914 ( .A(n3803), .ZN(n2303) );
  OR2_X1 U2915 ( .A1(n4651), .A2(n4697), .ZN(n2256) );
  OR2_X1 U2916 ( .A1(n4274), .A2(n3472), .ZN(n2257) );
  INV_X1 U2917 ( .A(n3600), .ZN(n3484) );
  NAND2_X1 U2918 ( .A1(n4368), .A2(n3694), .ZN(n2258) );
  OR2_X1 U2919 ( .A1(n3961), .A2(n3938), .ZN(n2259) );
  AND2_X1 U2920 ( .A1(n2843), .A2(n2301), .ZN(n2260) );
  INV_X1 U2921 ( .A(n3672), .ZN(n2431) );
  OR2_X1 U2922 ( .A1(n4271), .A2(n3713), .ZN(n2261) );
  AND2_X1 U2923 ( .A1(n4271), .A2(n4042), .ZN(n3827) );
  INV_X1 U2924 ( .A(n3827), .ZN(n2293) );
  MUX2_X1 U2925 ( .A(n4541), .B(DATAI_12_), .S(n2513), .Z(n4365) );
  NAND2_X1 U2926 ( .A1(n2318), .A2(n2316), .ZN(n2887) );
  INV_X1 U2927 ( .A(n4220), .ZN(n4482) );
  AND4_X1 U2928 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n4220)
         );
  INV_X1 U2929 ( .A(n2306), .ZN(n2305) );
  NAND2_X1 U2930 ( .A1(n2307), .A2(n3805), .ZN(n2306) );
  NAND2_X1 U2931 ( .A1(n2535), .A2(n2378), .ZN(n2377) );
  NAND2_X1 U2932 ( .A1(n3774), .A2(n3771), .ZN(n2754) );
  NAND2_X1 U2933 ( .A1(n3391), .A2(n2232), .ZN(n2262) );
  NAND2_X1 U2934 ( .A1(n2578), .A2(n2577), .ZN(n3409) );
  NAND2_X1 U2935 ( .A1(n3005), .A2(n3004), .ZN(n3103) );
  NAND2_X1 U2936 ( .A1(n3380), .A2(n3733), .ZN(n3379) );
  NAND2_X1 U2937 ( .A1(n3652), .A2(n3651), .ZN(n3650) );
  NOR2_X1 U2938 ( .A1(n3150), .A2(n3149), .ZN(n2263) );
  NAND2_X1 U2939 ( .A1(n2365), .A2(n2754), .ZN(n3173) );
  INV_X1 U2940 ( .A(n2287), .ZN(n4231) );
  NOR2_X1 U2941 ( .A1(n4229), .A2(n4228), .ZN(n2287) );
  INV_X1 U2942 ( .A(n2381), .ZN(n2617) );
  INV_X1 U2943 ( .A(n4211), .ZN(n4333) );
  AND2_X2 U2944 ( .A1(n2828), .A2(n2919), .ZN(n4699) );
  INV_X1 U2945 ( .A(n4699), .ZN(n4696) );
  NAND2_X1 U2946 ( .A1(n3173), .A2(n2485), .ZN(n3022) );
  INV_X1 U2947 ( .A(n4003), .ZN(n3839) );
  NAND2_X1 U2948 ( .A1(n2513), .A2(DATAI_24_), .ZN(n4074) );
  INV_X1 U2949 ( .A(n4056), .ZN(n3642) );
  NAND2_X1 U2950 ( .A1(n2513), .A2(DATAI_25_), .ZN(n4056) );
  INV_X1 U2951 ( .A(IR_REG_15__SCAN_IN), .ZN(n2626) );
  INV_X1 U2952 ( .A(n4541), .ZN(n2320) );
  INV_X1 U2953 ( .A(n4520), .ZN(n2319) );
  INV_X1 U2954 ( .A(IR_REG_17__SCAN_IN), .ZN(n2410) );
  INV_X1 U2955 ( .A(DATAI_1_), .ZN(n2359) );
  INV_X1 U2956 ( .A(IR_REG_2__SCAN_IN), .ZN(n2391) );
  OR2_X1 U2957 ( .A1(n3981), .A2(REG2_REG_17__SCAN_IN), .ZN(n2264) );
  NOR2_X1 U2958 ( .A1(n4643), .A2(n3983), .ZN(n2265) );
  INV_X1 U2959 ( .A(U4043), .ZN(n3903) );
  OAI21_X2 U2960 ( .B1(n2406), .B2(n2274), .A(n2272), .ZN(n2407) );
  INV_X2 U2961 ( .A(n3099), .ZN(n3562) );
  MUX2_X1 U2962 ( .A(n4960), .B(n2279), .S(n2513), .Z(n3086) );
  NAND3_X1 U2963 ( .A1(n2381), .A2(n2380), .A3(n2283), .ZN(n2793) );
  NAND3_X1 U2964 ( .A1(n2381), .A2(n2380), .A3(n2284), .ZN(n2286) );
  NAND3_X1 U2965 ( .A1(n3076), .A2(n2290), .A3(n2288), .ZN(n3206) );
  NAND2_X1 U2966 ( .A1(n2291), .A2(n3085), .ZN(n3768) );
  NAND2_X1 U2967 ( .A1(n2291), .A2(n3562), .ZN(n2433) );
  AOI21_X1 U2968 ( .B1(n4065), .B2(n2254), .A(n2292), .ZN(n4016) );
  OAI21_X1 U2969 ( .B1(n3245), .B2(n2306), .A(n2302), .ZN(n3419) );
  OAI21_X1 U2970 ( .B1(n3245), .B2(n3802), .A(n3787), .ZN(n3395) );
  NAND2_X1 U2971 ( .A1(n3802), .A2(n3787), .ZN(n2307) );
  OAI21_X1 U2972 ( .B1(n2752), .B2(n3767), .A(n2753), .ZN(n3181) );
  INV_X1 U2973 ( .A(n2740), .ZN(n2310) );
  NOR2_X1 U2974 ( .A1(n2740), .A2(n2312), .ZN(n2743) );
  NAND2_X1 U2975 ( .A1(n2310), .A2(n2311), .ZN(n2460) );
  MUX2_X1 U2976 ( .A(n2888), .B(REG2_REG_1__SCAN_IN), .S(n2887), .Z(n3908) );
  NAND2_X1 U2977 ( .A1(n2775), .A2(n3812), .ZN(n4199) );
  NAND2_X1 U2978 ( .A1(n3850), .A2(n3381), .ZN(n3447) );
  OAI22_X1 U2979 ( .A1(n4551), .A2(n4554), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3958), .ZN(n3947) );
  XNOR2_X1 U2980 ( .A(n4648), .B(n3947), .ZN(n4564) );
  NOR2_X1 U2981 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2326)
         );
  INV_X1 U2982 ( .A(n4081), .ZN(n2329) );
  NAND2_X1 U2983 ( .A1(n2353), .A2(n2354), .ZN(n4141) );
  NAND2_X1 U2984 ( .A1(n4183), .A2(n2355), .ZN(n2353) );
  MUX2_X1 U2985 ( .A(n2887), .B(n2359), .S(n2513), .Z(n3085) );
  NOR2_X1 U2986 ( .A1(n3072), .A2(n3194), .ZN(n2361) );
  INV_X1 U2987 ( .A(n3174), .ZN(n2365) );
  NAND2_X1 U2988 ( .A1(n2383), .A2(n2384), .ZN(n3986) );
  NAND2_X1 U2989 ( .A1(n4595), .A2(n2385), .ZN(n2383) );
  NOR2_X1 U2990 ( .A1(n4595), .A2(n4594), .ZN(n4596) );
  MUX2_X1 U2991 ( .A(REG1_REG_2__SCAN_IN), .B(n4690), .S(n4455), .Z(n3921) );
  OAI21_X2 U2992 ( .B1(n2399), .B2(n2396), .A(n2394), .ZN(n3231) );
  NAND2_X1 U2993 ( .A1(n3710), .A2(n3708), .ZN(n2402) );
  OAI211_X1 U2994 ( .C1(n2404), .C2(n3587), .A(n3586), .B(n2403), .ZN(U3217)
         );
  NAND2_X1 U2995 ( .A1(n2404), .A2(n3577), .ZN(n2403) );
  NAND2_X1 U2996 ( .A1(n3693), .A2(n2414), .ZN(n2411) );
  NAND2_X1 U2997 ( .A1(n2411), .A2(n2412), .ZN(n3492) );
  INV_X1 U2998 ( .A(n3691), .ZN(n2420) );
  INV_X1 U2999 ( .A(n3690), .ZN(n2421) );
  NAND2_X1 U3000 ( .A1(n3700), .A2(n3701), .ZN(n3607) );
  NAND2_X1 U3001 ( .A1(n2462), .A2(REG2_REG_1__SCAN_IN), .ZN(n2473) );
  OR2_X1 U3002 ( .A1(n3757), .A2(n2886), .ZN(n2481) );
  OR2_X1 U3003 ( .A1(n3757), .A2(n3051), .ZN(n2927) );
  NAND2_X1 U3004 ( .A1(n2469), .A2(n2466), .ZN(n2476) );
  INV_X1 U3005 ( .A(n2469), .ZN(n2465) );
  INV_X1 U3006 ( .A(n3679), .ZN(n4479) );
  AND2_X1 U3007 ( .A1(n4169), .A2(n4143), .ZN(n2439) );
  NAND2_X1 U3008 ( .A1(n3496), .A2(n3596), .ZN(n2440) );
  AND2_X1 U3009 ( .A1(n3628), .A2(n3627), .ZN(n2441) );
  AND2_X1 U3010 ( .A1(n4318), .A2(n4133), .ZN(n2442) );
  OR2_X1 U3011 ( .A1(n4135), .A2(n4116), .ZN(n2443) );
  OR2_X1 U3012 ( .A1(n4430), .A2(n4429), .ZN(U3499) );
  OR2_X1 U3013 ( .A1(n3466), .A2(n4443), .ZN(n2445) );
  OR2_X1 U3014 ( .A1(n3466), .A2(n4377), .ZN(n2446) );
  INV_X1 U3015 ( .A(IR_REG_14__SCAN_IN), .ZN(n2451) );
  NAND2_X1 U3016 ( .A1(n3557), .A2(n3088), .ZN(n2967) );
  INV_X1 U3017 ( .A(n3516), .ZN(n3517) );
  AND2_X1 U3018 ( .A1(n3753), .A2(n4031), .ZN(n3861) );
  AND2_X1 U3019 ( .A1(n4164), .A2(n2776), .ZN(n4084) );
  NOR2_X1 U3020 ( .A1(n3721), .A2(n4466), .ZN(n3504) );
  INV_X1 U3021 ( .A(n2984), .ZN(n3009) );
  OAI21_X1 U3022 ( .B1(n3426), .B2(n3425), .A(n3424), .ZN(n3428) );
  INV_X1 U3023 ( .A(REG3_REG_12__SCAN_IN), .ZN(n5047) );
  INV_X1 U3024 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2907) );
  INV_X1 U3025 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2549) );
  OR2_X1 U3026 ( .A1(n3499), .A2(n3498), .ZN(n3502) );
  AND2_X1 U3027 ( .A1(n3434), .A2(n3435), .ZN(n3477) );
  INV_X1 U3028 ( .A(n3529), .ZN(n3530) );
  OR2_X1 U3029 ( .A1(n2707), .A2(n2705), .ZN(n2715) );
  OR2_X1 U3030 ( .A1(n2692), .A2(n4940), .ZN(n2707) );
  INV_X1 U3031 ( .A(n3891), .ZN(n4035) );
  AND2_X1 U3032 ( .A1(n4037), .A2(n4056), .ZN(n3766) );
  AND2_X1 U3033 ( .A1(n4152), .A2(n2779), .ZN(n4087) );
  NOR2_X1 U3034 ( .A1(n4220), .A2(n4211), .ZN(n2643) );
  NOR2_X1 U3035 ( .A1(n2601), .A2(n4957), .ZN(n2610) );
  OR2_X1 U3036 ( .A1(n2591), .A2(n2590), .ZN(n2601) );
  NOR2_X1 U3037 ( .A1(n2550), .A2(n2549), .ZN(n2560) );
  NAND2_X1 U3038 ( .A1(n2525), .A2(REG3_REG_7__SCAN_IN), .ZN(n2536) );
  INV_X1 U3039 ( .A(n3372), .ZN(n3370) );
  INV_X1 U3040 ( .A(n2754), .ZN(n3180) );
  OR3_X1 U3041 ( .A1(n2556), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2567) );
  AND2_X1 U3042 ( .A1(n2560), .A2(REG3_REG_10__SCAN_IN), .ZN(n2570) );
  NOR2_X1 U3043 ( .A1(n3575), .A2(n3679), .ZN(n3576) );
  NOR2_X1 U3044 ( .A1(n2633), .A2(n2632), .ZN(n2645) );
  NOR2_X1 U3045 ( .A1(n2715), .A2(n4941), .ZN(n2724) );
  INV_X1 U3046 ( .A(REG3_REG_16__SCAN_IN), .ZN(n5041) );
  AND2_X1 U3047 ( .A1(n4005), .A2(n3472), .ZN(n3825) );
  AND2_X1 U3048 ( .A1(n2787), .A2(n2788), .ZN(n4015) );
  INV_X1 U3049 ( .A(n4037), .ZN(n4292) );
  OR2_X1 U3050 ( .A1(n2536), .A2(n4847), .ZN(n2550) );
  INV_X1 U3051 ( .A(n3026), .ZN(n3194) );
  AND2_X1 U3052 ( .A1(n2868), .A2(n2864), .ZN(n2821) );
  INV_X1 U3053 ( .A(n4074), .ZN(n4288) );
  MUX2_X1 U3054 ( .A(n3956), .B(DATAI_15_), .S(n2513), .Z(n4347) );
  INV_X1 U3055 ( .A(n4222), .ZN(n4242) );
  AND2_X1 U3056 ( .A1(n2683), .A2(REG3_REG_22__SCAN_IN), .ZN(n2687) );
  OR2_X1 U3057 ( .A1(n2716), .A2(n2724), .ZN(n4021) );
  AND4_X1 U3058 ( .A1(n2658), .A2(n2657), .A3(n2656), .A4(n2655), .ZN(n4151)
         );
  AND2_X1 U3059 ( .A1(n2882), .A2(n2881), .ZN(n4496) );
  AND2_X1 U3060 ( .A1(n4496), .A2(n3053), .ZN(n4606) );
  INV_X1 U3061 ( .A(n4317), .ZN(n4367) );
  NAND2_X1 U3062 ( .A1(n2790), .A2(n2789), .ZN(n4222) );
  INV_X1 U3063 ( .A(n4449), .ZN(n3989) );
  AND2_X1 U3064 ( .A1(n4256), .A2(n3047), .ZN(n4624) );
  AOI21_X1 U3065 ( .B1(n2823), .B2(n2822), .A(n2821), .ZN(n2919) );
  NAND2_X1 U3066 ( .A1(n2513), .A2(DATAI_22_), .ZN(n4116) );
  INV_X1 U3067 ( .A(n3694), .ZN(n4250) );
  INV_X1 U3068 ( .A(n3358), .ZN(n3396) );
  AND2_X1 U3069 ( .A1(n3034), .A2(n2943), .ZN(n4684) );
  INV_X1 U3070 ( .A(n3040), .ZN(n2949) );
  NAND2_X1 U3071 ( .A1(n2924), .A2(n2923), .ZN(n3679) );
  INV_X1 U3072 ( .A(n4274), .ZN(n4005) );
  NAND2_X1 U3073 ( .A1(n4496), .A2(n4457), .ZN(n4610) );
  INV_X1 U3074 ( .A(n4552), .ZN(n4600) );
  INV_X1 U3075 ( .A(n4256), .ZN(n4629) );
  INV_X1 U3076 ( .A(n4256), .ZN(n4489) );
  NAND2_X1 U3077 ( .A1(n4699), .A2(n4664), .ZN(n4377) );
  OR2_X1 U3078 ( .A1(n4008), .A2(n4443), .ZN(n2849) );
  NAND2_X1 U3079 ( .A1(n4687), .A2(n4664), .ZN(n4443) );
  INV_X1 U3080 ( .A(n4687), .ZN(n4685) );
  XNOR2_X1 U3081 ( .A(n2745), .B(n2744), .ZN(n4457) );
  NAND4_X1 U3082 ( .A1(n2450), .A2(n2449), .A3(n2448), .A4(n2447), .ZN(n2597)
         );
  NAND3_X1 U3083 ( .A1(n2451), .A2(n2510), .A3(n4793), .ZN(n2452) );
  NOR2_X1 U3084 ( .A1(n2597), .A2(n2452), .ZN(n2453) );
  INV_X1 U3085 ( .A(IR_REG_27__SCAN_IN), .ZN(n2457) );
  NOR2_X1 U3086 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2458)
         );
  NAND2_X1 U3087 ( .A1(n2743), .A2(n2458), .ZN(n2856) );
  NAND2_X4 U3088 ( .A1(n4445), .A2(n2465), .ZN(n3757) );
  INV_X1 U3089 ( .A(n3757), .ZN(n2462) );
  INV_X1 U3090 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2464) );
  OR2_X1 U3091 ( .A1(n2476), .A2(n2464), .ZN(n2468) );
  AND2_X2 U3092 ( .A1(n2466), .A2(n2465), .ZN(n2516) );
  NAND2_X1 U3093 ( .A1(n2516), .A2(REG0_REG_1__SCAN_IN), .ZN(n2467) );
  NAND2_X4 U3094 ( .A1(n2469), .A2(n4445), .ZN(n2486) );
  INV_X1 U3095 ( .A(n2486), .ZN(n2470) );
  NAND2_X1 U3096 ( .A1(n2470), .A2(REG3_REG_1__SCAN_IN), .ZN(n2471) );
  INV_X1 U3097 ( .A(n2887), .ZN(n4456) );
  NAND2_X1 U3098 ( .A1(n2838), .A2(n2744), .ZN(n2474) );
  NAND2_X1 U3099 ( .A1(n3184), .A2(n3088), .ZN(n2753) );
  NAND2_X1 U3100 ( .A1(n2753), .A2(n3768), .ZN(n2752) );
  INV_X1 U3101 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2475) );
  INV_X1 U3102 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3103 ( .A1(n2717), .A2(REG1_REG_0__SCAN_IN), .ZN(n2926) );
  NAND2_X1 U3104 ( .A1(n2631), .A2(REG0_REG_0__SCAN_IN), .ZN(n2925) );
  NOR2_X1 U3105 ( .A1(n2978), .A2(n3086), .ZN(n3081) );
  NAND2_X1 U3106 ( .A1(n2752), .A2(n3081), .ZN(n3083) );
  NAND2_X1 U3107 ( .A1(n2291), .A2(n3088), .ZN(n2477) );
  NAND2_X1 U3108 ( .A1(n3083), .A2(n2477), .ZN(n3174) );
  INV_X1 U3109 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2886) );
  INV_X1 U3110 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3179) );
  OR2_X1 U3111 ( .A1(n2486), .A2(n3179), .ZN(n2480) );
  NAND2_X1 U3112 ( .A1(n2516), .A2(REG0_REG_2__SCAN_IN), .ZN(n2479) );
  NAND2_X1 U3113 ( .A1(n2717), .A2(REG1_REG_2__SCAN_IN), .ZN(n2478) );
  INV_X1 U3114 ( .A(n3199), .ZN(n3902) );
  NOR2_X1 U3115 ( .A1(n2482), .A2(n2796), .ZN(n2483) );
  MUX2_X1 U3116 ( .A(n4455), .B(DATAI_2_), .S(n2513), .Z(n3182) );
  INV_X1 U3117 ( .A(n3182), .ZN(n2995) );
  NAND2_X1 U3118 ( .A1(n3902), .A2(n2995), .ZN(n3774) );
  NAND2_X1 U3119 ( .A1(n3199), .A2(n3182), .ZN(n3771) );
  NAND2_X1 U3120 ( .A1(n3199), .A2(n2995), .ZN(n2485) );
  OR2_X1 U3121 ( .A1(n2486), .A2(REG3_REG_3__SCAN_IN), .ZN(n2490) );
  INV_X1 U3122 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3929) );
  OR2_X1 U3123 ( .A1(n3757), .A2(n3929), .ZN(n2489) );
  NAND2_X1 U3124 ( .A1(n2717), .A2(REG1_REG_3__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U3125 ( .A1(n2631), .A2(REG0_REG_3__SCAN_IN), .ZN(n2487) );
  OR2_X1 U3126 ( .A1(n2484), .A2(n2796), .ZN(n2499) );
  XNOR2_X1 U3127 ( .A(n2499), .B(IR_REG_3__SCAN_IN), .ZN(n4454) );
  MUX2_X1 U3128 ( .A(n4454), .B(DATAI_3_), .S(n2513), .Z(n3026) );
  INV_X1 U3129 ( .A(n3901), .ZN(n3072) );
  NAND2_X1 U3130 ( .A1(n2717), .A2(REG1_REG_4__SCAN_IN), .ZN(n2497) );
  INV_X1 U3131 ( .A(n2505), .ZN(n2493) );
  INV_X1 U3132 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3017) );
  INV_X1 U3133 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U3134 ( .A1(n3017), .A2(n2491), .ZN(n2492) );
  NAND2_X1 U3135 ( .A1(n2493), .A2(n2492), .ZN(n3113) );
  OR2_X1 U3136 ( .A1(n2486), .A2(n3113), .ZN(n2496) );
  INV_X1 U3137 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2895) );
  OR2_X1 U3138 ( .A1(n3757), .A2(n2895), .ZN(n2495) );
  NAND2_X1 U3139 ( .A1(n2631), .A2(REG0_REG_4__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U3140 ( .A1(n2499), .A2(n2498), .ZN(n2500) );
  NAND2_X1 U3141 ( .A1(n2500), .A2(IR_REG_31__SCAN_IN), .ZN(n2501) );
  XNOR2_X1 U3142 ( .A(n2501), .B(IR_REG_4__SCAN_IN), .ZN(n4453) );
  MUX2_X1 U3143 ( .A(n4453), .B(DATAI_4_), .S(n2513), .Z(n3110) );
  NAND2_X1 U3144 ( .A1(n3282), .A2(n3110), .ZN(n3777) );
  NAND2_X1 U3145 ( .A1(n2502), .A2(n3101), .ZN(n3780) );
  NAND2_X1 U3146 ( .A1(n3777), .A2(n3780), .ZN(n3739) );
  NAND2_X1 U3147 ( .A1(n3069), .A2(n3739), .ZN(n2504) );
  NAND2_X1 U31480 ( .A1(n2502), .A2(n3110), .ZN(n2503) );
  NAND2_X1 U31490 ( .A1(n2504), .A2(n2503), .ZN(n3116) );
  INV_X1 U3150 ( .A(n3116), .ZN(n2522) );
  OAI21_X1 U3151 ( .B1(n2505), .B2(REG3_REG_5__SCAN_IN), .A(n2514), .ZN(n3655)
         );
  OR2_X1 U3152 ( .A1(n2486), .A2(n3655), .ZN(n2509) );
  INV_X1 U3153 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2885) );
  OR2_X1 U3154 ( .A1(n3757), .A2(n2885), .ZN(n2508) );
  NAND2_X1 U3155 ( .A1(n2631), .A2(REG0_REG_5__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3156 ( .A1(n2717), .A2(REG1_REG_5__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3157 ( .A1(n2511), .A2(n2510), .ZN(n2598) );
  NAND2_X1 U3158 ( .A1(n2598), .A2(IR_REG_31__SCAN_IN), .ZN(n2512) );
  XNOR2_X1 U3159 ( .A(n2512), .B(IR_REG_5__SCAN_IN), .ZN(n4452) );
  MUX2_X1 U3160 ( .A(n4452), .B(DATAI_5_), .S(n2513), .Z(n3654) );
  AND2_X1 U3161 ( .A1(n3900), .A2(n3654), .ZN(n3127) );
  AND2_X1 U3162 ( .A1(n2514), .A2(n2907), .ZN(n2515) );
  OR2_X1 U3163 ( .A1(n2515), .A2(n2525), .ZN(n3169) );
  OR2_X1 U3164 ( .A1(n2486), .A2(n3169), .ZN(n2520) );
  INV_X1 U3165 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3138) );
  OR2_X1 U3166 ( .A1(n3757), .A2(n3138), .ZN(n2519) );
  NAND2_X1 U3167 ( .A1(n2631), .A2(REG0_REG_6__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U3168 ( .A1(n2717), .A2(REG1_REG_6__SCAN_IN), .ZN(n2517) );
  OR2_X1 U3169 ( .A1(n2532), .A2(n2796), .ZN(n2521) );
  XNOR2_X1 U3170 ( .A(n2521), .B(IR_REG_6__SCAN_IN), .ZN(n4451) );
  MUX2_X1 U3171 ( .A(n4451), .B(DATAI_6_), .S(n2513), .Z(n3166) );
  AND2_X1 U3172 ( .A1(n3899), .A2(n3166), .ZN(n2524) );
  NAND2_X1 U3173 ( .A1(n2522), .A2(n2228), .ZN(n3213) );
  INV_X1 U3174 ( .A(n3900), .ZN(n2758) );
  INV_X1 U3175 ( .A(n3654), .ZN(n3154) );
  NAND2_X1 U3176 ( .A1(n2758), .A2(n3154), .ZN(n3128) );
  AND2_X1 U3177 ( .A1(n3128), .A2(n2252), .ZN(n2523) );
  OR2_X1 U3178 ( .A1(n2524), .A2(n2523), .ZN(n3212) );
  NAND2_X1 U3179 ( .A1(n2631), .A2(REG0_REG_7__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U3180 ( .A1(n2717), .A2(REG1_REG_7__SCAN_IN), .ZN(n2529) );
  OR2_X1 U3181 ( .A1(n2525), .A2(REG3_REG_7__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U3182 ( .A1(n2536), .A2(n2526), .ZN(n3240) );
  OR2_X1 U3183 ( .A1(n2486), .A2(n3240), .ZN(n2528) );
  INV_X1 U3184 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3938) );
  OR2_X1 U3185 ( .A1(n3757), .A2(n3938), .ZN(n2527) );
  INV_X1 U3186 ( .A(IR_REG_6__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U3187 ( .A1(n2532), .A2(n2531), .ZN(n2556) );
  NAND2_X1 U3188 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2544) );
  XNOR2_X1 U3189 ( .A(n2544), .B(IR_REG_7__SCAN_IN), .ZN(n4450) );
  MUX2_X1 U3190 ( .A(n4450), .B(DATAI_7_), .S(n2513), .Z(n3237) );
  NAND2_X1 U3191 ( .A1(n3321), .A2(n3237), .ZN(n2759) );
  NAND2_X1 U3192 ( .A1(n3898), .A2(n3235), .ZN(n3786) );
  NAND2_X1 U3193 ( .A1(n2759), .A2(n3786), .ZN(n3745) );
  AND2_X1 U3194 ( .A1(n3212), .A2(n3745), .ZN(n2533) );
  NAND2_X1 U3195 ( .A1(n3213), .A2(n2533), .ZN(n2535) );
  NAND2_X1 U3196 ( .A1(n3898), .A2(n3237), .ZN(n2534) );
  NAND2_X1 U3197 ( .A1(n2536), .A2(n4847), .ZN(n2537) );
  AND2_X1 U3198 ( .A1(n2550), .A2(n2537), .ZN(n4620) );
  INV_X1 U3199 ( .A(n4620), .ZN(n3277) );
  OR2_X1 U3200 ( .A1(n2486), .A2(n3277), .ZN(n2542) );
  INV_X1 U3201 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2538) );
  OR2_X1 U3202 ( .A1(n3757), .A2(n2538), .ZN(n2541) );
  NAND2_X1 U3203 ( .A1(n2717), .A2(REG1_REG_8__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U3204 ( .A1(n2631), .A2(REG0_REG_8__SCAN_IN), .ZN(n2539) );
  NAND4_X1 U3205 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(n3897)
         );
  INV_X1 U3206 ( .A(IR_REG_7__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U3207 ( .A1(n2544), .A2(n2543), .ZN(n2545) );
  NAND2_X1 U3208 ( .A1(n2545), .A2(IR_REG_31__SCAN_IN), .ZN(n2546) );
  XNOR2_X1 U3209 ( .A(n2546), .B(IR_REG_8__SCAN_IN), .ZN(n3964) );
  MUX2_X1 U32100 ( .A(n3964), .B(DATAI_8_), .S(n2513), .Z(n3274) );
  AND2_X1 U32110 ( .A1(n3897), .A2(n3274), .ZN(n2547) );
  INV_X1 U32120 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2548) );
  OR2_X1 U32130 ( .A1(n3757), .A2(n2548), .ZN(n2555) );
  AND2_X1 U32140 ( .A1(n2550), .A2(n2549), .ZN(n2551) );
  OR2_X1 U32150 ( .A1(n2551), .A2(n2560), .ZN(n3302) );
  OR2_X1 U32160 ( .A1(n2486), .A2(n3302), .ZN(n2554) );
  NAND2_X1 U32170 ( .A1(n2717), .A2(REG1_REG_9__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32180 ( .A1(n2631), .A2(REG0_REG_9__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32190 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2557) );
  XNOR2_X1 U32200 ( .A(n2557), .B(IR_REG_9__SCAN_IN), .ZN(n3960) );
  NOR2_X1 U32210 ( .A1(n3896), .A2(n3306), .ZN(n2559) );
  NAND2_X1 U32220 ( .A1(n3896), .A2(n3306), .ZN(n2558) );
  NOR2_X1 U32230 ( .A1(n2560), .A2(REG3_REG_10__SCAN_IN), .ZN(n2561) );
  OR2_X1 U32240 ( .A1(n2570), .A2(n2561), .ZN(n4611) );
  OR2_X1 U32250 ( .A1(n2486), .A2(n4611), .ZN(n2566) );
  INV_X1 U32260 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2562) );
  OR2_X1 U32270 ( .A1(n3757), .A2(n2562), .ZN(n2565) );
  NAND2_X1 U32280 ( .A1(n2717), .A2(REG1_REG_10__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U32290 ( .A1(n2631), .A2(REG0_REG_10__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32300 ( .A1(n2576), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  XNOR2_X1 U32310 ( .A(n2568), .B(IR_REG_10__SCAN_IN), .ZN(n4520) );
  MUX2_X1 U32320 ( .A(n4520), .B(DATAI_10_), .S(n2513), .Z(n3358) );
  INV_X1 U32330 ( .A(n3895), .ZN(n2762) );
  NAND2_X1 U32340 ( .A1(n2762), .A2(n3396), .ZN(n2569) );
  NAND2_X1 U32350 ( .A1(n2631), .A2(REG0_REG_11__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U32360 ( .A1(n2717), .A2(REG1_REG_11__SCAN_IN), .ZN(n2574) );
  OR2_X1 U32370 ( .A1(n2570), .A2(REG3_REG_11__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U32380 ( .A1(n2579), .A2(n2571), .ZN(n3375) );
  OR2_X1 U32390 ( .A1(n2486), .A2(n3375), .ZN(n2573) );
  INV_X1 U32400 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3338) );
  OR2_X1 U32410 ( .A1(n3757), .A2(n3338), .ZN(n2572) );
  OAI21_X1 U32420 ( .B1(n2576), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2586) );
  XNOR2_X1 U32430 ( .A(n2586), .B(IR_REG_11__SCAN_IN), .ZN(n3959) );
  MUX2_X1 U32440 ( .A(n3959), .B(DATAI_11_), .S(n2513), .Z(n3372) );
  NAND2_X1 U32450 ( .A1(n4372), .A2(n3372), .ZN(n3416) );
  NAND2_X1 U32460 ( .A1(n3894), .A2(n3370), .ZN(n3418) );
  NAND2_X1 U32470 ( .A1(n3416), .A2(n3418), .ZN(n3746) );
  NAND2_X1 U32480 ( .A1(n3332), .A2(n3746), .ZN(n2578) );
  NAND2_X1 U32490 ( .A1(n4372), .A2(n3370), .ZN(n2577) );
  NAND2_X1 U32500 ( .A1(n2579), .A2(n5047), .ZN(n2580) );
  NAND2_X1 U32510 ( .A1(n2591), .A2(n2580), .ZN(n3443) );
  OR2_X1 U32520 ( .A1(n2486), .A2(n3443), .ZN(n2584) );
  INV_X1 U32530 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3412) );
  OR2_X1 U32540 ( .A1(n3757), .A2(n3412), .ZN(n2583) );
  NAND2_X1 U32550 ( .A1(n2631), .A2(REG0_REG_12__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U32560 ( .A1(n2717), .A2(REG1_REG_12__SCAN_IN), .ZN(n2581) );
  INV_X1 U32570 ( .A(IR_REG_11__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U32580 ( .A1(n2586), .A2(n2585), .ZN(n2587) );
  NAND2_X1 U32590 ( .A1(n2587), .A2(IR_REG_31__SCAN_IN), .ZN(n2588) );
  XNOR2_X1 U32600 ( .A(n2588), .B(IR_REG_12__SCAN_IN), .ZN(n4541) );
  NOR2_X1 U32610 ( .A1(n4246), .A2(n4365), .ZN(n2589) );
  INV_X1 U32620 ( .A(n4365), .ZN(n2763) );
  INV_X1 U32630 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U32640 ( .A1(n2591), .A2(n2590), .ZN(n2592) );
  NAND2_X1 U32650 ( .A1(n2601), .A2(n2592), .ZN(n4254) );
  OR2_X1 U32660 ( .A1(n2486), .A2(n4254), .ZN(n2596) );
  INV_X1 U32670 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4255) );
  OR2_X1 U32680 ( .A1(n3757), .A2(n4255), .ZN(n2595) );
  NAND2_X1 U32690 ( .A1(n2631), .A2(REG0_REG_13__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U32700 ( .A1(n2717), .A2(REG1_REG_13__SCAN_IN), .ZN(n2593) );
  OR2_X1 U32710 ( .A1(n2598), .A2(n2597), .ZN(n2607) );
  NAND2_X1 U32720 ( .A1(n2607), .A2(IR_REG_31__SCAN_IN), .ZN(n2599) );
  XNOR2_X1 U32730 ( .A(n2599), .B(IR_REG_13__SCAN_IN), .ZN(n3958) );
  MUX2_X1 U32740 ( .A(n3958), .B(DATAI_13_), .S(n2513), .Z(n3694) );
  INV_X1 U32750 ( .A(n4368), .ZN(n3385) );
  NAND2_X1 U32760 ( .A1(n3385), .A2(n4250), .ZN(n2600) );
  NAND2_X1 U32770 ( .A1(n2631), .A2(REG0_REG_14__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U32780 ( .A1(n2717), .A2(REG1_REG_14__SCAN_IN), .ZN(n2605) );
  AND2_X1 U32790 ( .A1(n2601), .A2(n4957), .ZN(n2602) );
  OR2_X1 U32800 ( .A1(n2602), .A2(n2610), .ZN(n3603) );
  OR2_X1 U32810 ( .A1(n2486), .A2(n3603), .ZN(n2604) );
  INV_X1 U32820 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3387) );
  OR2_X1 U32830 ( .A1(n3757), .A2(n3387), .ZN(n2603) );
  OAI21_X1 U32840 ( .B1(n2607), .B2(IR_REG_13__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2608) );
  XNOR2_X1 U32850 ( .A(n2608), .B(IR_REG_14__SCAN_IN), .ZN(n3973) );
  MUX2_X1 U32860 ( .A(n3973), .B(DATAI_14_), .S(n2513), .Z(n3600) );
  NAND2_X1 U32870 ( .A1(n4351), .A2(n3600), .ZN(n3810) );
  INV_X1 U32880 ( .A(n4351), .ZN(n3893) );
  NAND2_X1 U32890 ( .A1(n3893), .A2(n3484), .ZN(n3791) );
  NAND2_X1 U32900 ( .A1(n3810), .A2(n3791), .ZN(n3733) );
  NAND2_X1 U32910 ( .A1(n4351), .A2(n3484), .ZN(n2609) );
  NAND2_X1 U32920 ( .A1(n3379), .A2(n2609), .ZN(n3451) );
  OR2_X1 U32930 ( .A1(n2610), .A2(REG3_REG_15__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U32940 ( .A1(n2620), .A2(n2611), .ZN(n3726) );
  OR2_X1 U32950 ( .A1(n2486), .A2(n3726), .ZN(n2616) );
  INV_X1 U32960 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2612) );
  OR2_X1 U32970 ( .A1(n3757), .A2(n2612), .ZN(n2615) );
  NAND2_X1 U32980 ( .A1(n2631), .A2(REG0_REG_15__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U32990 ( .A1(n2717), .A2(REG1_REG_15__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U33000 ( .A1(n2617), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  XNOR2_X1 U33010 ( .A(n2627), .B(IR_REG_15__SCAN_IN), .ZN(n3956) );
  NOR2_X1 U33020 ( .A1(n4217), .A2(n4347), .ZN(n2619) );
  NAND2_X1 U33030 ( .A1(n4217), .A2(n4347), .ZN(n2618) );
  NAND2_X1 U33040 ( .A1(n2717), .A2(REG1_REG_16__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U33050 ( .A1(n2631), .A2(REG0_REG_16__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U33060 ( .A1(n2620), .A2(n5041), .ZN(n2621) );
  NAND2_X1 U33070 ( .A1(n2633), .A2(n2621), .ZN(n4470) );
  OR2_X1 U33080 ( .A1(n2486), .A2(n4470), .ZN(n2623) );
  INV_X1 U33090 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4232) );
  OR2_X1 U33100 ( .A1(n3757), .A2(n4232), .ZN(n2622) );
  NAND2_X1 U33110 ( .A1(n2627), .A2(n2626), .ZN(n2628) );
  NAND2_X1 U33120 ( .A1(n2628), .A2(IR_REG_31__SCAN_IN), .ZN(n2629) );
  XNOR2_X1 U33130 ( .A(n2629), .B(IR_REG_16__SCAN_IN), .ZN(n3977) );
  MUX2_X1 U33140 ( .A(n3977), .B(DATAI_16_), .S(n2513), .Z(n4228) );
  NAND2_X1 U33150 ( .A1(n4337), .A2(n4228), .ZN(n3852) );
  NAND2_X1 U33160 ( .A1(n4348), .A2(n4460), .ZN(n3812) );
  NAND2_X1 U33170 ( .A1(n3852), .A2(n3812), .ZN(n4225) );
  NAND2_X1 U33180 ( .A1(n4226), .A2(n4225), .ZN(n4224) );
  NAND2_X1 U33190 ( .A1(n4224), .A2(n2630), .ZN(n4202) );
  NAND2_X1 U33200 ( .A1(n2717), .A2(REG1_REG_17__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U33210 ( .A1(n2631), .A2(REG0_REG_17__SCAN_IN), .ZN(n2638) );
  INV_X1 U33220 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2632) );
  AND2_X1 U33230 ( .A1(n2633), .A2(n2632), .ZN(n2634) );
  OR2_X1 U33240 ( .A1(n2634), .A2(n2645), .ZN(n4206) );
  OR2_X1 U33250 ( .A1(n2486), .A2(n4206), .ZN(n2637) );
  INV_X1 U33260 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2635) );
  OR2_X1 U33270 ( .A1(n3757), .A2(n2635), .ZN(n2636) );
  NAND2_X1 U33280 ( .A1(n2640), .A2(IR_REG_31__SCAN_IN), .ZN(n2641) );
  XNOR2_X1 U33290 ( .A(n2641), .B(IR_REG_17__SCAN_IN), .ZN(n3981) );
  INV_X1 U33300 ( .A(n3981), .ZN(n4644) );
  INV_X1 U33310 ( .A(DATAI_17_), .ZN(n2642) );
  MUX2_X1 U33320 ( .A(n4644), .B(n2642), .S(n2513), .Z(n4211) );
  NAND2_X1 U33330 ( .A1(n4220), .A2(n4211), .ZN(n2644) );
  AOI21_X1 U33340 ( .B1(n4202), .B2(n2644), .A(n2643), .ZN(n4183) );
  NAND2_X1 U33350 ( .A1(n2631), .A2(REG0_REG_18__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U33360 ( .A1(n2717), .A2(REG1_REG_18__SCAN_IN), .ZN(n2649) );
  NOR2_X1 U33370 ( .A1(n2645), .A2(REG3_REG_18__SCAN_IN), .ZN(n2646) );
  OR2_X1 U33380 ( .A1(n2653), .A2(n2646), .ZN(n4487) );
  OR2_X1 U33390 ( .A1(n2486), .A2(n4487), .ZN(n2648) );
  INV_X1 U33400 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4194) );
  OR2_X1 U33410 ( .A1(n3757), .A2(n4194), .ZN(n2647) );
  OR2_X1 U33420 ( .A1(n2651), .A2(n2796), .ZN(n2652) );
  XNOR2_X1 U33430 ( .A(n2652), .B(IR_REG_18__SCAN_IN), .ZN(n3954) );
  MUX2_X1 U33440 ( .A(n3954), .B(DATAI_18_), .S(n2513), .Z(n4483) );
  INV_X1 U33450 ( .A(n4483), .ZN(n4187) );
  NAND2_X1 U33460 ( .A1(n4334), .A2(n4187), .ZN(n4164) );
  NAND2_X1 U33470 ( .A1(n4172), .A2(n4483), .ZN(n4163) );
  NAND2_X1 U33480 ( .A1(n4164), .A2(n4163), .ZN(n4190) );
  NAND2_X1 U33490 ( .A1(n2631), .A2(REG0_REG_19__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U33500 ( .A1(n2717), .A2(REG1_REG_19__SCAN_IN), .ZN(n2657) );
  OR2_X1 U33510 ( .A1(n2653), .A2(REG3_REG_19__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U33520 ( .A1(n2663), .A2(n2654), .ZN(n4176) );
  OR2_X1 U3353 ( .A1(n2486), .A2(n4176), .ZN(n2656) );
  INV_X1 U33540 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4177) );
  OR2_X1 U3355 ( .A1(n3757), .A2(n4177), .ZN(n2655) );
  NAND2_X1 U3356 ( .A1(n2659), .A2(IR_REG_31__SCAN_IN), .ZN(n2736) );
  INV_X1 U3357 ( .A(DATAI_19_), .ZN(n2660) );
  MUX2_X1 U3358 ( .A(n3989), .B(n2660), .S(n2513), .Z(n4173) );
  INV_X1 U3359 ( .A(n4173), .ZN(n2661) );
  INV_X1 U3360 ( .A(n4141), .ZN(n2671) );
  INV_X1 U3361 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U3362 ( .A1(n2663), .A2(n4822), .ZN(n2664) );
  NAND2_X1 U3363 ( .A1(n2673), .A2(n2664), .ZN(n4146) );
  OR2_X1 U3364 ( .A1(n2486), .A2(n4146), .ZN(n2669) );
  INV_X1 U3365 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2665) );
  OR2_X1 U3366 ( .A1(n3757), .A2(n2665), .ZN(n2668) );
  NAND2_X1 U3367 ( .A1(n2631), .A2(REG0_REG_20__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3368 ( .A1(n2717), .A2(REG1_REG_20__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3369 ( .A1(n2513), .A2(DATAI_20_), .ZN(n4316) );
  NOR2_X1 U3370 ( .A1(n4169), .A2(n4143), .ZN(n3754) );
  INV_X1 U3371 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2672) );
  AND2_X1 U3372 ( .A1(n2673), .A2(n2672), .ZN(n2674) );
  OR2_X1 U3373 ( .A1(n2674), .A2(n2683), .ZN(n4130) );
  INV_X1 U3374 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2675) );
  OR2_X1 U3375 ( .A1(n3757), .A2(n2675), .ZN(n2676) );
  OAI21_X1 U3376 ( .B1(n4130), .B2(n2486), .A(n2676), .ZN(n2677) );
  INV_X1 U3377 ( .A(n2677), .ZN(n2681) );
  NAND2_X1 U3378 ( .A1(n2516), .A2(REG0_REG_21__SCAN_IN), .ZN(n2679) );
  NAND2_X1 U3379 ( .A1(n2717), .A2(REG1_REG_21__SCAN_IN), .ZN(n2678) );
  AND2_X1 U3380 ( .A1(n2679), .A2(n2678), .ZN(n2680) );
  NAND2_X1 U3381 ( .A1(n4145), .A2(n4306), .ZN(n2682) );
  AOI21_X1 U3382 ( .B1(n4124), .B2(n2682), .A(n2442), .ZN(n4107) );
  NOR2_X1 U3383 ( .A1(n2683), .A2(REG3_REG_22__SCAN_IN), .ZN(n2684) );
  OR2_X1 U3384 ( .A1(n2687), .A2(n2684), .ZN(n4117) );
  AOI22_X1 U3385 ( .A1(n2631), .A2(REG0_REG_22__SCAN_IN), .B1(n2717), .B2(
        REG1_REG_22__SCAN_IN), .ZN(n2686) );
  INV_X1 U3386 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4118) );
  OAI211_X1 U3387 ( .C1(n4117), .C2(n2486), .A(n2686), .B(n2685), .ZN(n4307)
         );
  NAND2_X1 U3388 ( .A1(n4307), .A2(n4116), .ZN(n2783) );
  NAND2_X1 U3389 ( .A1(n4090), .A2(n2783), .ZN(n4108) );
  NAND2_X1 U3390 ( .A1(n4107), .A2(n4108), .ZN(n4106) );
  NAND2_X1 U3391 ( .A1(n4106), .A2(n2443), .ZN(n4081) );
  OR2_X1 U3392 ( .A1(n2687), .A2(REG3_REG_23__SCAN_IN), .ZN(n2688) );
  NAND2_X1 U3393 ( .A1(n2692), .A2(n2688), .ZN(n4100) );
  AOI22_X1 U3394 ( .A1(n2631), .A2(REG0_REG_23__SCAN_IN), .B1(n2717), .B2(
        REG1_REG_23__SCAN_IN), .ZN(n2690) );
  INV_X1 U3395 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4101) );
  OR2_X1 U3396 ( .A1(n3757), .A2(n4101), .ZN(n2689) );
  INV_X1 U3397 ( .A(n4289), .ZN(n4075) );
  NAND2_X1 U3398 ( .A1(n4075), .A2(n4099), .ZN(n2691) );
  INV_X1 U3399 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U3400 ( .A1(n2692), .A2(n4940), .ZN(n2693) );
  NAND2_X1 U3401 ( .A1(n2707), .A2(n2693), .ZN(n3674) );
  OR2_X1 U3402 ( .A1(n3674), .A2(n2486), .ZN(n2697) );
  AOI22_X1 U3403 ( .A1(n2631), .A2(REG0_REG_24__SCAN_IN), .B1(n2717), .B2(
        REG1_REG_24__SCAN_IN), .ZN(n2696) );
  INV_X1 U3404 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2694) );
  OR2_X1 U3405 ( .A1(n3757), .A2(n2694), .ZN(n2695) );
  NAND2_X1 U3406 ( .A1(n3892), .A2(n4288), .ZN(n2699) );
  NOR2_X1 U3407 ( .A1(n3892), .A2(n4288), .ZN(n2698) );
  XNOR2_X1 U3408 ( .A(n2707), .B(REG3_REG_25__SCAN_IN), .ZN(n3641) );
  NAND2_X1 U3409 ( .A1(n3641), .A2(n2470), .ZN(n2704) );
  INV_X1 U3410 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4058) );
  NAND2_X1 U3411 ( .A1(n2717), .A2(REG1_REG_25__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U3412 ( .A1(n2631), .A2(REG0_REG_25__SCAN_IN), .ZN(n2700) );
  OAI211_X1 U3413 ( .C1(n4058), .C2(n3757), .A(n2701), .B(n2700), .ZN(n2702)
         );
  INV_X1 U3414 ( .A(n2702), .ZN(n2703) );
  NAND2_X1 U3415 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2705) );
  INV_X1 U3416 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3643) );
  INV_X1 U3417 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2706) );
  OAI21_X1 U3418 ( .B1(n2707), .B2(n3643), .A(n2706), .ZN(n2708) );
  NAND2_X1 U3419 ( .A1(n4043), .A2(n2470), .ZN(n2714) );
  INV_X1 U3420 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3421 ( .A1(n2631), .A2(REG0_REG_26__SCAN_IN), .ZN(n2710) );
  NAND2_X1 U3422 ( .A1(n2717), .A2(REG1_REG_26__SCAN_IN), .ZN(n2709) );
  OAI211_X1 U3423 ( .C1(n2711), .C2(n3757), .A(n2710), .B(n2709), .ZN(n2712)
         );
  INV_X1 U3424 ( .A(n2712), .ZN(n2713) );
  NAND2_X1 U3425 ( .A1(n2513), .A2(DATAI_26_), .ZN(n4042) );
  INV_X1 U3426 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4941) );
  AND2_X1 U3427 ( .A1(n2715), .A2(n4941), .ZN(n2716) );
  INV_X1 U3428 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4020) );
  NAND2_X1 U3429 ( .A1(n2717), .A2(REG1_REG_27__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U3430 ( .A1(n2516), .A2(REG0_REG_27__SCAN_IN), .ZN(n2718) );
  OAI211_X1 U3431 ( .C1(n4020), .C2(n3757), .A(n2719), .B(n2718), .ZN(n2720)
         );
  INV_X1 U3432 ( .A(n2720), .ZN(n2721) );
  OAI21_X1 U3433 ( .B1(n4021), .B2(n2486), .A(n2721), .ZN(n3891) );
  NAND2_X1 U3434 ( .A1(n2513), .A2(DATAI_27_), .ZN(n4019) );
  NAND2_X1 U3435 ( .A1(n4035), .A2(n4019), .ZN(n2723) );
  NOR2_X1 U3436 ( .A1(n4035), .A2(n4019), .ZN(n2722) );
  NAND2_X1 U3437 ( .A1(n2724), .A2(REG3_REG_28__SCAN_IN), .ZN(n4007) );
  INV_X1 U3438 ( .A(n2724), .ZN(n2726) );
  INV_X1 U3439 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2725) );
  NAND2_X1 U3440 ( .A1(n2726), .A2(n2725), .ZN(n2727) );
  NAND2_X1 U3441 ( .A1(n4007), .A2(n2727), .ZN(n3583) );
  OR2_X1 U3442 ( .A1(n3583), .A2(n2486), .ZN(n2732) );
  INV_X1 U3443 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3462) );
  NAND2_X1 U3444 ( .A1(n2717), .A2(REG1_REG_28__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U3445 ( .A1(n2516), .A2(REG0_REG_28__SCAN_IN), .ZN(n2728) );
  OAI211_X1 U3446 ( .C1(n3462), .C2(n3757), .A(n2729), .B(n2728), .ZN(n2730)
         );
  INV_X1 U3447 ( .A(n2730), .ZN(n2731) );
  NAND2_X1 U3448 ( .A1(n2513), .A2(DATAI_28_), .ZN(n3472) );
  INV_X1 U3449 ( .A(n3472), .ZN(n3580) );
  XNOR2_X1 U3450 ( .A(n2833), .B(n2832), .ZN(n3470) );
  NAND2_X1 U3451 ( .A1(n2244), .A2(IR_REG_31__SCAN_IN), .ZN(n2734) );
  NAND2_X1 U3452 ( .A1(n2736), .A2(n2735), .ZN(n2737) );
  NAND2_X1 U3453 ( .A1(n2737), .A2(IR_REG_31__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U3454 ( .A1(n2740), .A2(IR_REG_31__SCAN_IN), .ZN(n2741) );
  XNOR2_X1 U3455 ( .A(n4447), .B(n3046), .ZN(n2742) );
  NAND2_X1 U3456 ( .A1(n2742), .A2(n3989), .ZN(n3132) );
  AND2_X1 U3457 ( .A1(n3832), .A2(n4449), .ZN(n3034) );
  INV_X1 U34580 ( .A(n4684), .ZN(n4659) );
  NAND2_X1 U34590 ( .A1(n3132), .A2(n4659), .ZN(n4676) );
  INV_X1 U3460 ( .A(n4676), .ZN(n4341) );
  OR2_X1 U3461 ( .A1(n2743), .A2(n2796), .ZN(n2745) );
  NAND2_X1 U3462 ( .A1(n4447), .A2(n3874), .ZN(n2921) );
  NOR2_X2 U3463 ( .A1(n4457), .A2(n2921), .ZN(n4320) );
  OR2_X1 U3464 ( .A1(n4007), .A2(n2486), .ZN(n2750) );
  INV_X1 U3465 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2844) );
  NAND2_X1 U3466 ( .A1(n2516), .A2(REG0_REG_29__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U34670 ( .A1(n2462), .A2(REG2_REG_29__SCAN_IN), .ZN(n2746) );
  OAI211_X1 U3468 ( .C1(n2844), .C2(n2476), .A(n2747), .B(n2746), .ZN(n2748)
         );
  INV_X1 U34690 ( .A(n2748), .ZN(n2749) );
  NAND2_X1 U3470 ( .A1(n2750), .A2(n2749), .ZN(n3890) );
  INV_X1 U34710 ( .A(n3890), .ZN(n3840) );
  INV_X1 U3472 ( .A(n2921), .ZN(n2871) );
  NAND2_X1 U34730 ( .A1(n4457), .A2(n2871), .ZN(n4317) );
  NAND2_X1 U3474 ( .A1(n2943), .A2(n2807), .ZN(n3033) );
  OAI22_X1 U34750 ( .A1(n3840), .A2(n4317), .B1(n4315), .B2(n3472), .ZN(n2751)
         );
  AOI21_X1 U3476 ( .B1(n4320), .B2(n3891), .A(n2751), .ZN(n2792) );
  NAND2_X1 U34770 ( .A1(n2978), .A2(n2933), .ZN(n3767) );
  NAND2_X1 U3478 ( .A1(n3072), .A2(n3026), .ZN(n3776) );
  NAND2_X1 U34790 ( .A1(n3901), .A2(n3194), .ZN(n3773) );
  AND2_X1 U3480 ( .A1(n3776), .A2(n3773), .ZN(n3023) );
  NAND2_X1 U34810 ( .A1(n3024), .A2(n3023), .ZN(n2755) );
  NAND2_X1 U3482 ( .A1(n2755), .A2(n3776), .ZN(n3070) );
  INV_X1 U34830 ( .A(n3777), .ZN(n2756) );
  NAND2_X1 U3484 ( .A1(n2757), .A2(n3780), .ZN(n3118) );
  AND2_X1 U34850 ( .A1(n3900), .A2(n3154), .ZN(n3117) );
  NAND2_X1 U3486 ( .A1(n2758), .A2(n3654), .ZN(n3795) );
  NAND2_X1 U34870 ( .A1(n3899), .A2(n2289), .ZN(n3794) );
  INV_X1 U3488 ( .A(n3899), .ZN(n3281) );
  NAND2_X1 U34890 ( .A1(n3281), .A2(n3166), .ZN(n3782) );
  INV_X1 U3490 ( .A(n2759), .ZN(n2760) );
  NAND2_X1 U34910 ( .A1(n2375), .A2(n3274), .ZN(n3788) );
  NAND2_X1 U3492 ( .A1(n3320), .A2(n3788), .ZN(n2761) );
  NAND2_X1 U34930 ( .A1(n3897), .A2(n2376), .ZN(n3785) );
  NAND2_X1 U3494 ( .A1(n2761), .A2(n3785), .ZN(n3245) );
  INV_X1 U34950 ( .A(n3306), .ZN(n3298) );
  AND2_X1 U3496 ( .A1(n3896), .A2(n3298), .ZN(n3802) );
  INV_X1 U34970 ( .A(n3896), .ZN(n3397) );
  NAND2_X1 U3498 ( .A1(n3397), .A2(n3306), .ZN(n3787) );
  NAND2_X1 U34990 ( .A1(n3895), .A2(n3396), .ZN(n3805) );
  NAND2_X1 U3500 ( .A1(n2762), .A2(n3358), .ZN(n3803) );
  NAND2_X1 U35010 ( .A1(n4246), .A2(n2763), .ZN(n4237) );
  NAND2_X1 U3502 ( .A1(n4368), .A2(n4250), .ZN(n2764) );
  NAND2_X1 U35030 ( .A1(n4237), .A2(n2764), .ZN(n2766) );
  INV_X1 U3504 ( .A(n3418), .ZN(n2765) );
  NOR2_X1 U35050 ( .A1(n2766), .A2(n2765), .ZN(n3806) );
  NAND2_X1 U35060 ( .A1(n3419), .A2(n3806), .ZN(n2770) );
  NAND2_X1 U35070 ( .A1(n3333), .A2(n4365), .ZN(n4239) );
  NAND2_X1 U35080 ( .A1(n3416), .A2(n4239), .ZN(n2769) );
  INV_X1 U35090 ( .A(n2766), .ZN(n2768) );
  NOR2_X1 U35100 ( .A1(n4368), .A2(n4250), .ZN(n2767) );
  AOI21_X1 U35110 ( .B1(n2769), .B2(n2768), .A(n2767), .ZN(n3808) );
  NAND2_X1 U35120 ( .A1(n2770), .A2(n3808), .ZN(n3850) );
  INV_X1 U35130 ( .A(n3733), .ZN(n3381) );
  INV_X1 U35140 ( .A(n4217), .ZN(n4459) );
  NAND2_X1 U35150 ( .A1(n4459), .A2(n4347), .ZN(n3809) );
  NAND2_X1 U35160 ( .A1(n4217), .A2(n3456), .ZN(n3792) );
  NAND2_X1 U35170 ( .A1(n3809), .A2(n3792), .ZN(n3732) );
  INV_X1 U35180 ( .A(n3810), .ZN(n2771) );
  NOR2_X1 U35190 ( .A1(n3732), .A2(n2771), .ZN(n2772) );
  NAND2_X1 U35200 ( .A1(n3447), .A2(n2772), .ZN(n2773) );
  NAND2_X1 U35210 ( .A1(n2773), .A2(n3792), .ZN(n4216) );
  INV_X1 U35220 ( .A(n4225), .ZN(n2774) );
  NAND2_X1 U35230 ( .A1(n4216), .A2(n2774), .ZN(n2775) );
  NAND2_X1 U35240 ( .A1(n4220), .A2(n4333), .ZN(n4161) );
  NAND2_X1 U35250 ( .A1(n4163), .A2(n4161), .ZN(n2778) );
  NAND2_X1 U35260 ( .A1(n4472), .A2(n4173), .ZN(n2776) );
  NOR2_X1 U35270 ( .A1(n4472), .A2(n4173), .ZN(n2777) );
  AOI21_X1 U35280 ( .B1(n2778), .B2(n4084), .A(n2777), .ZN(n4152) );
  INV_X1 U35290 ( .A(n4169), .ZN(n4310) );
  NAND2_X1 U35300 ( .A1(n4310), .A2(n4143), .ZN(n2779) );
  NAND2_X1 U35310 ( .A1(n4199), .A2(n4087), .ZN(n2780) );
  NAND2_X1 U35320 ( .A1(n4482), .A2(n4211), .ZN(n4082) );
  NAND2_X1 U35330 ( .A1(n4084), .A2(n4082), .ZN(n3815) );
  AND2_X1 U35340 ( .A1(n4169), .A2(n4316), .ZN(n4086) );
  AOI21_X1 U35350 ( .B1(n4087), .B2(n3815), .A(n4086), .ZN(n3854) );
  NAND2_X1 U35360 ( .A1(n2780), .A2(n3854), .ZN(n2782) );
  NAND2_X1 U35370 ( .A1(n4318), .A2(n4306), .ZN(n3738) );
  NAND2_X1 U35380 ( .A1(n4090), .A2(n3738), .ZN(n3859) );
  INV_X1 U35390 ( .A(n3859), .ZN(n2781) );
  NAND2_X1 U35400 ( .A1(n2782), .A2(n2781), .ZN(n2786) );
  NOR2_X1 U35410 ( .A1(n4318), .A2(n4306), .ZN(n3819) );
  AND2_X1 U35420 ( .A1(n3819), .A2(n4090), .ZN(n2785) );
  NAND2_X1 U35430 ( .A1(n4289), .A2(n4099), .ZN(n2784) );
  NAND2_X1 U35440 ( .A1(n2784), .A2(n2783), .ZN(n3822) );
  NOR2_X1 U35450 ( .A1(n2785), .A2(n3822), .ZN(n3858) );
  NAND2_X1 U35460 ( .A1(n2786), .A2(n3858), .ZN(n4065) );
  NAND2_X1 U35470 ( .A1(n4097), .A2(n4288), .ZN(n3731) );
  OR2_X1 U35480 ( .A1(n4289), .A2(n4099), .ZN(n4064) );
  NAND2_X1 U35490 ( .A1(n3892), .A2(n4074), .ZN(n3765) );
  INV_X1 U35500 ( .A(n4271), .ZN(n4022) );
  NAND2_X1 U35510 ( .A1(n4022), .A2(n3713), .ZN(n3753) );
  OR2_X1 U35520 ( .A1(n4037), .A2(n4056), .ZN(n4031) );
  AND2_X1 U35530 ( .A1(n3891), .A2(n4019), .ZN(n3829) );
  INV_X1 U35540 ( .A(n3829), .ZN(n2787) );
  OR2_X1 U35550 ( .A1(n3891), .A2(n4019), .ZN(n2788) );
  INV_X1 U35560 ( .A(n2788), .ZN(n3867) );
  AOI21_X1 U35570 ( .B1(n4016), .B2(n4015), .A(n3867), .ZN(n2835) );
  INV_X1 U35580 ( .A(n2832), .ZN(n3737) );
  XNOR2_X1 U35590 ( .A(n2835), .B(n3737), .ZN(n2791) );
  NAND2_X1 U35600 ( .A1(n4447), .A2(n4449), .ZN(n2790) );
  INV_X1 U35610 ( .A(n3832), .ZN(n4448) );
  NAND2_X1 U35620 ( .A1(n4448), .A2(n3874), .ZN(n2789) );
  NAND2_X1 U35630 ( .A1(n2791), .A2(n4222), .ZN(n3461) );
  OAI211_X1 U35640 ( .C1(n3470), .C2(n4341), .A(n2792), .B(n3461), .ZN(n2829)
         );
  NAND2_X1 U35650 ( .A1(n2793), .A2(IR_REG_31__SCAN_IN), .ZN(n2794) );
  MUX2_X1 U35660 ( .A(IR_REG_31__SCAN_IN), .B(n2794), .S(IR_REG_25__SCAN_IN), 
        .Z(n2795) );
  NAND2_X1 U35670 ( .A1(n2795), .A2(n2237), .ZN(n2867) );
  NAND2_X1 U35680 ( .A1(n2867), .A2(B_REG_SCAN_IN), .ZN(n2800) );
  OR2_X1 U35690 ( .A1(n2797), .A2(n2796), .ZN(n2806) );
  INV_X1 U35700 ( .A(IR_REG_23__SCAN_IN), .ZN(n2805) );
  NAND2_X1 U35710 ( .A1(n2806), .A2(n2805), .ZN(n2798) );
  NAND2_X1 U35720 ( .A1(n2798), .A2(IR_REG_31__SCAN_IN), .ZN(n2799) );
  MUX2_X1 U35730 ( .A(n2800), .B(B_REG_SCAN_IN), .S(n4446), .Z(n2802) );
  NAND2_X1 U35740 ( .A1(n2802), .A2(n2804), .ZN(n2863) );
  INV_X1 U35750 ( .A(D_REG_1__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U35760 ( .A1(n2823), .A2(n2803), .ZN(n3041) );
  INV_X1 U35770 ( .A(n2804), .ZN(n2868) );
  NAND2_X1 U35780 ( .A1(n2868), .A2(n2867), .ZN(n2917) );
  NAND2_X1 U35790 ( .A1(n3041), .A2(n2917), .ZN(n2820) );
  INV_X1 U35800 ( .A(n2867), .ZN(n2853) );
  XNOR2_X1 U35810 ( .A(n2806), .B(n2805), .ZN(n3011) );
  NAND2_X1 U3582 ( .A1(n4684), .A2(n2807), .ZN(n2947) );
  AND2_X1 U3583 ( .A1(n3832), .A2(n3989), .ZN(n2920) );
  OR2_X1 U3584 ( .A1(n2921), .A2(n2920), .ZN(n3038) );
  NAND2_X1 U3585 ( .A1(n2947), .A2(n3038), .ZN(n2808) );
  NOR2_X1 U3586 ( .A1(n3040), .A2(n2808), .ZN(n2819) );
  NOR4_X1 U3587 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2812) );
  NOR4_X1 U3588 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2811) );
  NOR4_X1 U3589 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2810) );
  NOR4_X1 U3590 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2809) );
  NAND4_X1 U3591 ( .A1(n2812), .A2(n2811), .A3(n2810), .A4(n2809), .ZN(n2818)
         );
  NOR2_X1 U3592 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_29__SCAN_IN), .ZN(n2816)
         );
  NOR4_X1 U3593 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2815) );
  NOR4_X1 U3594 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2814) );
  NOR4_X1 U3595 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2813) );
  NAND4_X1 U3596 ( .A1(n2816), .A2(n2815), .A3(n2814), .A4(n2813), .ZN(n2817)
         );
  OAI21_X1 U3597 ( .B1(n2818), .B2(n2817), .A(n2823), .ZN(n2918) );
  INV_X1 U3598 ( .A(D_REG_0__SCAN_IN), .ZN(n2822) );
  INV_X1 U3599 ( .A(n4446), .ZN(n2864) );
  MUX2_X1 U3600 ( .A(REG1_REG_28__SCAN_IN), .B(n2829), .S(n4699), .Z(n2824) );
  INV_X1 U3601 ( .A(n2824), .ZN(n2827) );
  NAND2_X1 U3602 ( .A1(n3085), .A2(n3086), .ZN(n3177) );
  INV_X1 U3603 ( .A(n4018), .ZN(n2825) );
  INV_X1 U3604 ( .A(n3033), .ZN(n2826) );
  NAND2_X1 U3605 ( .A1(n2827), .A2(n2446), .ZN(U3546) );
  INV_X1 U3606 ( .A(n2919), .ZN(n3044) );
  MUX2_X1 U3607 ( .A(REG0_REG_28__SCAN_IN), .B(n2829), .S(n4687), .Z(n2830) );
  INV_X1 U3608 ( .A(n2830), .ZN(n2831) );
  NAND2_X1 U3609 ( .A1(n2831), .A2(n2445), .ZN(U3514) );
  NAND2_X1 U3610 ( .A1(n2513), .A2(DATAI_29_), .ZN(n4003) );
  XNOR2_X1 U3611 ( .A(n3890), .B(n3839), .ZN(n3763) );
  INV_X1 U3612 ( .A(n3763), .ZN(n2837) );
  INV_X1 U3613 ( .A(n3868), .ZN(n2834) );
  XOR2_X1 U3614 ( .A(n2837), .B(n2836), .Z(n2842) );
  XNOR2_X1 U3615 ( .A(n2838), .B(IR_REG_27__SCAN_IN), .ZN(n4494) );
  AOI21_X1 U3616 ( .B1(B_REG_SCAN_IN), .B2(n4494), .A(n4317), .ZN(n3995) );
  INV_X1 U3617 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2841) );
  NAND2_X1 U3618 ( .A1(n2717), .A2(REG1_REG_30__SCAN_IN), .ZN(n2840) );
  NAND2_X1 U3619 ( .A1(n2516), .A2(REG0_REG_30__SCAN_IN), .ZN(n2839) );
  OAI211_X1 U3620 ( .C1(n3757), .C2(n2841), .A(n2840), .B(n2839), .ZN(n3889)
         );
  AOI22_X1 U3621 ( .A1(n2842), .A2(n4222), .B1(n3995), .B2(n3889), .ZN(n4006)
         );
  NAND2_X1 U3622 ( .A1(n4005), .A2(n4320), .ZN(n2843) );
  INV_X1 U3623 ( .A(n2845), .ZN(n2846) );
  NAND2_X1 U3624 ( .A1(n2848), .A2(n2847), .ZN(U3547) );
  NAND2_X1 U3625 ( .A1(n2850), .A2(n2849), .ZN(U3515) );
  INV_X2 U3626 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3627 ( .A(n4641), .ZN(n2851) );
  NOR2_X2 U3628 ( .A1(n3012), .A2(n2851), .ZN(U4043) );
  INV_X1 U3629 ( .A(DATAI_21_), .ZN(n5044) );
  NAND2_X1 U3630 ( .A1(n3874), .A2(STATE_REG_SCAN_IN), .ZN(n2852) );
  OAI21_X1 U3631 ( .B1(STATE_REG_SCAN_IN), .B2(n5044), .A(n2852), .ZN(U3331)
         );
  INV_X1 U3632 ( .A(DATAI_25_), .ZN(n2855) );
  NAND2_X1 U3633 ( .A1(n2853), .A2(STATE_REG_SCAN_IN), .ZN(n2854) );
  OAI21_X1 U3634 ( .B1(STATE_REG_SCAN_IN), .B2(n2855), .A(n2854), .ZN(U3327)
         );
  INV_X1 U3635 ( .A(IR_REG_30__SCAN_IN), .ZN(n2857) );
  NAND3_X1 U3636 ( .A1(n2857), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n2859) );
  INV_X1 U3637 ( .A(DATAI_31_), .ZN(n2858) );
  OAI22_X1 U3638 ( .A1(n2856), .A2(n2859), .B1(STATE_REG_SCAN_IN), .B2(n2858), 
        .ZN(U3321) );
  INV_X1 U3639 ( .A(DATAI_27_), .ZN(n4943) );
  NAND2_X1 U3640 ( .A1(n4494), .A2(STATE_REG_SCAN_IN), .ZN(n2860) );
  OAI21_X1 U3641 ( .B1(STATE_REG_SCAN_IN), .B2(n4943), .A(n2860), .ZN(U3325)
         );
  INV_X1 U3642 ( .A(DATAI_29_), .ZN(n2862) );
  NAND2_X1 U3643 ( .A1(n2469), .A2(STATE_REG_SCAN_IN), .ZN(n2861) );
  OAI21_X1 U3644 ( .B1(STATE_REG_SCAN_IN), .B2(n2862), .A(n2861), .ZN(U3323)
         );
  AND2_X2 U3645 ( .A1(n2863), .A2(n2949), .ZN(n4640) );
  NAND3_X1 U3646 ( .A1(n2868), .A2(n4641), .A3(n2864), .ZN(n2865) );
  OAI21_X1 U3647 ( .B1(n4640), .B2(D_REG_0__SCAN_IN), .A(n2865), .ZN(n2866) );
  INV_X1 U3648 ( .A(n2866), .ZN(U3458) );
  NAND3_X1 U3649 ( .A1(n2868), .A2(n4641), .A3(n2867), .ZN(n2869) );
  OAI21_X1 U3650 ( .B1(n4640), .B2(D_REG_1__SCAN_IN), .A(n2869), .ZN(n2870) );
  INV_X1 U3651 ( .A(n2870), .ZN(U3459) );
  NAND2_X1 U3652 ( .A1(n3011), .A2(n2871), .ZN(n2872) );
  NAND2_X1 U3653 ( .A1(n2513), .A2(n2872), .ZN(n2880) );
  INV_X1 U3654 ( .A(n3011), .ZN(n2874) );
  NAND2_X1 U3655 ( .A1(n2874), .A2(STATE_REG_SCAN_IN), .ZN(n3887) );
  NAND2_X1 U3656 ( .A1(n3040), .A2(n3887), .ZN(n2881) );
  NOR2_X1 U3657 ( .A1(n4604), .A2(U4043), .ZN(U3148) );
  INV_X1 U3658 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4690) );
  XNOR2_X1 U3659 ( .A(n2887), .B(REG1_REG_1__SCAN_IN), .ZN(n3906) );
  AND2_X1 U3660 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3905)
         );
  NAND2_X1 U3661 ( .A1(n3906), .A2(n3905), .ZN(n3904) );
  NAND2_X1 U3662 ( .A1(n4456), .A2(REG1_REG_1__SCAN_IN), .ZN(n2875) );
  NAND2_X1 U3663 ( .A1(n3904), .A2(n2875), .ZN(n3920) );
  NAND2_X1 U3664 ( .A1(n4455), .A2(REG1_REG_2__SCAN_IN), .ZN(n2876) );
  NAND2_X1 U3665 ( .A1(n3919), .A2(n2876), .ZN(n2877) );
  INV_X1 U3666 ( .A(n4454), .ZN(n2891) );
  XNOR2_X1 U3667 ( .A(n2877), .B(n2891), .ZN(n3928) );
  NAND2_X1 U3668 ( .A1(n3928), .A2(REG1_REG_3__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U3669 ( .A1(n2877), .A2(n4454), .ZN(n2878) );
  NAND2_X1 U3670 ( .A1(n3927), .A2(n2878), .ZN(n2879) );
  INV_X1 U3671 ( .A(n4453), .ZN(n3065) );
  XNOR2_X1 U3672 ( .A(n4452), .B(REG1_REG_5__SCAN_IN), .ZN(n2883) );
  NOR2_X1 U3673 ( .A1(n2884), .A2(n2883), .ZN(n2910) );
  INV_X1 U3674 ( .A(n2880), .ZN(n2882) );
  INV_X1 U3675 ( .A(n4494), .ZN(n3053) );
  INV_X1 U3676 ( .A(n4606), .ZN(n2911) );
  AOI211_X1 U3677 ( .C1(n2884), .C2(n2883), .A(n2910), .B(n2911), .ZN(n2904)
         );
  INV_X1 U3678 ( .A(n4452), .ZN(n2902) );
  MUX2_X1 U3679 ( .A(REG2_REG_5__SCAN_IN), .B(n2885), .S(n4452), .Z(n2899) );
  MUX2_X1 U3680 ( .A(REG2_REG_2__SCAN_IN), .B(n2886), .S(n4455), .Z(n3918) );
  INV_X1 U3681 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2888) );
  AND2_X1 U3682 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3909)
         );
  NAND2_X1 U3683 ( .A1(n4456), .A2(REG2_REG_1__SCAN_IN), .ZN(n2889) );
  NAND2_X1 U3684 ( .A1(n3907), .A2(n2889), .ZN(n3917) );
  NAND2_X1 U3685 ( .A1(n4455), .A2(REG2_REG_2__SCAN_IN), .ZN(n2890) );
  NAND2_X1 U3686 ( .A1(n3916), .A2(n2890), .ZN(n2892) );
  XNOR2_X1 U3687 ( .A(n2892), .B(n2891), .ZN(n3930) );
  NAND2_X1 U3688 ( .A1(n3930), .A2(REG2_REG_3__SCAN_IN), .ZN(n2894) );
  NAND2_X1 U3689 ( .A1(n2892), .A2(n4454), .ZN(n2893) );
  NAND2_X1 U3690 ( .A1(n2896), .A2(n4453), .ZN(n2897) );
  NOR2_X1 U3691 ( .A1(n4457), .A2(n3053), .ZN(n3884) );
  NAND2_X1 U3692 ( .A1(n2898), .A2(n2899), .ZN(n2906) );
  OAI211_X1 U3693 ( .C1(n2899), .C2(n2898), .A(n4552), .B(n2906), .ZN(n2901)
         );
  INV_X1 U3694 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4831) );
  NOR2_X1 U3695 ( .A1(STATE_REG_SCAN_IN), .A2(n4831), .ZN(n3653) );
  AOI21_X1 U3696 ( .B1(n4604), .B2(ADDR_REG_5__SCAN_IN), .A(n3653), .ZN(n2900)
         );
  OAI211_X1 U3697 ( .C1(n4610), .C2(n2902), .A(n2901), .B(n2900), .ZN(n2903)
         );
  OR2_X1 U3698 ( .A1(n2904), .A2(n2903), .ZN(U3245) );
  NAND2_X1 U3699 ( .A1(n4452), .A2(REG2_REG_5__SCAN_IN), .ZN(n2905) );
  NAND2_X1 U3700 ( .A1(n2906), .A2(n2905), .ZN(n2957) );
  INV_X1 U3701 ( .A(n4451), .ZN(n2909) );
  XNOR2_X1 U3702 ( .A(n2957), .B(n2909), .ZN(n2959) );
  XNOR2_X1 U3703 ( .A(n2959), .B(n3138), .ZN(n2915) );
  NOR2_X1 U3704 ( .A1(STATE_REG_SCAN_IN), .A2(n2907), .ZN(n3165) );
  AOI21_X1 U3705 ( .B1(n4604), .B2(ADDR_REG_6__SCAN_IN), .A(n3165), .ZN(n2908)
         );
  OAI21_X1 U3706 ( .B1(n4610), .B2(n2909), .A(n2908), .ZN(n2914) );
  INV_X1 U3707 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3228) );
  NOR2_X1 U3708 ( .A1(n2912), .A2(n3228), .ZN(n2954) );
  AOI211_X1 U3709 ( .C1(n3228), .C2(n2912), .A(n2911), .B(n2954), .ZN(n2913)
         );
  AOI211_X1 U3710 ( .C1(n4552), .C2(n2915), .A(n2914), .B(n2913), .ZN(n2916)
         );
  INV_X1 U3711 ( .A(n2916), .ZN(U3246) );
  AND2_X1 U3712 ( .A1(n2918), .A2(n2917), .ZN(n3043) );
  NAND3_X1 U3713 ( .A1(n3043), .A2(n2919), .A3(n3041), .ZN(n2977) );
  INV_X1 U3714 ( .A(n2977), .ZN(n2924) );
  OR2_X1 U3715 ( .A1(n3033), .A2(n2920), .ZN(n2922) );
  NAND2_X1 U3716 ( .A1(n2922), .A2(n2921), .ZN(n2940) );
  NOR2_X1 U3717 ( .A1(n3040), .A2(n2940), .ZN(n2923) );
  NAND4_X1 U3718 ( .A1(n2928), .A2(n2927), .A3(n2926), .A4(n2925), .ZN(n3035)
         );
  INV_X1 U3719 ( .A(n3569), .ZN(n2929) );
  NAND2_X2 U3720 ( .A1(n2929), .A2(n4679), .ZN(n2984) );
  NAND2_X1 U3721 ( .A1(n3035), .A2(n3009), .ZN(n2932) );
  INV_X1 U3722 ( .A(n3012), .ZN(n2930) );
  AOI22_X1 U3723 ( .A1(n2933), .A2(n3562), .B1(IR_REG_0__SCAN_IN), .B2(n2930), 
        .ZN(n2931) );
  NAND2_X1 U3724 ( .A1(n2932), .A2(n2931), .ZN(n2938) );
  NAND2_X1 U3725 ( .A1(n3035), .A2(n3562), .ZN(n2937) );
  INV_X1 U3726 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2934) );
  NAND2_X1 U3727 ( .A1(n2933), .A2(n3557), .ZN(n2971) );
  OAI21_X1 U3728 ( .B1(n3012), .B2(n2934), .A(n2971), .ZN(n2935) );
  INV_X1 U3729 ( .A(n2935), .ZN(n2936) );
  NAND2_X1 U3730 ( .A1(n2937), .A2(n2936), .ZN(n2939) );
  NAND2_X1 U3731 ( .A1(n2939), .A2(n2938), .ZN(n2973) );
  OAI21_X1 U3732 ( .B1(n2938), .B2(n2939), .A(n2973), .ZN(n3055) );
  NAND2_X1 U3733 ( .A1(n2940), .A2(n4315), .ZN(n2941) );
  NAND2_X1 U3734 ( .A1(n2977), .A2(n2941), .ZN(n2942) );
  NAND2_X1 U3735 ( .A1(n2942), .A2(n3038), .ZN(n3014) );
  INV_X1 U3736 ( .A(n3014), .ZN(n2945) );
  NOR2_X1 U3737 ( .A1(n2943), .A2(n4449), .ZN(n2968) );
  AND2_X1 U3738 ( .A1(n4641), .A2(n2968), .ZN(n2944) );
  AND2_X1 U3739 ( .A1(n3562), .A2(n2944), .ZN(n3883) );
  NAND2_X1 U3740 ( .A1(n2977), .A2(n3883), .ZN(n3015) );
  NAND3_X1 U3741 ( .A1(n2945), .A2(n2949), .A3(n3015), .ZN(n2997) );
  NAND2_X1 U3742 ( .A1(n2949), .A2(n4366), .ZN(n2946) );
  OR2_X1 U3743 ( .A1(n2977), .A2(n2946), .ZN(n2950) );
  INV_X1 U3744 ( .A(n2947), .ZN(n2948) );
  NAND2_X2 U3745 ( .A1(n2949), .A2(n2948), .ZN(n4253) );
  NAND2_X1 U3746 ( .A1(n2950), .A2(n4253), .ZN(n4484) );
  INV_X1 U3747 ( .A(n4484), .ZN(n4461) );
  NAND2_X1 U3748 ( .A1(n3883), .A2(n4457), .ZN(n2951) );
  OR2_X1 U3749 ( .A1(n2977), .A2(n2951), .ZN(n3703) );
  OAI22_X1 U3750 ( .A1(n4461), .A2(n3086), .B1(n3184), .B2(n3703), .ZN(n2952)
         );
  AOI21_X1 U3751 ( .B1(REG3_REG_0__SCAN_IN), .B2(n2997), .A(n2952), .ZN(n2953)
         );
  OAI21_X1 U3752 ( .B1(n3679), .B2(n3055), .A(n2953), .ZN(U3229) );
  AOI21_X1 U3753 ( .B1(n4451), .B2(n2955), .A(n2954), .ZN(n3963) );
  INV_X1 U3754 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4694) );
  MUX2_X1 U3755 ( .A(REG1_REG_7__SCAN_IN), .B(n4694), .S(n4450), .Z(n2956) );
  XNOR2_X1 U3756 ( .A(n3963), .B(n2956), .ZN(n2965) );
  AND2_X1 U3757 ( .A1(n2957), .A2(n4451), .ZN(n2958) );
  AOI21_X1 U3758 ( .B1(n2959), .B2(REG2_REG_6__SCAN_IN), .A(n2958), .ZN(n2961)
         );
  MUX2_X1 U3759 ( .A(n3938), .B(REG2_REG_7__SCAN_IN), .S(n4450), .Z(n2960) );
  AOI211_X1 U3760 ( .C1(n2961), .C2(n2960), .A(n3937), .B(n4600), .ZN(n2964)
         );
  INV_X1 U3761 ( .A(n4450), .ZN(n3961) );
  INV_X1 U3762 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4969) );
  NOR2_X1 U3763 ( .A1(STATE_REG_SCAN_IN), .A2(n4969), .ZN(n3236) );
  AOI21_X1 U3764 ( .B1(n4604), .B2(ADDR_REG_7__SCAN_IN), .A(n3236), .ZN(n2962)
         );
  OAI21_X1 U3765 ( .B1(n4610), .B2(n3961), .A(n2962), .ZN(n2963) );
  AOI211_X1 U3766 ( .C1(n2965), .C2(n4606), .A(n2964), .B(n2963), .ZN(n2966)
         );
  INV_X1 U3767 ( .A(n2966), .ZN(U3247) );
  INV_X1 U3768 ( .A(n2997), .ZN(n2982) );
  INV_X1 U3769 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3087) );
  INV_X1 U3770 ( .A(n2968), .ZN(n2969) );
  NAND2_X1 U3771 ( .A1(n2971), .A2(n3552), .ZN(n2972) );
  NAND2_X1 U3772 ( .A1(n2973), .A2(n2972), .ZN(n2975) );
  NAND2_X1 U3773 ( .A1(n2974), .A2(n2975), .ZN(n2988) );
  OAI211_X1 U3774 ( .C1(n2974), .C2(n2975), .A(n2988), .B(n4479), .ZN(n2981)
         );
  INV_X1 U3775 ( .A(n4457), .ZN(n3054) );
  NAND2_X1 U3776 ( .A1(n3054), .A2(n3883), .ZN(n2976) );
  OR2_X1 U3777 ( .A1(n2977), .A2(n2976), .ZN(n4458) );
  OAI22_X1 U3778 ( .A1(n2978), .A2(n4458), .B1(n3199), .B2(n3703), .ZN(n2979)
         );
  AOI21_X1 U3779 ( .B1(n3088), .B2(n4484), .A(n2979), .ZN(n2980) );
  OAI211_X1 U3780 ( .C1(n2982), .C2(n3087), .A(n2981), .B(n2980), .ZN(U3219)
         );
  OAI22_X1 U3781 ( .A1(n3199), .A2(n3099), .B1(n2995), .B2(n3569), .ZN(n2983)
         );
  XNOR2_X1 U3782 ( .A(n2983), .B(n3570), .ZN(n3000) );
  OAI22_X1 U3783 ( .A1(n3199), .A2(n2984), .B1(n2995), .B2(n3572), .ZN(n3001)
         );
  XNOR2_X1 U3784 ( .A(n3000), .B(n3001), .ZN(n2993) );
  INV_X1 U3785 ( .A(n2985), .ZN(n2986) );
  NAND2_X1 U3786 ( .A1(n2988), .A2(n2987), .ZN(n2992) );
  INV_X1 U3787 ( .A(n2992), .ZN(n2990) );
  INV_X1 U3788 ( .A(n3005), .ZN(n2991) );
  AOI21_X1 U3789 ( .B1(n2993), .B2(n2992), .A(n2991), .ZN(n2999) );
  INV_X2 U3790 ( .A(n3703), .ZN(n4471) );
  AOI22_X1 U3791 ( .A1(n2291), .A2(n4481), .B1(n4471), .B2(n3901), .ZN(n2994)
         );
  OAI21_X1 U3792 ( .B1(n4461), .B2(n2995), .A(n2994), .ZN(n2996) );
  AOI21_X1 U3793 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2997), .A(n2996), .ZN(n2998)
         );
  OAI21_X1 U3794 ( .B1(n2999), .B2(n3679), .A(n2998), .ZN(U3234) );
  INV_X1 U3795 ( .A(n3000), .ZN(n3003) );
  INV_X1 U3796 ( .A(n3001), .ZN(n3002) );
  NAND2_X1 U3797 ( .A1(n3003), .A2(n3002), .ZN(n3004) );
  NAND2_X1 U3798 ( .A1(n3901), .A2(n3562), .ZN(n3007) );
  NAND2_X1 U3799 ( .A1(n3026), .A2(n3557), .ZN(n3006) );
  NAND2_X1 U3800 ( .A1(n3007), .A2(n3006), .ZN(n3008) );
  NOR2_X1 U3801 ( .A1(n3194), .A2(n3572), .ZN(n3010) );
  AOI21_X1 U3802 ( .B1(n3901), .B2(n3561), .A(n3010), .ZN(n3105) );
  XNOR2_X1 U3803 ( .A(n3104), .B(n3105), .ZN(n3102) );
  XOR2_X1 U3804 ( .A(n3103), .B(n3102), .Z(n3021) );
  OAI22_X1 U3805 ( .A1(n3282), .A2(n3703), .B1(n3199), .B2(n4458), .ZN(n3019)
         );
  NAND2_X1 U3806 ( .A1(n3012), .A2(n3011), .ZN(n3013) );
  OAI21_X1 U3807 ( .B1(n3014), .B2(n3013), .A(STATE_REG_SCAN_IN), .ZN(n3016)
         );
  INV_X1 U3808 ( .A(n4488), .ZN(n3712) );
  MUX2_X1 U3809 ( .A(U3149), .B(n3712), .S(n3017), .Z(n3018) );
  AOI211_X1 U3810 ( .C1(n3026), .C2(n4484), .A(n3019), .B(n3018), .ZN(n3020)
         );
  OAI21_X1 U3811 ( .B1(n3021), .B2(n3679), .A(n3020), .ZN(U3215) );
  INV_X1 U3812 ( .A(n3023), .ZN(n3740) );
  XNOR2_X1 U3813 ( .A(n3022), .B(n3740), .ZN(n3192) );
  XNOR2_X1 U3814 ( .A(n3024), .B(n3023), .ZN(n3025) );
  NAND2_X1 U3815 ( .A1(n3025), .A2(n4222), .ZN(n3193) );
  AOI22_X1 U3816 ( .A1(n2502), .A2(n4367), .B1(n3026), .B2(n4366), .ZN(n3027)
         );
  OAI211_X1 U3817 ( .C1(n3199), .C2(n4371), .A(n3193), .B(n3027), .ZN(n3028)
         );
  AOI21_X1 U3818 ( .B1(n4676), .B2(n3192), .A(n3028), .ZN(n3032) );
  NOR2_X1 U3819 ( .A1(n3176), .A2(n3194), .ZN(n3029) );
  NOR2_X1 U3820 ( .A1(n3029), .A2(n3076), .ZN(n3195) );
  INV_X1 U3821 ( .A(n4443), .ZN(n4415) );
  AOI22_X1 U3822 ( .A1(n3195), .A2(n4415), .B1(REG0_REG_3__SCAN_IN), .B2(n4685), .ZN(n3030) );
  OAI21_X1 U3823 ( .B1(n3032), .B2(n4685), .A(n3030), .ZN(U3473) );
  INV_X1 U3824 ( .A(n4377), .ZN(n4325) );
  AOI22_X1 U3825 ( .A1(n3195), .A2(n4325), .B1(REG1_REG_3__SCAN_IN), .B2(n4696), .ZN(n3031) );
  OAI21_X1 U3826 ( .B1(n3032), .B2(n4696), .A(n3031), .ZN(U3521) );
  NOR2_X1 U3827 ( .A1(n3086), .A2(n3033), .ZN(n4655) );
  INV_X1 U3828 ( .A(n3034), .ZN(n3037) );
  INV_X1 U3829 ( .A(n3132), .ZN(n3402) );
  NAND2_X1 U3830 ( .A1(n3035), .A2(n3086), .ZN(n3769) );
  NAND2_X1 U3831 ( .A1(n3767), .A2(n3769), .ZN(n4656) );
  OAI21_X1 U3832 ( .B1(n3402), .B2(n4222), .A(n4656), .ZN(n3036) );
  OAI21_X1 U3833 ( .B1(n3184), .B2(n4317), .A(n3036), .ZN(n4654) );
  AOI21_X1 U3834 ( .B1(n4655), .B2(n3037), .A(n4654), .ZN(n3050) );
  INV_X1 U3835 ( .A(n3038), .ZN(n3039) );
  NOR2_X1 U3836 ( .A1(n3040), .A2(n3039), .ZN(n3042) );
  NAND4_X1 U3837 ( .A1(n3044), .A2(n3043), .A3(n3042), .A4(n3041), .ZN(n3045)
         );
  NAND2_X2 U3838 ( .A1(n3045), .A2(n4253), .ZN(n4256) );
  INV_X1 U3839 ( .A(n4253), .ZN(n4619) );
  AOI22_X1 U3840 ( .A1(n4489), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4619), .ZN(n3049) );
  OR2_X1 U3841 ( .A1(n3046), .A2(n3989), .ZN(n3131) );
  INV_X1 U3842 ( .A(n3131), .ZN(n3047) );
  NAND2_X1 U3843 ( .A1(n4656), .A2(n4624), .ZN(n3048) );
  OAI211_X1 U3844 ( .C1(n3050), .C2(n4489), .A(n3049), .B(n3048), .ZN(U3290)
         );
  NAND2_X1 U3845 ( .A1(n4494), .A2(n3051), .ZN(n3052) );
  NAND2_X1 U3846 ( .A1(n3054), .A2(n3052), .ZN(n4495) );
  INV_X1 U3847 ( .A(n4495), .ZN(n4493) );
  INV_X1 U3848 ( .A(IR_REG_0__SCAN_IN), .ZN(n4960) );
  NAND3_X1 U3849 ( .A1(n3055), .A2(n3054), .A3(n3053), .ZN(n3057) );
  AOI21_X1 U3850 ( .B1(n3884), .B2(n3909), .A(n3903), .ZN(n3056) );
  OAI211_X1 U3851 ( .C1(n4493), .C2(IR_REG_0__SCAN_IN), .A(n3057), .B(n3056), 
        .ZN(n3925) );
  XNOR2_X1 U3852 ( .A(n3058), .B(REG2_REG_4__SCAN_IN), .ZN(n3067) );
  INV_X1 U3853 ( .A(n3059), .ZN(n3060) );
  INV_X1 U3854 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4692) );
  NAND2_X1 U3855 ( .A1(n3060), .A2(n4692), .ZN(n3061) );
  NAND3_X1 U3856 ( .A1(n4606), .A2(n3062), .A3(n3061), .ZN(n3064) );
  AND2_X1 U3857 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3109) );
  AOI21_X1 U3858 ( .B1(n4604), .B2(ADDR_REG_4__SCAN_IN), .A(n3109), .ZN(n3063)
         );
  OAI211_X1 U3859 ( .C1(n4610), .C2(n3065), .A(n3064), .B(n3063), .ZN(n3066)
         );
  AOI21_X1 U3860 ( .B1(n4552), .B2(n3067), .A(n3066), .ZN(n3068) );
  NAND2_X1 U3861 ( .A1(n3925), .A2(n3068), .ZN(U3244) );
  XNOR2_X1 U3862 ( .A(n3069), .B(n3739), .ZN(n3078) );
  XOR2_X1 U3863 ( .A(n3739), .B(n3070), .Z(n3074) );
  AOI22_X1 U3864 ( .A1(n3900), .A2(n4367), .B1(n4366), .B2(n3110), .ZN(n3071)
         );
  OAI21_X1 U3865 ( .B1(n3072), .B2(n4371), .A(n3071), .ZN(n3073) );
  AOI21_X1 U3866 ( .B1(n3074), .B2(n4222), .A(n3073), .ZN(n3075) );
  OAI21_X1 U3867 ( .B1(n3078), .B2(n3132), .A(n3075), .ZN(n4670) );
  OAI211_X1 U3868 ( .C1(n3076), .C2(n3101), .A(n4664), .B(n3123), .ZN(n4669)
         );
  OAI22_X1 U3869 ( .A1(n4669), .A2(n4449), .B1(n4253), .B2(n3113), .ZN(n3077)
         );
  OAI21_X1 U3870 ( .B1(n4670), .B2(n3077), .A(n4256), .ZN(n3080) );
  INV_X1 U3871 ( .A(n3078), .ZN(n4672) );
  AOI22_X1 U3872 ( .A1(n4672), .A2(n4624), .B1(REG2_REG_4__SCAN_IN), .B2(n4489), .ZN(n3079) );
  NAND2_X1 U3873 ( .A1(n3080), .A2(n3079), .ZN(U3286) );
  OR2_X1 U3874 ( .A1(n3081), .A2(n2752), .ZN(n3082) );
  NAND2_X1 U3875 ( .A1(n3083), .A2(n3082), .ZN(n4660) );
  INV_X1 U3876 ( .A(n4660), .ZN(n3097) );
  AND2_X1 U3877 ( .A1(n4664), .A2(n3989), .ZN(n3084) );
  OAI21_X1 U3878 ( .B1(n3086), .B2(n3085), .A(n3177), .ZN(n4658) );
  OAI22_X1 U3879 ( .A1(n4252), .A2(n4658), .B1(n3087), .B2(n4253), .ZN(n3096)
         );
  NAND2_X1 U3880 ( .A1(n3088), .A2(n4366), .ZN(n3090) );
  NAND2_X1 U3881 ( .A1(n3035), .A2(n4320), .ZN(n3089) );
  OAI211_X1 U3882 ( .C1(n3199), .C2(n4317), .A(n3090), .B(n3089), .ZN(n3091)
         );
  INV_X1 U3883 ( .A(n3091), .ZN(n3094) );
  XNOR2_X1 U3884 ( .A(n2752), .B(n3767), .ZN(n3092) );
  NAND2_X1 U3885 ( .A1(n3092), .A2(n4222), .ZN(n3093) );
  OAI211_X1 U3886 ( .C1(n4660), .C2(n3132), .A(n3094), .B(n3093), .ZN(n4662)
         );
  MUX2_X1 U3887 ( .A(n4662), .B(REG2_REG_1__SCAN_IN), .S(n4629), .Z(n3095) );
  AOI211_X1 U3888 ( .C1(n3097), .C2(n4624), .A(n3096), .B(n3095), .ZN(n3098)
         );
  INV_X1 U3889 ( .A(n3098), .ZN(U3289) );
  XNOR2_X1 U3890 ( .A(n3100), .B(n3570), .ZN(n3147) );
  OAI22_X1 U3891 ( .A1(n3282), .A2(n2984), .B1(n3572), .B2(n3101), .ZN(n3146)
         );
  XNOR2_X1 U3892 ( .A(n3147), .B(n3146), .ZN(n3149) );
  INV_X1 U3893 ( .A(n3104), .ZN(n3106) );
  NAND2_X1 U3894 ( .A1(n3106), .A2(n3105), .ZN(n3107) );
  AOI211_X1 U3895 ( .C1(n3149), .C2(n3150), .A(n3679), .B(n2263), .ZN(n3115)
         );
  AOI21_X1 U3896 ( .B1(n4471), .B2(n3900), .A(n3109), .ZN(n3112) );
  AOI22_X1 U3897 ( .A1(n4481), .A2(n3901), .B1(n4484), .B2(n3110), .ZN(n3111)
         );
  OAI211_X1 U3898 ( .C1(n4488), .C2(n3113), .A(n3112), .B(n3111), .ZN(n3114)
         );
  OR2_X1 U3899 ( .A1(n3115), .A2(n3114), .ZN(U3227) );
  INV_X1 U3900 ( .A(n3117), .ZN(n3779) );
  NAND2_X1 U3901 ( .A1(n3779), .A2(n3795), .ZN(n3743) );
  XOR2_X1 U3902 ( .A(n3116), .B(n3743), .Z(n3290) );
  XNOR2_X1 U3903 ( .A(n3118), .B(n3743), .ZN(n3119) );
  NAND2_X1 U3904 ( .A1(n3119), .A2(n4222), .ZN(n3288) );
  AOI22_X1 U3905 ( .A1(n3899), .A2(n4367), .B1(n4366), .B2(n3654), .ZN(n3120)
         );
  OAI211_X1 U3906 ( .C1(n3282), .C2(n4371), .A(n3288), .B(n3120), .ZN(n3121)
         );
  AOI21_X1 U3907 ( .B1(n3290), .B2(n4676), .A(n3121), .ZN(n3126) );
  INV_X1 U3908 ( .A(n3136), .ZN(n3122) );
  AOI21_X1 U3909 ( .B1(n3654), .B2(n3123), .A(n3122), .ZN(n3285) );
  AOI22_X1 U3910 ( .A1(n3285), .A2(n4325), .B1(REG1_REG_5__SCAN_IN), .B2(n4696), .ZN(n3124) );
  OAI21_X1 U3911 ( .B1(n3126), .B2(n4696), .A(n3124), .ZN(U3523) );
  AOI22_X1 U3912 ( .A1(n3285), .A2(n4415), .B1(REG0_REG_5__SCAN_IN), .B2(n4685), .ZN(n3125) );
  OAI21_X1 U3913 ( .B1(n3126), .B2(n4685), .A(n3125), .ZN(U3477) );
  NAND2_X1 U3914 ( .A1(n3782), .A2(n3794), .ZN(n3747) );
  OR2_X1 U3915 ( .A1(n3116), .A2(n3127), .ZN(n3129) );
  NAND2_X1 U3916 ( .A1(n3129), .A2(n3128), .ZN(n3130) );
  XOR2_X1 U3917 ( .A(n3747), .B(n3130), .Z(n3221) );
  NAND2_X1 U3918 ( .A1(n3132), .A2(n3131), .ZN(n3133) );
  NAND2_X1 U3919 ( .A1(n4256), .A2(n3133), .ZN(n4227) );
  XNOR2_X1 U3920 ( .A(n3134), .B(n3747), .ZN(n3135) );
  NOR2_X1 U3921 ( .A1(n3135), .A2(n4242), .ZN(n3218) );
  AND2_X1 U3922 ( .A1(n3136), .A2(n3166), .ZN(n3137) );
  NOR2_X1 U3923 ( .A1(n3205), .A2(n3137), .ZN(n3225) );
  NAND2_X1 U3924 ( .A1(n3225), .A2(n4623), .ZN(n3143) );
  AND2_X1 U3925 ( .A1(n4256), .A2(n4320), .ZN(n4204) );
  OAI22_X1 U3926 ( .A1(n4256), .A2(n3138), .B1(n3169), .B2(n4253), .ZN(n3139)
         );
  AOI21_X1 U3927 ( .B1(n4204), .B2(n3900), .A(n3139), .ZN(n3142) );
  NAND2_X1 U3928 ( .A1(n4256), .A2(n4367), .ZN(n4134) );
  NAND2_X1 U3929 ( .A1(n4256), .A2(n4366), .ZN(n4210) );
  OAI22_X1 U3930 ( .A1(n3321), .A2(n4134), .B1(n4210), .B2(n2289), .ZN(n3140)
         );
  INV_X1 U3931 ( .A(n3140), .ZN(n3141) );
  NAND3_X1 U3932 ( .A1(n3143), .A2(n3142), .A3(n3141), .ZN(n3144) );
  AOI21_X1 U3933 ( .B1(n3218), .B2(n4256), .A(n3144), .ZN(n3145) );
  OAI21_X1 U3934 ( .B1(n3221), .B2(n4227), .A(n3145), .ZN(U3284) );
  NAND2_X1 U3935 ( .A1(n3147), .A2(n3146), .ZN(n3148) );
  NAND2_X1 U3936 ( .A1(n3900), .A2(n3562), .ZN(n3152) );
  NAND2_X1 U3937 ( .A1(n3654), .A2(n3557), .ZN(n3151) );
  NAND2_X1 U3938 ( .A1(n3152), .A2(n3151), .ZN(n3153) );
  XNOR2_X1 U3939 ( .A(n3153), .B(n3570), .ZN(n3158) );
  NOR2_X1 U3940 ( .A1(n3154), .A2(n3572), .ZN(n3155) );
  AOI21_X1 U3941 ( .B1(n3900), .B2(n3561), .A(n3155), .ZN(n3156) );
  XNOR2_X1 U3942 ( .A(n3158), .B(n3156), .ZN(n3651) );
  INV_X1 U3943 ( .A(n3156), .ZN(n3157) );
  NAND2_X1 U3944 ( .A1(n3899), .A2(n3562), .ZN(n3160) );
  NAND2_X1 U3945 ( .A1(n3166), .A2(n3557), .ZN(n3159) );
  NAND2_X1 U3946 ( .A1(n3160), .A2(n3159), .ZN(n3161) );
  XNOR2_X1 U3947 ( .A(n3161), .B(n3570), .ZN(n3229) );
  NAND2_X1 U3948 ( .A1(n3899), .A2(n3561), .ZN(n3163) );
  NAND2_X1 U3949 ( .A1(n3166), .A2(n3562), .ZN(n3162) );
  NAND2_X1 U3950 ( .A1(n3163), .A2(n3162), .ZN(n3230) );
  XNOR2_X1 U3951 ( .A(n3229), .B(n3230), .ZN(n3164) );
  XNOR2_X1 U3952 ( .A(n3231), .B(n3164), .ZN(n3171) );
  AOI21_X1 U3953 ( .B1(n3898), .B2(n4471), .A(n3165), .ZN(n3168) );
  AOI22_X1 U3954 ( .A1(n4481), .A2(n3900), .B1(n4484), .B2(n3166), .ZN(n3167)
         );
  OAI211_X1 U3955 ( .C1(n4488), .C2(n3169), .A(n3168), .B(n3167), .ZN(n3170)
         );
  AOI21_X1 U3956 ( .B1(n3171), .B2(n4479), .A(n3170), .ZN(n3172) );
  INV_X1 U3957 ( .A(n3172), .ZN(U3236) );
  NAND2_X1 U3958 ( .A1(n3174), .A2(n3180), .ZN(n3175) );
  NAND2_X1 U3959 ( .A1(n3173), .A2(n3175), .ZN(n4668) );
  INV_X1 U3960 ( .A(n3176), .ZN(n4665) );
  NAND2_X1 U3961 ( .A1(n3177), .A2(n3182), .ZN(n4663) );
  NAND3_X1 U3962 ( .A1(n4623), .A2(n4665), .A3(n4663), .ZN(n3178) );
  OAI21_X1 U3963 ( .B1(n4253), .B2(n3179), .A(n3178), .ZN(n3190) );
  XNOR2_X1 U3964 ( .A(n3181), .B(n2754), .ZN(n3188) );
  NAND2_X1 U3965 ( .A1(n4668), .A2(n3402), .ZN(n3187) );
  AOI22_X1 U3966 ( .A1(n3901), .A2(n4367), .B1(n4366), .B2(n3182), .ZN(n3183)
         );
  OAI21_X1 U3967 ( .B1(n3184), .B2(n4371), .A(n3183), .ZN(n3185) );
  INV_X1 U3968 ( .A(n3185), .ZN(n3186) );
  OAI211_X1 U3969 ( .C1(n3188), .C2(n4242), .A(n3187), .B(n3186), .ZN(n4666)
         );
  MUX2_X1 U3970 ( .A(n4666), .B(REG2_REG_2__SCAN_IN), .S(n4489), .Z(n3189) );
  AOI211_X1 U3971 ( .C1(n4624), .C2(n4668), .A(n3190), .B(n3189), .ZN(n3191)
         );
  INV_X1 U3972 ( .A(n3191), .ZN(U3288) );
  INV_X1 U3973 ( .A(n3192), .ZN(n3204) );
  INV_X1 U3974 ( .A(n3193), .ZN(n3202) );
  OAI22_X1 U3975 ( .A1(n3282), .A2(n4134), .B1(n4210), .B2(n3194), .ZN(n3201)
         );
  INV_X1 U3976 ( .A(n4204), .ZN(n4150) );
  NAND2_X1 U3977 ( .A1(n3195), .A2(n4623), .ZN(n3198) );
  OAI22_X1 U3978 ( .A1(n4256), .A2(n3929), .B1(REG3_REG_3__SCAN_IN), .B2(n4253), .ZN(n3196) );
  INV_X1 U3979 ( .A(n3196), .ZN(n3197) );
  OAI211_X1 U3980 ( .C1(n3199), .C2(n4150), .A(n3198), .B(n3197), .ZN(n3200)
         );
  AOI211_X1 U3981 ( .C1(n3202), .C2(n4256), .A(n3201), .B(n3200), .ZN(n3203)
         );
  OAI21_X1 U3982 ( .B1(n3204), .B2(n4227), .A(n3203), .ZN(U3287) );
  INV_X1 U3983 ( .A(n3205), .ZN(n3207) );
  INV_X1 U3984 ( .A(n3206), .ZN(n3318) );
  AOI211_X1 U3985 ( .C1(n3237), .C2(n3207), .A(n4679), .B(n3318), .ZN(n4675)
         );
  INV_X1 U3986 ( .A(n3745), .ZN(n3783) );
  XNOR2_X1 U3987 ( .A(n3208), .B(n3783), .ZN(n3209) );
  NAND2_X1 U3988 ( .A1(n3209), .A2(n4222), .ZN(n3211) );
  AOI22_X1 U3989 ( .A1(n3897), .A2(n4367), .B1(n4366), .B2(n3237), .ZN(n3210)
         );
  OAI211_X1 U3990 ( .C1(n3281), .C2(n4371), .A(n3211), .B(n3210), .ZN(n4674)
         );
  AOI21_X1 U3991 ( .B1(n4675), .B2(n3989), .A(n4674), .ZN(n3217) );
  AND2_X1 U3992 ( .A1(n3213), .A2(n3212), .ZN(n3214) );
  XOR2_X1 U3993 ( .A(n3745), .B(n3214), .Z(n4677) );
  OAI22_X1 U3994 ( .A1(n4256), .A2(n3938), .B1(n3240), .B2(n4253), .ZN(n3215)
         );
  AOI21_X1 U3995 ( .B1(n4677), .B2(n4259), .A(n3215), .ZN(n3216) );
  OAI21_X1 U3996 ( .B1(n3217), .B2(n4489), .A(n3216), .ZN(U3283) );
  INV_X1 U3997 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4980) );
  OAI22_X1 U3998 ( .A1(n3321), .A2(n4317), .B1(n4315), .B2(n2289), .ZN(n3219)
         );
  AOI211_X1 U3999 ( .C1(n4320), .C2(n3900), .A(n3219), .B(n3218), .ZN(n3220)
         );
  OAI21_X1 U4000 ( .B1(n4341), .B2(n3221), .A(n3220), .ZN(n3224) );
  NAND2_X1 U4001 ( .A1(n3224), .A2(n4687), .ZN(n3223) );
  NAND2_X1 U4002 ( .A1(n3225), .A2(n4415), .ZN(n3222) );
  OAI211_X1 U4003 ( .C1(n4687), .C2(n4980), .A(n3223), .B(n3222), .ZN(U3479)
         );
  NAND2_X1 U4004 ( .A1(n3224), .A2(n4699), .ZN(n3227) );
  NAND2_X1 U4005 ( .A1(n3225), .A2(n4325), .ZN(n3226) );
  OAI211_X1 U4006 ( .C1(n4699), .C2(n3228), .A(n3227), .B(n3226), .ZN(U3524)
         );
  OAI21_X1 U4007 ( .B1(n3231), .B2(n3230), .A(n3229), .ZN(n3233) );
  NAND2_X1 U4008 ( .A1(n3231), .A2(n3230), .ZN(n3232) );
  NAND2_X1 U4009 ( .A1(n3233), .A2(n3232), .ZN(n3257) );
  OAI22_X1 U4010 ( .A1(n3321), .A2(n3572), .B1(n3569), .B2(n3235), .ZN(n3234)
         );
  XNOR2_X1 U4011 ( .A(n3234), .B(n3552), .ZN(n3258) );
  OAI22_X1 U4012 ( .A1(n3321), .A2(n2984), .B1(n3572), .B2(n3235), .ZN(n3259)
         );
  XNOR2_X1 U4013 ( .A(n3258), .B(n3259), .ZN(n3256) );
  XOR2_X1 U4014 ( .A(n3257), .B(n3256), .Z(n3242) );
  AOI21_X1 U4015 ( .B1(n4471), .B2(n3897), .A(n3236), .ZN(n3239) );
  AOI22_X1 U4016 ( .A1(n4481), .A2(n3899), .B1(n4484), .B2(n3237), .ZN(n3238)
         );
  OAI211_X1 U4017 ( .C1(n4488), .C2(n3240), .A(n3239), .B(n3238), .ZN(n3241)
         );
  AOI21_X1 U4018 ( .B1(n3242), .B2(n4479), .A(n3241), .ZN(n3243) );
  INV_X1 U4019 ( .A(n3243), .ZN(U3210) );
  INV_X1 U4020 ( .A(n3802), .ZN(n3244) );
  NAND2_X1 U4021 ( .A1(n3244), .A2(n3787), .ZN(n3744) );
  XNOR2_X1 U4022 ( .A(n3245), .B(n3744), .ZN(n3246) );
  NAND2_X1 U4023 ( .A1(n3246), .A2(n4222), .ZN(n3308) );
  XNOR2_X1 U4024 ( .A(n3247), .B(n3744), .ZN(n3310) );
  NAND2_X1 U4025 ( .A1(n3310), .A2(n4259), .ZN(n3255) );
  INV_X1 U4026 ( .A(n3317), .ZN(n3249) );
  INV_X1 U4027 ( .A(n3393), .ZN(n3248) );
  OAI21_X1 U4028 ( .B1(n3249), .B2(n3298), .A(n3248), .ZN(n3316) );
  INV_X1 U4029 ( .A(n3316), .ZN(n3253) );
  OAI22_X1 U4030 ( .A1(n3302), .A2(n4253), .B1(n2548), .B2(n4256), .ZN(n3252)
         );
  INV_X1 U4031 ( .A(n4210), .ZN(n4144) );
  INV_X1 U4032 ( .A(n4134), .ZN(n4205) );
  AOI22_X1 U4033 ( .A1(n4144), .A2(n3306), .B1(n4205), .B2(n3895), .ZN(n3250)
         );
  OAI21_X1 U4034 ( .B1(n2375), .B2(n4150), .A(n3250), .ZN(n3251) );
  AOI211_X1 U4035 ( .C1(n3253), .C2(n4623), .A(n3252), .B(n3251), .ZN(n3254)
         );
  OAI211_X1 U4036 ( .C1(n4489), .C2(n3308), .A(n3255), .B(n3254), .ZN(U3281)
         );
  INV_X1 U4037 ( .A(n3258), .ZN(n3260) );
  NAND2_X1 U4038 ( .A1(n3260), .A2(n3259), .ZN(n3261) );
  NAND2_X1 U4039 ( .A1(n3897), .A2(n3562), .ZN(n3263) );
  NAND2_X1 U4040 ( .A1(n3274), .A2(n3557), .ZN(n3262) );
  NAND2_X1 U4041 ( .A1(n3263), .A2(n3262), .ZN(n3264) );
  XNOR2_X1 U4042 ( .A(n3264), .B(n3570), .ZN(n3267) );
  NAND2_X1 U40430 ( .A1(n3897), .A2(n3561), .ZN(n3266) );
  NAND2_X1 U4044 ( .A1(n3274), .A2(n3562), .ZN(n3265) );
  NAND2_X1 U4045 ( .A1(n3266), .A2(n3265), .ZN(n3268) );
  AND2_X1 U4046 ( .A1(n3267), .A2(n3268), .ZN(n3293) );
  INV_X1 U4047 ( .A(n3293), .ZN(n3271) );
  INV_X1 U4048 ( .A(n3267), .ZN(n3270) );
  INV_X1 U4049 ( .A(n3268), .ZN(n3269) );
  NAND2_X1 U4050 ( .A1(n3270), .A2(n3269), .ZN(n3294) );
  NAND2_X1 U4051 ( .A1(n3271), .A2(n3294), .ZN(n3272) );
  XNOR2_X1 U4052 ( .A(n3292), .B(n3272), .ZN(n3279) );
  NAND2_X1 U4053 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4502) );
  INV_X1 U4054 ( .A(n4502), .ZN(n3273) );
  AOI21_X1 U4055 ( .B1(n4471), .B2(n3896), .A(n3273), .ZN(n3276) );
  AOI22_X1 U4056 ( .A1(n3898), .A2(n4481), .B1(n3274), .B2(n4484), .ZN(n3275)
         );
  OAI211_X1 U4057 ( .C1(n4488), .C2(n3277), .A(n3276), .B(n3275), .ZN(n3278)
         );
  AOI21_X1 U4058 ( .B1(n3279), .B2(n4479), .A(n3278), .ZN(n3280) );
  INV_X1 U4059 ( .A(n3280), .ZN(U3218) );
  OAI22_X1 U4060 ( .A1(n4256), .A2(n2885), .B1(n3655), .B2(n4253), .ZN(n3284)
         );
  OAI22_X1 U4061 ( .A1(n4150), .A2(n3282), .B1(n3281), .B2(n4134), .ZN(n3283)
         );
  AOI211_X1 U4062 ( .C1(n3654), .C2(n4144), .A(n3284), .B(n3283), .ZN(n3287)
         );
  NAND2_X1 U4063 ( .A1(n3285), .A2(n4623), .ZN(n3286) );
  OAI211_X1 U4064 ( .C1(n3288), .C2(n4489), .A(n3287), .B(n3286), .ZN(n3289)
         );
  AOI21_X1 U4065 ( .B1(n3290), .B2(n4259), .A(n3289), .ZN(n3291) );
  INV_X1 U4066 ( .A(n3291), .ZN(U3285) );
  NAND2_X1 U4067 ( .A1(n3896), .A2(n3562), .ZN(n3296) );
  NAND2_X1 U4068 ( .A1(n3306), .A2(n3557), .ZN(n3295) );
  NAND2_X1 U4069 ( .A1(n3296), .A2(n3295), .ZN(n3297) );
  XNOR2_X1 U4070 ( .A(n3297), .B(n3570), .ZN(n3349) );
  NOR2_X1 U4071 ( .A1(n3298), .A2(n3572), .ZN(n3299) );
  AOI21_X1 U4072 ( .B1(n3896), .B2(n3561), .A(n3299), .ZN(n3350) );
  XNOR2_X1 U4073 ( .A(n3349), .B(n3350), .ZN(n3347) );
  XNOR2_X1 U4074 ( .A(n3348), .B(n3347), .ZN(n3304) );
  NOR2_X1 U4075 ( .A1(STATE_REG_SCAN_IN), .A2(n2549), .ZN(n4518) );
  AOI21_X1 U4076 ( .B1(n4471), .B2(n3895), .A(n4518), .ZN(n3301) );
  AOI22_X1 U4077 ( .A1(n4481), .A2(n3897), .B1(n4484), .B2(n3306), .ZN(n3300)
         );
  OAI211_X1 U4078 ( .C1(n4488), .C2(n3302), .A(n3301), .B(n3300), .ZN(n3303)
         );
  AOI21_X1 U4079 ( .B1(n3304), .B2(n4479), .A(n3303), .ZN(n3305) );
  INV_X1 U4080 ( .A(n3305), .ZN(U3228) );
  INV_X1 U4081 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4082 ( .A1(n3895), .A2(n4367), .B1(n4366), .B2(n3306), .ZN(n3307)
         );
  OAI211_X1 U4083 ( .C1(n2375), .C2(n4371), .A(n3308), .B(n3307), .ZN(n3309)
         );
  AOI21_X1 U4084 ( .B1(n4676), .B2(n3310), .A(n3309), .ZN(n3313) );
  MUX2_X1 U4085 ( .A(n3311), .B(n3313), .S(n4687), .Z(n3312) );
  OAI21_X1 U4086 ( .B1(n3316), .B2(n4443), .A(n3312), .ZN(U3485) );
  INV_X1 U4087 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3314) );
  MUX2_X1 U4088 ( .A(n3314), .B(n3313), .S(n4699), .Z(n3315) );
  OAI21_X1 U4089 ( .B1(n4377), .B2(n3316), .A(n3315), .ZN(U3527) );
  OAI21_X1 U4090 ( .B1(n3318), .B2(n2376), .A(n3317), .ZN(n4621) );
  INV_X1 U4091 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4092 ( .A1(n3788), .A2(n3785), .ZN(n3741) );
  XOR2_X1 U4093 ( .A(n3741), .B(n3319), .Z(n4625) );
  XOR2_X1 U4094 ( .A(n3320), .B(n3741), .Z(n3324) );
  OAI22_X1 U4095 ( .A1(n3321), .A2(n4371), .B1(n2376), .B2(n4315), .ZN(n3322)
         );
  AOI21_X1 U4096 ( .B1(n4367), .B2(n3896), .A(n3322), .ZN(n3323) );
  OAI21_X1 U4097 ( .B1(n3324), .B2(n4242), .A(n3323), .ZN(n3325) );
  AOI21_X1 U4098 ( .B1(n3402), .B2(n4625), .A(n3325), .ZN(n4628) );
  INV_X1 U4099 ( .A(n4628), .ZN(n3326) );
  AOI21_X1 U4100 ( .B1(n4684), .B2(n4625), .A(n3326), .ZN(n3329) );
  MUX2_X1 U4101 ( .A(n3327), .B(n3329), .S(n4699), .Z(n3328) );
  OAI21_X1 U4102 ( .B1(n4621), .B2(n4377), .A(n3328), .ZN(U3526) );
  INV_X1 U4103 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3330) );
  MUX2_X1 U4104 ( .A(n3330), .B(n3329), .S(n4687), .Z(n3331) );
  OAI21_X1 U4105 ( .B1(n4621), .B2(n4443), .A(n3331), .ZN(U3483) );
  XNOR2_X1 U4106 ( .A(n3419), .B(n3746), .ZN(n3337) );
  XNOR2_X1 U4107 ( .A(n3332), .B(n3746), .ZN(n4683) );
  NAND2_X1 U4108 ( .A1(n4683), .A2(n3402), .ZN(n3336) );
  OAI22_X1 U4109 ( .A1(n3333), .A2(n4317), .B1(n4315), .B2(n3370), .ZN(n3334)
         );
  AOI21_X1 U4110 ( .B1(n4320), .B2(n3895), .A(n3334), .ZN(n3335) );
  OAI211_X1 U4111 ( .C1(n4242), .C2(n3337), .A(n3336), .B(n3335), .ZN(n4681)
         );
  INV_X1 U4112 ( .A(n4681), .ZN(n3342) );
  OAI21_X1 U4113 ( .B1(n3391), .B2(n3370), .A(n3410), .ZN(n4680) );
  NOR2_X1 U4114 ( .A1(n4680), .A2(n4252), .ZN(n3340) );
  OAI22_X1 U4115 ( .A1(n4256), .A2(n3338), .B1(n3375), .B2(n4253), .ZN(n3339)
         );
  AOI211_X1 U4116 ( .C1(n4683), .C2(n4624), .A(n3340), .B(n3339), .ZN(n3341)
         );
  OAI21_X1 U4117 ( .B1(n3342), .B2(n4629), .A(n3341), .ZN(U3279) );
  NAND2_X1 U4118 ( .A1(n3895), .A2(n3562), .ZN(n3344) );
  NAND2_X1 U4119 ( .A1(n3358), .A2(n3557), .ZN(n3343) );
  NAND2_X1 U4120 ( .A1(n3344), .A2(n3343), .ZN(n3345) );
  XNOR2_X1 U4121 ( .A(n3345), .B(n3552), .ZN(n3363) );
  NOR2_X1 U4122 ( .A1(n3396), .A2(n3572), .ZN(n3346) );
  AOI21_X1 U4123 ( .B1(n3895), .B2(n3561), .A(n3346), .ZN(n3364) );
  XNOR2_X1 U4124 ( .A(n3363), .B(n3364), .ZN(n3356) );
  INV_X1 U4125 ( .A(n3349), .ZN(n3351) );
  NAND2_X1 U4126 ( .A1(n3351), .A2(n3350), .ZN(n3352) );
  INV_X1 U4127 ( .A(n3356), .ZN(n3353) );
  INV_X1 U4128 ( .A(n3368), .ZN(n3354) );
  AOI211_X1 U4129 ( .C1(n3356), .C2(n3355), .A(n3679), .B(n3354), .ZN(n3362)
         );
  NAND2_X1 U4130 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4523) );
  INV_X1 U4131 ( .A(n4523), .ZN(n3357) );
  AOI21_X1 U4132 ( .B1(n4481), .B2(n3896), .A(n3357), .ZN(n3360) );
  AOI22_X1 U4133 ( .A1(n3894), .A2(n4471), .B1(n3358), .B2(n4484), .ZN(n3359)
         );
  OAI211_X1 U4134 ( .C1(n4488), .C2(n4611), .A(n3360), .B(n3359), .ZN(n3361)
         );
  OR2_X1 U4135 ( .A1(n3362), .A2(n3361), .ZN(U3214) );
  INV_X1 U4136 ( .A(n3363), .ZN(n3366) );
  INV_X1 U4137 ( .A(n3364), .ZN(n3365) );
  NAND2_X1 U4138 ( .A1(n3366), .A2(n3365), .ZN(n3367) );
  NAND2_X1 U4139 ( .A1(n3368), .A2(n3367), .ZN(n3426) );
  OAI22_X1 U4140 ( .A1(n4372), .A2(n3572), .B1(n3569), .B2(n3370), .ZN(n3369)
         );
  XNOR2_X1 U4141 ( .A(n3369), .B(n3570), .ZN(n3424) );
  OAI22_X1 U4142 ( .A1(n4372), .A2(n2984), .B1(n3572), .B2(n3370), .ZN(n3425)
         );
  XNOR2_X1 U4143 ( .A(n3424), .B(n3425), .ZN(n3371) );
  XNOR2_X1 U4144 ( .A(n3426), .B(n3371), .ZN(n3377) );
  AND2_X1 U4145 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4539) );
  AOI21_X1 U4146 ( .B1(n4481), .B2(n3895), .A(n4539), .ZN(n3374) );
  AOI22_X1 U4147 ( .A1(n4471), .A2(n4246), .B1(n4484), .B2(n3372), .ZN(n3373)
         );
  OAI211_X1 U4148 ( .C1(n4488), .C2(n3375), .A(n3374), .B(n3373), .ZN(n3376)
         );
  AOI21_X1 U4149 ( .B1(n3377), .B2(n4479), .A(n3376), .ZN(n3378) );
  INV_X1 U4150 ( .A(n3378), .ZN(U3233) );
  OAI21_X1 U4151 ( .B1(n3380), .B2(n3733), .A(n3379), .ZN(n4355) );
  OAI21_X1 U4152 ( .B1(n3381), .B2(n3850), .A(n3447), .ZN(n3382) );
  NAND2_X1 U4153 ( .A1(n3382), .A2(n4222), .ZN(n3384) );
  AOI22_X1 U4154 ( .A1(n4217), .A2(n4367), .B1(n4366), .B2(n3600), .ZN(n3383)
         );
  OAI211_X1 U4155 ( .C1(n3385), .C2(n4371), .A(n3384), .B(n3383), .ZN(n3386)
         );
  AOI21_X1 U4156 ( .B1(n4355), .B2(n3402), .A(n3386), .ZN(n4359) );
  INV_X1 U4157 ( .A(n3452), .ZN(n4357) );
  NAND2_X1 U4158 ( .A1(n2262), .A2(n3600), .ZN(n4356) );
  AND3_X1 U4159 ( .A1(n4357), .A2(n4623), .A3(n4356), .ZN(n3389) );
  OAI22_X1 U4160 ( .A1(n4256), .A2(n3387), .B1(n3603), .B2(n4253), .ZN(n3388)
         );
  AOI211_X1 U4161 ( .C1(n4355), .C2(n4624), .A(n3389), .B(n3388), .ZN(n3390)
         );
  OAI21_X1 U4162 ( .B1(n4359), .B2(n4629), .A(n3390), .ZN(U3276) );
  INV_X1 U4163 ( .A(n3391), .ZN(n3392) );
  OAI21_X1 U4164 ( .B1(n3393), .B2(n3396), .A(n3392), .ZN(n4613) );
  INV_X1 U4165 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U4166 ( .A1(n3803), .A2(n3805), .ZN(n3748) );
  XOR2_X1 U4167 ( .A(n3748), .B(n3394), .Z(n4615) );
  XNOR2_X1 U4168 ( .A(n3395), .B(n3748), .ZN(n3400) );
  OAI22_X1 U4169 ( .A1(n3397), .A2(n4371), .B1(n3396), .B2(n4315), .ZN(n3398)
         );
  AOI21_X1 U4170 ( .B1(n4367), .B2(n3894), .A(n3398), .ZN(n3399) );
  OAI21_X1 U4171 ( .B1(n3400), .B2(n4242), .A(n3399), .ZN(n3401) );
  AOI21_X1 U4172 ( .B1(n4615), .B2(n3402), .A(n3401), .ZN(n4618) );
  INV_X1 U4173 ( .A(n4618), .ZN(n3403) );
  AOI21_X1 U4174 ( .B1(n4684), .B2(n4615), .A(n3403), .ZN(n3406) );
  MUX2_X1 U4175 ( .A(n3404), .B(n3406), .S(n4687), .Z(n3405) );
  OAI21_X1 U4176 ( .B1(n4613), .B2(n4443), .A(n3405), .ZN(U3487) );
  INV_X1 U4177 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3407) );
  MUX2_X1 U4178 ( .A(n3407), .B(n3406), .S(n4699), .Z(n3408) );
  OAI21_X1 U4179 ( .B1(n4613), .B2(n4377), .A(n3408), .ZN(U3528) );
  NAND2_X1 U4180 ( .A1(n4239), .A2(n4237), .ZN(n3742) );
  XNOR2_X1 U4181 ( .A(n3409), .B(n3742), .ZN(n4374) );
  NAND2_X1 U4182 ( .A1(n3410), .A2(n4365), .ZN(n3411) );
  NAND2_X1 U4183 ( .A1(n4249), .A2(n3411), .ZN(n4444) );
  OAI22_X1 U4184 ( .A1(n4256), .A2(n3412), .B1(n3443), .B2(n4253), .ZN(n3413)
         );
  AOI21_X1 U4185 ( .B1(n4365), .B2(n4144), .A(n3413), .ZN(n3415) );
  AOI22_X1 U4186 ( .A1(n4205), .A2(n4368), .B1(n3894), .B2(n4204), .ZN(n3414)
         );
  OAI211_X1 U4187 ( .C1(n4444), .C2(n4252), .A(n3415), .B(n3414), .ZN(n3422)
         );
  INV_X1 U4188 ( .A(n3416), .ZN(n3417) );
  AOI21_X1 U4189 ( .B1(n3419), .B2(n3418), .A(n3417), .ZN(n4240) );
  XNOR2_X1 U4190 ( .A(n4240), .B(n3742), .ZN(n3420) );
  NAND2_X1 U4191 ( .A1(n3420), .A2(n4222), .ZN(n4370) );
  NOR2_X1 U4192 ( .A1(n4370), .A2(n4489), .ZN(n3421) );
  AOI211_X1 U4193 ( .C1(n4259), .C2(n4374), .A(n3422), .B(n3421), .ZN(n3423)
         );
  INV_X1 U4194 ( .A(n3423), .ZN(U3278) );
  NAND2_X1 U4195 ( .A1(n3426), .A2(n3425), .ZN(n3427) );
  NAND2_X1 U4196 ( .A1(n3428), .A2(n3427), .ZN(n3478) );
  NAND2_X1 U4197 ( .A1(n4246), .A2(n3562), .ZN(n3430) );
  NAND2_X1 U4198 ( .A1(n4365), .A2(n3557), .ZN(n3429) );
  NAND2_X1 U4199 ( .A1(n3430), .A2(n3429), .ZN(n3431) );
  XNOR2_X1 U4200 ( .A(n3431), .B(n3570), .ZN(n3434) );
  NAND2_X1 U4201 ( .A1(n4246), .A2(n3561), .ZN(n3433) );
  NAND2_X1 U4202 ( .A1(n4365), .A2(n3562), .ZN(n3432) );
  NAND2_X1 U4203 ( .A1(n3433), .A2(n3432), .ZN(n3435) );
  INV_X1 U4204 ( .A(n3477), .ZN(n3438) );
  INV_X1 U4205 ( .A(n3434), .ZN(n3437) );
  INV_X1 U4206 ( .A(n3435), .ZN(n3436) );
  NAND2_X1 U4207 ( .A1(n3437), .A2(n3436), .ZN(n3476) );
  NAND2_X1 U4208 ( .A1(n3438), .A2(n3476), .ZN(n3439) );
  XNOR2_X1 U4209 ( .A(n3478), .B(n3439), .ZN(n3445) );
  NAND2_X1 U4210 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4544) );
  OAI21_X1 U4211 ( .B1(n4372), .B2(n4458), .A(n4544), .ZN(n3440) );
  INV_X1 U4212 ( .A(n3440), .ZN(n3442) );
  AOI22_X1 U4213 ( .A1(n4471), .A2(n4368), .B1(n4484), .B2(n4365), .ZN(n3441)
         );
  OAI211_X1 U4214 ( .C1(n4488), .C2(n3443), .A(n3442), .B(n3441), .ZN(n3444)
         );
  AOI21_X1 U4215 ( .B1(n3445), .B2(n4479), .A(n3444), .ZN(n3446) );
  INV_X1 U4216 ( .A(n3446), .ZN(U3221) );
  NAND2_X1 U4217 ( .A1(n3447), .A2(n3810), .ZN(n3449) );
  INV_X1 U4218 ( .A(n3732), .ZN(n3448) );
  XNOR2_X1 U4219 ( .A(n3449), .B(n3448), .ZN(n3450) );
  NAND2_X1 U4220 ( .A1(n3450), .A2(n4222), .ZN(n4350) );
  XNOR2_X1 U4221 ( .A(n3451), .B(n3732), .ZN(n4353) );
  NAND2_X1 U4222 ( .A1(n4353), .A2(n4259), .ZN(n3460) );
  OAI21_X1 U4223 ( .B1(n3452), .B2(n3456), .A(n4229), .ZN(n4434) );
  INV_X1 U4224 ( .A(n4434), .ZN(n3458) );
  AOI22_X1 U4225 ( .A1(n4205), .A2(n4348), .B1(n3893), .B2(n4204), .ZN(n3455)
         );
  INV_X1 U4226 ( .A(n3726), .ZN(n3453) );
  AOI22_X1 U4227 ( .A1(n4489), .A2(REG2_REG_15__SCAN_IN), .B1(n3453), .B2(
        n4619), .ZN(n3454) );
  OAI211_X1 U4228 ( .C1(n3456), .C2(n4210), .A(n3455), .B(n3454), .ZN(n3457)
         );
  AOI21_X1 U4229 ( .B1(n3458), .B2(n4623), .A(n3457), .ZN(n3459) );
  OAI211_X1 U4230 ( .C1(n4489), .C2(n4350), .A(n3460), .B(n3459), .ZN(U3275)
         );
  INV_X1 U4231 ( .A(n3461), .ZN(n3468) );
  OAI22_X1 U4232 ( .A1(n3583), .A2(n4253), .B1(n3462), .B2(n4256), .ZN(n3464)
         );
  OAI22_X1 U4233 ( .A1(n4035), .A2(n4150), .B1(n3840), .B2(n4134), .ZN(n3463)
         );
  AOI211_X1 U4234 ( .C1(n3580), .C2(n4144), .A(n3464), .B(n3463), .ZN(n3465)
         );
  OAI21_X1 U4235 ( .B1(n3466), .B2(n4252), .A(n3465), .ZN(n3467) );
  AOI21_X1 U4236 ( .B1(n3468), .B2(n4256), .A(n3467), .ZN(n3469) );
  OAI21_X1 U4237 ( .B1(n3470), .B2(n4227), .A(n3469), .ZN(U3262) );
  OAI22_X1 U4238 ( .A1(n4274), .A2(n2984), .B1(n3472), .B2(n3099), .ZN(n3471)
         );
  XNOR2_X1 U4239 ( .A(n3471), .B(n3552), .ZN(n3474) );
  OAI22_X1 U4240 ( .A1(n4274), .A2(n3099), .B1(n3472), .B2(n3569), .ZN(n3473)
         );
  XNOR2_X1 U4241 ( .A(n3474), .B(n3473), .ZN(n3579) );
  INV_X1 U4242 ( .A(n3579), .ZN(n3475) );
  NAND2_X1 U4243 ( .A1(n3475), .A2(n4479), .ZN(n3587) );
  NAND2_X1 U4244 ( .A1(n4368), .A2(n3562), .ZN(n3480) );
  NAND2_X1 U4245 ( .A1(n3694), .A2(n3557), .ZN(n3479) );
  NAND2_X1 U4246 ( .A1(n3480), .A2(n3479), .ZN(n3481) );
  XNOR2_X1 U4247 ( .A(n3481), .B(n3552), .ZN(n3690) );
  NOR2_X1 U4248 ( .A1(n4250), .A2(n3572), .ZN(n3482) );
  AOI21_X1 U4249 ( .B1(n4368), .B2(n3561), .A(n3482), .ZN(n3691) );
  OAI22_X1 U4250 ( .A1(n4351), .A2(n3572), .B1(n3484), .B2(n3569), .ZN(n3483)
         );
  XNOR2_X1 U4251 ( .A(n3483), .B(n3570), .ZN(n3485) );
  OAI22_X1 U4252 ( .A1(n4351), .A2(n2984), .B1(n3484), .B2(n3572), .ZN(n3486)
         );
  NAND2_X1 U4253 ( .A1(n3485), .A2(n3486), .ZN(n3597) );
  INV_X1 U4254 ( .A(n3485), .ZN(n3488) );
  INV_X1 U4255 ( .A(n3486), .ZN(n3487) );
  NAND2_X1 U4256 ( .A1(n3488), .A2(n3487), .ZN(n3596) );
  NAND2_X1 U4257 ( .A1(n4217), .A2(n3562), .ZN(n3490) );
  NAND2_X1 U4258 ( .A1(n4347), .A2(n3557), .ZN(n3489) );
  NAND2_X1 U4259 ( .A1(n3490), .A2(n3489), .ZN(n3491) );
  XNOR2_X1 U4260 ( .A(n3491), .B(n3552), .ZN(n3495) );
  NAND2_X1 U4261 ( .A1(n3492), .A2(n3495), .ZN(n3722) );
  NAND2_X1 U4262 ( .A1(n4217), .A2(n3561), .ZN(n3494) );
  NAND2_X1 U4263 ( .A1(n4347), .A2(n3562), .ZN(n3493) );
  NAND2_X1 U4264 ( .A1(n3494), .A2(n3493), .ZN(n4464) );
  NAND2_X1 U4265 ( .A1(n3722), .A2(n4464), .ZN(n3505) );
  INV_X1 U4266 ( .A(n3495), .ZN(n3496) );
  OAI22_X1 U4267 ( .A1(n4337), .A2(n3572), .B1(n4460), .B2(n3569), .ZN(n3497)
         );
  XNOR2_X1 U4268 ( .A(n3497), .B(n3570), .ZN(n3499) );
  INV_X1 U4269 ( .A(n3499), .ZN(n3501) );
  OAI22_X1 U4270 ( .A1(n4337), .A2(n2984), .B1(n4460), .B2(n3572), .ZN(n3498)
         );
  INV_X1 U4271 ( .A(n3498), .ZN(n3500) );
  OAI21_X1 U4272 ( .B1(n3501), .B2(n3500), .A(n3502), .ZN(n4466) );
  INV_X1 U4273 ( .A(n3502), .ZN(n3503) );
  OAI22_X1 U4274 ( .A1(n4220), .A2(n3572), .B1(n4211), .B2(n3569), .ZN(n3506)
         );
  XNOR2_X1 U4275 ( .A(n3506), .B(n3570), .ZN(n3508) );
  OAI22_X1 U4276 ( .A1(n4220), .A2(n2984), .B1(n4211), .B2(n3572), .ZN(n3507)
         );
  AND2_X1 U4277 ( .A1(n3508), .A2(n3507), .ZN(n3661) );
  OR2_X1 U4278 ( .A1(n3508), .A2(n3507), .ZN(n3662) );
  OAI22_X1 U4279 ( .A1(n4172), .A2(n3572), .B1(n3569), .B2(n4187), .ZN(n3509)
         );
  XNOR2_X1 U4280 ( .A(n3509), .B(n3570), .ZN(n3510) );
  OAI22_X1 U4281 ( .A1(n4172), .A2(n2984), .B1(n3572), .B2(n4187), .ZN(n3511)
         );
  NAND2_X1 U4282 ( .A1(n3510), .A2(n3511), .ZN(n4473) );
  INV_X1 U4283 ( .A(n3510), .ZN(n3513) );
  INV_X1 U4284 ( .A(n3511), .ZN(n3512) );
  NAND2_X1 U4285 ( .A1(n3513), .A2(n3512), .ZN(n4474) );
  OAI22_X1 U4286 ( .A1(n4151), .A2(n2984), .B1(n4173), .B2(n3572), .ZN(n3516)
         );
  OAI22_X1 U4287 ( .A1(n4151), .A2(n3572), .B1(n4173), .B2(n3569), .ZN(n3514)
         );
  XNOR2_X1 U4288 ( .A(n3514), .B(n3570), .ZN(n3515) );
  XOR2_X1 U4289 ( .A(n3516), .B(n3515), .Z(n3618) );
  NAND2_X1 U4290 ( .A1(n3617), .A2(n3618), .ZN(n3616) );
  NAND2_X1 U4291 ( .A1(n3616), .A2(n3519), .ZN(n3625) );
  NAND2_X1 U4292 ( .A1(n4169), .A2(n3562), .ZN(n3521) );
  NAND2_X1 U4293 ( .A1(n4143), .A2(n3557), .ZN(n3520) );
  NAND2_X1 U4294 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  XNOR2_X1 U4295 ( .A(n3522), .B(n3552), .ZN(n3528) );
  INV_X1 U4296 ( .A(n3528), .ZN(n3525) );
  NOR2_X1 U4297 ( .A1(n4316), .A2(n3572), .ZN(n3523) );
  AOI21_X1 U4298 ( .B1(n4169), .B2(n3561), .A(n3523), .ZN(n3527) );
  INV_X1 U4299 ( .A(n3527), .ZN(n3524) );
  NAND2_X1 U4300 ( .A1(n3525), .A2(n3524), .ZN(n3682) );
  NAND2_X1 U4301 ( .A1(n3625), .A2(n3682), .ZN(n3531) );
  OAI22_X1 U4302 ( .A1(n4318), .A2(n3099), .B1(n4133), .B2(n3569), .ZN(n3526)
         );
  XNOR2_X1 U4303 ( .A(n3526), .B(n3570), .ZN(n3628) );
  OAI22_X1 U4304 ( .A1(n4318), .A2(n2984), .B1(n4133), .B2(n3099), .ZN(n3627)
         );
  NAND2_X1 U4305 ( .A1(n3528), .A2(n3527), .ZN(n3681) );
  OAI21_X1 U4306 ( .B1(n3628), .B2(n3627), .A(n3681), .ZN(n3529) );
  AOI21_X2 U4307 ( .B1(n3531), .B2(n3530), .A(n2441), .ZN(n3700) );
  OAI22_X1 U4308 ( .A1(n4135), .A2(n2984), .B1(n4116), .B2(n3572), .ZN(n3538)
         );
  OAI22_X1 U4309 ( .A1(n4135), .A2(n3572), .B1(n4116), .B2(n3569), .ZN(n3532)
         );
  XNOR2_X1 U4310 ( .A(n3532), .B(n3570), .ZN(n3537) );
  XOR2_X1 U4311 ( .A(n3538), .B(n3537), .Z(n3701) );
  NAND2_X1 U4312 ( .A1(n4289), .A2(n3562), .ZN(n3534) );
  NAND2_X1 U4313 ( .A1(n4094), .A2(n3557), .ZN(n3533) );
  NAND2_X1 U4314 ( .A1(n3534), .A2(n3533), .ZN(n3535) );
  XNOR2_X1 U4315 ( .A(n3535), .B(n3570), .ZN(n3542) );
  NOR2_X1 U4316 ( .A1(n4099), .A2(n3572), .ZN(n3536) );
  AOI21_X1 U4317 ( .B1(n4289), .B2(n3561), .A(n3536), .ZN(n3543) );
  XNOR2_X1 U4318 ( .A(n3542), .B(n3543), .ZN(n3608) );
  INV_X1 U4319 ( .A(n3537), .ZN(n3540) );
  INV_X1 U4320 ( .A(n3538), .ZN(n3539) );
  NAND2_X1 U4321 ( .A1(n3540), .A2(n3539), .ZN(n3609) );
  OAI22_X1 U4322 ( .A1(n4097), .A2(n2984), .B1(n4074), .B2(n3572), .ZN(n3548)
         );
  INV_X1 U4323 ( .A(n3548), .ZN(n3546) );
  INV_X1 U4324 ( .A(n3542), .ZN(n3544) );
  NOR2_X1 U4325 ( .A1(n3544), .A2(n3543), .ZN(n3549) );
  INV_X1 U4326 ( .A(n3549), .ZN(n3545) );
  OAI22_X1 U4327 ( .A1(n4097), .A2(n3572), .B1(n4074), .B2(n3569), .ZN(n3547)
         );
  XOR2_X1 U4328 ( .A(n3570), .B(n3547), .Z(n3672) );
  NAND2_X1 U4329 ( .A1(n4037), .A2(n3562), .ZN(n3551) );
  NAND2_X1 U4330 ( .A1(n3642), .A2(n3557), .ZN(n3550) );
  NAND2_X1 U4331 ( .A1(n3551), .A2(n3550), .ZN(n3553) );
  XNOR2_X1 U4332 ( .A(n3553), .B(n3552), .ZN(n3556) );
  NOR2_X1 U4333 ( .A1(n4056), .A2(n3572), .ZN(n3554) );
  AOI21_X1 U4334 ( .B1(n4037), .B2(n3561), .A(n3554), .ZN(n3555) );
  NAND2_X1 U4335 ( .A1(n3556), .A2(n3555), .ZN(n3637) );
  NOR2_X1 U4336 ( .A1(n3556), .A2(n3555), .ZN(n3636) );
  NAND2_X1 U4337 ( .A1(n4271), .A2(n3562), .ZN(n3559) );
  NAND2_X1 U4338 ( .A1(n3713), .A2(n3557), .ZN(n3558) );
  NAND2_X1 U4339 ( .A1(n3559), .A2(n3558), .ZN(n3560) );
  XNOR2_X1 U4340 ( .A(n3560), .B(n3570), .ZN(n3565) );
  NAND2_X1 U4341 ( .A1(n4271), .A2(n3561), .ZN(n3564) );
  NAND2_X1 U4342 ( .A1(n3713), .A2(n3562), .ZN(n3563) );
  NAND2_X1 U4343 ( .A1(n3564), .A2(n3563), .ZN(n3566) );
  NAND2_X1 U4344 ( .A1(n3565), .A2(n3566), .ZN(n3708) );
  INV_X1 U4345 ( .A(n3565), .ZN(n3568) );
  INV_X1 U4346 ( .A(n3566), .ZN(n3567) );
  NAND2_X1 U4347 ( .A1(n3568), .A2(n3567), .ZN(n3709) );
  OAI22_X1 U4348 ( .A1(n4035), .A2(n3099), .B1(n3569), .B2(n4019), .ZN(n3571)
         );
  XNOR2_X1 U4349 ( .A(n3571), .B(n3570), .ZN(n3574) );
  OAI22_X1 U4350 ( .A1(n4035), .A2(n2984), .B1(n3572), .B2(n4019), .ZN(n3573)
         );
  XNOR2_X1 U4351 ( .A(n3574), .B(n3573), .ZN(n3588) );
  NAND2_X1 U4352 ( .A1(n3574), .A2(n3573), .ZN(n3578) );
  INV_X1 U4353 ( .A(n3578), .ZN(n3575) );
  AND2_X1 U4354 ( .A1(n3579), .A2(n3576), .ZN(n3577) );
  NOR3_X1 U4355 ( .A1(n3579), .A2(n3578), .A3(n3679), .ZN(n3585) );
  AOI22_X1 U4356 ( .A1(n3891), .A2(n4481), .B1(n3580), .B2(n4484), .ZN(n3582)
         );
  AOI22_X1 U4357 ( .A1(n3890), .A2(n4471), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3581) );
  OAI211_X1 U4358 ( .C1(n4488), .C2(n3583), .A(n3582), .B(n3581), .ZN(n3584)
         );
  NOR2_X1 U4359 ( .A1(n3585), .A2(n3584), .ZN(n3586) );
  XNOR2_X1 U4360 ( .A(n3589), .B(n3588), .ZN(n3594) );
  NOR2_X1 U4361 ( .A1(n4021), .A2(n4488), .ZN(n3592) );
  AOI22_X1 U4362 ( .A1(n4271), .A2(n4481), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3590) );
  OAI21_X1 U4363 ( .B1(n4461), .B2(n4019), .A(n3590), .ZN(n3591) );
  AOI211_X1 U4364 ( .C1(n4471), .C2(n4005), .A(n3592), .B(n3591), .ZN(n3593)
         );
  OAI21_X1 U4365 ( .B1(n3594), .B2(n3679), .A(n3593), .ZN(U3211) );
  INV_X1 U4366 ( .A(n3595), .ZN(n3599) );
  NAND2_X1 U4367 ( .A1(n3597), .A2(n3596), .ZN(n3598) );
  XNOR2_X1 U4368 ( .A(n3599), .B(n3598), .ZN(n3605) );
  AND2_X1 U4369 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4566) );
  AOI21_X1 U4370 ( .B1(n4471), .B2(n4217), .A(n4566), .ZN(n3602) );
  AOI22_X1 U4371 ( .A1(n4481), .A2(n4368), .B1(n4484), .B2(n3600), .ZN(n3601)
         );
  OAI211_X1 U4372 ( .C1(n4488), .C2(n3603), .A(n3602), .B(n3601), .ZN(n3604)
         );
  AOI21_X1 U4373 ( .B1(n3605), .B2(n4479), .A(n3604), .ZN(n3606) );
  INV_X1 U4374 ( .A(n3606), .ZN(U3212) );
  AOI21_X1 U4375 ( .B1(n3607), .B2(n3609), .A(n3608), .ZN(n3610) );
  NOR3_X1 U4376 ( .A1(n3611), .A2(n3610), .A3(n3679), .ZN(n3615) );
  AOI22_X1 U4377 ( .A1(n3892), .A2(n4471), .B1(n4094), .B2(n4484), .ZN(n3613)
         );
  AOI22_X1 U4378 ( .A1(n4307), .A2(n4481), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3612) );
  OAI211_X1 U4379 ( .C1(n4488), .C2(n4100), .A(n3613), .B(n3612), .ZN(n3614)
         );
  OR2_X1 U4380 ( .A1(n3615), .A2(n3614), .ZN(U3213) );
  OAI21_X1 U4381 ( .B1(n3618), .B2(n3617), .A(n3616), .ZN(n3623) );
  NAND2_X1 U4382 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3988) );
  OAI21_X1 U4383 ( .B1(n4172), .B2(n4458), .A(n3988), .ZN(n3619) );
  INV_X1 U4384 ( .A(n3619), .ZN(n3621) );
  AOI22_X1 U4385 ( .A1(n4471), .A2(n4169), .B1(n4484), .B2(n2661), .ZN(n3620)
         );
  OAI211_X1 U4386 ( .C1(n4488), .C2(n4176), .A(n3621), .B(n3620), .ZN(n3622)
         );
  AOI21_X1 U4387 ( .B1(n3623), .B2(n4479), .A(n3622), .ZN(n3624) );
  INV_X1 U4388 ( .A(n3624), .ZN(U3216) );
  INV_X1 U4389 ( .A(n3681), .ZN(n3626) );
  OAI21_X1 U4390 ( .B1(n3625), .B2(n3626), .A(n3682), .ZN(n3630) );
  XNOR2_X1 U4391 ( .A(n3628), .B(n3627), .ZN(n3629) );
  XNOR2_X1 U4392 ( .A(n3630), .B(n3629), .ZN(n3634) );
  AOI22_X1 U4393 ( .A1(n4307), .A2(n4471), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3632) );
  AOI22_X1 U4394 ( .A1(n4481), .A2(n4169), .B1(n4484), .B2(n4306), .ZN(n3631)
         );
  OAI211_X1 U4395 ( .C1(n4488), .C2(n4130), .A(n3632), .B(n3631), .ZN(n3633)
         );
  AOI21_X1 U4396 ( .B1(n3634), .B2(n4479), .A(n3633), .ZN(n3635) );
  INV_X1 U4397 ( .A(n3635), .ZN(U3220) );
  INV_X1 U4398 ( .A(n3636), .ZN(n3638) );
  NAND2_X1 U4399 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  XNOR2_X1 U4400 ( .A(n3640), .B(n3639), .ZN(n3648) );
  INV_X1 U4401 ( .A(n3641), .ZN(n4059) );
  AOI22_X1 U4402 ( .A1(n4271), .A2(n4471), .B1(n3642), .B2(n4484), .ZN(n3646)
         );
  OAI22_X1 U4403 ( .A1(n4097), .A2(n4458), .B1(STATE_REG_SCAN_IN), .B2(n3643), 
        .ZN(n3644) );
  INV_X1 U4404 ( .A(n3644), .ZN(n3645) );
  OAI211_X1 U4405 ( .C1(n4488), .C2(n4059), .A(n3646), .B(n3645), .ZN(n3647)
         );
  AOI21_X1 U4406 ( .B1(n3648), .B2(n4479), .A(n3647), .ZN(n3649) );
  INV_X1 U4407 ( .A(n3649), .ZN(U3222) );
  OAI211_X1 U4408 ( .C1(n3652), .C2(n3651), .A(n3650), .B(n4479), .ZN(n3659)
         );
  AOI21_X1 U4409 ( .B1(n2502), .B2(n4481), .A(n3653), .ZN(n3658) );
  AOI22_X1 U4410 ( .A1(n4471), .A2(n3899), .B1(n4484), .B2(n3654), .ZN(n3657)
         );
  OR2_X1 U4411 ( .A1(n4488), .A2(n3655), .ZN(n3656) );
  NAND4_X1 U4412 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(U3224)
         );
  INV_X1 U4413 ( .A(n3661), .ZN(n3663) );
  NAND2_X1 U4414 ( .A1(n3663), .A2(n3662), .ZN(n3664) );
  XNOR2_X1 U4415 ( .A(n3660), .B(n3664), .ZN(n3668) );
  NOR2_X1 U4416 ( .A1(STATE_REG_SCAN_IN), .A2(n2632), .ZN(n4593) );
  AOI21_X1 U4417 ( .B1(n4348), .B2(n4481), .A(n4593), .ZN(n3666) );
  AOI22_X1 U4418 ( .A1(n4334), .A2(n4471), .B1(n4333), .B2(n4484), .ZN(n3665)
         );
  OAI211_X1 U4419 ( .C1(n4488), .C2(n4206), .A(n3666), .B(n3665), .ZN(n3667)
         );
  AOI21_X1 U4420 ( .B1(n3668), .B2(n4479), .A(n3667), .ZN(n3669) );
  INV_X1 U4421 ( .A(n3669), .ZN(U3225) );
  NAND2_X1 U4422 ( .A1(n3671), .A2(n3670), .ZN(n3673) );
  XNOR2_X1 U4423 ( .A(n3673), .B(n3672), .ZN(n3680) );
  INV_X1 U4424 ( .A(n3674), .ZN(n4072) );
  NAND2_X1 U4425 ( .A1(n4037), .A2(n4471), .ZN(n3676) );
  AOI22_X1 U4426 ( .A1(n4289), .A2(n4481), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3675) );
  OAI211_X1 U4427 ( .C1(n4461), .C2(n4074), .A(n3676), .B(n3675), .ZN(n3677)
         );
  AOI21_X1 U4428 ( .B1(n4072), .B2(n3712), .A(n3677), .ZN(n3678) );
  OAI21_X1 U4429 ( .B1(n3680), .B2(n3679), .A(n3678), .ZN(U3226) );
  NAND2_X1 U4430 ( .A1(n3682), .A2(n3681), .ZN(n3683) );
  XOR2_X1 U4431 ( .A(n3683), .B(n3625), .Z(n3688) );
  OAI22_X1 U4432 ( .A1(n4151), .A2(n4458), .B1(STATE_REG_SCAN_IN), .B2(n4822), 
        .ZN(n3684) );
  INV_X1 U4433 ( .A(n3684), .ZN(n3686) );
  AOI22_X1 U4434 ( .A1(n4145), .A2(n4471), .B1(n4143), .B2(n4484), .ZN(n3685)
         );
  OAI211_X1 U4435 ( .C1(n4488), .C2(n4146), .A(n3686), .B(n3685), .ZN(n3687)
         );
  AOI21_X1 U4436 ( .B1(n3688), .B2(n4479), .A(n3687), .ZN(n3689) );
  INV_X1 U4437 ( .A(n3689), .ZN(U3230) );
  XOR2_X1 U4438 ( .A(n3691), .B(n3690), .Z(n3692) );
  XNOR2_X1 U4439 ( .A(n3693), .B(n3692), .ZN(n3698) );
  AND2_X1 U4440 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4557) );
  AOI21_X1 U4441 ( .B1(n4481), .B2(n4246), .A(n4557), .ZN(n3696) );
  AOI22_X1 U4442 ( .A1(n3893), .A2(n4471), .B1(n3694), .B2(n4484), .ZN(n3695)
         );
  OAI211_X1 U4443 ( .C1(n4488), .C2(n4254), .A(n3696), .B(n3695), .ZN(n3697)
         );
  AOI21_X1 U4444 ( .B1(n3698), .B2(n4479), .A(n3697), .ZN(n3699) );
  INV_X1 U4445 ( .A(n3699), .ZN(U3231) );
  OAI21_X1 U4446 ( .B1(n3701), .B2(n3700), .A(n3607), .ZN(n3702) );
  NAND2_X1 U4447 ( .A1(n3702), .A2(n4479), .ZN(n3707) );
  NOR2_X1 U4448 ( .A1(n4318), .A2(n4458), .ZN(n3705) );
  OAI22_X1 U4449 ( .A1(n4075), .A2(n3703), .B1(n4461), .B2(n4116), .ZN(n3704)
         );
  AOI211_X1 U4450 ( .C1(REG3_REG_22__SCAN_IN), .C2(U3149), .A(n3705), .B(n3704), .ZN(n3706) );
  OAI211_X1 U4451 ( .C1(n4488), .C2(n4117), .A(n3707), .B(n3706), .ZN(U3232)
         );
  NAND2_X1 U4452 ( .A1(n3709), .A2(n3708), .ZN(n3711) );
  XOR2_X1 U4453 ( .A(n3711), .B(n3710), .Z(n3719) );
  AOI22_X1 U4454 ( .A1(n3891), .A2(n4471), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3717) );
  NAND2_X1 U4455 ( .A1(n3712), .A2(n4043), .ZN(n3716) );
  NAND2_X1 U4456 ( .A1(n4037), .A2(n4481), .ZN(n3715) );
  NAND2_X1 U4457 ( .A1(n4484), .A2(n3713), .ZN(n3714) );
  NAND4_X1 U4458 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3718)
         );
  AOI21_X1 U4459 ( .B1(n3719), .B2(n4479), .A(n3718), .ZN(n3720) );
  INV_X1 U4460 ( .A(n3720), .ZN(U3237) );
  INV_X1 U4461 ( .A(n3721), .ZN(n4463) );
  NAND2_X1 U4462 ( .A1(n4463), .A2(n3722), .ZN(n3723) );
  XNOR2_X1 U4463 ( .A(n3723), .B(n4464), .ZN(n3728) );
  AND2_X1 U4464 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4575) );
  AOI21_X1 U4465 ( .B1(n4348), .B2(n4471), .A(n4575), .ZN(n3725) );
  AOI22_X1 U4466 ( .A1(n3893), .A2(n4481), .B1(n4347), .B2(n4484), .ZN(n3724)
         );
  OAI211_X1 U4467 ( .C1(n4488), .C2(n3726), .A(n3725), .B(n3724), .ZN(n3727)
         );
  AOI21_X1 U4468 ( .B1(n3728), .B2(n4479), .A(n3727), .ZN(n3729) );
  INV_X1 U4469 ( .A(n3729), .ZN(U3238) );
  INV_X1 U4470 ( .A(n4031), .ZN(n3730) );
  NOR2_X1 U4471 ( .A1(n3730), .A2(n3766), .ZN(n4052) );
  NAND2_X1 U4472 ( .A1(n3731), .A2(n3765), .ZN(n4069) );
  NOR4_X1 U4473 ( .A1(n4069), .A2(n3733), .A3(n3732), .A4(n4656), .ZN(n3734)
         );
  NAND3_X1 U4474 ( .A1(n4015), .A2(n4052), .A3(n3734), .ZN(n3736) );
  XNOR2_X1 U4475 ( .A(n4289), .B(n4094), .ZN(n4091) );
  INV_X1 U4476 ( .A(n4091), .ZN(n3735) );
  XNOR2_X1 U4477 ( .A(n4151), .B(n2661), .ZN(n4166) );
  NOR4_X1 U4478 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n4166), .ZN(n3764)
         );
  INV_X1 U4479 ( .A(n3738), .ZN(n4089) );
  OR2_X1 U4480 ( .A1(n4089), .A2(n3819), .ZN(n4088) );
  NOR4_X1 U4481 ( .A1(n3740), .A2(n4088), .A3(n2752), .A4(n3739), .ZN(n3752)
         );
  NOR4_X1 U4482 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3751)
         );
  NOR4_X1 U4483 ( .A1(n2754), .A2(n4190), .A3(n3746), .A4(n3745), .ZN(n3750)
         );
  NOR4_X1 U4484 ( .A1(n4108), .A2(n4225), .A3(n3748), .A4(n3747), .ZN(n3749)
         );
  NAND4_X1 U4485 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3761)
         );
  NAND2_X1 U4486 ( .A1(n2293), .A2(n3753), .ZN(n4033) );
  XNOR2_X1 U4487 ( .A(n4368), .B(n4250), .ZN(n4248) );
  OR2_X1 U4488 ( .A1(n2439), .A2(n3754), .ZN(n4154) );
  INV_X1 U4489 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3998) );
  NAND2_X1 U4490 ( .A1(n2717), .A2(REG1_REG_31__SCAN_IN), .ZN(n3756) );
  NAND2_X1 U4491 ( .A1(n2516), .A2(REG0_REG_31__SCAN_IN), .ZN(n3755) );
  OAI211_X1 U4492 ( .C1(n3757), .C2(n3998), .A(n3756), .B(n3755), .ZN(n3996)
         );
  NAND2_X1 U4493 ( .A1(n2513), .A2(DATAI_31_), .ZN(n3997) );
  NAND2_X1 U4494 ( .A1(n3996), .A2(n3997), .ZN(n3837) );
  NAND2_X1 U4495 ( .A1(n2513), .A2(DATAI_30_), .ZN(n3994) );
  OR2_X1 U4496 ( .A1(n3889), .A2(n3994), .ZN(n3758) );
  NAND2_X1 U4497 ( .A1(n3837), .A2(n3758), .ZN(n3838) );
  NOR2_X1 U4498 ( .A1(n3838), .A2(n3874), .ZN(n3759) );
  AND2_X1 U4499 ( .A1(n4161), .A2(n4082), .ZN(n4201) );
  NAND3_X1 U4500 ( .A1(n4154), .A2(n3759), .A3(n4201), .ZN(n3760) );
  NOR4_X1 U4501 ( .A1(n3761), .A2(n4033), .A3(n4248), .A4(n3760), .ZN(n3762)
         );
  NAND3_X1 U4502 ( .A1(n3764), .A2(n3763), .A3(n3762), .ZN(n3834) );
  NOR2_X1 U4503 ( .A1(n3766), .A2(n2296), .ZN(n3847) );
  INV_X1 U4504 ( .A(n3767), .ZN(n3770) );
  OAI211_X1 U4505 ( .C1(n3770), .C2(n3874), .A(n3769), .B(n3768), .ZN(n3772)
         );
  NAND3_X1 U4506 ( .A1(n3772), .A2(n3771), .A3(n2753), .ZN(n3775) );
  NAND3_X1 U4507 ( .A1(n3775), .A2(n3774), .A3(n3773), .ZN(n3778) );
  NAND3_X1 U4508 ( .A1(n3778), .A2(n3777), .A3(n3776), .ZN(n3781) );
  NAND4_X1 U4509 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3794), .ZN(n3784)
         );
  NAND3_X1 U4510 ( .A1(n3784), .A2(n3783), .A3(n3782), .ZN(n3790) );
  AND2_X1 U4511 ( .A1(n3786), .A2(n3785), .ZN(n3793) );
  INV_X1 U4512 ( .A(n3788), .ZN(n3789) );
  AOI211_X1 U4513 ( .C1(n3790), .C2(n3793), .A(n2304), .B(n3789), .ZN(n3801)
         );
  NAND2_X1 U4514 ( .A1(n3792), .A2(n3791), .ZN(n3800) );
  INV_X1 U4515 ( .A(n3793), .ZN(n3797) );
  INV_X1 U4516 ( .A(n3794), .ZN(n3796) );
  NOR3_X1 U4517 ( .A1(n3797), .A2(n3796), .A3(n3795), .ZN(n3798) );
  NAND2_X1 U4518 ( .A1(n3800), .A2(n3809), .ZN(n3848) );
  OAI21_X1 U4519 ( .B1(n3798), .B2(n2303), .A(n3848), .ZN(n3799) );
  OAI21_X1 U4520 ( .B1(n3801), .B2(n3800), .A(n3799), .ZN(n3807) );
  NAND2_X1 U4521 ( .A1(n3803), .A2(n3802), .ZN(n3804) );
  NAND4_X1 U4522 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3814)
         );
  INV_X1 U4523 ( .A(n3808), .ZN(n3811) );
  NAND2_X1 U4524 ( .A1(n3810), .A2(n3809), .ZN(n3849) );
  OAI21_X1 U4525 ( .B1(n3811), .B2(n3849), .A(n3848), .ZN(n3813) );
  INV_X1 U4526 ( .A(n3812), .ZN(n3851) );
  AOI21_X1 U4527 ( .B1(n3814), .B2(n3813), .A(n3851), .ZN(n3818) );
  INV_X1 U4528 ( .A(n3852), .ZN(n3817) );
  INV_X1 U4529 ( .A(n3815), .ZN(n3816) );
  OAI21_X1 U4530 ( .B1(n3818), .B2(n3817), .A(n3816), .ZN(n3820) );
  AOI211_X1 U4531 ( .C1(n3820), .C2(n4087), .A(n3819), .B(n4086), .ZN(n3821)
         );
  NOR2_X1 U4532 ( .A1(n3821), .A2(n3859), .ZN(n3823) );
  OAI21_X1 U4533 ( .B1(n3823), .B2(n3822), .A(n3863), .ZN(n3824) );
  NAND2_X1 U4534 ( .A1(n3847), .A2(n3824), .ZN(n3830) );
  INV_X1 U4535 ( .A(n3825), .ZN(n3826) );
  OAI21_X1 U4536 ( .B1(n3840), .B2(n3839), .A(n3826), .ZN(n3841) );
  NOR2_X1 U4537 ( .A1(n3827), .A2(n3841), .ZN(n3871) );
  INV_X1 U4538 ( .A(n3871), .ZN(n3828) );
  AOI211_X1 U4539 ( .C1(n3861), .C2(n3830), .A(n3829), .B(n3828), .ZN(n3831)
         );
  INV_X1 U4540 ( .A(n3831), .ZN(n3833) );
  MUX2_X1 U4541 ( .A(n3834), .B(n3833), .S(n3832), .Z(n3881) );
  OR2_X1 U4542 ( .A1(n3996), .A2(n3997), .ZN(n3836) );
  AND2_X1 U4543 ( .A1(n3889), .A2(n3994), .ZN(n3846) );
  INV_X1 U4544 ( .A(n3846), .ZN(n3835) );
  AND2_X1 U4545 ( .A1(n3836), .A2(n3835), .ZN(n3843) );
  INV_X1 U4546 ( .A(n3843), .ZN(n3880) );
  INV_X1 U4547 ( .A(n3837), .ZN(n3844) );
  NOR2_X1 U4548 ( .A1(n3868), .A2(n3867), .ZN(n3842) );
  AOI21_X1 U4549 ( .B1(n3840), .B2(n3839), .A(n3838), .ZN(n3865) );
  OAI21_X1 U4550 ( .B1(n3842), .B2(n3841), .A(n3865), .ZN(n3870) );
  OAI21_X1 U4551 ( .B1(n3844), .B2(n3843), .A(n3870), .ZN(n3878) );
  INV_X1 U4552 ( .A(n3996), .ZN(n3845) );
  NOR2_X1 U4553 ( .A1(n3846), .A2(n3845), .ZN(n3876) );
  INV_X1 U4554 ( .A(n3847), .ZN(n3864) );
  OAI21_X1 U4555 ( .B1(n3850), .B2(n3849), .A(n3848), .ZN(n3853) );
  AOI21_X1 U4556 ( .B1(n3853), .B2(n3852), .A(n3851), .ZN(n3856) );
  INV_X1 U4557 ( .A(n4087), .ZN(n3855) );
  OAI21_X1 U4558 ( .B1(n3856), .B2(n3855), .A(n3854), .ZN(n3857) );
  INV_X1 U4559 ( .A(n3857), .ZN(n3860) );
  OAI21_X1 U4560 ( .B1(n3860), .B2(n3859), .A(n3858), .ZN(n3862) );
  OAI221_X1 U4561 ( .B1(n3864), .B2(n3863), .C1(n3864), .C2(n3862), .A(n3861), 
        .ZN(n3869) );
  INV_X1 U4562 ( .A(n3865), .ZN(n3866) );
  NOR4_X1 U4563 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3873)
         );
  AOI21_X1 U4564 ( .B1(n4015), .B2(n3871), .A(n3870), .ZN(n3872) );
  OAI22_X1 U4565 ( .A1(n3873), .A2(n3872), .B1(n3996), .B2(n3994), .ZN(n3875)
         );
  OAI211_X1 U4566 ( .C1(n3876), .C2(n3997), .A(n3875), .B(n3874), .ZN(n3877)
         );
  MUX2_X1 U4567 ( .A(n3878), .B(n3877), .S(n4448), .Z(n3879) );
  OAI21_X1 U4568 ( .B1(n3881), .B2(n3880), .A(n3879), .ZN(n3882) );
  XNOR2_X1 U4569 ( .A(n3882), .B(n4449), .ZN(n3888) );
  NAND2_X1 U4570 ( .A1(n3884), .A2(n3883), .ZN(n3885) );
  OAI211_X1 U4571 ( .C1(n4447), .C2(n3887), .A(n3885), .B(B_REG_SCAN_IN), .ZN(
        n3886) );
  OAI21_X1 U4572 ( .B1(n3888), .B2(n3887), .A(n3886), .ZN(U3239) );
  MUX2_X1 U4573 ( .A(DATAO_REG_31__SCAN_IN), .B(n3996), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4574 ( .A(DATAO_REG_30__SCAN_IN), .B(n3889), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4575 ( .A(DATAO_REG_29__SCAN_IN), .B(n3890), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4576 ( .A(DATAO_REG_28__SCAN_IN), .B(n4005), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4577 ( .A(DATAO_REG_27__SCAN_IN), .B(n3891), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4578 ( .A(n4271), .B(DATAO_REG_26__SCAN_IN), .S(n3903), .Z(U3576)
         );
  MUX2_X1 U4579 ( .A(n4037), .B(DATAO_REG_25__SCAN_IN), .S(n3903), .Z(U3575)
         );
  MUX2_X1 U4580 ( .A(n3892), .B(DATAO_REG_24__SCAN_IN), .S(n3903), .Z(U3574)
         );
  MUX2_X1 U4581 ( .A(n4289), .B(DATAO_REG_23__SCAN_IN), .S(n3903), .Z(U3573)
         );
  MUX2_X1 U4582 ( .A(n4307), .B(DATAO_REG_22__SCAN_IN), .S(n3903), .Z(U3572)
         );
  MUX2_X1 U4583 ( .A(DATAO_REG_21__SCAN_IN), .B(n4145), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4584 ( .A(n4169), .B(DATAO_REG_20__SCAN_IN), .S(n3903), .Z(U3570)
         );
  MUX2_X1 U4585 ( .A(DATAO_REG_19__SCAN_IN), .B(n4472), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4586 ( .A(DATAO_REG_18__SCAN_IN), .B(n4334), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4587 ( .A(DATAO_REG_17__SCAN_IN), .B(n4482), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4588 ( .A(DATAO_REG_16__SCAN_IN), .B(n4348), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4589 ( .A(n4217), .B(DATAO_REG_15__SCAN_IN), .S(n3903), .Z(U3565)
         );
  MUX2_X1 U4590 ( .A(DATAO_REG_14__SCAN_IN), .B(n3893), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4591 ( .A(n4368), .B(DATAO_REG_13__SCAN_IN), .S(n3903), .Z(U3563)
         );
  MUX2_X1 U4592 ( .A(n4246), .B(DATAO_REG_12__SCAN_IN), .S(n3903), .Z(U3562)
         );
  MUX2_X1 U4593 ( .A(DATAO_REG_11__SCAN_IN), .B(n3894), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4594 ( .A(n3895), .B(DATAO_REG_10__SCAN_IN), .S(n3903), .Z(U3560)
         );
  MUX2_X1 U4595 ( .A(n3896), .B(DATAO_REG_9__SCAN_IN), .S(n3903), .Z(U3559) );
  MUX2_X1 U4596 ( .A(n3897), .B(DATAO_REG_8__SCAN_IN), .S(n3903), .Z(U3558) );
  MUX2_X1 U4597 ( .A(DATAO_REG_7__SCAN_IN), .B(n3898), .S(U4043), .Z(U3557) );
  MUX2_X1 U4598 ( .A(n3899), .B(DATAO_REG_6__SCAN_IN), .S(n3903), .Z(U3556) );
  MUX2_X1 U4599 ( .A(n3900), .B(DATAO_REG_5__SCAN_IN), .S(n3903), .Z(U3555) );
  MUX2_X1 U4600 ( .A(DATAO_REG_4__SCAN_IN), .B(n2502), .S(U4043), .Z(U3554) );
  MUX2_X1 U4601 ( .A(n3901), .B(DATAO_REG_3__SCAN_IN), .S(n3903), .Z(U3553) );
  MUX2_X1 U4602 ( .A(DATAO_REG_2__SCAN_IN), .B(n3902), .S(U4043), .Z(U3552) );
  MUX2_X1 U4603 ( .A(DATAO_REG_1__SCAN_IN), .B(n2291), .S(U4043), .Z(U3551) );
  MUX2_X1 U4604 ( .A(n3035), .B(DATAO_REG_0__SCAN_IN), .S(n3903), .Z(U3550) );
  INV_X1 U4605 ( .A(n4610), .ZN(n3926) );
  NAND2_X1 U4606 ( .A1(n3926), .A2(n4456), .ZN(n3913) );
  OAI211_X1 U4607 ( .C1(n3906), .C2(n3905), .A(n4606), .B(n3904), .ZN(n3912)
         );
  OAI211_X1 U4608 ( .C1(n3909), .C2(n3908), .A(n4552), .B(n3907), .ZN(n3911)
         );
  AOI22_X1 U4609 ( .A1(n4604), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3910) );
  NAND4_X1 U4610 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(U3241)
         );
  AOI22_X1 U4611 ( .A1(n4604), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3914) );
  INV_X1 U4612 ( .A(n3914), .ZN(n3915) );
  AOI21_X1 U4613 ( .B1(n3926), .B2(n4455), .A(n3915), .ZN(n3924) );
  OAI211_X1 U4614 ( .C1(n3918), .C2(n3917), .A(n4552), .B(n3916), .ZN(n3923)
         );
  OAI211_X1 U4615 ( .C1(n3921), .C2(n3920), .A(n4606), .B(n3919), .ZN(n3922)
         );
  NAND4_X1 U4616 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(U3242)
         );
  NAND2_X1 U4617 ( .A1(n3926), .A2(n4454), .ZN(n3935) );
  OAI211_X1 U4618 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3928), .A(n4606), .B(n3927), 
        .ZN(n3934) );
  AOI22_X1 U4619 ( .A1(n4604), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3933) );
  XNOR2_X1 U4620 ( .A(n3930), .B(n3929), .ZN(n3931) );
  NAND2_X1 U4621 ( .A1(n4552), .A2(n3931), .ZN(n3932) );
  NAND4_X1 U4622 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(U3243)
         );
  MUX2_X1 U4623 ( .A(REG2_REG_19__SCAN_IN), .B(n4177), .S(n4449), .Z(n3953) );
  INV_X1 U4624 ( .A(n3954), .ZN(n4643) );
  AOI22_X1 U4625 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4643), .B1(n3954), .B2(
        n4194), .ZN(n4602) );
  NOR2_X1 U4626 ( .A1(n3981), .A2(REG2_REG_17__SCAN_IN), .ZN(n3936) );
  AOI21_X1 U4627 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3981), .A(n3936), .ZN(n4591) );
  INV_X1 U4628 ( .A(n3973), .ZN(n4648) );
  INV_X1 U4629 ( .A(n3958), .ZN(n4649) );
  NOR2_X1 U4630 ( .A1(n4255), .A2(n4649), .ZN(n4551) );
  NAND2_X1 U4631 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3959), .ZN(n3944) );
  INV_X1 U4632 ( .A(n3959), .ZN(n4651) );
  AOI22_X1 U4633 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3959), .B1(n4651), .B2(
        n3338), .ZN(n4535) );
  NAND2_X1 U4634 ( .A1(n3960), .A2(REG2_REG_9__SCAN_IN), .ZN(n3941) );
  INV_X1 U4635 ( .A(n3960), .ZN(n4653) );
  AOI22_X1 U4636 ( .A1(n3960), .A2(REG2_REG_9__SCAN_IN), .B1(n2548), .B2(n4653), .ZN(n4514) );
  NAND2_X1 U4637 ( .A1(n3964), .A2(n3939), .ZN(n3940) );
  NAND2_X1 U4638 ( .A1(n3940), .A2(n4500), .ZN(n4513) );
  NAND2_X1 U4639 ( .A1(n4514), .A2(n4513), .ZN(n4512) );
  NAND2_X1 U4640 ( .A1(n4520), .A2(n3942), .ZN(n3943) );
  NAND2_X1 U4641 ( .A1(n4535), .A2(n4534), .ZN(n4533) );
  NAND2_X1 U4642 ( .A1(n4541), .A2(n3945), .ZN(n3946) );
  NOR2_X1 U4643 ( .A1(n4648), .A2(n3947), .ZN(n3948) );
  NOR2_X1 U4644 ( .A1(n3387), .A2(n4564), .ZN(n4563) );
  NOR2_X1 U4645 ( .A1(n3948), .A2(n4563), .ZN(n4573) );
  NAND2_X1 U4646 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3956), .ZN(n3949) );
  OAI21_X1 U4647 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3956), .A(n3949), .ZN(n4572) );
  NOR2_X1 U4648 ( .A1(n4573), .A2(n4572), .ZN(n4571) );
  AOI21_X1 U4649 ( .B1(n3956), .B2(REG2_REG_15__SCAN_IN), .A(n4571), .ZN(n3950) );
  INV_X1 U4650 ( .A(n3977), .ZN(n4645) );
  NAND2_X1 U4651 ( .A1(n3950), .A2(n4645), .ZN(n3951) );
  XOR2_X1 U4652 ( .A(n3950), .B(n4645), .Z(n4582) );
  NAND2_X1 U4653 ( .A1(n4582), .A2(n4232), .ZN(n4581) );
  NAND2_X1 U4654 ( .A1(n3951), .A2(n4581), .ZN(n4589) );
  NAND2_X1 U4655 ( .A1(n4591), .A2(n4589), .ZN(n4590) );
  AOI21_X1 U4656 ( .B1(n3954), .B2(REG2_REG_18__SCAN_IN), .A(n4601), .ZN(n3952) );
  XOR2_X1 U4657 ( .A(n3953), .B(n3952), .Z(n3993) );
  INV_X1 U4658 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4659 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3954), .B1(n4643), .B2(
        n3983), .ZN(n4607) );
  NOR2_X1 U4660 ( .A1(n3981), .A2(REG1_REG_17__SCAN_IN), .ZN(n3982) );
  NAND2_X1 U4661 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3956), .ZN(n3976) );
  INV_X1 U4662 ( .A(n3956), .ZN(n4646) );
  INV_X1 U4663 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4664 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3956), .B1(n4646), .B2(
        n3955), .ZN(n4578) );
  NAND2_X1 U4665 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3958), .ZN(n3972) );
  INV_X1 U4666 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4667 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3958), .B1(n4649), .B2(
        n3957), .ZN(n4560) );
  INV_X1 U4668 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U4669 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3959), .B1(n4651), .B2(
        n4697), .ZN(n4532) );
  NAND2_X1 U4670 ( .A1(n3960), .A2(REG1_REG_9__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4671 ( .A1(n3960), .A2(REG1_REG_9__SCAN_IN), .B1(n3314), .B2(n4653), .ZN(n4511) );
  NOR2_X1 U4672 ( .A1(n4450), .A2(REG1_REG_7__SCAN_IN), .ZN(n3962) );
  OAI22_X1 U4673 ( .A1(n3963), .A2(n3962), .B1(n4694), .B2(n3961), .ZN(n3965)
         );
  NAND2_X1 U4674 ( .A1(n3965), .A2(n3964), .ZN(n3966) );
  XNOR2_X1 U4675 ( .A(n3965), .B(n2314), .ZN(n4506) );
  NAND2_X1 U4676 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4506), .ZN(n4505) );
  NAND2_X1 U4677 ( .A1(n4520), .A2(n3968), .ZN(n3969) );
  NAND2_X1 U4678 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4527), .ZN(n4526) );
  NAND2_X1 U4679 ( .A1(n4541), .A2(n3970), .ZN(n3971) );
  NAND2_X1 U4680 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4548), .ZN(n4547) );
  NAND2_X1 U4681 ( .A1(n3973), .A2(n3974), .ZN(n3975) );
  NAND2_X1 U4682 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4568), .ZN(n4567) );
  NAND2_X1 U4683 ( .A1(n3975), .A2(n4567), .ZN(n4577) );
  NAND2_X1 U4684 ( .A1(n4578), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U4685 ( .A1(n3976), .A2(n4576), .ZN(n3978) );
  NOR2_X1 U4686 ( .A1(n3977), .A2(n3978), .ZN(n3979) );
  XNOR2_X1 U4687 ( .A(n3978), .B(n3977), .ZN(n4585) );
  NOR2_X1 U4688 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4585), .ZN(n4586) );
  NOR2_X1 U4689 ( .A1(n3979), .A2(n4586), .ZN(n4595) );
  INV_X1 U4690 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4691 ( .A1(n3981), .A2(n3980), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4644), .ZN(n4594) );
  INV_X1 U4692 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3984) );
  MUX2_X1 U4693 ( .A(n3984), .B(REG1_REG_19__SCAN_IN), .S(n4449), .Z(n3985) );
  XNOR2_X1 U4694 ( .A(n3986), .B(n3985), .ZN(n3991) );
  NAND2_X1 U4695 ( .A1(n4604), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3987) );
  OAI211_X1 U4696 ( .C1(n4610), .C2(n3989), .A(n3988), .B(n3987), .ZN(n3990)
         );
  AOI21_X1 U4697 ( .B1(n3991), .B2(n4606), .A(n3990), .ZN(n3992) );
  OAI21_X1 U4698 ( .B1(n3993), .B2(n4600), .A(n3992), .ZN(U3259) );
  INV_X1 U4699 ( .A(n3994), .ZN(n4267) );
  XNOR2_X1 U4700 ( .A(n4263), .B(n3997), .ZN(n4381) );
  NAND2_X1 U4701 ( .A1(n3996), .A2(n3995), .ZN(n4265) );
  OAI21_X1 U4702 ( .B1(n3997), .B2(n4315), .A(n4265), .ZN(n4378) );
  NOR2_X1 U4703 ( .A1(n4256), .A2(n3998), .ZN(n3999) );
  AOI21_X1 U4704 ( .B1(n4256), .B2(n4378), .A(n3999), .ZN(n4000) );
  OAI21_X1 U4705 ( .B1(n4381), .B2(n4252), .A(n4000), .ZN(U3260) );
  INV_X1 U4706 ( .A(n4001), .ZN(n4013) );
  INV_X1 U4707 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4002) );
  OAI22_X1 U4708 ( .A1(n4210), .A2(n4003), .B1(n4002), .B2(n4256), .ZN(n4004)
         );
  AOI21_X1 U4709 ( .B1(n4005), .B2(n4204), .A(n4004), .ZN(n4012) );
  INV_X1 U4710 ( .A(n4006), .ZN(n4010) );
  OAI22_X1 U4711 ( .A1(n4008), .A2(n4252), .B1(n4007), .B2(n4253), .ZN(n4009)
         );
  OAI21_X1 U4712 ( .B1(n4010), .B2(n4009), .A(n4256), .ZN(n4011) );
  OAI211_X1 U4713 ( .C1(n4013), .C2(n4227), .A(n4012), .B(n4011), .ZN(U3354)
         );
  XNOR2_X1 U4714 ( .A(n4014), .B(n4015), .ZN(n4276) );
  INV_X1 U4715 ( .A(n4276), .ZN(n4029) );
  XNOR2_X1 U4716 ( .A(n4016), .B(n4015), .ZN(n4017) );
  NAND2_X1 U4717 ( .A1(n4017), .A2(n4222), .ZN(n4273) );
  INV_X1 U4718 ( .A(n4273), .ZN(n4027) );
  OAI21_X1 U4719 ( .B1(n4040), .B2(n4019), .A(n4018), .ZN(n4388) );
  INV_X1 U4720 ( .A(n4019), .ZN(n4270) );
  OAI22_X1 U4721 ( .A1(n4021), .A2(n4253), .B1(n4020), .B2(n4256), .ZN(n4024)
         );
  OAI22_X1 U4722 ( .A1(n4274), .A2(n4134), .B1(n4022), .B2(n4150), .ZN(n4023)
         );
  AOI211_X1 U4723 ( .C1(n4270), .C2(n4144), .A(n4024), .B(n4023), .ZN(n4025)
         );
  OAI21_X1 U4724 ( .B1(n4388), .B2(n4252), .A(n4025), .ZN(n4026) );
  AOI21_X1 U4725 ( .B1(n4027), .B2(n4256), .A(n4026), .ZN(n4028) );
  OAI21_X1 U4726 ( .B1(n4029), .B2(n4227), .A(n4028), .ZN(U3263) );
  XNOR2_X1 U4727 ( .A(n4030), .B(n4033), .ZN(n4280) );
  INV_X1 U4728 ( .A(n4280), .ZN(n4047) );
  NAND2_X1 U4729 ( .A1(n4032), .A2(n4031), .ZN(n4034) );
  XNOR2_X1 U4730 ( .A(n4034), .B(n4033), .ZN(n4039) );
  OAI22_X1 U4731 ( .A1(n4035), .A2(n4317), .B1(n4315), .B2(n4042), .ZN(n4036)
         );
  AOI21_X1 U4732 ( .B1(n4320), .B2(n4037), .A(n4036), .ZN(n4038) );
  OAI21_X1 U4733 ( .B1(n4039), .B2(n4242), .A(n4038), .ZN(n4279) );
  INV_X1 U4734 ( .A(n4040), .ZN(n4041) );
  OAI21_X1 U4735 ( .B1(n4054), .B2(n4042), .A(n4041), .ZN(n4392) );
  AOI22_X1 U4736 ( .A1(n4043), .A2(n4619), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4489), .ZN(n4044) );
  OAI21_X1 U4737 ( .B1(n4392), .B2(n4252), .A(n4044), .ZN(n4045) );
  AOI21_X1 U4738 ( .B1(n4256), .B2(n4279), .A(n4045), .ZN(n4046) );
  OAI21_X1 U4739 ( .B1(n4047), .B2(n4227), .A(n4046), .ZN(U3264) );
  OAI22_X1 U4740 ( .A1(n4097), .A2(n4371), .B1(n4056), .B2(n4315), .ZN(n4051)
         );
  XNOR2_X1 U4741 ( .A(n4048), .B(n4052), .ZN(n4049) );
  NOR2_X1 U4742 ( .A1(n4049), .A2(n4242), .ZN(n4050) );
  AOI211_X1 U4743 ( .C1(n4367), .C2(n4271), .A(n4051), .B(n4050), .ZN(n4283)
         );
  XNOR2_X1 U4744 ( .A(n4053), .B(n4052), .ZN(n4285) );
  NAND2_X1 U4745 ( .A1(n4285), .A2(n4259), .ZN(n4063) );
  INV_X1 U4746 ( .A(n4070), .ZN(n4057) );
  INV_X1 U4747 ( .A(n4054), .ZN(n4055) );
  OAI21_X1 U4748 ( .B1(n4057), .B2(n4056), .A(n4055), .ZN(n4396) );
  INV_X1 U4749 ( .A(n4396), .ZN(n4061) );
  OAI22_X1 U4750 ( .A1(n4059), .A2(n4253), .B1(n4058), .B2(n4256), .ZN(n4060)
         );
  AOI21_X1 U4751 ( .B1(n4061), .B2(n4623), .A(n4060), .ZN(n4062) );
  OAI211_X1 U4752 ( .C1(n4629), .C2(n4283), .A(n4063), .B(n4062), .ZN(U3265)
         );
  NAND2_X1 U4753 ( .A1(n4065), .A2(n4064), .ZN(n4067) );
  INV_X1 U4754 ( .A(n4069), .ZN(n4066) );
  XNOR2_X1 U4755 ( .A(n4067), .B(n4066), .ZN(n4068) );
  NAND2_X1 U4756 ( .A1(n4068), .A2(n4222), .ZN(n4291) );
  XNOR2_X1 U4757 ( .A(n2253), .B(n4069), .ZN(n4294) );
  NAND2_X1 U4758 ( .A1(n4294), .A2(n4259), .ZN(n4080) );
  INV_X1 U4759 ( .A(n4098), .ZN(n4071) );
  OAI21_X1 U4760 ( .B1(n4071), .B2(n4074), .A(n4070), .ZN(n4400) );
  INV_X1 U4761 ( .A(n4400), .ZN(n4078) );
  AOI22_X1 U4762 ( .A1(n4072), .A2(n4619), .B1(n4489), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n4073) );
  OAI21_X1 U4763 ( .B1(n4074), .B2(n4210), .A(n4073), .ZN(n4077) );
  OAI22_X1 U4764 ( .A1(n4292), .A2(n4134), .B1(n4075), .B2(n4150), .ZN(n4076)
         );
  AOI211_X1 U4765 ( .C1(n4078), .C2(n4623), .A(n4077), .B(n4076), .ZN(n4079)
         );
  OAI211_X1 U4766 ( .C1(n4489), .C2(n4291), .A(n4080), .B(n4079), .ZN(U3266)
         );
  XNOR2_X1 U4767 ( .A(n4081), .B(n4091), .ZN(n4298) );
  INV_X1 U4768 ( .A(n4298), .ZN(n4105) );
  INV_X1 U4769 ( .A(n4082), .ZN(n4083) );
  INV_X1 U4770 ( .A(n4084), .ZN(n4085) );
  AOI21_X1 U4771 ( .B1(n4153), .B2(n4087), .A(n4086), .ZN(n4122) );
  INV_X1 U4772 ( .A(n4088), .ZN(n4125) );
  AOI21_X1 U4773 ( .B1(n4122), .B2(n4125), .A(n4089), .ZN(n4109) );
  OAI21_X1 U4774 ( .B1(n4109), .B2(n4108), .A(n4090), .ZN(n4092) );
  XNOR2_X1 U4775 ( .A(n4092), .B(n4091), .ZN(n4093) );
  NAND2_X1 U4776 ( .A1(n4093), .A2(n4222), .ZN(n4096) );
  AOI22_X1 U4777 ( .A1(n4307), .A2(n4320), .B1(n4366), .B2(n4094), .ZN(n4095)
         );
  OAI211_X1 U4778 ( .C1(n4097), .C2(n4317), .A(n4096), .B(n4095), .ZN(n4297)
         );
  OAI21_X1 U4779 ( .B1(n4114), .B2(n4099), .A(n4098), .ZN(n4404) );
  NOR2_X1 U4780 ( .A1(n4404), .A2(n4252), .ZN(n4103) );
  OAI22_X1 U4781 ( .A1(n4256), .A2(n4101), .B1(n4100), .B2(n4253), .ZN(n4102)
         );
  AOI211_X1 U4782 ( .C1(n4297), .C2(n4256), .A(n4103), .B(n4102), .ZN(n4104)
         );
  OAI21_X1 U4783 ( .B1(n4105), .B2(n4227), .A(n4104), .ZN(U3267) );
  OAI21_X1 U4784 ( .B1(n4107), .B2(n4108), .A(n4106), .ZN(n4301) );
  XNOR2_X1 U4785 ( .A(n4109), .B(n4108), .ZN(n4110) );
  NAND2_X1 U4786 ( .A1(n4110), .A2(n4222), .ZN(n4113) );
  NOR2_X1 U4787 ( .A1(n4116), .A2(n4315), .ZN(n4111) );
  AOI21_X1 U4788 ( .B1(n4289), .B2(n4367), .A(n4111), .ZN(n4112) );
  OAI211_X1 U4789 ( .C1(n4318), .C2(n4371), .A(n4113), .B(n4112), .ZN(n4302)
         );
  INV_X1 U4790 ( .A(n4114), .ZN(n4115) );
  OAI21_X1 U4791 ( .B1(n4128), .B2(n4116), .A(n4115), .ZN(n4408) );
  NOR2_X1 U4792 ( .A1(n4408), .A2(n4252), .ZN(n4120) );
  OAI22_X1 U4793 ( .A1(n4256), .A2(n4118), .B1(n4117), .B2(n4253), .ZN(n4119)
         );
  AOI211_X1 U4794 ( .C1(n4302), .C2(n4256), .A(n4120), .B(n4119), .ZN(n4121)
         );
  OAI21_X1 U4795 ( .B1(n4301), .B2(n4227), .A(n4121), .ZN(U3268) );
  XNOR2_X1 U4796 ( .A(n4122), .B(n4125), .ZN(n4123) );
  NAND2_X1 U4797 ( .A1(n4123), .A2(n4222), .ZN(n4309) );
  INV_X1 U4798 ( .A(n4124), .ZN(n4126) );
  XNOR2_X1 U4799 ( .A(n4126), .B(n4125), .ZN(n4312) );
  NAND2_X1 U4800 ( .A1(n4312), .A2(n4259), .ZN(n4140) );
  INV_X1 U4801 ( .A(n4127), .ZN(n4142) );
  INV_X1 U4802 ( .A(n4128), .ZN(n4129) );
  OAI21_X1 U4803 ( .B1(n4142), .B2(n4133), .A(n4129), .ZN(n4412) );
  INV_X1 U4804 ( .A(n4412), .ZN(n4138) );
  INV_X1 U4805 ( .A(n4130), .ZN(n4131) );
  AOI22_X1 U4806 ( .A1(n4489), .A2(REG2_REG_21__SCAN_IN), .B1(n4131), .B2(
        n4619), .ZN(n4132) );
  OAI21_X1 U4807 ( .B1(n4133), .B2(n4210), .A(n4132), .ZN(n4137) );
  OAI22_X1 U4808 ( .A1(n4310), .A2(n4150), .B1(n4135), .B2(n4134), .ZN(n4136)
         );
  AOI211_X1 U4809 ( .C1(n4138), .C2(n4623), .A(n4137), .B(n4136), .ZN(n4139)
         );
  OAI211_X1 U4810 ( .C1(n4629), .C2(n4309), .A(n4140), .B(n4139), .ZN(U3269)
         );
  XNOR2_X1 U4811 ( .A(n4141), .B(n4154), .ZN(n4323) );
  AOI21_X1 U4812 ( .B1(n4143), .B2(n4175), .A(n4142), .ZN(n4416) );
  AOI22_X1 U4813 ( .A1(n4205), .A2(n4145), .B1(n4144), .B2(n4143), .ZN(n4149)
         );
  INV_X1 U4814 ( .A(n4146), .ZN(n4147) );
  AOI22_X1 U4815 ( .A1(n4489), .A2(REG2_REG_20__SCAN_IN), .B1(n4147), .B2(
        n4619), .ZN(n4148) );
  OAI211_X1 U4816 ( .C1(n4151), .C2(n4150), .A(n4149), .B(n4148), .ZN(n4158)
         );
  NAND2_X1 U4817 ( .A1(n4153), .A2(n4152), .ZN(n4155) );
  XNOR2_X1 U4818 ( .A(n4155), .B(n4154), .ZN(n4156) );
  NAND2_X1 U4819 ( .A1(n4156), .A2(n4222), .ZN(n4321) );
  NOR2_X1 U4820 ( .A1(n4321), .A2(n4489), .ZN(n4157) );
  AOI211_X1 U4821 ( .C1(n4416), .C2(n4623), .A(n4158), .B(n4157), .ZN(n4159)
         );
  OAI21_X1 U4822 ( .B1(n4323), .B2(n4227), .A(n4159), .ZN(U3270) );
  XNOR2_X1 U4823 ( .A(n4160), .B(n4166), .ZN(n4328) );
  INV_X1 U4824 ( .A(n4328), .ZN(n4181) );
  NAND2_X1 U4825 ( .A1(n4162), .A2(n4161), .ZN(n4189) );
  INV_X1 U4826 ( .A(n4163), .ZN(n4165) );
  OAI21_X1 U4827 ( .B1(n4189), .B2(n4165), .A(n4164), .ZN(n4167) );
  XNOR2_X1 U4828 ( .A(n4167), .B(n4166), .ZN(n4168) );
  NAND2_X1 U4829 ( .A1(n4168), .A2(n4222), .ZN(n4171) );
  AOI22_X1 U4830 ( .A1(n4169), .A2(n4367), .B1(n4366), .B2(n2661), .ZN(n4170)
         );
  OAI211_X1 U4831 ( .C1(n4172), .C2(n4371), .A(n4171), .B(n4170), .ZN(n4327)
         );
  OR2_X1 U4832 ( .A1(n4185), .A2(n4173), .ZN(n4174) );
  NAND2_X1 U4833 ( .A1(n4175), .A2(n4174), .ZN(n4421) );
  NOR2_X1 U4834 ( .A1(n4421), .A2(n4252), .ZN(n4179) );
  OAI22_X1 U4835 ( .A1(n4256), .A2(n4177), .B1(n4176), .B2(n4253), .ZN(n4178)
         );
  AOI211_X1 U4836 ( .C1(n4327), .C2(n4256), .A(n4179), .B(n4178), .ZN(n4180)
         );
  OAI21_X1 U4837 ( .B1(n4181), .B2(n4227), .A(n4180), .ZN(U3271) );
  OAI21_X1 U4838 ( .B1(n4183), .B2(n4190), .A(n4182), .ZN(n4184) );
  INV_X1 U4839 ( .A(n4184), .ZN(n4332) );
  INV_X1 U4840 ( .A(n4203), .ZN(n4188) );
  INV_X1 U4841 ( .A(n4185), .ZN(n4186) );
  OAI211_X1 U4842 ( .C1(n4188), .C2(n4187), .A(n4186), .B(n4664), .ZN(n4330)
         );
  XOR2_X1 U4843 ( .A(n4190), .B(n4189), .Z(n4193) );
  AOI22_X1 U4844 ( .A1(n4472), .A2(n4367), .B1(n4483), .B2(n4366), .ZN(n4191)
         );
  OAI21_X1 U4845 ( .B1(n4220), .B2(n4371), .A(n4191), .ZN(n4192) );
  AOI21_X1 U4846 ( .B1(n4193), .B2(n4222), .A(n4192), .ZN(n4331) );
  OAI21_X1 U4847 ( .B1(n4449), .B2(n4330), .A(n4331), .ZN(n4196) );
  OAI22_X1 U4848 ( .A1(n4256), .A2(n4194), .B1(n4487), .B2(n4253), .ZN(n4195)
         );
  AOI21_X1 U4849 ( .B1(n4196), .B2(n4256), .A(n4195), .ZN(n4197) );
  OAI21_X1 U4850 ( .B1(n4332), .B2(n4227), .A(n4197), .ZN(U3272) );
  INV_X1 U4851 ( .A(n4201), .ZN(n4198) );
  XNOR2_X1 U4852 ( .A(n4199), .B(n4198), .ZN(n4200) );
  NAND2_X1 U4853 ( .A1(n4200), .A2(n4222), .ZN(n4336) );
  XNOR2_X1 U4854 ( .A(n4202), .B(n4201), .ZN(n4339) );
  NAND2_X1 U4855 ( .A1(n4339), .A2(n4259), .ZN(n4215) );
  OAI21_X1 U4856 ( .B1(n2287), .B2(n4211), .A(n4203), .ZN(n4426) );
  INV_X1 U4857 ( .A(n4426), .ZN(n4213) );
  AOI22_X1 U4858 ( .A1(n4205), .A2(n4334), .B1(n4348), .B2(n4204), .ZN(n4209)
         );
  INV_X1 U4859 ( .A(n4206), .ZN(n4207) );
  AOI22_X1 U4860 ( .A1(n4489), .A2(REG2_REG_17__SCAN_IN), .B1(n4207), .B2(
        n4619), .ZN(n4208) );
  OAI211_X1 U4861 ( .C1(n4211), .C2(n4210), .A(n4209), .B(n4208), .ZN(n4212)
         );
  AOI21_X1 U4862 ( .B1(n4213), .B2(n4623), .A(n4212), .ZN(n4214) );
  OAI211_X1 U4863 ( .C1(n4629), .C2(n4336), .A(n4215), .B(n4214), .ZN(U3273)
         );
  XNOR2_X1 U4864 ( .A(n4216), .B(n4225), .ZN(n4223) );
  NAND2_X1 U4865 ( .A1(n4228), .A2(n4366), .ZN(n4219) );
  NAND2_X1 U4866 ( .A1(n4217), .A2(n4320), .ZN(n4218) );
  OAI211_X1 U4867 ( .C1(n4220), .C2(n4317), .A(n4219), .B(n4218), .ZN(n4221)
         );
  AOI21_X1 U4868 ( .B1(n4223), .B2(n4222), .A(n4221), .ZN(n4343) );
  OAI21_X1 U4869 ( .B1(n4226), .B2(n4225), .A(n4224), .ZN(n4342) );
  OR2_X1 U4870 ( .A1(n4342), .A2(n4227), .ZN(n4236) );
  NAND2_X1 U4871 ( .A1(n4229), .A2(n4228), .ZN(n4230) );
  NAND2_X1 U4872 ( .A1(n4231), .A2(n4230), .ZN(n4428) );
  INV_X1 U4873 ( .A(n4428), .ZN(n4234) );
  OAI22_X1 U4874 ( .A1(n4256), .A2(n4232), .B1(n4470), .B2(n4253), .ZN(n4233)
         );
  AOI21_X1 U4875 ( .B1(n4234), .B2(n4623), .A(n4233), .ZN(n4235) );
  OAI211_X1 U4876 ( .C1(n4629), .C2(n4343), .A(n4236), .B(n4235), .ZN(U3274)
         );
  OAI22_X1 U4877 ( .A1(n4351), .A2(n4317), .B1(n4315), .B2(n4250), .ZN(n4245)
         );
  INV_X1 U4878 ( .A(n4237), .ZN(n4238) );
  AOI21_X1 U4879 ( .B1(n4240), .B2(n4239), .A(n4238), .ZN(n4241) );
  XNOR2_X1 U4880 ( .A(n4241), .B(n4248), .ZN(n4243) );
  NOR2_X1 U4881 ( .A1(n4243), .A2(n4242), .ZN(n4244) );
  AOI211_X1 U4882 ( .C1(n4320), .C2(n4246), .A(n4245), .B(n4244), .ZN(n4361)
         );
  XOR2_X1 U4883 ( .A(n4248), .B(n4247), .Z(n4363) );
  INV_X1 U4884 ( .A(n4249), .ZN(n4251) );
  OAI21_X1 U4885 ( .B1(n4251), .B2(n4250), .A(n2262), .ZN(n4439) );
  NOR2_X1 U4886 ( .A1(n4439), .A2(n4252), .ZN(n4258) );
  OAI22_X1 U4887 ( .A1(n4256), .A2(n4255), .B1(n4254), .B2(n4253), .ZN(n4257)
         );
  AOI211_X1 U4888 ( .C1(n4363), .C2(n4259), .A(n4258), .B(n4257), .ZN(n4260)
         );
  OAI21_X1 U4889 ( .B1(n4361), .B2(n4489), .A(n4260), .ZN(U3277) );
  NAND2_X1 U4890 ( .A1(n4378), .A2(n4699), .ZN(n4262) );
  NAND2_X1 U4891 ( .A1(n4696), .A2(REG1_REG_31__SCAN_IN), .ZN(n4261) );
  OAI211_X1 U4892 ( .C1(n4381), .C2(n4377), .A(n4262), .B(n4261), .ZN(U3549)
         );
  AOI21_X1 U4893 ( .B1(n4267), .B2(n4264), .A(n4263), .ZN(n4490) );
  INV_X1 U4894 ( .A(n4490), .ZN(n4384) );
  INV_X1 U4895 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4268) );
  INV_X1 U4896 ( .A(n4265), .ZN(n4266) );
  AOI21_X1 U4897 ( .B1(n4267), .B2(n4366), .A(n4266), .ZN(n4492) );
  MUX2_X1 U4898 ( .A(n4268), .B(n4492), .S(n4699), .Z(n4269) );
  OAI21_X1 U4899 ( .B1(n4384), .B2(n4377), .A(n4269), .ZN(U3548) );
  INV_X1 U4900 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U4901 ( .A1(n4271), .A2(n4320), .B1(n4270), .B2(n4366), .ZN(n4272)
         );
  OAI211_X1 U4902 ( .C1(n4274), .C2(n4317), .A(n4273), .B(n4272), .ZN(n4275)
         );
  AOI21_X1 U4903 ( .B1(n4276), .B2(n4676), .A(n4275), .ZN(n4385) );
  MUX2_X1 U4904 ( .A(n4277), .B(n4385), .S(n4699), .Z(n4278) );
  OAI21_X1 U4905 ( .B1(n4377), .B2(n4388), .A(n4278), .ZN(U3545) );
  INV_X1 U4906 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4281) );
  AOI21_X1 U4907 ( .B1(n4280), .B2(n4676), .A(n4279), .ZN(n4389) );
  MUX2_X1 U4908 ( .A(n4281), .B(n4389), .S(n4699), .Z(n4282) );
  OAI21_X1 U4909 ( .B1(n4377), .B2(n4392), .A(n4282), .ZN(U3544) );
  INV_X1 U4910 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4286) );
  INV_X1 U4911 ( .A(n4283), .ZN(n4284) );
  AOI21_X1 U4912 ( .B1(n4285), .B2(n4676), .A(n4284), .ZN(n4393) );
  MUX2_X1 U4913 ( .A(n4286), .B(n4393), .S(n4699), .Z(n4287) );
  OAI21_X1 U4914 ( .B1(n4377), .B2(n4396), .A(n4287), .ZN(U3543) );
  INV_X1 U4915 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U4916 ( .A1(n4289), .A2(n4320), .B1(n4288), .B2(n4366), .ZN(n4290)
         );
  OAI211_X1 U4917 ( .C1(n4292), .C2(n4317), .A(n4291), .B(n4290), .ZN(n4293)
         );
  AOI21_X1 U4918 ( .B1(n4294), .B2(n4676), .A(n4293), .ZN(n4397) );
  MUX2_X1 U4919 ( .A(n4295), .B(n4397), .S(n4699), .Z(n4296) );
  OAI21_X1 U4920 ( .B1(n4377), .B2(n4400), .A(n4296), .ZN(U3542) );
  INV_X1 U4921 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4299) );
  AOI21_X1 U4922 ( .B1(n4298), .B2(n4676), .A(n4297), .ZN(n4401) );
  MUX2_X1 U4923 ( .A(n4299), .B(n4401), .S(n4699), .Z(n4300) );
  OAI21_X1 U4924 ( .B1(n4377), .B2(n4404), .A(n4300), .ZN(U3541) );
  INV_X1 U4925 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4304) );
  INV_X1 U4926 ( .A(n4301), .ZN(n4303) );
  AOI21_X1 U4927 ( .B1(n4303), .B2(n4676), .A(n4302), .ZN(n4405) );
  MUX2_X1 U4928 ( .A(n4304), .B(n4405), .S(n4699), .Z(n4305) );
  OAI21_X1 U4929 ( .B1(n4377), .B2(n4408), .A(n4305), .ZN(U3540) );
  INV_X1 U4930 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4313) );
  AOI22_X1 U4931 ( .A1(n4307), .A2(n4367), .B1(n4366), .B2(n4306), .ZN(n4308)
         );
  OAI211_X1 U4932 ( .C1(n4310), .C2(n4371), .A(n4309), .B(n4308), .ZN(n4311)
         );
  AOI21_X1 U4933 ( .B1(n4312), .B2(n4676), .A(n4311), .ZN(n4409) );
  MUX2_X1 U4934 ( .A(n4313), .B(n4409), .S(n4699), .Z(n4314) );
  OAI21_X1 U4935 ( .B1(n4377), .B2(n4412), .A(n4314), .ZN(U3539) );
  OAI22_X1 U4936 ( .A1(n4318), .A2(n4317), .B1(n4316), .B2(n4315), .ZN(n4319)
         );
  AOI21_X1 U4937 ( .B1(n4320), .B2(n4472), .A(n4319), .ZN(n4322) );
  OAI211_X1 U4938 ( .C1(n4323), .C2(n4341), .A(n4322), .B(n4321), .ZN(n4413)
         );
  MUX2_X1 U4939 ( .A(REG1_REG_20__SCAN_IN), .B(n4413), .S(n4699), .Z(n4324) );
  AOI21_X1 U4940 ( .B1(n4325), .B2(n4416), .A(n4324), .ZN(n4326) );
  INV_X1 U4941 ( .A(n4326), .ZN(U3538) );
  AOI21_X1 U4942 ( .B1(n4328), .B2(n4676), .A(n4327), .ZN(n4418) );
  MUX2_X1 U4943 ( .A(n3984), .B(n4418), .S(n4699), .Z(n4329) );
  OAI21_X1 U4944 ( .B1(n4377), .B2(n4421), .A(n4329), .ZN(U3537) );
  OAI211_X1 U4945 ( .C1(n4332), .C2(n4341), .A(n4331), .B(n4330), .ZN(n4422)
         );
  MUX2_X1 U4946 ( .A(REG1_REG_18__SCAN_IN), .B(n4422), .S(n4699), .Z(U3536) );
  AOI22_X1 U4947 ( .A1(n4334), .A2(n4367), .B1(n4366), .B2(n4333), .ZN(n4335)
         );
  OAI211_X1 U4948 ( .C1(n4337), .C2(n4371), .A(n4336), .B(n4335), .ZN(n4338)
         );
  AOI21_X1 U4949 ( .B1(n4339), .B2(n4676), .A(n4338), .ZN(n4423) );
  MUX2_X1 U4950 ( .A(n3980), .B(n4423), .S(n4699), .Z(n4340) );
  OAI21_X1 U4951 ( .B1(n4377), .B2(n4426), .A(n4340), .ZN(U3535) );
  OR2_X1 U4952 ( .A1(n4342), .A2(n4341), .ZN(n4344) );
  NAND2_X1 U4953 ( .A1(n4344), .A2(n4343), .ZN(n4427) );
  MUX2_X1 U4954 ( .A(REG1_REG_16__SCAN_IN), .B(n4427), .S(n4699), .Z(n4345) );
  INV_X1 U4955 ( .A(n4345), .ZN(n4346) );
  OAI21_X1 U4956 ( .B1(n4377), .B2(n4428), .A(n4346), .ZN(U3534) );
  AOI22_X1 U4957 ( .A1(n4348), .A2(n4367), .B1(n4366), .B2(n4347), .ZN(n4349)
         );
  OAI211_X1 U4958 ( .C1(n4351), .C2(n4371), .A(n4350), .B(n4349), .ZN(n4352)
         );
  AOI21_X1 U4959 ( .B1(n4353), .B2(n4676), .A(n4352), .ZN(n4431) );
  MUX2_X1 U4960 ( .A(n3955), .B(n4431), .S(n4699), .Z(n4354) );
  OAI21_X1 U4961 ( .B1(n4377), .B2(n4434), .A(n4354), .ZN(U3533) );
  INV_X1 U4962 ( .A(n4355), .ZN(n4360) );
  NAND3_X1 U4963 ( .A1(n4357), .A2(n4664), .A3(n4356), .ZN(n4358) );
  OAI211_X1 U4964 ( .C1(n4360), .C2(n4659), .A(n4359), .B(n4358), .ZN(n4435)
         );
  MUX2_X1 U4965 ( .A(REG1_REG_14__SCAN_IN), .B(n4435), .S(n4699), .Z(U3532) );
  INV_X1 U4966 ( .A(n4361), .ZN(n4362) );
  AOI21_X1 U4967 ( .B1(n4363), .B2(n4676), .A(n4362), .ZN(n4436) );
  MUX2_X1 U4968 ( .A(n3957), .B(n4436), .S(n4699), .Z(n4364) );
  OAI21_X1 U4969 ( .B1(n4377), .B2(n4439), .A(n4364), .ZN(U3531) );
  INV_X1 U4970 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U4971 ( .A1(n4368), .A2(n4367), .B1(n4366), .B2(n4365), .ZN(n4369)
         );
  OAI211_X1 U4972 ( .C1(n4372), .C2(n4371), .A(n4370), .B(n4369), .ZN(n4373)
         );
  AOI21_X1 U4973 ( .B1(n4676), .B2(n4374), .A(n4373), .ZN(n4440) );
  MUX2_X1 U4974 ( .A(n4375), .B(n4440), .S(n4699), .Z(n4376) );
  OAI21_X1 U4975 ( .B1(n4444), .B2(n4377), .A(n4376), .ZN(U3530) );
  NAND2_X1 U4976 ( .A1(n4378), .A2(n4687), .ZN(n4380) );
  NAND2_X1 U4977 ( .A1(n4685), .A2(REG0_REG_31__SCAN_IN), .ZN(n4379) );
  OAI211_X1 U4978 ( .C1(n4381), .C2(n4443), .A(n4380), .B(n4379), .ZN(U3517)
         );
  INV_X1 U4979 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4382) );
  MUX2_X1 U4980 ( .A(n4382), .B(n4492), .S(n4687), .Z(n4383) );
  OAI21_X1 U4981 ( .B1(n4384), .B2(n4443), .A(n4383), .ZN(U3516) );
  INV_X1 U4982 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4386) );
  MUX2_X1 U4983 ( .A(n4386), .B(n4385), .S(n4687), .Z(n4387) );
  OAI21_X1 U4984 ( .B1(n4388), .B2(n4443), .A(n4387), .ZN(U3513) );
  INV_X1 U4985 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4390) );
  MUX2_X1 U4986 ( .A(n4390), .B(n4389), .S(n4687), .Z(n4391) );
  OAI21_X1 U4987 ( .B1(n4392), .B2(n4443), .A(n4391), .ZN(U3512) );
  INV_X1 U4988 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4394) );
  MUX2_X1 U4989 ( .A(n4394), .B(n4393), .S(n4687), .Z(n4395) );
  OAI21_X1 U4990 ( .B1(n4396), .B2(n4443), .A(n4395), .ZN(U3511) );
  INV_X1 U4991 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4398) );
  MUX2_X1 U4992 ( .A(n4398), .B(n4397), .S(n4687), .Z(n4399) );
  OAI21_X1 U4993 ( .B1(n4400), .B2(n4443), .A(n4399), .ZN(U3510) );
  INV_X1 U4994 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4402) );
  MUX2_X1 U4995 ( .A(n4402), .B(n4401), .S(n4687), .Z(n4403) );
  OAI21_X1 U4996 ( .B1(n4404), .B2(n4443), .A(n4403), .ZN(U3509) );
  INV_X1 U4997 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4406) );
  MUX2_X1 U4998 ( .A(n4406), .B(n4405), .S(n4687), .Z(n4407) );
  OAI21_X1 U4999 ( .B1(n4408), .B2(n4443), .A(n4407), .ZN(U3508) );
  INV_X1 U5000 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4410) );
  MUX2_X1 U5001 ( .A(n4410), .B(n4409), .S(n4687), .Z(n4411) );
  OAI21_X1 U5002 ( .B1(n4412), .B2(n4443), .A(n4411), .ZN(U3507) );
  MUX2_X1 U5003 ( .A(REG0_REG_20__SCAN_IN), .B(n4413), .S(n4687), .Z(n4414) );
  AOI21_X1 U5004 ( .B1(n4416), .B2(n4415), .A(n4414), .ZN(n4417) );
  INV_X1 U5005 ( .A(n4417), .ZN(U3506) );
  INV_X1 U5006 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4419) );
  MUX2_X1 U5007 ( .A(n4419), .B(n4418), .S(n4687), .Z(n4420) );
  OAI21_X1 U5008 ( .B1(n4421), .B2(n4443), .A(n4420), .ZN(U3505) );
  MUX2_X1 U5009 ( .A(REG0_REG_18__SCAN_IN), .B(n4422), .S(n4687), .Z(U3503) );
  INV_X1 U5010 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4424) );
  MUX2_X1 U5011 ( .A(n4424), .B(n4423), .S(n4687), .Z(n4425) );
  OAI21_X1 U5012 ( .B1(n4426), .B2(n4443), .A(n4425), .ZN(U3501) );
  MUX2_X1 U5013 ( .A(REG0_REG_16__SCAN_IN), .B(n4427), .S(n4687), .Z(n4430) );
  NOR2_X1 U5014 ( .A1(n4428), .A2(n4443), .ZN(n4429) );
  INV_X1 U5015 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4432) );
  MUX2_X1 U5016 ( .A(n4432), .B(n4431), .S(n4687), .Z(n4433) );
  OAI21_X1 U5017 ( .B1(n4434), .B2(n4443), .A(n4433), .ZN(U3497) );
  MUX2_X1 U5018 ( .A(REG0_REG_14__SCAN_IN), .B(n4435), .S(n4687), .Z(U3495) );
  INV_X1 U5019 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4437) );
  MUX2_X1 U5020 ( .A(n4437), .B(n4436), .S(n4687), .Z(n4438) );
  OAI21_X1 U5021 ( .B1(n4439), .B2(n4443), .A(n4438), .ZN(U3493) );
  INV_X1 U5022 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4441) );
  MUX2_X1 U5023 ( .A(n4441), .B(n4440), .S(n4687), .Z(n4442) );
  OAI21_X1 U5024 ( .B1(n4444), .B2(n4443), .A(n4442), .ZN(U3491) );
  MUX2_X1 U5025 ( .A(n4445), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5026 ( .A(n2804), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5027 ( .A(n4446), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5028 ( .A(DATAI_22_), .B(n4447), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5029 ( .A(DATAI_20_), .B(n4448), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5030 ( .A(DATAI_19_), .B(n4449), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5031 ( .A(DATAI_7_), .B(n4450), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5032 ( .A(DATAI_6_), .B(n4451), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U5033 ( .A(DATAI_5_), .B(n4452), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U5034 ( .A(n4453), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U5035 ( .A(n4454), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5036 ( .A(DATAI_2_), .B(n4455), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5037 ( .A(n4456), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5038 ( .A(DATAI_28_), .ZN(n4944) );
  AOI22_X1 U5039 ( .A1(STATE_REG_SCAN_IN), .A2(n4457), .B1(n4944), .B2(U3149), 
        .ZN(U3324) );
  NOR2_X1 U5040 ( .A1(STATE_REG_SCAN_IN), .A2(n5041), .ZN(n4584) );
  OAI22_X1 U5041 ( .A1(n4461), .A2(n4460), .B1(n4459), .B2(n4458), .ZN(n4462)
         );
  AOI211_X1 U5042 ( .C1(n4471), .C2(n4482), .A(n4584), .B(n4462), .ZN(n4469)
         );
  OAI21_X1 U5043 ( .B1(n3721), .B2(n4464), .A(n3722), .ZN(n4465) );
  XOR2_X1 U5044 ( .A(n4466), .B(n4465), .Z(n4467) );
  NAND2_X1 U5045 ( .A1(n4467), .A2(n4479), .ZN(n4468) );
  OAI211_X1 U5046 ( .C1(n4488), .C2(n4470), .A(n4469), .B(n4468), .ZN(U3223)
         );
  AOI22_X1 U5047 ( .A1(n4472), .A2(n4471), .B1(REG3_REG_18__SCAN_IN), .B2(
        U3149), .ZN(n4486) );
  INV_X1 U5048 ( .A(n4474), .ZN(n4477) );
  AND2_X1 U5049 ( .A1(n4474), .A2(n4473), .ZN(n4476) );
  OAI22_X1 U5050 ( .A1(n4478), .A2(n4477), .B1(n4476), .B2(n4475), .ZN(n4480)
         );
  AOI222_X1 U5051 ( .A1(n4484), .A2(n4483), .B1(n4482), .B2(n4481), .C1(n4480), 
        .C2(n4479), .ZN(n4485) );
  OAI211_X1 U5052 ( .C1(n4488), .C2(n4487), .A(n4486), .B(n4485), .ZN(U3235)
         );
  AOI22_X1 U5053 ( .A1(n4490), .A2(n4623), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4489), .ZN(n4491) );
  OAI21_X1 U5054 ( .B1(n4629), .B2(n4492), .A(n4491), .ZN(U3261) );
  OAI211_X1 U5055 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4494), .A(n4493), .B(n4496), 
        .ZN(n4499) );
  AOI22_X1 U5056 ( .A1(n4496), .A2(n4495), .B1(n4606), .B2(n2934), .ZN(n4498)
         );
  AOI22_X1 U5057 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4604), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4497) );
  OAI221_X1 U5058 ( .B1(IR_REG_0__SCAN_IN), .B2(n4499), .C1(n4960), .C2(n4498), 
        .A(n4497), .ZN(U3240) );
  OAI211_X1 U5059 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4501), .A(n4552), .B(n4500), 
        .ZN(n4503) );
  NAND2_X1 U5060 ( .A1(n4503), .A2(n4502), .ZN(n4504) );
  AOI21_X1 U5061 ( .B1(n4604), .B2(ADDR_REG_8__SCAN_IN), .A(n4504), .ZN(n4508)
         );
  OAI211_X1 U5062 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4506), .A(n4606), .B(n4505), 
        .ZN(n4507) );
  OAI211_X1 U5063 ( .C1(n4610), .C2(n2314), .A(n4508), .B(n4507), .ZN(U3248)
         );
  OAI211_X1 U5064 ( .C1(n4511), .C2(n4510), .A(n4606), .B(n4509), .ZN(n4516)
         );
  OAI211_X1 U5065 ( .C1(n4514), .C2(n4513), .A(n4552), .B(n4512), .ZN(n4515)
         );
  OAI211_X1 U5066 ( .C1(n4610), .C2(n4653), .A(n4516), .B(n4515), .ZN(n4517)
         );
  AOI211_X1 U5067 ( .C1(n4604), .C2(ADDR_REG_9__SCAN_IN), .A(n4518), .B(n4517), 
        .ZN(n4519) );
  INV_X1 U5068 ( .A(n4519), .ZN(U3249) );
  OAI211_X1 U5069 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4522), .A(n4552), .B(n4521), .ZN(n4524) );
  NAND2_X1 U5070 ( .A1(n4524), .A2(n4523), .ZN(n4525) );
  AOI21_X1 U5071 ( .B1(n4604), .B2(ADDR_REG_10__SCAN_IN), .A(n4525), .ZN(n4529) );
  OAI211_X1 U5072 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4527), .A(n4606), .B(n4526), .ZN(n4528) );
  OAI211_X1 U5073 ( .C1(n4610), .C2(n2319), .A(n4529), .B(n4528), .ZN(U3250)
         );
  OAI211_X1 U5074 ( .C1(n4532), .C2(n4531), .A(n4606), .B(n4530), .ZN(n4537)
         );
  OAI211_X1 U5075 ( .C1(n4535), .C2(n4534), .A(n4552), .B(n4533), .ZN(n4536)
         );
  OAI211_X1 U5076 ( .C1(n4610), .C2(n4651), .A(n4537), .B(n4536), .ZN(n4538)
         );
  AOI211_X1 U5077 ( .C1(n4604), .C2(ADDR_REG_11__SCAN_IN), .A(n4539), .B(n4538), .ZN(n4540) );
  INV_X1 U5078 ( .A(n4540), .ZN(U3251) );
  OAI211_X1 U5079 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4543), .A(n4552), .B(n4542), .ZN(n4545) );
  NAND2_X1 U5080 ( .A1(n4545), .A2(n4544), .ZN(n4546) );
  AOI21_X1 U5081 ( .B1(n4604), .B2(ADDR_REG_12__SCAN_IN), .A(n4546), .ZN(n4550) );
  OAI211_X1 U5082 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4548), .A(n4606), .B(n4547), .ZN(n4549) );
  OAI211_X1 U5083 ( .C1(n4610), .C2(n2320), .A(n4550), .B(n4549), .ZN(U3252)
         );
  AOI21_X1 U5084 ( .B1(n4255), .B2(n4649), .A(n4551), .ZN(n4555) );
  OAI21_X1 U5085 ( .B1(n4555), .B2(n4554), .A(n4552), .ZN(n4553) );
  AOI21_X1 U5086 ( .B1(n4555), .B2(n4554), .A(n4553), .ZN(n4556) );
  AOI211_X1 U5087 ( .C1(n4604), .C2(ADDR_REG_13__SCAN_IN), .A(n4557), .B(n4556), .ZN(n4562) );
  OAI211_X1 U5088 ( .C1(n4560), .C2(n4559), .A(n4606), .B(n4558), .ZN(n4561)
         );
  OAI211_X1 U5089 ( .C1(n4610), .C2(n4649), .A(n4562), .B(n4561), .ZN(U3253)
         );
  AOI211_X1 U5090 ( .C1(n3387), .C2(n4564), .A(n4563), .B(n4600), .ZN(n4565)
         );
  AOI211_X1 U5091 ( .C1(n4604), .C2(ADDR_REG_14__SCAN_IN), .A(n4566), .B(n4565), .ZN(n4570) );
  OAI211_X1 U5092 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4568), .A(n4606), .B(n4567), .ZN(n4569) );
  OAI211_X1 U5093 ( .C1(n4610), .C2(n4648), .A(n4570), .B(n4569), .ZN(U3254)
         );
  AOI211_X1 U5094 ( .C1(n4573), .C2(n4572), .A(n4571), .B(n4600), .ZN(n4574)
         );
  AOI211_X1 U5095 ( .C1(n4604), .C2(ADDR_REG_15__SCAN_IN), .A(n4575), .B(n4574), .ZN(n4580) );
  OAI211_X1 U5096 ( .C1(n4578), .C2(n4577), .A(n4606), .B(n4576), .ZN(n4579)
         );
  OAI211_X1 U5097 ( .C1(n4610), .C2(n4646), .A(n4580), .B(n4579), .ZN(U3255)
         );
  AOI221_X1 U5098 ( .B1(n4582), .B2(n4581), .C1(n4232), .C2(n4581), .A(n4600), 
        .ZN(n4583) );
  AOI211_X1 U5099 ( .C1(n4604), .C2(ADDR_REG_16__SCAN_IN), .A(n4584), .B(n4583), .ZN(n4588) );
  OAI221_X1 U5100 ( .B1(n4586), .B2(REG1_REG_16__SCAN_IN), .C1(n4586), .C2(
        n4585), .A(n4606), .ZN(n4587) );
  OAI211_X1 U5101 ( .C1(n4610), .C2(n4645), .A(n4588), .B(n4587), .ZN(U3256)
         );
  AOI221_X1 U5102 ( .B1(n4591), .B2(n4590), .C1(n4589), .C2(n4590), .A(n4600), 
        .ZN(n4592) );
  AOI211_X1 U5103 ( .C1(n4604), .C2(ADDR_REG_17__SCAN_IN), .A(n4593), .B(n4592), .ZN(n4598) );
  OAI221_X1 U5104 ( .B1(n4596), .B2(n4595), .C1(n4596), .C2(n4594), .A(n4606), 
        .ZN(n4597) );
  OAI211_X1 U5105 ( .C1(n4610), .C2(n4644), .A(n4598), .B(n4597), .ZN(U3257)
         );
  INV_X1 U5106 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4599) );
  NOR2_X1 U5107 ( .A1(STATE_REG_SCAN_IN), .A2(n4599), .ZN(n4603) );
  OAI211_X1 U5108 ( .C1(n4607), .C2(n2255), .A(n4606), .B(n4605), .ZN(n4608)
         );
  OAI211_X1 U5109 ( .C1(n4610), .C2(n4643), .A(n4609), .B(n4608), .ZN(U3258)
         );
  INV_X1 U5110 ( .A(n4611), .ZN(n4612) );
  AOI22_X1 U5111 ( .A1(n4612), .A2(n4619), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4629), .ZN(n4617) );
  INV_X1 U5112 ( .A(n4613), .ZN(n4614) );
  AOI22_X1 U5113 ( .A1(n4615), .A2(n4624), .B1(n4623), .B2(n4614), .ZN(n4616)
         );
  OAI211_X1 U5114 ( .C1(n4629), .C2(n4618), .A(n4617), .B(n4616), .ZN(U3280)
         );
  AOI22_X1 U5115 ( .A1(n4620), .A2(n4619), .B1(REG2_REG_8__SCAN_IN), .B2(n4629), .ZN(n4627) );
  INV_X1 U5116 ( .A(n4621), .ZN(n4622) );
  AOI22_X1 U5117 ( .A1(n4625), .A2(n4624), .B1(n4623), .B2(n4622), .ZN(n4626)
         );
  OAI211_X1 U5118 ( .C1(n4629), .C2(n4628), .A(n4627), .B(n4626), .ZN(U3282)
         );
  INV_X1 U5119 ( .A(D_REG_31__SCAN_IN), .ZN(n4630) );
  NOR2_X1 U5120 ( .A1(n4640), .A2(n4630), .ZN(U3291) );
  INV_X1 U5121 ( .A(D_REG_30__SCAN_IN), .ZN(n4805) );
  NOR2_X1 U5122 ( .A1(n4640), .A2(n4805), .ZN(U3292) );
  INV_X1 U5123 ( .A(D_REG_29__SCAN_IN), .ZN(n4631) );
  NOR2_X1 U5124 ( .A1(n4640), .A2(n4631), .ZN(U3293) );
  INV_X1 U5125 ( .A(D_REG_28__SCAN_IN), .ZN(n4792) );
  NOR2_X1 U5126 ( .A1(n4640), .A2(n4792), .ZN(U3294) );
  INV_X1 U5127 ( .A(D_REG_27__SCAN_IN), .ZN(n4632) );
  NOR2_X1 U5128 ( .A1(n4640), .A2(n4632), .ZN(U3295) );
  INV_X1 U5129 ( .A(D_REG_26__SCAN_IN), .ZN(n5024) );
  NOR2_X1 U5130 ( .A1(n4640), .A2(n5024), .ZN(U3296) );
  INV_X1 U5131 ( .A(D_REG_25__SCAN_IN), .ZN(n5033) );
  NOR2_X1 U5132 ( .A1(n4640), .A2(n5033), .ZN(U3297) );
  INV_X1 U5133 ( .A(D_REG_24__SCAN_IN), .ZN(n5017) );
  NOR2_X1 U5134 ( .A1(n4640), .A2(n5017), .ZN(U3298) );
  INV_X1 U5135 ( .A(D_REG_23__SCAN_IN), .ZN(n5014) );
  NOR2_X1 U5136 ( .A1(n4640), .A2(n5014), .ZN(U3299) );
  INV_X1 U5137 ( .A(D_REG_22__SCAN_IN), .ZN(n4633) );
  NOR2_X1 U5138 ( .A1(n4640), .A2(n4633), .ZN(U3300) );
  INV_X1 U5139 ( .A(D_REG_21__SCAN_IN), .ZN(n4634) );
  NOR2_X1 U5140 ( .A1(n4640), .A2(n4634), .ZN(U3301) );
  INV_X1 U5141 ( .A(D_REG_20__SCAN_IN), .ZN(n5027) );
  NOR2_X1 U5142 ( .A1(n4640), .A2(n5027), .ZN(U3302) );
  INV_X1 U5143 ( .A(D_REG_19__SCAN_IN), .ZN(n5026) );
  NOR2_X1 U5144 ( .A1(n4640), .A2(n5026), .ZN(U3303) );
  INV_X1 U5145 ( .A(D_REG_18__SCAN_IN), .ZN(n5011) );
  NOR2_X1 U5146 ( .A1(n4640), .A2(n5011), .ZN(U3304) );
  INV_X1 U5147 ( .A(D_REG_17__SCAN_IN), .ZN(n4635) );
  NOR2_X1 U5148 ( .A1(n4640), .A2(n4635), .ZN(U3305) );
  INV_X1 U5149 ( .A(D_REG_16__SCAN_IN), .ZN(n4636) );
  NOR2_X1 U5150 ( .A1(n4640), .A2(n4636), .ZN(U3306) );
  INV_X1 U5151 ( .A(D_REG_15__SCAN_IN), .ZN(n4637) );
  NOR2_X1 U5152 ( .A1(n4640), .A2(n4637), .ZN(U3307) );
  INV_X1 U5153 ( .A(D_REG_14__SCAN_IN), .ZN(n4783) );
  NOR2_X1 U5154 ( .A1(n4640), .A2(n4783), .ZN(U3308) );
  INV_X1 U5155 ( .A(D_REG_13__SCAN_IN), .ZN(n5029) );
  NOR2_X1 U5156 ( .A1(n4640), .A2(n5029), .ZN(U3309) );
  INV_X1 U5157 ( .A(D_REG_12__SCAN_IN), .ZN(n5032) );
  NOR2_X1 U5158 ( .A1(n4640), .A2(n5032), .ZN(U3310) );
  INV_X1 U5159 ( .A(D_REG_11__SCAN_IN), .ZN(n5016) );
  NOR2_X1 U5160 ( .A1(n4640), .A2(n5016), .ZN(U3311) );
  INV_X1 U5161 ( .A(D_REG_10__SCAN_IN), .ZN(n5007) );
  NOR2_X1 U5162 ( .A1(n4640), .A2(n5007), .ZN(U3312) );
  INV_X1 U5163 ( .A(D_REG_9__SCAN_IN), .ZN(n5008) );
  NOR2_X1 U5164 ( .A1(n4640), .A2(n5008), .ZN(U3313) );
  INV_X1 U5165 ( .A(D_REG_8__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U5166 ( .A1(n4640), .A2(n4638), .ZN(U3314) );
  INV_X1 U5167 ( .A(D_REG_7__SCAN_IN), .ZN(n4639) );
  NOR2_X1 U5168 ( .A1(n4640), .A2(n4639), .ZN(U3315) );
  INV_X1 U5169 ( .A(D_REG_6__SCAN_IN), .ZN(n4780) );
  NOR2_X1 U5170 ( .A1(n4640), .A2(n4780), .ZN(U3316) );
  INV_X1 U5171 ( .A(D_REG_5__SCAN_IN), .ZN(n5023) );
  NOR2_X1 U5172 ( .A1(n4640), .A2(n5023), .ZN(U3317) );
  INV_X1 U5173 ( .A(D_REG_4__SCAN_IN), .ZN(n5030) );
  NOR2_X1 U5174 ( .A1(n4640), .A2(n5030), .ZN(U3318) );
  INV_X1 U5175 ( .A(D_REG_3__SCAN_IN), .ZN(n5010) );
  NOR2_X1 U5176 ( .A1(n4640), .A2(n5010), .ZN(U3319) );
  INV_X1 U5177 ( .A(D_REG_2__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U5178 ( .A1(n4640), .A2(n5013), .ZN(U3320) );
  INV_X1 U5179 ( .A(DATAI_23_), .ZN(n4946) );
  AOI21_X1 U5180 ( .B1(U3149), .B2(n4946), .A(n4641), .ZN(U3329) );
  INV_X1 U5181 ( .A(DATAI_18_), .ZN(n4642) );
  AOI22_X1 U5182 ( .A1(STATE_REG_SCAN_IN), .A2(n4643), .B1(n4642), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5183 ( .A1(STATE_REG_SCAN_IN), .A2(n4644), .B1(n2642), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5184 ( .A(DATAI_16_), .ZN(n5039) );
  AOI22_X1 U5185 ( .A1(STATE_REG_SCAN_IN), .A2(n4645), .B1(n5039), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5186 ( .A(DATAI_15_), .ZN(n4956) );
  AOI22_X1 U5187 ( .A1(STATE_REG_SCAN_IN), .A2(n4646), .B1(n4956), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5188 ( .A(DATAI_14_), .ZN(n4647) );
  AOI22_X1 U5189 ( .A1(STATE_REG_SCAN_IN), .A2(n4648), .B1(n4647), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5190 ( .A(DATAI_13_), .ZN(n4808) );
  AOI22_X1 U5191 ( .A1(STATE_REG_SCAN_IN), .A2(n4649), .B1(n4808), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5192 ( .A(DATAI_12_), .ZN(n4650) );
  AOI22_X1 U5193 ( .A1(STATE_REG_SCAN_IN), .A2(n2320), .B1(n4650), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5194 ( .A(DATAI_11_), .ZN(n4995) );
  AOI22_X1 U5195 ( .A1(STATE_REG_SCAN_IN), .A2(n4651), .B1(n4995), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5196 ( .A(DATAI_10_), .ZN(n4807) );
  AOI22_X1 U5197 ( .A1(STATE_REG_SCAN_IN), .A2(n2319), .B1(n4807), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5198 ( .A(DATAI_9_), .ZN(n4652) );
  AOI22_X1 U5199 ( .A1(STATE_REG_SCAN_IN), .A2(n4653), .B1(n4652), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5200 ( .A(DATAI_8_), .ZN(n4998) );
  AOI22_X1 U5201 ( .A1(STATE_REG_SCAN_IN), .A2(n2314), .B1(n4998), .B2(U3149), 
        .ZN(U3344) );
  AOI211_X1 U5202 ( .C1(n4684), .C2(n4656), .A(n4655), .B(n4654), .ZN(n4688)
         );
  INV_X1 U5203 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5204 ( .A1(n4687), .A2(n4688), .B1(n4657), .B2(n4685), .ZN(U3467)
         );
  OAI22_X1 U5205 ( .A1(n4660), .A2(n4659), .B1(n4679), .B2(n4658), .ZN(n4661)
         );
  NOR2_X1 U5206 ( .A1(n4662), .A2(n4661), .ZN(n4689) );
  INV_X1 U5207 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4782) );
  AOI22_X1 U5208 ( .A1(n4687), .A2(n4689), .B1(n4782), .B2(n4685), .ZN(U3469)
         );
  AND3_X1 U5209 ( .A1(n4665), .A2(n4664), .A3(n4663), .ZN(n4667) );
  AOI211_X1 U5210 ( .C1(n4684), .C2(n4668), .A(n4667), .B(n4666), .ZN(n4691)
         );
  INV_X1 U5211 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5045) );
  AOI22_X1 U5212 ( .A1(n4687), .A2(n4691), .B1(n5045), .B2(n4685), .ZN(U3471)
         );
  INV_X1 U5213 ( .A(n4669), .ZN(n4671) );
  AOI211_X1 U5214 ( .C1(n4672), .C2(n4684), .A(n4671), .B(n4670), .ZN(n4693)
         );
  INV_X1 U5215 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5216 ( .A1(n4687), .A2(n4693), .B1(n4673), .B2(n4685), .ZN(U3475)
         );
  AOI211_X1 U5217 ( .C1(n4677), .C2(n4676), .A(n4675), .B(n4674), .ZN(n4695)
         );
  INV_X1 U5218 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5219 ( .A1(n4687), .A2(n4695), .B1(n4678), .B2(n4685), .ZN(U3481)
         );
  NOR2_X1 U5220 ( .A1(n4680), .A2(n4679), .ZN(n4682) );
  AOI211_X1 U5221 ( .C1(n4684), .C2(n4683), .A(n4682), .B(n4681), .ZN(n4698)
         );
  INV_X1 U5222 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U5223 ( .A1(n4687), .A2(n4698), .B1(n4686), .B2(n4685), .ZN(U3489)
         );
  AOI22_X1 U5224 ( .A1(n4699), .A2(n4688), .B1(n2934), .B2(n4696), .ZN(U3518)
         );
  AOI22_X1 U5225 ( .A1(n4699), .A2(n4689), .B1(n2464), .B2(n4696), .ZN(U3519)
         );
  AOI22_X1 U5226 ( .A1(n4699), .A2(n4691), .B1(n4690), .B2(n4696), .ZN(U3520)
         );
  AOI22_X1 U5227 ( .A1(n4699), .A2(n4693), .B1(n4692), .B2(n4696), .ZN(U3522)
         );
  AOI22_X1 U5228 ( .A1(n4699), .A2(n4695), .B1(n4694), .B2(n4696), .ZN(U3525)
         );
  AOI22_X1 U5229 ( .A1(n4699), .A2(n4698), .B1(n4697), .B2(n4696), .ZN(U3529)
         );
  OAI22_X1 U5230 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput_g81), .B1(
        keyinput_g84), .B2(IR_REG_29__SCAN_IN), .ZN(n4700) );
  AOI221_X1 U5231 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput_g81), .C1(
        IR_REG_29__SCAN_IN), .C2(keyinput_g84), .A(n4700), .ZN(n4707) );
  OAI22_X1 U5232 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput_g95), .B1(keyinput_g11), 
        .B2(DATAI_20_), .ZN(n4701) );
  AOI221_X1 U5233 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput_g95), .C1(DATAI_20_), 
        .C2(keyinput_g11), .A(n4701), .ZN(n4706) );
  OAI22_X1 U5234 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_g85), .B1(
        REG0_REG_8__SCAN_IN), .B2(keyinput_g127), .ZN(n4702) );
  AOI221_X1 U5235 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_g85), .C1(
        keyinput_g127), .C2(REG0_REG_8__SCAN_IN), .A(n4702), .ZN(n4705) );
  OAI22_X1 U5236 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput_g75), .B1(
        keyinput_g56), .B2(IR_REG_1__SCAN_IN), .ZN(n4703) );
  AOI221_X1 U5237 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput_g75), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput_g56), .A(n4703), .ZN(n4704) );
  NAND4_X1 U5238 ( .A1(n4707), .A2(n4706), .A3(n4705), .A4(n4704), .ZN(n4735)
         );
  OAI22_X1 U5239 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput_g79), .B1(
        keyinput_g112), .B2(D_REG_25__SCAN_IN), .ZN(n4708) );
  AOI221_X1 U5240 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput_g79), .C1(
        D_REG_25__SCAN_IN), .C2(keyinput_g112), .A(n4708), .ZN(n4715) );
  OAI22_X1 U5241 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_g45), .B1(DATAI_28_), .B2(keyinput_g3), .ZN(n4709) );
  AOI221_X1 U5242 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_g45), .C1(
        keyinput_g3), .C2(DATAI_28_), .A(n4709), .ZN(n4714) );
  OAI22_X1 U5243 ( .A1(DATAI_27_), .A2(keyinput_g4), .B1(DATAI_26_), .B2(
        keyinput_g5), .ZN(n4710) );
  AOI221_X1 U5244 ( .B1(DATAI_27_), .B2(keyinput_g4), .C1(keyinput_g5), .C2(
        DATAI_26_), .A(n4710), .ZN(n4713) );
  OAI22_X1 U5245 ( .A1(DATAI_23_), .A2(keyinput_g8), .B1(DATAI_19_), .B2(
        keyinput_g12), .ZN(n4711) );
  AOI221_X1 U5246 ( .B1(DATAI_23_), .B2(keyinput_g8), .C1(keyinput_g12), .C2(
        DATAI_19_), .A(n4711), .ZN(n4712) );
  NAND4_X1 U5247 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4734)
         );
  OAI22_X1 U5248 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_g54), .B1(
        keyinput_g13), .B2(DATAI_18_), .ZN(n4716) );
  AOI221_X1 U5249 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_g54), .C1(
        DATAI_18_), .C2(keyinput_g13), .A(n4716), .ZN(n4723) );
  OAI22_X1 U5250 ( .A1(D_REG_29__SCAN_IN), .A2(keyinput_g116), .B1(
        D_REG_21__SCAN_IN), .B2(keyinput_g108), .ZN(n4717) );
  AOI221_X1 U5251 ( .B1(D_REG_29__SCAN_IN), .B2(keyinput_g116), .C1(
        keyinput_g108), .C2(D_REG_21__SCAN_IN), .A(n4717), .ZN(n4722) );
  OAI22_X1 U5252 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput_g86), .B1(
        keyinput_g94), .B2(D_REG_7__SCAN_IN), .ZN(n4718) );
  AOI221_X1 U5253 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput_g86), .C1(
        D_REG_7__SCAN_IN), .C2(keyinput_g94), .A(n4718), .ZN(n4721) );
  OAI22_X1 U5254 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput_g83), .B1(
        keyinput_g119), .B2(REG0_REG_0__SCAN_IN), .ZN(n4719) );
  AOI221_X1 U5255 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput_g83), .C1(
        REG0_REG_0__SCAN_IN), .C2(keyinput_g119), .A(n4719), .ZN(n4720) );
  NAND4_X1 U5256 ( .A1(n4723), .A2(n4722), .A3(n4721), .A4(n4720), .ZN(n4733)
         );
  OAI22_X1 U5257 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput_g67), .B1(
        REG0_REG_6__SCAN_IN), .B2(keyinput_g125), .ZN(n4724) );
  AOI221_X1 U5258 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput_g67), .C1(
        keyinput_g125), .C2(REG0_REG_6__SCAN_IN), .A(n4724), .ZN(n4731) );
  OAI22_X1 U5259 ( .A1(IR_REG_22__SCAN_IN), .A2(keyinput_g77), .B1(
        keyinput_g60), .B2(IR_REG_5__SCAN_IN), .ZN(n4725) );
  AOI221_X1 U5260 ( .B1(IR_REG_22__SCAN_IN), .B2(keyinput_g77), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_g60), .A(n4725), .ZN(n4730) );
  OAI22_X1 U5261 ( .A1(D_REG_3__SCAN_IN), .A2(keyinput_g90), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_g48), .ZN(n4726) );
  AOI221_X1 U5262 ( .B1(D_REG_3__SCAN_IN), .B2(keyinput_g90), .C1(keyinput_g48), .C2(REG3_REG_17__SCAN_IN), .A(n4726), .ZN(n4729) );
  OAI22_X1 U5263 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput_g44), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .ZN(n4727) );
  AOI221_X1 U5264 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .C1(
        keyinput_g37), .C2(REG3_REG_10__SCAN_IN), .A(n4727), .ZN(n4728) );
  NAND4_X1 U5265 ( .A1(n4731), .A2(n4730), .A3(n4729), .A4(n4728), .ZN(n4732)
         );
  NOR4_X1 U5266 ( .A1(n4735), .A2(n4734), .A3(n4733), .A4(n4732), .ZN(n5069)
         );
  OAI22_X1 U5267 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_g88), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput_g113), .ZN(n4736) );
  AOI221_X1 U5268 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_g88), .C1(
        keyinput_g113), .C2(D_REG_26__SCAN_IN), .A(n4736), .ZN(n4743) );
  OAI22_X1 U5269 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_g32), .B1(DATAI_29_), 
        .B2(keyinput_g2), .ZN(n4737) );
  AOI221_X1 U5270 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_g32), .C1(keyinput_g2), .C2(DATAI_29_), .A(n4737), .ZN(n4742) );
  OAI22_X1 U5271 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput_g114), .B1(
        REG0_REG_4__SCAN_IN), .B2(keyinput_g123), .ZN(n4738) );
  AOI221_X1 U5272 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput_g114), .C1(
        keyinput_g123), .C2(REG0_REG_4__SCAN_IN), .A(n4738), .ZN(n4741) );
  OAI22_X1 U5273 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_g33), .B1(DATAI_0_), 
        .B2(keyinput_g31), .ZN(n4739) );
  AOI221_X1 U5274 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_g33), .C1(
        keyinput_g31), .C2(DATAI_0_), .A(n4739), .ZN(n4740) );
  NAND4_X1 U5275 ( .A1(n4743), .A2(n4742), .A3(n4741), .A4(n4740), .ZN(n4868)
         );
  AOI22_X1 U5276 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_g36), .ZN(n4744) );
  OAI221_X1 U5277 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_g36), .A(n4744), .ZN(n4751) );
  AOI22_X1 U5278 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(REG3_REG_28__SCAN_IN), 
        .B2(keyinput_g40), .ZN(n4745) );
  OAI221_X1 U5279 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(REG3_REG_28__SCAN_IN), .C2(keyinput_g40), .A(n4745), .ZN(n4750) );
  AOI22_X1 U5280 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_g39), .B1(
        D_REG_22__SCAN_IN), .B2(keyinput_g109), .ZN(n4746) );
  OAI221_X1 U5281 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .C1(
        D_REG_22__SCAN_IN), .C2(keyinput_g109), .A(n4746), .ZN(n4749) );
  AOI22_X1 U5282 ( .A1(DATAI_31_), .A2(keyinput_g0), .B1(D_REG_15__SCAN_IN), 
        .B2(keyinput_g102), .ZN(n4747) );
  OAI221_X1 U5283 ( .B1(DATAI_31_), .B2(keyinput_g0), .C1(D_REG_15__SCAN_IN), 
        .C2(keyinput_g102), .A(n4747), .ZN(n4748) );
  NOR4_X1 U5284 ( .A1(n4751), .A2(n4750), .A3(n4749), .A4(n4748), .ZN(n4769)
         );
  AOI22_X1 U5285 ( .A1(REG0_REG_7__SCAN_IN), .A2(keyinput_g126), .B1(
        IR_REG_11__SCAN_IN), .B2(keyinput_g66), .ZN(n4752) );
  OAI221_X1 U5286 ( .B1(REG0_REG_7__SCAN_IN), .B2(keyinput_g126), .C1(
        IR_REG_11__SCAN_IN), .C2(keyinput_g66), .A(n4752), .ZN(n4759) );
  AOI22_X1 U5287 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(D_REG_31__SCAN_IN), 
        .B2(keyinput_g118), .ZN(n4753) );
  OAI221_X1 U5288 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(D_REG_31__SCAN_IN), 
        .C2(keyinput_g118), .A(n4753), .ZN(n4758) );
  AOI22_X1 U5289 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_g122), .B1(
        IR_REG_7__SCAN_IN), .B2(keyinput_g62), .ZN(n4754) );
  OAI221_X1 U5290 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_g122), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput_g62), .A(n4754), .ZN(n4757) );
  AOI22_X1 U5291 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(REG3_REG_4__SCAN_IN), 
        .B2(keyinput_g50), .ZN(n4755) );
  OAI221_X1 U5292 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(REG3_REG_4__SCAN_IN), 
        .C2(keyinput_g50), .A(n4755), .ZN(n4756) );
  NOR4_X1 U5293 ( .A1(n4759), .A2(n4758), .A3(n4757), .A4(n4756), .ZN(n4768)
         );
  OAI22_X1 U5294 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput_g63), .B1(keyinput_g29), .B2(DATAI_2_), .ZN(n4760) );
  AOI221_X1 U5295 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput_g63), .C1(DATAI_2_), 
        .C2(keyinput_g29), .A(n4760), .ZN(n4766) );
  OAI22_X1 U5296 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_g34), .B1(
        keyinput_g6), .B2(DATAI_25_), .ZN(n4761) );
  AOI221_X1 U5297 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .C1(
        DATAI_25_), .C2(keyinput_g6), .A(n4761), .ZN(n4765) );
  OAI22_X1 U5298 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_g55), .B1(
        D_REG_16__SCAN_IN), .B2(keyinput_g103), .ZN(n4762) );
  AOI221_X1 U5299 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_g55), .C1(
        keyinput_g103), .C2(D_REG_16__SCAN_IN), .A(n4762), .ZN(n4764) );
  XNOR2_X1 U5300 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_g76), .ZN(n4763) );
  AND4_X1 U5301 ( .A1(n4766), .A2(n4765), .A3(n4764), .A4(n4763), .ZN(n4767)
         );
  NAND3_X1 U5302 ( .A1(n4769), .A2(n4768), .A3(n4767), .ZN(n4867) );
  AOI22_X1 U5303 ( .A1(REG0_REG_2__SCAN_IN), .A2(keyinput_g121), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput_g104), .ZN(n4770) );
  OAI221_X1 U5304 ( .B1(REG0_REG_2__SCAN_IN), .B2(keyinput_g121), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput_g104), .A(n4770), .ZN(n4778) );
  INV_X1 U5305 ( .A(DATAI_30_), .ZN(n4772) );
  AOI22_X1 U5306 ( .A1(n4772), .A2(keyinput_g1), .B1(n5023), .B2(keyinput_g92), 
        .ZN(n4771) );
  OAI221_X1 U5307 ( .B1(n4772), .B2(keyinput_g1), .C1(n5023), .C2(keyinput_g92), .A(n4771), .ZN(n4777) );
  AOI22_X1 U5308 ( .A1(n5027), .A2(keyinput_g107), .B1(keyinput_g43), .B2(
        n2672), .ZN(n4773) );
  OAI221_X1 U5309 ( .B1(n5027), .B2(keyinput_g107), .C1(n2672), .C2(
        keyinput_g43), .A(n4773), .ZN(n4776) );
  INV_X1 U5310 ( .A(DATAI_22_), .ZN(n4950) );
  AOI22_X1 U5311 ( .A1(n2822), .A2(keyinput_g87), .B1(keyinput_g9), .B2(n4950), 
        .ZN(n4774) );
  OAI221_X1 U5312 ( .B1(n2822), .B2(keyinput_g87), .C1(n4950), .C2(keyinput_g9), .A(n4774), .ZN(n4775) );
  NOR4_X1 U5313 ( .A1(n4778), .A2(n4777), .A3(n4776), .A4(n4775), .ZN(n4818)
         );
  AOI22_X1 U5314 ( .A1(n5032), .A2(keyinput_g99), .B1(keyinput_g93), .B2(n4780), .ZN(n4779) );
  OAI221_X1 U5315 ( .B1(n5032), .B2(keyinput_g99), .C1(n4780), .C2(
        keyinput_g93), .A(n4779), .ZN(n4790) );
  AOI22_X1 U5316 ( .A1(n4783), .A2(keyinput_g101), .B1(keyinput_g120), .B2(
        n4782), .ZN(n4781) );
  OAI221_X1 U5317 ( .B1(n4783), .B2(keyinput_g101), .C1(n4782), .C2(
        keyinput_g120), .A(n4781), .ZN(n4789) );
  XNOR2_X1 U5318 ( .A(DATAI_12_), .B(keyinput_g19), .ZN(n4787) );
  XNOR2_X1 U5319 ( .A(DATAI_4_), .B(keyinput_g27), .ZN(n4786) );
  XNOR2_X1 U5320 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n4785) );
  XNOR2_X1 U5321 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4784) );
  NAND4_X1 U5322 ( .A1(n4787), .A2(n4786), .A3(n4785), .A4(n4784), .ZN(n4788)
         );
  NOR3_X1 U5323 ( .A1(n4790), .A2(n4789), .A3(n4788), .ZN(n4817) );
  AOI22_X1 U5324 ( .A1(n4792), .A2(keyinput_g115), .B1(keyinput_g35), .B2(
        n4957), .ZN(n4791) );
  OAI221_X1 U5325 ( .B1(n4792), .B2(keyinput_g115), .C1(n4957), .C2(
        keyinput_g35), .A(n4791), .ZN(n4796) );
  XNOR2_X1 U5326 ( .A(n5029), .B(keyinput_g100), .ZN(n4795) );
  XNOR2_X1 U5327 ( .A(n4793), .B(keyinput_g68), .ZN(n4794) );
  OR3_X1 U5328 ( .A1(n4796), .A2(n4795), .A3(n4794), .ZN(n4801) );
  AOI22_X1 U5329 ( .A1(n5026), .A2(keyinput_g106), .B1(keyinput_g91), .B2(
        n5030), .ZN(n4797) );
  OAI221_X1 U5330 ( .B1(n5026), .B2(keyinput_g106), .C1(n5030), .C2(
        keyinput_g91), .A(n4797), .ZN(n4800) );
  AOI22_X1 U5331 ( .A1(n5044), .A2(keyinput_g10), .B1(n2626), .B2(keyinput_g70), .ZN(n4798) );
  OAI221_X1 U5332 ( .B1(n5044), .B2(keyinput_g10), .C1(n2626), .C2(
        keyinput_g70), .A(n4798), .ZN(n4799) );
  NOR3_X1 U5333 ( .A1(n4801), .A2(n4800), .A3(n4799), .ZN(n4816) );
  INV_X1 U5334 ( .A(IR_REG_10__SCAN_IN), .ZN(n4803) );
  AOI22_X1 U5335 ( .A1(n5011), .A2(keyinput_g105), .B1(n4803), .B2(
        keyinput_g65), .ZN(n4802) );
  OAI221_X1 U5336 ( .B1(n5011), .B2(keyinput_g105), .C1(n4803), .C2(
        keyinput_g65), .A(n4802), .ZN(n4814) );
  AOI22_X1 U5337 ( .A1(n5014), .A2(keyinput_g110), .B1(n4805), .B2(
        keyinput_g117), .ZN(n4804) );
  OAI221_X1 U5338 ( .B1(n5014), .B2(keyinput_g110), .C1(n4805), .C2(
        keyinput_g117), .A(n4804), .ZN(n4813) );
  AOI22_X1 U5339 ( .A1(n5007), .A2(keyinput_g97), .B1(keyinput_g21), .B2(n4807), .ZN(n4806) );
  OAI221_X1 U5340 ( .B1(n5007), .B2(keyinput_g97), .C1(n4807), .C2(
        keyinput_g21), .A(n4806), .ZN(n4812) );
  XOR2_X1 U5341 ( .A(n4808), .B(keyinput_g18), .Z(n4810) );
  XNOR2_X1 U5342 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_g73), .ZN(n4809) );
  NAND2_X1 U5343 ( .A1(n4810), .A2(n4809), .ZN(n4811) );
  NOR4_X1 U5344 ( .A1(n4814), .A2(n4813), .A3(n4812), .A4(n4811), .ZN(n4815)
         );
  NAND4_X1 U5345 ( .A1(n4818), .A2(n4817), .A3(n4816), .A4(n4815), .ZN(n4866)
         );
  INV_X1 U5346 ( .A(DATAI_3_), .ZN(n4820) );
  AOI22_X1 U5347 ( .A1(n5041), .A2(keyinput_g46), .B1(keyinput_g28), .B2(n4820), .ZN(n4819) );
  OAI221_X1 U5348 ( .B1(n5041), .B2(keyinput_g46), .C1(n4820), .C2(
        keyinput_g28), .A(n4819), .ZN(n4829) );
  AOI22_X1 U5349 ( .A1(n2451), .A2(keyinput_g69), .B1(keyinput_g53), .B2(n4822), .ZN(n4821) );
  OAI221_X1 U5350 ( .B1(n2451), .B2(keyinput_g69), .C1(n4822), .C2(
        keyinput_g53), .A(n4821), .ZN(n4828) );
  AOI22_X1 U5351 ( .A1(n4998), .A2(keyinput_g23), .B1(n4968), .B2(keyinput_g71), .ZN(n4823) );
  OAI221_X1 U5352 ( .B1(n4998), .B2(keyinput_g23), .C1(n4968), .C2(
        keyinput_g71), .A(n4823), .ZN(n4827) );
  XOR2_X1 U5353 ( .A(n2410), .B(keyinput_g72), .Z(n4825) );
  XNOR2_X1 U5354 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_g59), .ZN(n4824) );
  NAND2_X1 U5355 ( .A1(n4825), .A2(n4824), .ZN(n4826) );
  NOR4_X1 U5356 ( .A1(n4829), .A2(n4828), .A3(n4827), .A4(n4826), .ZN(n4864)
         );
  INV_X1 U5357 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4979) );
  AOI22_X1 U5358 ( .A1(n4979), .A2(keyinput_g124), .B1(n4831), .B2(
        keyinput_g47), .ZN(n4830) );
  OAI221_X1 U5359 ( .B1(n4979), .B2(keyinput_g124), .C1(n4831), .C2(
        keyinput_g47), .A(n4830), .ZN(n4840) );
  AOI22_X1 U5360 ( .A1(n2391), .A2(keyinput_g57), .B1(keyinput_g14), .B2(n2642), .ZN(n4832) );
  OAI221_X1 U5361 ( .B1(n2391), .B2(keyinput_g57), .C1(n2642), .C2(
        keyinput_g14), .A(n4832), .ZN(n4839) );
  INV_X1 U5362 ( .A(DATAI_6_), .ZN(n4834) );
  AOI22_X1 U5363 ( .A1(n5008), .A2(keyinput_g96), .B1(keyinput_g25), .B2(n4834), .ZN(n4833) );
  OAI221_X1 U5364 ( .B1(n5008), .B2(keyinput_g96), .C1(n4834), .C2(
        keyinput_g25), .A(n4833), .ZN(n4838) );
  XNOR2_X1 U5365 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_g82), .ZN(n4836) );
  XNOR2_X1 U5366 ( .A(keyinput_g24), .B(DATAI_7_), .ZN(n4835) );
  NAND2_X1 U5367 ( .A1(n4836), .A2(n4835), .ZN(n4837) );
  NOR4_X1 U5368 ( .A1(n4840), .A2(n4839), .A3(n4838), .A4(n4837), .ZN(n4863)
         );
  AOI22_X1 U5369 ( .A1(n5013), .A2(keyinput_g89), .B1(keyinput_g49), .B2(n4940), .ZN(n4841) );
  OAI221_X1 U5370 ( .B1(n5013), .B2(keyinput_g89), .C1(n4940), .C2(
        keyinput_g49), .A(n4841), .ZN(n4844) );
  XNOR2_X1 U5371 ( .A(n5017), .B(keyinput_g111), .ZN(n4843) );
  XOR2_X1 U5372 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_g64), .Z(n4842) );
  OR3_X1 U5373 ( .A1(n4844), .A2(n4843), .A3(n4842), .ZN(n4850) );
  AOI22_X1 U5374 ( .A1(n4956), .A2(keyinput_g16), .B1(n3087), .B2(keyinput_g42), .ZN(n4845) );
  OAI221_X1 U5375 ( .B1(n4956), .B2(keyinput_g16), .C1(n3087), .C2(
        keyinput_g42), .A(n4845), .ZN(n4849) );
  AOI22_X1 U5376 ( .A1(n4847), .A2(keyinput_g41), .B1(keyinput_g52), .B2(n2475), .ZN(n4846) );
  OAI221_X1 U5377 ( .B1(n4847), .B2(keyinput_g41), .C1(n2475), .C2(
        keyinput_g52), .A(n4846), .ZN(n4848) );
  NOR3_X1 U5378 ( .A1(n4850), .A2(n4849), .A3(n4848), .ZN(n4862) );
  INV_X1 U5379 ( .A(DATAI_5_), .ZN(n4852) );
  AOI22_X1 U5380 ( .A1(n5016), .A2(keyinput_g98), .B1(keyinput_g26), .B2(n4852), .ZN(n4851) );
  OAI221_X1 U5381 ( .B1(n5016), .B2(keyinput_g98), .C1(n4852), .C2(
        keyinput_g26), .A(n4851), .ZN(n4860) );
  AOI22_X1 U5382 ( .A1(n2735), .A2(keyinput_g74), .B1(keyinput_g51), .B2(n2549), .ZN(n4853) );
  OAI221_X1 U5383 ( .B1(n2735), .B2(keyinput_g74), .C1(n2549), .C2(
        keyinput_g51), .A(n4853), .ZN(n4859) );
  XOR2_X1 U5384 ( .A(n4995), .B(keyinput_g20), .Z(n4857) );
  XNOR2_X1 U5385 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_g58), .ZN(n4856) );
  XNOR2_X1 U5386 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_g80), .ZN(n4855) );
  XNOR2_X1 U5387 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_g78), .ZN(n4854) );
  NAND4_X1 U5388 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n4858)
         );
  NOR3_X1 U5389 ( .A1(n4860), .A2(n4859), .A3(n4858), .ZN(n4861) );
  NAND4_X1 U5390 ( .A1(n4864), .A2(n4863), .A3(n4862), .A4(n4861), .ZN(n4865)
         );
  NOR4_X1 U5391 ( .A1(n4868), .A2(n4867), .A3(n4866), .A4(n4865), .ZN(n5068)
         );
  OAI22_X1 U5392 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput_f67), .B1(
        keyinput_f83), .B2(IR_REG_28__SCAN_IN), .ZN(n4869) );
  AOI221_X1 U5393 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput_f67), .C1(
        IR_REG_28__SCAN_IN), .C2(keyinput_f83), .A(n4869), .ZN(n4876) );
  OAI22_X1 U5394 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput_f66), .B1(DATAI_10_), 
        .B2(keyinput_f21), .ZN(n4870) );
  AOI221_X1 U5395 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput_f66), .C1(
        keyinput_f21), .C2(DATAI_10_), .A(n4870), .ZN(n4875) );
  OAI22_X1 U5396 ( .A1(IR_REG_10__SCAN_IN), .A2(keyinput_f65), .B1(DATAI_7_), 
        .B2(keyinput_f24), .ZN(n4871) );
  AOI221_X1 U5397 ( .B1(IR_REG_10__SCAN_IN), .B2(keyinput_f65), .C1(
        keyinput_f24), .C2(DATAI_7_), .A(n4871), .ZN(n4874) );
  OAI22_X1 U5398 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_f62), .B1(DATAI_6_), 
        .B2(keyinput_f25), .ZN(n4872) );
  AOI221_X1 U5399 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_f62), .C1(
        keyinput_f25), .C2(DATAI_6_), .A(n4872), .ZN(n4873) );
  NAND4_X1 U5400 ( .A1(n4876), .A2(n4875), .A3(n4874), .A4(n4873), .ZN(n4904)
         );
  OAI22_X1 U5401 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_f60), .B1(keyinput_f47), .B2(REG3_REG_5__SCAN_IN), .ZN(n4877) );
  AOI221_X1 U5402 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_f60), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput_f47), .A(n4877), .ZN(n4884) );
  OAI22_X1 U5403 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput_f120), .B1(
        keyinput_f31), .B2(DATAI_0_), .ZN(n4878) );
  AOI221_X1 U5404 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput_f120), .C1(DATAI_0_), .C2(keyinput_f31), .A(n4878), .ZN(n4883) );
  OAI22_X1 U5405 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput_f64), .B1(keyinput_f28), .B2(DATAI_3_), .ZN(n4879) );
  AOI221_X1 U5406 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput_f64), .C1(DATAI_3_), 
        .C2(keyinput_f28), .A(n4879), .ZN(n4882) );
  OAI22_X1 U5407 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_f88), .B1(keyinput_f51), 
        .B2(REG3_REG_9__SCAN_IN), .ZN(n4880) );
  AOI221_X1 U5408 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_f88), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_f51), .A(n4880), .ZN(n4881) );
  NAND4_X1 U5409 ( .A1(n4884), .A2(n4883), .A3(n4882), .A4(n4881), .ZN(n4903)
         );
  OAI22_X1 U5410 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput_f75), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput_f93), .ZN(n4885) );
  AOI221_X1 U5411 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput_f75), .C1(
        keyinput_f93), .C2(D_REG_6__SCAN_IN), .A(n4885), .ZN(n4892) );
  OAI22_X1 U5412 ( .A1(D_REG_30__SCAN_IN), .A2(keyinput_f117), .B1(
        D_REG_28__SCAN_IN), .B2(keyinput_f115), .ZN(n4886) );
  AOI221_X1 U5413 ( .B1(D_REG_30__SCAN_IN), .B2(keyinput_f117), .C1(
        keyinput_f115), .C2(D_REG_28__SCAN_IN), .A(n4886), .ZN(n4891) );
  OAI22_X1 U5414 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .ZN(n4887) );
  AOI221_X1 U5415 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f43), .C2(REG3_REG_21__SCAN_IN), .A(n4887), .ZN(n4890) );
  OAI22_X1 U5416 ( .A1(IR_REG_29__SCAN_IN), .A2(keyinput_f84), .B1(
        keyinput_f36), .B2(REG3_REG_23__SCAN_IN), .ZN(n4888) );
  AOI221_X1 U5417 ( .B1(IR_REG_29__SCAN_IN), .B2(keyinput_f84), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_f36), .A(n4888), .ZN(n4889) );
  NAND4_X1 U5418 ( .A1(n4892), .A2(n4891), .A3(n4890), .A4(n4889), .ZN(n4902)
         );
  OAI22_X1 U5419 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput_f80), .B1(
        IR_REG_23__SCAN_IN), .B2(keyinput_f78), .ZN(n4893) );
  AOI221_X1 U5420 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput_f80), .C1(
        keyinput_f78), .C2(IR_REG_23__SCAN_IN), .A(n4893), .ZN(n4900) );
  OAI22_X1 U5421 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(keyinput_f1), .B2(
        DATAI_30_), .ZN(n4894) );
  AOI221_X1 U5422 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(DATAI_30_), .C2(
        keyinput_f1), .A(n4894), .ZN(n4899) );
  OAI22_X1 U5423 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput_f87), .B1(keyinput_f27), 
        .B2(DATAI_4_), .ZN(n4895) );
  AOI221_X1 U5424 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput_f87), .C1(DATAI_4_), 
        .C2(keyinput_f27), .A(n4895), .ZN(n4898) );
  OAI22_X1 U5425 ( .A1(U3149), .A2(keyinput_f32), .B1(keyinput_f41), .B2(
        REG3_REG_8__SCAN_IN), .ZN(n4896) );
  AOI221_X1 U5426 ( .B1(U3149), .B2(keyinput_f32), .C1(REG3_REG_8__SCAN_IN), 
        .C2(keyinput_f41), .A(n4896), .ZN(n4897) );
  NAND4_X1 U5427 ( .A1(n4900), .A2(n4899), .A3(n4898), .A4(n4897), .ZN(n4901)
         );
  NOR4_X1 U5428 ( .A1(n4904), .A2(n4903), .A3(n4902), .A4(n4901), .ZN(n5062)
         );
  OAI22_X1 U5429 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_f53), .B1(DATAI_29_), .B2(keyinput_f2), .ZN(n4905) );
  AOI221_X1 U5430 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_f53), .C1(
        keyinput_f2), .C2(DATAI_29_), .A(n4905), .ZN(n4912) );
  OAI22_X1 U5431 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput_f38), .B1(
        keyinput_f13), .B2(DATAI_18_), .ZN(n4906) );
  AOI221_X1 U5432 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_f38), .C1(DATAI_18_), .C2(keyinput_f13), .A(n4906), .ZN(n4911) );
  OAI22_X1 U5433 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput_f82), .B1(
        keyinput_f54), .B2(REG3_REG_13__SCAN_IN), .ZN(n4907) );
  AOI221_X1 U5434 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput_f82), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput_f54), .A(n4907), .ZN(n4910) );
  OAI22_X1 U5435 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput_f118), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput_f116), .ZN(n4908) );
  AOI221_X1 U5436 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput_f118), .C1(
        keyinput_f116), .C2(D_REG_29__SCAN_IN), .A(n4908), .ZN(n4909) );
  NAND4_X1 U5437 ( .A1(n4912), .A2(n4911), .A3(n4910), .A4(n4909), .ZN(n5060)
         );
  AOI22_X1 U5438 ( .A1(D_REG_22__SCAN_IN), .A2(keyinput_f109), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput_f114), .ZN(n4913) );
  OAI221_X1 U5439 ( .B1(D_REG_22__SCAN_IN), .B2(keyinput_f109), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput_f114), .A(n4913), .ZN(n4920) );
  AOI22_X1 U5440 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput_f104), .B1(
        D_REG_21__SCAN_IN), .B2(keyinput_f108), .ZN(n4914) );
  OAI221_X1 U5441 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput_f104), .C1(
        D_REG_21__SCAN_IN), .C2(keyinput_f108), .A(n4914), .ZN(n4919) );
  AOI22_X1 U5442 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput_f102), .B1(
        D_REG_16__SCAN_IN), .B2(keyinput_f103), .ZN(n4915) );
  OAI221_X1 U5443 ( .B1(D_REG_15__SCAN_IN), .B2(keyinput_f102), .C1(
        D_REG_16__SCAN_IN), .C2(keyinput_f103), .A(n4915), .ZN(n4918) );
  AOI22_X1 U5444 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput_f94), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput_f95), .ZN(n4916) );
  OAI221_X1 U5445 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput_f94), .C1(
        D_REG_8__SCAN_IN), .C2(keyinput_f95), .A(n4916), .ZN(n4917) );
  NOR4_X1 U5446 ( .A1(n4920), .A2(n4919), .A3(n4918), .A4(n4917), .ZN(n4938)
         );
  AOI22_X1 U5447 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(IR_REG_14__SCAN_IN), 
        .B2(keyinput_f69), .ZN(n4921) );
  OAI221_X1 U5448 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(IR_REG_14__SCAN_IN), 
        .C2(keyinput_f69), .A(n4921), .ZN(n4928) );
  AOI22_X1 U5449 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput_f119), .B1(DATAI_14_), .B2(keyinput_f17), .ZN(n4922) );
  OAI221_X1 U5450 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput_f119), .C1(
        DATAI_14_), .C2(keyinput_f17), .A(n4922), .ZN(n4927) );
  AOI22_X1 U5451 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput_f123), .B1(
        REG0_REG_3__SCAN_IN), .B2(keyinput_f122), .ZN(n4923) );
  OAI221_X1 U5452 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput_f123), .C1(
        REG0_REG_3__SCAN_IN), .C2(keyinput_f122), .A(n4923), .ZN(n4926) );
  AOI22_X1 U5453 ( .A1(REG0_REG_7__SCAN_IN), .A2(keyinput_f126), .B1(
        REG0_REG_8__SCAN_IN), .B2(keyinput_f127), .ZN(n4924) );
  OAI221_X1 U5454 ( .B1(REG0_REG_7__SCAN_IN), .B2(keyinput_f126), .C1(
        REG0_REG_8__SCAN_IN), .C2(keyinput_f127), .A(n4924), .ZN(n4925) );
  NOR4_X1 U5455 ( .A1(n4928), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(n4937)
         );
  OAI22_X1 U5456 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput_f40), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput_f39), .ZN(n4929) );
  AOI221_X1 U5457 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .C1(
        keyinput_f39), .C2(REG3_REG_19__SCAN_IN), .A(n4929), .ZN(n4935) );
  OAI22_X1 U5458 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(
        keyinput_f7), .B2(DATAI_24_), .ZN(n4930) );
  AOI221_X1 U5459 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(DATAI_24_), .C2(keyinput_f7), .A(n4930), .ZN(n4934) );
  OAI22_X1 U5460 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_f45), .B1(DATAI_25_), .B2(keyinput_f6), .ZN(n4931) );
  AOI221_X1 U5461 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_f45), .C1(
        keyinput_f6), .C2(DATAI_25_), .A(n4931), .ZN(n4933) );
  XNOR2_X1 U5462 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_f79), .ZN(n4932) );
  AND4_X1 U5463 ( .A1(n4935), .A2(n4934), .A3(n4933), .A4(n4932), .ZN(n4936)
         );
  NAND3_X1 U5464 ( .A1(n4938), .A2(n4937), .A3(n4936), .ZN(n5059) );
  AOI22_X1 U5465 ( .A1(n4941), .A2(keyinput_f34), .B1(keyinput_f49), .B2(n4940), .ZN(n4939) );
  OAI221_X1 U5466 ( .B1(n4941), .B2(keyinput_f34), .C1(n4940), .C2(
        keyinput_f49), .A(n4939), .ZN(n4954) );
  AOI22_X1 U5467 ( .A1(n4944), .A2(keyinput_f3), .B1(keyinput_f4), .B2(n4943), 
        .ZN(n4942) );
  OAI221_X1 U5468 ( .B1(n4944), .B2(keyinput_f3), .C1(n4943), .C2(keyinput_f4), 
        .A(n4942), .ZN(n4953) );
  INV_X1 U5469 ( .A(DATAI_26_), .ZN(n4947) );
  AOI22_X1 U5470 ( .A1(n4947), .A2(keyinput_f5), .B1(n4946), .B2(keyinput_f8), 
        .ZN(n4945) );
  OAI221_X1 U5471 ( .B1(n4947), .B2(keyinput_f5), .C1(n4946), .C2(keyinput_f8), 
        .A(n4945), .ZN(n4952) );
  INV_X1 U5472 ( .A(DATAI_20_), .ZN(n4949) );
  AOI22_X1 U5473 ( .A1(n4950), .A2(keyinput_f9), .B1(keyinput_f11), .B2(n4949), 
        .ZN(n4948) );
  OAI221_X1 U5474 ( .B1(n4950), .B2(keyinput_f9), .C1(n4949), .C2(keyinput_f11), .A(n4948), .ZN(n4951) );
  NOR4_X1 U5475 ( .A1(n4954), .A2(n4953), .A3(n4952), .A4(n4951), .ZN(n4993)
         );
  AOI22_X1 U5476 ( .A1(n4957), .A2(keyinput_f35), .B1(keyinput_f16), .B2(n4956), .ZN(n4955) );
  OAI221_X1 U5477 ( .B1(n4957), .B2(keyinput_f35), .C1(n4956), .C2(
        keyinput_f16), .A(n4955), .ZN(n4966) );
  AOI22_X1 U5478 ( .A1(n2660), .A2(keyinput_f12), .B1(keyinput_f14), .B2(n2642), .ZN(n4958) );
  OAI221_X1 U5479 ( .B1(n2660), .B2(keyinput_f12), .C1(n2642), .C2(
        keyinput_f14), .A(n4958), .ZN(n4965) );
  AOI22_X1 U5480 ( .A1(n3087), .A2(keyinput_f42), .B1(n4960), .B2(keyinput_f55), .ZN(n4959) );
  OAI221_X1 U5481 ( .B1(n3087), .B2(keyinput_f42), .C1(n4960), .C2(
        keyinput_f55), .A(n4959), .ZN(n4964) );
  XOR2_X1 U5482 ( .A(n2857), .B(keyinput_f85), .Z(n4962) );
  XNOR2_X1 U5483 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_f86), .ZN(n4961) );
  NAND2_X1 U5484 ( .A1(n4962), .A2(n4961), .ZN(n4963) );
  NOR4_X1 U5485 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n4992)
         );
  AOI22_X1 U5486 ( .A1(n4968), .A2(keyinput_f71), .B1(keyinput_f70), .B2(n2626), .ZN(n4967) );
  OAI221_X1 U5487 ( .B1(n4968), .B2(keyinput_f71), .C1(n2626), .C2(
        keyinput_f70), .A(n4967), .ZN(n4977) );
  XNOR2_X1 U5488 ( .A(keyinput_f72), .B(n2410), .ZN(n4976) );
  XNOR2_X1 U5489 ( .A(keyinput_f33), .B(n4969), .ZN(n4975) );
  XNOR2_X1 U5490 ( .A(DATAI_12_), .B(keyinput_f19), .ZN(n4973) );
  XNOR2_X1 U5491 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_f73), .ZN(n4972) );
  XNOR2_X1 U5492 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n4971) );
  XNOR2_X1 U5493 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_f68), .ZN(n4970) );
  NAND4_X1 U5494 ( .A1(n4973), .A2(n4972), .A3(n4971), .A4(n4970), .ZN(n4974)
         );
  NOR4_X1 U5495 ( .A1(n4977), .A2(n4976), .A3(n4975), .A4(n4974), .ZN(n4991)
         );
  AOI22_X1 U5496 ( .A1(n4980), .A2(keyinput_f125), .B1(keyinput_f124), .B2(
        n4979), .ZN(n4978) );
  OAI221_X1 U5497 ( .B1(n4980), .B2(keyinput_f125), .C1(n4979), .C2(
        keyinput_f124), .A(n4978), .ZN(n4989) );
  INV_X1 U5498 ( .A(IR_REG_1__SCAN_IN), .ZN(n4982) );
  AOI22_X1 U5499 ( .A1(n2359), .A2(keyinput_f30), .B1(n4982), .B2(keyinput_f56), .ZN(n4981) );
  OAI221_X1 U5500 ( .B1(n2359), .B2(keyinput_f30), .C1(n4982), .C2(
        keyinput_f56), .A(n4981), .ZN(n4988) );
  XNOR2_X1 U5501 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4986) );
  XNOR2_X1 U5502 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4985) );
  XNOR2_X1 U5503 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n4984) );
  XNOR2_X1 U5504 ( .A(keyinput_f26), .B(DATAI_5_), .ZN(n4983) );
  NAND4_X1 U5505 ( .A1(n4986), .A2(n4985), .A3(n4984), .A4(n4983), .ZN(n4987)
         );
  NOR3_X1 U5506 ( .A1(n4989), .A2(n4988), .A3(n4987), .ZN(n4990) );
  NAND4_X1 U5507 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(n5058)
         );
  AOI22_X1 U5508 ( .A1(n4995), .A2(keyinput_f20), .B1(n2735), .B2(keyinput_f74), .ZN(n4994) );
  OAI221_X1 U5509 ( .B1(n4995), .B2(keyinput_f20), .C1(n2735), .C2(
        keyinput_f74), .A(n4994), .ZN(n5005) );
  INV_X1 U5510 ( .A(IR_REG_8__SCAN_IN), .ZN(n4997) );
  AOI22_X1 U5511 ( .A1(n4998), .A2(keyinput_f23), .B1(n4997), .B2(keyinput_f63), .ZN(n4996) );
  OAI221_X1 U5512 ( .B1(n4998), .B2(keyinput_f23), .C1(n4997), .C2(
        keyinput_f63), .A(n4996), .ZN(n5004) );
  XOR2_X1 U5513 ( .A(n2391), .B(keyinput_f57), .Z(n5002) );
  XOR2_X1 U5514 ( .A(n2733), .B(keyinput_f77), .Z(n5001) );
  XNOR2_X1 U5515 ( .A(DATAI_2_), .B(keyinput_f29), .ZN(n5000) );
  XNOR2_X1 U5516 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_f76), .ZN(n4999) );
  NAND4_X1 U5517 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n5003)
         );
  NOR3_X1 U5518 ( .A1(n5005), .A2(n5004), .A3(n5003), .ZN(n5056) );
  AOI22_X1 U5519 ( .A1(n5008), .A2(keyinput_f96), .B1(keyinput_f97), .B2(n5007), .ZN(n5006) );
  OAI221_X1 U5520 ( .B1(n5008), .B2(keyinput_f96), .C1(n5007), .C2(
        keyinput_f97), .A(n5006), .ZN(n5021) );
  AOI22_X1 U5521 ( .A1(n5011), .A2(keyinput_f105), .B1(keyinput_f90), .B2(
        n5010), .ZN(n5009) );
  OAI221_X1 U5522 ( .B1(n5011), .B2(keyinput_f105), .C1(n5010), .C2(
        keyinput_f90), .A(n5009), .ZN(n5020) );
  AOI22_X1 U5523 ( .A1(n5014), .A2(keyinput_f110), .B1(keyinput_f89), .B2(
        n5013), .ZN(n5012) );
  OAI221_X1 U5524 ( .B1(n5014), .B2(keyinput_f110), .C1(n5013), .C2(
        keyinput_f89), .A(n5012), .ZN(n5019) );
  AOI22_X1 U5525 ( .A1(n5017), .A2(keyinput_f111), .B1(keyinput_f98), .B2(
        n5016), .ZN(n5015) );
  OAI221_X1 U5526 ( .B1(n5017), .B2(keyinput_f111), .C1(n5016), .C2(
        keyinput_f98), .A(n5015), .ZN(n5018) );
  NOR4_X1 U5527 ( .A1(n5021), .A2(n5020), .A3(n5019), .A4(n5018), .ZN(n5055)
         );
  AOI22_X1 U5528 ( .A1(n5024), .A2(keyinput_f113), .B1(keyinput_f92), .B2(
        n5023), .ZN(n5022) );
  OAI221_X1 U5529 ( .B1(n5024), .B2(keyinput_f113), .C1(n5023), .C2(
        keyinput_f92), .A(n5022), .ZN(n5037) );
  AOI22_X1 U5530 ( .A1(n5027), .A2(keyinput_f107), .B1(keyinput_f106), .B2(
        n5026), .ZN(n5025) );
  OAI221_X1 U5531 ( .B1(n5027), .B2(keyinput_f107), .C1(n5026), .C2(
        keyinput_f106), .A(n5025), .ZN(n5036) );
  AOI22_X1 U5532 ( .A1(n5030), .A2(keyinput_f91), .B1(keyinput_f100), .B2(
        n5029), .ZN(n5028) );
  OAI221_X1 U5533 ( .B1(n5030), .B2(keyinput_f91), .C1(n5029), .C2(
        keyinput_f100), .A(n5028), .ZN(n5035) );
  AOI22_X1 U5534 ( .A1(n5033), .A2(keyinput_f112), .B1(keyinput_f99), .B2(
        n5032), .ZN(n5031) );
  OAI221_X1 U5535 ( .B1(n5033), .B2(keyinput_f112), .C1(n5032), .C2(
        keyinput_f99), .A(n5031), .ZN(n5034) );
  NOR4_X1 U5536 ( .A1(n5037), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n5054)
         );
  AOI22_X1 U5537 ( .A1(n2632), .A2(keyinput_f48), .B1(keyinput_f15), .B2(n5039), .ZN(n5038) );
  OAI221_X1 U5538 ( .B1(n2632), .B2(keyinput_f48), .C1(n5039), .C2(
        keyinput_f15), .A(n5038), .ZN(n5052) );
  AOI22_X1 U5539 ( .A1(n5042), .A2(keyinput_f81), .B1(keyinput_f46), .B2(n5041), .ZN(n5040) );
  OAI221_X1 U5540 ( .B1(n5042), .B2(keyinput_f81), .C1(n5041), .C2(
        keyinput_f46), .A(n5040), .ZN(n5051) );
  AOI22_X1 U5541 ( .A1(n5045), .A2(keyinput_f121), .B1(n5044), .B2(
        keyinput_f10), .ZN(n5043) );
  OAI221_X1 U5542 ( .B1(n5045), .B2(keyinput_f121), .C1(n5044), .C2(
        keyinput_f10), .A(n5043), .ZN(n5050) );
  INV_X1 U5543 ( .A(REG3_REG_10__SCAN_IN), .ZN(n5048) );
  AOI22_X1 U5544 ( .A1(n5048), .A2(keyinput_f37), .B1(n5047), .B2(keyinput_f44), .ZN(n5046) );
  OAI221_X1 U5545 ( .B1(n5048), .B2(keyinput_f37), .C1(n5047), .C2(
        keyinput_f44), .A(n5046), .ZN(n5049) );
  NOR4_X1 U5546 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n5053)
         );
  NAND4_X1 U5547 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n5057)
         );
  NOR4_X1 U5548 ( .A1(n5060), .A2(n5059), .A3(n5058), .A4(n5057), .ZN(n5061)
         );
  NAND2_X1 U5549 ( .A1(n5062), .A2(n5061), .ZN(n5064) );
  AOI21_X1 U5550 ( .B1(keyinput_f22), .B2(n5064), .A(DATAI_9_), .ZN(n5066) );
  INV_X1 U5551 ( .A(keyinput_f22), .ZN(n5063) );
  AOI21_X1 U5552 ( .B1(n5064), .B2(n5063), .A(keyinput_g22), .ZN(n5065) );
  AOI22_X1 U5553 ( .A1(keyinput_g22), .A2(n5066), .B1(DATAI_9_), .B2(n5065), 
        .ZN(n5067) );
  AOI21_X1 U5554 ( .B1(n5069), .B2(n5068), .A(n5067), .ZN(n5071) );
  AOI22_X1 U5555 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5070) );
  XNOR2_X1 U5556 ( .A(n5071), .B(n5070), .ZN(U3352) );
endmodule

