

module b20_C_AntiSAT_k_128_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235;

  OR2_X1 U4821 ( .A1(n8592), .A2(n8591), .ZN(n8593) );
  OAI211_X1 U4822 ( .C1(n7822), .C2(n6476), .A(n6475), .B(n6474), .ZN(n8525)
         );
  OR2_X1 U4823 ( .A1(n6938), .A2(n7487), .ZN(n7207) );
  CLKBUF_X2 U4824 ( .A(n5122), .Z(n5695) );
  BUF_X1 U4825 ( .A(n7247), .Z(n4321) );
  INV_X4 U4826 ( .A(n6508), .ZN(n5846) );
  INV_X1 U4827 ( .A(n7060), .ZN(n8756) );
  INV_X1 U4828 ( .A(n6133), .ZN(n6229) );
  BUF_X2 U4829 ( .A(n5122), .Z(n5281) );
  INV_X1 U4830 ( .A(n6004), .ZN(n6180) );
  CLKBUF_X1 U4831 ( .A(n5966), .Z(n6614) );
  NAND4_X1 U4832 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n6526)
         );
  AND2_X1 U4833 ( .A1(n5462), .A2(n8394), .ZN(n8451) );
  INV_X2 U4834 ( .A(n5515), .ZN(n4324) );
  INV_X1 U4835 ( .A(n4317), .ZN(n4319) );
  INV_X4 U4836 ( .A(n6632), .ZN(n6631) );
  NAND2_X1 U4837 ( .A1(n5727), .A2(n9796), .ZN(n5125) );
  CLKBUF_X1 U4838 ( .A(n9052), .Z(n4315) );
  NOR2_X1 U4839 ( .A1(n6970), .A2(n8937), .ZN(n9052) );
  OR2_X1 U4840 ( .A1(n6902), .A2(n7098), .ZN(n4338) );
  NOR2_X1 U4842 ( .A1(n6270), .A2(n6269), .ZN(n6291) );
  INV_X1 U4843 ( .A(n5125), .ZN(n5151) );
  INV_X1 U4844 ( .A(n7064), .ZN(n8564) );
  INV_X1 U4845 ( .A(n8589), .ZN(n4802) );
  AND2_X1 U4846 ( .A1(n5125), .A2(n6632), .ZN(n5146) );
  INV_X1 U4847 ( .A(n4317), .ZN(n4320) );
  INV_X1 U4848 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5243) );
  INV_X1 U4849 ( .A(n8924), .ZN(n8713) );
  INV_X1 U4850 ( .A(n6614), .ZN(n6880) );
  NAND2_X1 U4851 ( .A1(n5812), .A2(n5811), .ZN(n6234) );
  AND3_X1 U4852 ( .A1(n5990), .A2(n5992), .A3(n5991), .ZN(n9926) );
  OR2_X2 U4853 ( .A1(n5987), .A2(n4325), .ZN(n5989) );
  NAND2_X1 U4854 ( .A1(n5436), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5021) );
  AND2_X1 U4855 ( .A1(n5208), .A2(n5207), .ZN(n7326) );
  INV_X1 U4856 ( .A(n4936), .ZN(n6632) );
  AND2_X1 U4857 ( .A1(n5859), .A2(n5858), .ZN(n8718) );
  NOR2_X1 U4858 ( .A1(n7772), .A2(n6102), .ZN(n7933) );
  NAND2_X1 U4859 ( .A1(n4460), .A2(n6077), .ZN(n7436) );
  NAND2_X1 U4860 ( .A1(n5547), .A2(n9198), .ZN(n9197) );
  AOI211_X1 U4861 ( .C1(n6700), .C2(n6699), .A(n9387), .B(n6722), .ZN(n6709)
         );
  INV_X1 U4862 ( .A(n7379), .ZN(n5178) );
  OAI22_X1 U4863 ( .A1(n9513), .A2(n6553), .B1(n9270), .B2(n9518), .ZN(n9496)
         );
  AOI21_X1 U4864 ( .B1(n9589), .B2(n9328), .A(n6550), .ZN(n9560) );
  INV_X1 U4865 ( .A(n9624), .ZN(n9620) );
  XNOR2_X1 U4866 ( .A(n6234), .B(P2_REG3_REG_26__SCAN_IN), .ZN(n8917) );
  AND3_X1 U4867 ( .A1(n5973), .A2(n5972), .A3(n5971), .ZN(n4316) );
  NAND2_X2 U4868 ( .A1(n7867), .A2(n7868), .ZN(n7866) );
  NAND2_X2 U4869 ( .A1(n7923), .A2(n5339), .ZN(n7867) );
  AOI21_X2 U4870 ( .B1(n4671), .B2(n4670), .A(n4667), .ZN(n8662) );
  NOR2_X2 U4871 ( .A1(n5035), .A2(n5034), .ZN(n5119) );
  NOR2_X2 U4872 ( .A1(n7689), .A2(n7699), .ZN(n7688) );
  OAI21_X2 U4874 ( .B1(n5575), .B2(n4597), .A(n9249), .ZN(n9250) );
  INV_X1 U4875 ( .A(n5151), .ZN(n4317) );
  INV_X1 U4876 ( .A(n4317), .ZN(n4318) );
  NAND3_X2 U4877 ( .A1(n5121), .A2(n4915), .A3(n5120), .ZN(n6524) );
  AND2_X2 U4878 ( .A1(n8068), .A2(n8067), .ZN(n8469) );
  NAND2_X2 U4879 ( .A1(n5092), .A2(n5091), .ZN(n7524) );
  XNOR2_X2 U4880 ( .A(n8479), .B(n9582), .ZN(n8491) );
  OR2_X2 U4881 ( .A1(n9388), .A2(n8478), .ZN(n8479) );
  AOI21_X2 U4882 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6727), .A(n6722), .ZN(
        n6726) );
  NOR2_X2 U4883 ( .A1(n6700), .A2(n6699), .ZN(n6722) );
  AOI21_X2 U4884 ( .B1(n8012), .B2(n9331), .A(n6547), .ZN(n8161) );
  INV_X2 U4885 ( .A(n5515), .ZN(n4322) );
  XNOR2_X2 U4886 ( .A(n5989), .B(n5988), .ZN(n6895) );
  XNOR2_X2 U4887 ( .A(n5965), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6897) );
  OAI21_X2 U4889 ( .B1(n5012), .B2(n5000), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5001) );
  AND2_X2 U4890 ( .A1(n8464), .A2(n5462), .ZN(n6562) );
  OR2_X1 U4891 ( .A1(n9546), .A2(n9545), .ZN(n9548) );
  OR2_X2 U4892 ( .A1(n9122), .A2(n8713), .ZN(n6375) );
  AND2_X1 U4893 ( .A1(n6749), .A2(n5134), .ZN(n6771) );
  INV_X1 U4894 ( .A(n7243), .ZN(n9940) );
  CLKBUF_X1 U4895 ( .A(n5303), .Z(n5697) );
  INV_X1 U4896 ( .A(n6185), .ZN(n6237) );
  CLKBUF_X2 U4897 ( .A(n5065), .Z(n5640) );
  CLKBUF_X1 U4898 ( .A(n5065), .Z(n5619) );
  CLKBUF_X2 U4899 ( .A(n5996), .Z(n6141) );
  AND3_X1 U4900 ( .A1(n5969), .A2(n5968), .A3(n5967), .ZN(n7267) );
  INV_X1 U4901 ( .A(n7321), .ZN(n6525) );
  CLKBUF_X3 U4902 ( .A(n5980), .Z(n6282) );
  OR2_X2 U4903 ( .A1(n5128), .A2(n5022), .ZN(n5690) );
  OR2_X1 U4905 ( .A1(n6409), .A2(n5723), .ZN(n5753) );
  OR3_X1 U4906 ( .A1(n8903), .A2(n9007), .A3(n8902), .ZN(n8906) );
  NOR2_X1 U4907 ( .A1(n4482), .A2(n9432), .ZN(n4481) );
  NAND2_X1 U4908 ( .A1(n4657), .A2(n4661), .ZN(n8574) );
  OAI21_X1 U4909 ( .B1(n4480), .B2(n4479), .A(n8458), .ZN(n4478) );
  NAND2_X1 U4910 ( .A1(n4630), .A2(n4352), .ZN(n9454) );
  AND2_X1 U4911 ( .A1(n9469), .A2(n9470), .ZN(n9471) );
  NAND2_X1 U4912 ( .A1(n4581), .A2(n4584), .ZN(n9280) );
  NAND2_X1 U4913 ( .A1(n5872), .A2(n5871), .ZN(n9122) );
  AND2_X1 U4914 ( .A1(n9479), .A2(n8366), .ZN(n9504) );
  NAND2_X1 U4915 ( .A1(n6231), .A2(n6230), .ZN(n9127) );
  NAND2_X1 U4916 ( .A1(n5851), .A2(n5850), .ZN(n9116) );
  NAND2_X1 U4917 ( .A1(n6219), .A2(n6218), .ZN(n9133) );
  NAND2_X1 U4918 ( .A1(n5586), .A2(n5585), .ZN(n6564) );
  AND2_X1 U4919 ( .A1(n4620), .A2(n4619), .ZN(n8797) );
  AND2_X1 U4920 ( .A1(n6583), .A2(n8265), .ZN(n8162) );
  NAND2_X1 U4921 ( .A1(n5557), .A2(n5556), .ZN(n6589) );
  OAI21_X1 U4922 ( .B1(n7896), .B2(n6443), .A(n6442), .ZN(n8100) );
  AND3_X1 U4923 ( .A1(n4691), .A2(n4692), .A3(n4402), .ZN(n8782) );
  NAND2_X1 U4924 ( .A1(n6206), .A2(n6205), .ZN(n9085) );
  OR2_X1 U4925 ( .A1(n7908), .A2(n7909), .ZN(n8003) );
  OAI21_X1 U4926 ( .B1(n5550), .B2(n5549), .A(n5548), .ZN(n5577) );
  NAND2_X1 U4927 ( .A1(n8052), .A2(n4617), .ZN(n8119) );
  NAND2_X1 U4928 ( .A1(n7683), .A2(n7684), .ZN(n7792) );
  NAND2_X1 U4929 ( .A1(n5911), .A2(n5910), .ZN(n9168) );
  INV_X1 U4930 ( .A(n9318), .ZN(n8012) );
  OR2_X1 U4931 ( .A1(n6348), .A2(n6147), .ZN(n8147) );
  XNOR2_X1 U4932 ( .A(n4689), .B(n7938), .ZN(n7772) );
  AND2_X1 U4933 ( .A1(n5365), .A2(n5364), .ZN(n9318) );
  NAND2_X1 U4934 ( .A1(n5927), .A2(n5926), .ZN(n8542) );
  INV_X1 U4935 ( .A(n8257), .ZN(n8414) );
  OR2_X1 U4936 ( .A1(n7699), .A2(n6541), .ZN(n8247) );
  AND2_X1 U4937 ( .A1(n7813), .A2(n6544), .ZN(n8257) );
  NAND2_X1 U4938 ( .A1(n5320), .A2(n5319), .ZN(n7699) );
  NAND2_X1 U4939 ( .A1(n5930), .A2(n5929), .ZN(n8537) );
  NAND2_X1 U4940 ( .A1(n5350), .A2(n5349), .ZN(n9702) );
  NAND2_X1 U4941 ( .A1(n4996), .A2(n4995), .ZN(n7813) );
  NAND2_X1 U4942 ( .A1(n6136), .A2(n6135), .ZN(n8111) );
  AND2_X1 U4943 ( .A1(n8220), .A2(n8333), .ZN(n8223) );
  NAND2_X1 U4944 ( .A1(n4972), .A2(n4971), .ZN(n5343) );
  NAND2_X1 U4945 ( .A1(n5074), .A2(n5073), .ZN(n7889) );
  NAND2_X1 U4946 ( .A1(n6058), .A2(n6057), .ZN(n9969) );
  AND3_X1 U4947 ( .A1(n5958), .A2(n5957), .A3(n5956), .ZN(n9951) );
  NAND2_X1 U4948 ( .A1(n5133), .A2(n4912), .ZN(n6751) );
  OR2_X1 U4949 ( .A1(n7455), .A2(n7454), .ZN(n7581) );
  NOR2_X1 U4950 ( .A1(n4654), .A2(n4652), .ZN(n4651) );
  AND2_X1 U4951 ( .A1(n5224), .A2(n5223), .ZN(n6955) );
  AND2_X1 U4952 ( .A1(n5127), .A2(n5126), .ZN(n5133) );
  NAND2_X1 U4953 ( .A1(n5240), .A2(n5239), .ZN(n5242) );
  AND4_X1 U4954 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n7253)
         );
  INV_X1 U4955 ( .A(n7254), .ZN(n8759) );
  NAND4_X1 U4956 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n9343)
         );
  NAND4_X1 U4957 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), .ZN(n9342)
         );
  NAND4_X2 U4958 ( .A1(n5986), .A2(n5985), .A3(n5984), .A4(n5983), .ZN(n8758)
         );
  NAND4_X1 U4959 ( .A1(n5144), .A2(n5143), .A3(n5142), .A4(n5141), .ZN(n9344)
         );
  INV_X1 U4960 ( .A(n9835), .ZN(n6963) );
  AND2_X1 U4961 ( .A1(n5118), .A2(n5117), .ZN(n4915) );
  NAND2_X1 U4962 ( .A1(n5041), .A2(n5040), .ZN(n5065) );
  AND3_X2 U4963 ( .A1(n5156), .A2(n5155), .A3(n5154), .ZN(n9835) );
  AND3_X2 U4964 ( .A1(n6617), .A2(P1_STATE_REG_SCAN_IN), .A3(n5128), .ZN(
        P1_U3973) );
  CLKBUF_X1 U4965 ( .A(n5469), .Z(n5731) );
  INV_X4 U4966 ( .A(n5442), .ZN(n5140) );
  NAND3_X1 U4967 ( .A1(n5112), .A2(n5113), .A3(n4521), .ZN(n7321) );
  INV_X1 U4968 ( .A(n5690), .ZN(n5122) );
  NAND2_X1 U4969 ( .A1(n5966), .A2(n6632), .ZN(n6133) );
  BUF_X4 U4970 ( .A(n5146), .Z(n4326) );
  INV_X4 U4971 ( .A(n5469), .ZN(n4323) );
  NAND2_X1 U4972 ( .A1(n9176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U4973 ( .A1(n5125), .A2(n6631), .ZN(n5316) );
  AND2_X2 U4974 ( .A1(n5700), .A2(n5005), .ZN(n5128) );
  NAND2_X1 U4975 ( .A1(n5820), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5822) );
  AND2_X1 U4976 ( .A1(n5015), .A2(n5717), .ZN(n8464) );
  NAND2_X1 U4977 ( .A1(n5031), .A2(n5030), .ZN(n5035) );
  XNOR2_X1 U4978 ( .A(n5002), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8197) );
  XNOR2_X1 U4979 ( .A(n5004), .B(P1_IR_REG_25__SCAN_IN), .ZN(n8175) );
  XNOR2_X1 U4980 ( .A(n5007), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5719) );
  AND2_X1 U4981 ( .A1(n5817), .A2(n5776), .ZN(n4854) );
  NAND2_X1 U4982 ( .A1(n4987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U4983 ( .A1(n5006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U4984 ( .A1(n5017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5415) );
  NAND2_X2 U4985 ( .A1(n6631), .A2(P1_U3086), .ZN(n9792) );
  AND2_X1 U4986 ( .A1(n5016), .A2(n4997), .ZN(n5008) );
  AND2_X1 U4987 ( .A1(n5780), .A2(n5779), .ZN(n5815) );
  CLKBUF_X1 U4988 ( .A(n4990), .Z(n5199) );
  AND2_X1 U4989 ( .A1(n5778), .A2(n5777), .ZN(n5779) );
  BUF_X2 U4990 ( .A(n6895), .Z(n7026) );
  AND3_X1 U4991 ( .A1(n4723), .A2(n4330), .A3(n4722), .ZN(n5016) );
  NOR2_X1 U4992 ( .A1(n5898), .A2(n5773), .ZN(n5774) );
  NAND4_X1 U4993 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n5898)
         );
  AND2_X1 U4994 ( .A1(n5152), .A2(n4514), .ZN(n4990) );
  AND4_X1 U4995 ( .A1(n5152), .A2(n4976), .A3(n4977), .A4(n4721), .ZN(n4722)
         );
  AND2_X1 U4996 ( .A1(n4976), .A2(n4977), .ZN(n4514) );
  AND2_X1 U4997 ( .A1(n6390), .A2(n5782), .ZN(n5780) );
  NAND3_X1 U4998 ( .A1(n8497), .A2(n4408), .A3(n4407), .ZN(n4754) );
  AND4_X1 U4999 ( .A1(n5346), .A2(n4975), .A3(n4992), .A4(n4974), .ZN(n4330)
         );
  AND3_X1 U5000 ( .A1(n4711), .A2(n4710), .A3(n4709), .ZN(n5770) );
  NAND3_X1 U5001 ( .A1(n4753), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4752) );
  INV_X1 U5002 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5018) );
  INV_X1 U5003 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8497) );
  INV_X1 U5004 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4753) );
  INV_X1 U5005 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4407) );
  INV_X1 U5006 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4992) );
  NOR2_X1 U5007 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4517) );
  INV_X1 U5008 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4998) );
  NOR2_X1 U5009 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4516) );
  NOR2_X1 U5010 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4518) );
  INV_X1 U5011 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4999) );
  INV_X1 U5012 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5346) );
  BUF_X1 U5013 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9798) );
  NOR2_X1 U5014 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5767) );
  NOR2_X1 U5015 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5768) );
  NOR2_X1 U5016 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5769) );
  INV_X1 U5017 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4709) );
  INV_X1 U5018 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4710) );
  INV_X1 U5019 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4711) );
  INV_X1 U5020 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10173) );
  INV_X1 U5021 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5818) );
  INV_X4 U5022 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X2 U5023 ( .A1(n9535), .A2(n6589), .ZN(n9516) );
  OAI21_X1 U5024 ( .B1(n4549), .B2(n4546), .A(n6354), .ZN(n6157) );
  NAND2_X2 U5025 ( .A1(n9122), .A2(n8713), .ZN(n6374) );
  NAND2_X1 U5026 ( .A1(n5034), .A2(n5035), .ZN(n5515) );
  XNOR2_X2 U5027 ( .A(n6418), .B(n6467), .ZN(n6476) );
  INV_X1 U5028 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4325) );
  OAI21_X2 U5029 ( .B1(n9280), .B2(n9276), .A(n9277), .ZN(n8514) );
  NOR2_X2 U5030 ( .A1(n7207), .A2(n9818), .ZN(n7500) );
  OAI22_X2 U5031 ( .A1(n9197), .A2(n5574), .B1(n9198), .B2(n5573), .ZN(n5575)
         );
  INV_X1 U5032 ( .A(n5119), .ZN(n5469) );
  NAND2_X1 U5033 ( .A1(n8279), .A2(n8427), .ZN(n8272) );
  INV_X1 U5034 ( .A(n8295), .ZN(n8298) );
  INV_X1 U5035 ( .A(n5406), .ZN(n5407) );
  OR2_X1 U5036 ( .A1(n9156), .A2(n9011), .ZN(n6358) );
  OR2_X1 U5037 ( .A1(n6714), .A2(n6493), .ZN(n6510) );
  AND2_X1 U5038 ( .A1(n8448), .A2(n8321), .ZN(n4773) );
  INV_X1 U5039 ( .A(n8322), .ZN(n4772) );
  CLKBUF_X1 U5040 ( .A(n5442), .Z(n5728) );
  OR2_X1 U5041 ( .A1(n9554), .A2(n9269), .ZN(n8436) );
  AOI21_X1 U5042 ( .B1(n4872), .B2(n4870), .A(n4373), .ZN(n4869) );
  INV_X1 U5043 ( .A(n4873), .ZN(n4870) );
  OAI21_X1 U5044 ( .B1(n5453), .B2(n4783), .A(n5456), .ZN(n5483) );
  INV_X1 U5045 ( .A(n5454), .ZN(n4783) );
  NAND2_X1 U5046 ( .A1(n4545), .A2(n4351), .ZN(n4412) );
  INV_X1 U5047 ( .A(n5288), .ZN(n4413) );
  OAI211_X1 U5048 ( .C1(n4476), .C2(n4475), .A(n6340), .B(n4474), .ZN(n6341)
         );
  NAND2_X1 U5049 ( .A1(n4477), .A2(n4826), .ZN(n4476) );
  AND3_X1 U5050 ( .A1(n5423), .A2(n5422), .A3(n5421), .ZN(n9282) );
  INV_X1 U5051 ( .A(n5034), .ZN(n4563) );
  NAND2_X1 U5052 ( .A1(n4856), .A2(n4855), .ZN(n9513) );
  AOI21_X1 U5053 ( .B1(n4858), .B2(n4860), .A(n4372), .ZN(n4855) );
  AOI21_X1 U5054 ( .B1(n8279), .B2(n8430), .A(n8278), .ZN(n8280) );
  AOI21_X1 U5055 ( .B1(n6204), .B2(n5846), .A(n6215), .ZN(n4554) );
  NAND2_X1 U5056 ( .A1(n6203), .A2(n6508), .ZN(n4555) );
  NOR2_X1 U5057 ( .A1(n4503), .A2(n4502), .ZN(n8295) );
  INV_X1 U5058 ( .A(n8294), .ZN(n4502) );
  AOI21_X1 U5059 ( .B1(n8291), .B2(n8290), .A(n4504), .ZN(n4503) );
  OR2_X1 U5060 ( .A1(n6250), .A2(n8900), .ZN(n4562) );
  INV_X1 U5061 ( .A(n5783), .ZN(n5788) );
  AND2_X1 U5062 ( .A1(n5836), .A2(n5782), .ZN(n5839) );
  INV_X1 U5063 ( .A(n5338), .ZN(n4716) );
  AOI21_X1 U5064 ( .B1(n4572), .B2(n5358), .A(n9187), .ZN(n4571) );
  INV_X1 U5065 ( .A(n4788), .ZN(n4787) );
  OAI21_X1 U5066 ( .B1(n5675), .B2(n4789), .A(n5754), .ZN(n4788) );
  AOI21_X1 U5067 ( .B1(n4775), .B2(n4779), .A(n4427), .ZN(n4426) );
  INV_X1 U5068 ( .A(n5648), .ZN(n4427) );
  NAND2_X1 U5069 ( .A1(n5343), .A2(n4396), .ZN(n4794) );
  NAND2_X1 U5070 ( .A1(n5359), .A2(SI_14_), .ZN(n4796) );
  INV_X1 U5071 ( .A(n9184), .ZN(n5823) );
  OAI21_X1 U5072 ( .B1(n4847), .B2(n4846), .A(n7417), .ZN(n4844) );
  AND2_X1 U5073 ( .A1(n9138), .A2(n8935), .ZN(n6367) );
  OR2_X1 U5074 ( .A1(n9085), .A2(n8985), .ZN(n6362) );
  OR2_X1 U5075 ( .A1(n8700), .A2(n8997), .ZN(n6357) );
  NAND2_X1 U5076 ( .A1(n9174), .A2(n6967), .ZN(n6821) );
  INV_X1 U5077 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5988) );
  INV_X1 U5078 ( .A(n4720), .ZN(n4592) );
  NAND2_X1 U5079 ( .A1(n4719), .A2(n4718), .ZN(n4717) );
  NAND2_X1 U5080 ( .A1(n7748), .A2(n5308), .ZN(n4718) );
  OAI21_X1 U5081 ( .B1(n9610), .B2(n4633), .A(n4631), .ZN(n6586) );
  INV_X1 U5082 ( .A(n4632), .ZN(n4631) );
  OAI21_X1 U5083 ( .B1(n4329), .B2(n4633), .A(n9579), .ZN(n4632) );
  OR2_X1 U5084 ( .A1(n9404), .A2(n8309), .ZN(n8354) );
  AND2_X1 U5085 ( .A1(n4438), .A2(n4437), .ZN(n6275) );
  NAND2_X1 U5086 ( .A1(n5759), .A2(n5760), .ZN(n4437) );
  NAND2_X1 U5087 ( .A1(n4441), .A2(n4439), .ZN(n4438) );
  OAI21_X1 U5088 ( .B1(n5483), .B2(n5482), .A(n5481), .ZN(n5505) );
  NOR2_X1 U5089 ( .A1(n5430), .A2(n4800), .ZN(n4799) );
  INV_X1 U5090 ( .A(n5408), .ZN(n4800) );
  AND2_X1 U5091 ( .A1(n4450), .A2(n4922), .ZN(n5109) );
  NAND2_X1 U5092 ( .A1(n4936), .A2(n5123), .ZN(n4922) );
  INV_X1 U5093 ( .A(n4451), .ZN(n4450) );
  OR2_X1 U5094 ( .A1(n7045), .A2(n7044), .ZN(n7047) );
  OR2_X1 U5095 ( .A1(n5845), .A2(n8741), .ZN(n6383) );
  INV_X1 U5096 ( .A(n6141), .ZN(n6235) );
  NAND2_X1 U5098 ( .A1(n7590), .A2(n7591), .ZN(n9901) );
  NAND2_X1 U5099 ( .A1(n7939), .A2(n7940), .ZN(n7941) );
  NAND2_X1 U5100 ( .A1(n7941), .A2(n7942), .ZN(n8052) );
  XNOR2_X1 U5101 ( .A(n8119), .B(n8124), .ZN(n8054) );
  NAND2_X1 U5102 ( .A1(n8054), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8120) );
  INV_X1 U5103 ( .A(n6232), .ZN(n5812) );
  INV_X1 U5104 ( .A(n8750), .ZN(n7900) );
  NAND2_X1 U5105 ( .A1(n7428), .A2(n7424), .ZN(n4744) );
  AND4_X1 U5106 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n7429)
         );
  OAI21_X1 U5107 ( .B1(n8944), .B2(n6460), .A(n6459), .ZN(n8933) );
  OR2_X1 U5108 ( .A1(n6457), .A2(n8968), .ZN(n6365) );
  OR2_X1 U5109 ( .A1(n9089), .A2(n8998), .ZN(n6360) );
  NAND2_X1 U5110 ( .A1(n8994), .A2(n6452), .ZN(n9000) );
  AOI21_X1 U5111 ( .B1(n4815), .B2(n4817), .A(n4813), .ZN(n4812) );
  INV_X1 U5112 ( .A(n4816), .ZN(n4815) );
  NAND2_X1 U5113 ( .A1(n6481), .A2(n6480), .ZN(n6714) );
  INV_X1 U5114 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U5115 ( .A1(n5558), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5610) );
  AND2_X1 U5116 ( .A1(n9293), .A2(n9290), .ZN(n5647) );
  OR2_X1 U5117 ( .A1(n4327), .A2(n8388), .ZN(n4436) );
  INV_X1 U5118 ( .A(n8324), .ZN(n4501) );
  AND2_X1 U5119 ( .A1(n5616), .A2(n5615), .ZN(n9254) );
  AND2_X1 U5120 ( .A1(n5518), .A2(n5517), .ZN(n9269) );
  AND2_X1 U5121 ( .A1(n5495), .A2(n5494), .ZN(n9211) );
  OR2_X1 U5122 ( .A1(n9361), .A2(n9360), .ZN(n4601) );
  NAND2_X1 U5123 ( .A1(n9462), .A2(n4522), .ZN(n9439) );
  NOR2_X1 U5124 ( .A1(n9404), .A2(n4523), .ZN(n4522) );
  INV_X1 U5125 ( .A(n4524), .ZN(n4523) );
  AOI21_X1 U5126 ( .B1(n4873), .B2(n6584), .A(n4374), .ZN(n4872) );
  INV_X1 U5127 ( .A(n9584), .ZN(n9616) );
  AOI21_X1 U5128 ( .B1(n4897), .B2(n4894), .A(n4332), .ZN(n4893) );
  INV_X1 U5129 ( .A(n4902), .ZN(n4894) );
  AOI21_X1 U5130 ( .B1(n9754), .B2(n9283), .A(n9578), .ZN(n6550) );
  INV_X2 U5131 ( .A(n5316), .ZN(n8313) );
  INV_X1 U5132 ( .A(n9609), .ZN(n9846) );
  INV_X1 U5133 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U5134 ( .A1(n9780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5025) );
  OAI21_X1 U5135 ( .B1(n4412), .B2(n4411), .A(n4375), .ZN(n5048) );
  INV_X1 U5136 ( .A(n5087), .ZN(n4411) );
  AND2_X1 U5137 ( .A1(n4962), .A2(n4960), .ZN(n4797) );
  OR3_X1 U5138 ( .A1(n8095), .A2(n8178), .A3(n8200), .ZN(n6884) );
  INV_X1 U5139 ( .A(n8753), .ZN(n7758) );
  INV_X1 U5140 ( .A(P2_U3893), .ZN(n8841) );
  INV_X1 U5141 ( .A(n9902), .ZN(n8840) );
  OR2_X1 U5142 ( .A1(n7936), .A2(n7935), .ZN(n4540) );
  NAND2_X1 U5143 ( .A1(n4559), .A2(n4558), .ZN(n6065) );
  NAND2_X1 U5144 ( .A1(n6339), .A2(n5846), .ZN(n4558) );
  AOI21_X1 U5145 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n4493) );
  AND2_X1 U5146 ( .A1(n8248), .A2(n8249), .ZN(n4492) );
  NAND2_X1 U5147 ( .A1(n8270), .A2(n9318), .ZN(n8262) );
  OAI21_X1 U5148 ( .B1(n8258), .B2(n8257), .A(n8419), .ZN(n8260) );
  OAI21_X1 U5149 ( .B1(n6548), .B2(n8164), .A(n4781), .ZN(n8270) );
  INV_X1 U5150 ( .A(n4782), .ZN(n4781) );
  OAI21_X1 U5151 ( .B1(n9242), .B2(n8164), .A(n8458), .ZN(n4782) );
  NAND2_X1 U5152 ( .A1(n8264), .A2(n8319), .ZN(n4509) );
  INV_X1 U5153 ( .A(n6156), .ZN(n4548) );
  AOI21_X1 U5154 ( .B1(n4790), .B2(n4791), .A(n8285), .ZN(n4513) );
  AOI21_X1 U5155 ( .B1(n8280), .B2(n8458), .A(n8282), .ZN(n4790) );
  NAND2_X1 U5156 ( .A1(n4792), .A2(n8319), .ZN(n4791) );
  INV_X1 U5157 ( .A(n8284), .ZN(n4512) );
  INV_X1 U5158 ( .A(n6214), .ZN(n4553) );
  AOI21_X1 U5159 ( .B1(n8306), .B2(n9431), .A(n8458), .ZN(n4482) );
  NOR2_X1 U5160 ( .A1(n8297), .A2(n8379), .ZN(n4480) );
  OR2_X1 U5161 ( .A1(n8900), .A2(n6256), .ZN(n6257) );
  OR2_X1 U5162 ( .A1(n6246), .A2(n8900), .ZN(n4561) );
  NOR2_X1 U5163 ( .A1(n6075), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6056) );
  INV_X1 U5164 ( .A(n4651), .ZN(n4485) );
  NOR2_X1 U5165 ( .A1(n6588), .A2(n4643), .ZN(n4642) );
  INV_X1 U5166 ( .A(n8283), .ZN(n4643) );
  INV_X1 U5167 ( .A(n5677), .ZN(n4789) );
  NAND2_X1 U5168 ( .A1(n5459), .A2(n5458), .ZN(n5481) );
  NAND2_X1 U5169 ( .A1(n8652), .A2(n4669), .ZN(n4668) );
  INV_X1 U5170 ( .A(n8545), .ZN(n4669) );
  AND2_X1 U5171 ( .A1(n4662), .A2(n8571), .ZN(n4661) );
  NAND2_X1 U5172 ( .A1(n6898), .A2(n6900), .ZN(n9882) );
  NAND2_X1 U5173 ( .A1(n4533), .A2(n4368), .ZN(n4532) );
  NOR2_X1 U5174 ( .A1(n8809), .A2(n4621), .ZN(n8845) );
  NOR2_X1 U5175 ( .A1(n8806), .A2(n9048), .ZN(n4621) );
  NOR2_X1 U5176 ( .A1(n8817), .A2(n4530), .ZN(n8830) );
  NOR2_X1 U5177 ( .A1(n8806), .A2(n9104), .ZN(n4530) );
  AOI21_X1 U5178 ( .B1(n4728), .B2(n4730), .A(n4377), .ZN(n4727) );
  INV_X1 U5179 ( .A(n4728), .ZN(n4725) );
  INV_X1 U5180 ( .A(n4731), .ZN(n4730) );
  AOI21_X1 U5181 ( .B1(n4731), .B2(n4729), .A(n4734), .ZN(n4728) );
  INV_X1 U5182 ( .A(n6465), .ZN(n4729) );
  AND2_X1 U5183 ( .A1(n9116), .A2(n8914), .ZN(n4734) );
  INV_X1 U5184 ( .A(n4707), .ZN(n4706) );
  OAI21_X1 U5185 ( .B1(n9040), .B2(n4708), .A(n6449), .ZN(n4707) );
  INV_X1 U5186 ( .A(n6448), .ZN(n4708) );
  NOR2_X1 U5187 ( .A1(n4845), .A2(n4846), .ZN(n4842) );
  NAND2_X1 U5188 ( .A1(n7254), .A2(n7267), .ZN(n6420) );
  AND2_X1 U5189 ( .A1(n8900), .A2(n4346), .ZN(n4731) );
  NAND2_X1 U5190 ( .A1(n9116), .A2(n8718), .ZN(n6376) );
  OR2_X1 U5191 ( .A1(n9116), .A2(n8718), .ZN(n6377) );
  NAND2_X1 U5192 ( .A1(n6366), .A2(n4831), .ZN(n4473) );
  NAND2_X1 U5193 ( .A1(n4831), .A2(n4829), .ZN(n4472) );
  AND2_X1 U5194 ( .A1(n4830), .A2(n6368), .ZN(n4834) );
  OR2_X1 U5195 ( .A1(n8955), .A2(n8953), .ZN(n6456) );
  NAND2_X1 U5196 ( .A1(n8101), .A2(n6444), .ZN(n4742) );
  OR2_X1 U5197 ( .A1(n8111), .A2(n8532), .ZN(n6347) );
  INV_X1 U5198 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U5199 ( .A1(n5776), .A2(n4686), .ZN(n4750) );
  NAND2_X1 U5200 ( .A1(n5790), .A2(n5789), .ZN(n6404) );
  NOR2_X1 U5201 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  NOR2_X1 U5202 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  INV_X1 U5203 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6390) );
  INV_X1 U5204 ( .A(n5839), .ZN(n6389) );
  INV_X1 U5205 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U5206 ( .A1(n4590), .A2(n4716), .ZN(n4587) );
  NAND2_X1 U5207 ( .A1(n4716), .A2(n5307), .ZN(n4588) );
  AND2_X1 U5208 ( .A1(n9262), .A2(n4713), .ZN(n4712) );
  NAND2_X1 U5209 ( .A1(n8517), .A2(n8515), .ZN(n4713) );
  NAND2_X1 U5210 ( .A1(n5719), .A2(n8394), .ZN(n5022) );
  NAND2_X1 U5211 ( .A1(n7474), .A2(n5306), .ZN(n4720) );
  NAND2_X1 U5212 ( .A1(n4571), .A2(n4573), .ZN(n4569) );
  OR2_X1 U5213 ( .A1(n8320), .A2(n8382), .ZN(n8448) );
  NOR2_X1 U5214 ( .A1(n9720), .A2(n9648), .ZN(n4526) );
  NOR2_X1 U5215 ( .A1(n5631), .A2(n9298), .ZN(n5683) );
  INV_X1 U5216 ( .A(n4642), .ZN(n4636) );
  AND2_X1 U5217 ( .A1(n6537), .A2(n8236), .ZN(n8335) );
  OAI21_X1 U5218 ( .B1(n7498), .B2(n4883), .A(n4882), .ZN(n4881) );
  INV_X1 U5219 ( .A(n4881), .ZN(n4880) );
  INV_X1 U5220 ( .A(n9451), .ZN(n4891) );
  NOR2_X1 U5221 ( .A1(n4898), .A2(n4900), .ZN(n4897) );
  OR2_X1 U5222 ( .A1(n6557), .A2(n4901), .ZN(n4898) );
  OR2_X1 U5223 ( .A1(n9493), .A2(n9254), .ZN(n8359) );
  NAND2_X1 U5224 ( .A1(n9532), .A2(n8289), .ZN(n4641) );
  INV_X1 U5225 ( .A(n4872), .ZN(n4871) );
  NOR2_X1 U5226 ( .A1(n4888), .A2(n8342), .ZN(n4885) );
  INV_X1 U5227 ( .A(n4906), .ZN(n4888) );
  OR2_X1 U5228 ( .A1(n9191), .A2(n8253), .ZN(n4906) );
  INV_X1 U5229 ( .A(n6546), .ZN(n4887) );
  NAND2_X1 U5230 ( .A1(n4424), .A2(n4422), .ZN(n5676) );
  AOI21_X1 U5231 ( .B1(n4426), .B2(n4428), .A(n4423), .ZN(n4422) );
  INV_X1 U5232 ( .A(n5650), .ZN(n4423) );
  AND2_X1 U5233 ( .A1(n5677), .A2(n5654), .ZN(n5675) );
  NAND2_X1 U5234 ( .A1(n5503), .A2(n5504), .ZN(n4420) );
  OR2_X1 U5235 ( .A1(n5503), .A2(n5504), .ZN(n4421) );
  AND3_X1 U5236 ( .A1(n5018), .A2(n5433), .A3(n5020), .ZN(n4997) );
  INV_X1 U5237 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U5238 ( .A1(n4794), .A2(n4395), .ZN(n5384) );
  NAND2_X1 U5239 ( .A1(n4794), .A2(n4793), .ZN(n5380) );
  INV_X1 U5240 ( .A(n4795), .ZN(n4793) );
  NAND2_X1 U5241 ( .A1(n4967), .A2(SI_13_), .ZN(n5342) );
  NOR2_X1 U5242 ( .A1(n4964), .A2(SI_11_), .ZN(n4760) );
  AOI21_X1 U5243 ( .B1(n5262), .B2(n4767), .A(n4766), .ZN(n4765) );
  INV_X1 U5244 ( .A(n4952), .ZN(n4766) );
  AND2_X1 U5245 ( .A1(n5262), .A2(n5239), .ZN(n4764) );
  NAND2_X1 U5246 ( .A1(n7042), .A2(n7051), .ZN(n7050) );
  INV_X1 U5247 ( .A(n8760), .ZN(n7042) );
  NAND2_X1 U5248 ( .A1(n8568), .A2(n8567), .ZN(n8643) );
  NOR2_X1 U5249 ( .A1(n7367), .A2(n4678), .ZN(n4677) );
  INV_X1 U5250 ( .A(n7364), .ZN(n4678) );
  NOR2_X1 U5251 ( .A1(n7836), .A2(n4676), .ZN(n4675) );
  INV_X1 U5252 ( .A(n7224), .ZN(n4676) );
  NAND2_X1 U5253 ( .A1(n8549), .A2(n8701), .ZN(n8704) );
  INV_X1 U5254 ( .A(n8934), .ZN(n8717) );
  AND2_X1 U5255 ( .A1(n6496), .A2(n6516), .ZN(n6826) );
  AND4_X1 U5256 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n7219)
         );
  OR2_X1 U5257 ( .A1(n6240), .A2(n5970), .ZN(n5973) );
  NOR2_X1 U5258 ( .A1(n7167), .A2(n4531), .ZN(n7137) );
  NOR2_X1 U5259 ( .A1(n4532), .A2(n7155), .ZN(n4531) );
  AND2_X1 U5260 ( .A1(n4532), .A2(n7155), .ZN(n7167) );
  NAND2_X1 U5261 ( .A1(n9901), .A2(n9900), .ZN(n9899) );
  XNOR2_X1 U5262 ( .A(n7723), .B(n7718), .ZN(n7593) );
  NAND2_X1 U5263 ( .A1(n4535), .A2(n4534), .ZN(n7717) );
  NAND2_X1 U5264 ( .A1(n9907), .A2(n7584), .ZN(n4534) );
  AND2_X1 U5265 ( .A1(n4540), .A2(n4539), .ZN(n8123) );
  NAND2_X1 U5266 ( .A1(n8050), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4539) );
  OR2_X1 U5267 ( .A1(n8051), .A2(n4694), .ZN(n4691) );
  OR2_X1 U5268 ( .A1(n8127), .A2(n8107), .ZN(n4694) );
  NAND2_X1 U5269 ( .A1(n8126), .A2(n4693), .ZN(n4692) );
  INV_X1 U5270 ( .A(n8127), .ZN(n4693) );
  OR2_X1 U5271 ( .A1(n8053), .A2(n7948), .ZN(n4617) );
  NAND2_X1 U5272 ( .A1(n8769), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4619) );
  NOR2_X1 U5273 ( .A1(n6073), .A2(n5898), .ZN(n5908) );
  NAND2_X1 U5274 ( .A1(n8892), .A2(n6379), .ZN(n6418) );
  OR2_X1 U5275 ( .A1(n8894), .A2(n8895), .ZN(n8892) );
  XNOR2_X1 U5276 ( .A(n9062), .B(n8596), .ZN(n8895) );
  NAND2_X1 U5277 ( .A1(n5810), .A2(n5809), .ZN(n6232) );
  INV_X1 U5278 ( .A(n6220), .ZN(n5810) );
  OR2_X1 U5279 ( .A1(n5889), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U5280 ( .A1(n4818), .A2(n4821), .ZN(n6363) );
  NOR2_X1 U5281 ( .A1(n4823), .A2(n4361), .ZN(n4821) );
  NAND2_X1 U5282 ( .A1(n9014), .A2(n4465), .ZN(n4818) );
  AND3_X1 U5283 ( .A1(n6212), .A2(n6211), .A3(n6210), .ZN(n8985) );
  NAND2_X1 U5284 ( .A1(n9000), .A2(n4735), .ZN(n8980) );
  NOR2_X1 U5285 ( .A1(n8983), .A2(n4736), .ZN(n4735) );
  INV_X1 U5286 ( .A(n6453), .ZN(n4736) );
  AND4_X1 U5287 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n9009)
         );
  INV_X1 U5288 ( .A(n6449), .ZN(n9027) );
  OR2_X1 U5289 ( .A1(n6087), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U5290 ( .A1(n6438), .A2(n6437), .ZN(n7896) );
  OR2_X1 U5291 ( .A1(n6068), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6059) );
  AND2_X1 U5292 ( .A1(n6310), .A2(n6434), .ZN(n4743) );
  AND2_X1 U5293 ( .A1(n6309), .A2(n6339), .ZN(n7561) );
  OAI21_X1 U5294 ( .B1(n7416), .B2(n7429), .A(n9951), .ZN(n6433) );
  NOR2_X1 U5295 ( .A1(n6023), .A2(n6335), .ZN(n4847) );
  INV_X1 U5296 ( .A(n4849), .ZN(n4845) );
  INV_X1 U5297 ( .A(n6334), .ZN(n4846) );
  AND2_X1 U5298 ( .A1(n6336), .A2(n6306), .ZN(n7417) );
  NOR2_X1 U5299 ( .A1(n6332), .A2(n4850), .ZN(n4849) );
  NAND3_X1 U5300 ( .A1(n6429), .A2(n6430), .A3(n7285), .ZN(n7284) );
  OR2_X1 U5301 ( .A1(n5982), .A2(n5995), .ZN(n6000) );
  AND2_X1 U5302 ( .A1(n6821), .A2(n6511), .ZN(n6968) );
  AND2_X1 U5303 ( .A1(n4732), .A2(n4346), .ZN(n8901) );
  AND2_X1 U5304 ( .A1(n4732), .A2(n4731), .ZN(n8902) );
  INV_X1 U5305 ( .A(n6375), .ZN(n4810) );
  NAND2_X2 U5306 ( .A1(n6377), .A2(n6376), .ZN(n8900) );
  INV_X1 U5307 ( .A(n4834), .ZN(n4829) );
  AOI21_X1 U5308 ( .B1(n4833), .B2(n4834), .A(n4832), .ZN(n4831) );
  INV_X1 U5309 ( .A(n4837), .ZN(n4833) );
  NOR2_X1 U5310 ( .A1(n6367), .A2(n4838), .ZN(n4837) );
  INV_X1 U5311 ( .A(n6365), .ZN(n4838) );
  INV_X1 U5312 ( .A(n8923), .ZN(n8946) );
  NOR2_X1 U5313 ( .A1(n6367), .A2(n4835), .ZN(n4914) );
  NAND2_X1 U5314 ( .A1(n8959), .A2(n6364), .ZN(n6366) );
  NAND2_X1 U5315 ( .A1(n5879), .A2(n5878), .ZN(n6457) );
  NAND2_X1 U5316 ( .A1(n4825), .A2(n6359), .ZN(n8979) );
  NAND2_X1 U5317 ( .A1(n8992), .A2(n6358), .ZN(n4825) );
  AND3_X1 U5318 ( .A1(n6198), .A2(n6197), .A3(n6196), .ZN(n8998) );
  NAND2_X1 U5319 ( .A1(n6450), .A2(n4908), .ZN(n8994) );
  INV_X1 U5320 ( .A(n9041), .ZN(n9010) );
  NAND2_X1 U5321 ( .A1(n5902), .A2(n5901), .ZN(n9100) );
  OR2_X1 U5322 ( .A1(n8148), .A2(n6348), .ZN(n6350) );
  INV_X1 U5323 ( .A(n9012), .ZN(n9043) );
  AND2_X1 U5324 ( .A1(n7040), .A2(n6508), .ZN(n9041) );
  AND2_X1 U5325 ( .A1(n6347), .A2(n6346), .ZN(n8101) );
  OR2_X1 U5326 ( .A1(n4458), .A2(n6342), .ZN(n4457) );
  INV_X1 U5327 ( .A(n7436), .ZN(n9956) );
  NAND2_X1 U5328 ( .A1(n6497), .A2(n7046), .ZN(n9046) );
  AND2_X1 U5329 ( .A1(n6884), .A2(n6717), .ZN(n6841) );
  XNOR2_X1 U5330 ( .A(n5842), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7044) );
  AND2_X1 U5331 ( .A1(n6076), .A2(n6075), .ZN(n7598) );
  INV_X1 U5332 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6036) );
  INV_X1 U5333 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4679) );
  NOR2_X1 U5334 ( .A1(n5358), .A2(n4572), .ZN(n4570) );
  AND2_X1 U5335 ( .A1(n4580), .A2(n9210), .ZN(n4579) );
  OR2_X1 U5336 ( .A1(n4712), .A2(n5500), .ZN(n4580) );
  NAND2_X1 U5337 ( .A1(n9229), .A2(n9230), .ZN(n9228) );
  NAND2_X1 U5338 ( .A1(n4714), .A2(n4712), .ZN(n9260) );
  XNOR2_X1 U5339 ( .A(n5116), .B(n5640), .ZN(n5135) );
  NAND2_X1 U5340 ( .A1(n5145), .A2(n7321), .ZN(n5114) );
  NOR2_X1 U5341 ( .A1(n4585), .A2(n4583), .ZN(n4582) );
  INV_X1 U5342 ( .A(n9240), .ZN(n4585) );
  INV_X1 U5343 ( .A(n9230), .ZN(n4583) );
  OR3_X1 U5344 ( .A1(n6618), .A2(n5128), .A3(P1_U3086), .ZN(n8463) );
  AND2_X1 U5345 ( .A1(n5565), .A2(n5564), .ZN(n9270) );
  OR2_X1 U5346 ( .A1(n6664), .A2(n6663), .ZN(n4608) );
  NAND2_X1 U5347 ( .A1(n4608), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U5348 ( .A1(n6685), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4607) );
  AND2_X1 U5349 ( .A1(n4606), .A2(n4605), .ZN(n6743) );
  INV_X1 U5350 ( .A(n6744), .ZN(n4605) );
  AND2_X1 U5351 ( .A1(n4603), .A2(n4602), .ZN(n7991) );
  NAND2_X1 U5352 ( .A1(n7996), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4602) );
  NAND2_X1 U5353 ( .A1(n4343), .A2(n9374), .ZN(n8475) );
  OR2_X1 U5354 ( .A1(n9720), .A2(n9295), .ZN(n9429) );
  OR2_X1 U5355 ( .A1(n6564), .A2(n9221), .ZN(n9479) );
  NAND2_X1 U5356 ( .A1(n9610), .A2(n4329), .ZN(n9593) );
  NOR2_X1 U5357 ( .A1(n4876), .A2(n6549), .ZN(n4873) );
  AND2_X1 U5358 ( .A1(n8210), .A2(n8237), .ZN(n8341) );
  OR2_X1 U5359 ( .A1(n7351), .A2(n7356), .ZN(n7349) );
  OR2_X1 U5360 ( .A1(n7524), .A2(n9337), .ZN(n6535) );
  NAND2_X1 U5361 ( .A1(n7499), .A2(n7498), .ZN(n7497) );
  NOR2_X1 U5362 ( .A1(n6575), .A2(n4656), .ZN(n4655) );
  INV_X1 U5363 ( .A(n6573), .ZN(n4656) );
  NAND2_X1 U5364 ( .A1(n6860), .A2(n8400), .ZN(n6574) );
  OR2_X1 U5365 ( .A1(n8323), .A2(n6593), .ZN(n9609) );
  INV_X1 U5366 ( .A(n4897), .ZN(n4895) );
  AND2_X1 U5367 ( .A1(n8373), .A2(n8375), .ZN(n9470) );
  NOR2_X1 U5368 ( .A1(n6556), .A2(n4903), .ZN(n4902) );
  INV_X1 U5369 ( .A(n6554), .ZN(n4903) );
  AND2_X1 U5370 ( .A1(n4902), .A2(n6555), .ZN(n4900) );
  NOR2_X1 U5371 ( .A1(n9731), .A2(n9254), .ZN(n4901) );
  NOR2_X1 U5372 ( .A1(n4344), .A2(n4863), .ZN(n4862) );
  INV_X1 U5373 ( .A(n6551), .ZN(n4863) );
  OR2_X1 U5374 ( .A1(n4864), .A2(n4344), .ZN(n4861) );
  AND2_X1 U5375 ( .A1(n6552), .A2(n4347), .ZN(n4864) );
  NAND2_X1 U5376 ( .A1(n5509), .A2(n5508), .ZN(n9554) );
  NAND2_X1 U5377 ( .A1(n5486), .A2(n5485), .ZN(n9673) );
  AND2_X1 U5378 ( .A1(n8281), .A2(n8432), .ZN(n9579) );
  NAND2_X1 U5379 ( .A1(n5417), .A2(n5416), .ZN(n9618) );
  AND2_X1 U5380 ( .A1(n8275), .A2(n8271), .ZN(n9612) );
  NAND2_X1 U5381 ( .A1(n7791), .A2(n7793), .ZN(n7790) );
  NAND2_X1 U5382 ( .A1(n5702), .A2(n8197), .ZN(n9777) );
  OR2_X1 U5383 ( .A1(n8175), .A2(n9407), .ZN(n5701) );
  AND2_X1 U5384 ( .A1(n4913), .A2(n4983), .ZN(n4599) );
  INV_X1 U5385 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4985) );
  XNOR2_X1 U5386 ( .A(n6280), .B(n6279), .ZN(n9175) );
  OAI21_X1 U5387 ( .B1(n6275), .B2(n6274), .A(n6273), .ZN(n6280) );
  XNOR2_X1 U5388 ( .A(n6275), .B(n6274), .ZN(n8588) );
  INV_X1 U5389 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4986) );
  AND2_X1 U5390 ( .A1(n4988), .A2(n5243), .ZN(n4645) );
  AND2_X1 U5391 ( .A1(n4982), .A2(n4647), .ZN(n4646) );
  XNOR2_X1 U5392 ( .A(n5676), .B(n5675), .ZN(n8202) );
  INV_X1 U5393 ( .A(n5389), .ZN(n4904) );
  NAND2_X1 U5394 ( .A1(n4777), .A2(n5602), .ZN(n5622) );
  NAND2_X1 U5395 ( .A1(n5601), .A2(n5600), .ZN(n4777) );
  NAND2_X1 U5396 ( .A1(n4763), .A2(n4762), .ZN(n4761) );
  INV_X1 U5397 ( .A(n4760), .ZN(n4758) );
  NAND2_X1 U5398 ( .A1(n4412), .A2(n4956), .ZN(n5088) );
  NAND2_X1 U5399 ( .A1(n5220), .A2(n4946), .ZN(n5240) );
  AND2_X1 U5400 ( .A1(n5152), .A2(n4976), .ZN(n5153) );
  NAND2_X1 U5401 ( .A1(n4447), .A2(n4923), .ZN(n5110) );
  AND2_X1 U5402 ( .A1(n5885), .A2(n5884), .ZN(n8968) );
  AND4_X1 U5403 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n7060)
         );
  AND2_X1 U5404 ( .A1(n6288), .A2(n5835), .ZN(n8741) );
  INV_X1 U5405 ( .A(n8935), .ZN(n8958) );
  AND3_X1 U5406 ( .A1(n6191), .A2(n6190), .A3(n6189), .ZN(n9011) );
  AND4_X1 U5407 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n8732)
         );
  NAND2_X1 U5408 ( .A1(n7044), .A2(n7234), .ZN(n7046) );
  INV_X1 U5409 ( .A(n8732), .ZN(n9023) );
  NAND2_X1 U5410 ( .A1(n4462), .A2(n4461), .ZN(n8753) );
  AND2_X1 U5411 ( .A1(n4389), .A2(n6071), .ZN(n4461) );
  NAND2_X1 U5412 ( .A1(n6237), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4462) );
  INV_X1 U5413 ( .A(n7429), .ZN(n8754) );
  NAND2_X1 U5414 ( .A1(n6983), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9891) );
  OR2_X1 U5415 ( .A1(n7456), .A2(n9997), .ZN(n4538) );
  XNOR2_X1 U5416 ( .A(n7581), .B(n7589), .ZN(n7456) );
  XNOR2_X1 U5417 ( .A(n6048), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9903) );
  OR2_X1 U5418 ( .A1(n7585), .A2(n7601), .ZN(n4529) );
  NOR2_X1 U5419 ( .A1(n7933), .A2(n7934), .ZN(n7936) );
  INV_X1 U5420 ( .A(n4689), .ZN(n7932) );
  OR2_X1 U5421 ( .A1(n8051), .A2(n8107), .ZN(n4696) );
  XNOR2_X1 U5422 ( .A(n8123), .B(n8124), .ZN(n8051) );
  NOR2_X1 U5423 ( .A1(n6881), .A2(n6880), .ZN(n9902) );
  OAI21_X1 U5424 ( .B1(n8880), .B2(n9908), .A(n4624), .ZN(n4623) );
  AOI21_X1 U5425 ( .B1(n8879), .B2(n9892), .A(n8878), .ZN(n4624) );
  NAND2_X1 U5426 ( .A1(n5888), .A2(n5887), .ZN(n8950) );
  NAND2_X1 U5427 ( .A1(n6193), .A2(n6192), .ZN(n9089) );
  NAND2_X1 U5428 ( .A1(n6121), .A2(n6120), .ZN(n9986) );
  NAND2_X1 U5429 ( .A1(n6086), .A2(n6085), .ZN(n9975) );
  INV_X2 U5430 ( .A(n9990), .ZN(n9988) );
  INV_X1 U5431 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U5432 ( .A1(n5783), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5781) );
  INV_X1 U5433 ( .A(n6480), .ZN(n8200) );
  NAND2_X1 U5434 ( .A1(n6395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U5435 ( .A1(n6395), .A2(n6394), .ZN(n8095) );
  INV_X1 U5436 ( .A(n8053), .ZN(n8050) );
  NAND2_X1 U5437 ( .A1(n5674), .A2(n4747), .ZN(n4746) );
  INV_X1 U5438 ( .A(n5647), .ZN(n4747) );
  INV_X1 U5439 ( .A(n9673), .ZN(n9563) );
  NAND2_X1 U5440 ( .A1(n5438), .A2(n5437), .ZN(n9684) );
  AND2_X1 U5441 ( .A1(n5744), .A2(n5721), .ZN(n9307) );
  NAND2_X1 U5442 ( .A1(n4436), .A2(n4435), .ZN(n4434) );
  NAND2_X1 U5443 ( .A1(n4323), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5142) );
  NOR2_X1 U5444 ( .A1(n8470), .A2(n8471), .ZN(n9361) );
  OAI21_X1 U5445 ( .B1(n9437), .B2(n9846), .A(n9436), .ZN(n9636) );
  AND2_X1 U5446 ( .A1(n9440), .A2(n9439), .ZN(n9635) );
  NAND2_X1 U5447 ( .A1(n5534), .A2(n5533), .ZN(n9540) );
  NAND2_X1 U5448 ( .A1(n5464), .A2(n5463), .ZN(n9589) );
  NAND2_X1 U5449 ( .A1(n6600), .A2(n9776), .ZN(n9601) );
  INV_X1 U5450 ( .A(n9699), .ZN(n9640) );
  INV_X1 U5451 ( .A(n9874), .ZN(n9876) );
  NOR2_X1 U5452 ( .A1(n9867), .A2(n9845), .ZN(n9763) );
  NAND2_X1 U5453 ( .A1(n9869), .A2(n9860), .ZN(n9773) );
  OAI21_X1 U5454 ( .B1(n6114), .B2(n4557), .A(n4556), .ZN(n6109) );
  AND2_X1 U5455 ( .A1(n6344), .A2(n6342), .ZN(n4556) );
  NAND2_X1 U5456 ( .A1(n4491), .A2(n8458), .ZN(n4490) );
  NAND2_X1 U5457 ( .A1(n8250), .A2(n8319), .ZN(n4494) );
  NAND2_X1 U5458 ( .A1(n8263), .A2(n8458), .ZN(n4510) );
  NAND2_X1 U5459 ( .A1(n6155), .A2(n4547), .ZN(n4546) );
  AOI21_X1 U5460 ( .B1(n6146), .B2(n8101), .A(n4550), .ZN(n4549) );
  NAND2_X1 U5461 ( .A1(n6301), .A2(n4548), .ZN(n4547) );
  NAND2_X1 U5462 ( .A1(n4511), .A2(n8287), .ZN(n8288) );
  NAND2_X1 U5463 ( .A1(n9504), .A2(n8293), .ZN(n4504) );
  OAI21_X1 U5464 ( .B1(n4552), .B2(n4551), .A(n6217), .ZN(n6247) );
  NAND2_X1 U5465 ( .A1(n8955), .A2(n6216), .ZN(n4551) );
  AOI21_X1 U5466 ( .B1(n4555), .B2(n4554), .A(n4553), .ZN(n4552) );
  INV_X1 U5467 ( .A(n5524), .ZN(n5525) );
  NOR2_X1 U5468 ( .A1(n4664), .A2(n4659), .ZN(n4658) );
  INV_X1 U5469 ( .A(n8645), .ZN(n4664) );
  INV_X1 U5470 ( .A(n8567), .ZN(n4659) );
  NAND2_X1 U5471 ( .A1(n8645), .A2(n4663), .ZN(n4662) );
  INV_X1 U5472 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U5473 ( .A1(n4481), .A2(n4478), .ZN(n4774) );
  INV_X1 U5474 ( .A(n8353), .ZN(n4479) );
  MUX2_X1 U5475 ( .A(n8384), .B(n8354), .S(n8319), .Z(n8310) );
  INV_X1 U5476 ( .A(n8277), .ZN(n4633) );
  NAND2_X1 U5477 ( .A1(n4440), .A2(SI_29_), .ZN(n4439) );
  INV_X1 U5478 ( .A(n5759), .ZN(n4440) );
  INV_X1 U5479 ( .A(n4775), .ZN(n4428) );
  INV_X1 U5480 ( .A(n5602), .ZN(n4780) );
  INV_X1 U5481 ( .A(n4420), .ZN(n4418) );
  INV_X1 U5482 ( .A(n4421), .ZN(n4415) );
  INV_X1 U5483 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5457) );
  INV_X1 U5484 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5410) );
  NOR2_X1 U5485 ( .A1(n5359), .A2(SI_14_), .ZN(n4795) );
  NOR2_X1 U5486 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4515) );
  INV_X1 U5487 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4977) );
  OAI21_X1 U5488 ( .B1(n4936), .B2(n4921), .A(n4449), .ZN(n4448) );
  NAND2_X1 U5489 ( .A1(n4936), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U5490 ( .A1(n7012), .A2(n6890), .ZN(n7089) );
  NOR2_X1 U5491 ( .A1(n4810), .A2(n4806), .ZN(n4805) );
  INV_X1 U5492 ( .A(n6372), .ZN(n4806) );
  NAND2_X1 U5493 ( .A1(n6375), .A2(n4809), .ZN(n4808) );
  INV_X1 U5494 ( .A(n6374), .ZN(n4809) );
  AND2_X1 U5495 ( .A1(n4819), .A2(n6357), .ZN(n4465) );
  NOR2_X1 U5496 ( .A1(n4824), .A2(n4820), .ZN(n4819) );
  INV_X1 U5497 ( .A(n6358), .ZN(n4820) );
  INV_X1 U5498 ( .A(n6360), .ZN(n4824) );
  INV_X1 U5499 ( .A(n6361), .ZN(n4823) );
  INV_X1 U5500 ( .A(n6359), .ZN(n4822) );
  INV_X1 U5501 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7953) );
  INV_X1 U5502 ( .A(n7705), .ZN(n4477) );
  INV_X1 U5503 ( .A(n9969), .ZN(n4560) );
  INV_X1 U5504 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5792) );
  OAI21_X1 U5505 ( .B1(n7981), .B2(n4817), .A(n6346), .ZN(n4816) );
  INV_X1 U5506 ( .A(n6345), .ZN(n4817) );
  INV_X1 U5507 ( .A(n6347), .ZN(n4813) );
  XOR2_X1 U5508 ( .A(n8758), .B(n9926), .Z(n7247) );
  OAI21_X1 U5509 ( .B1(n7050), .B2(n4803), .A(n6420), .ZN(n7248) );
  INV_X1 U5510 ( .A(SI_18_), .ZN(n10197) );
  INV_X1 U5511 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10068) );
  INV_X1 U5512 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U5513 ( .A1(n5839), .A2(n6390), .ZN(n6392) );
  OR2_X1 U5514 ( .A1(n6118), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5920) );
  AND2_X1 U5515 ( .A1(n6056), .A2(n5918), .ZN(n6096) );
  AND2_X1 U5516 ( .A1(n5057), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5075) );
  NOR2_X1 U5517 ( .A1(n5535), .A2(n9271), .ZN(n5558) );
  NAND2_X1 U5518 ( .A1(n4342), .A2(n5023), .ZN(n4702) );
  AND2_X1 U5519 ( .A1(n5193), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5225) );
  NOR2_X1 U5520 ( .A1(n5366), .A2(n9309), .ZN(n5394) );
  NOR2_X1 U5521 ( .A1(n6560), .A2(n4525), .ZN(n4524) );
  INV_X1 U5522 ( .A(n4526), .ZN(n4525) );
  NAND2_X1 U5523 ( .A1(n6559), .A2(n6558), .ZN(n8353) );
  NAND2_X1 U5524 ( .A1(n9516), .A2(n9499), .ZN(n9489) );
  AOI21_X1 U5525 ( .B1(n4861), .B2(n4859), .A(n4367), .ZN(n4858) );
  INV_X1 U5526 ( .A(n4862), .ZN(n4859) );
  INV_X1 U5527 ( .A(n4861), .ZN(n4860) );
  NOR2_X1 U5528 ( .A1(n9551), .A2(n9554), .ZN(n9534) );
  AND2_X1 U5529 ( .A1(n5465), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5487) );
  NOR2_X1 U5530 ( .A1(n5440), .A2(n5439), .ZN(n5465) );
  NAND2_X1 U5531 ( .A1(n6548), .A2(n9242), .ZN(n8424) );
  OR2_X1 U5532 ( .A1(n6548), .A2(n9242), .ZN(n8267) );
  NOR2_X1 U5533 ( .A1(n5095), .A2(n7749), .ZN(n5057) );
  NOR2_X1 U5534 ( .A1(n7524), .A2(n9861), .ZN(n4528) );
  AND2_X1 U5535 ( .A1(n8213), .A2(n8332), .ZN(n8407) );
  INV_X1 U5536 ( .A(n8403), .ZN(n4652) );
  INV_X1 U5537 ( .A(n5022), .ZN(n7314) );
  NAND2_X1 U5538 ( .A1(n9548), .A2(n4642), .ZN(n4640) );
  OR2_X1 U5539 ( .A1(n9673), .A2(n9211), .ZN(n8360) );
  OR2_X1 U5540 ( .A1(n6548), .A2(n8168), .ZN(n9617) );
  NAND2_X1 U5541 ( .A1(n7688), .A2(n6545), .ZN(n7914) );
  AND2_X1 U5542 ( .A1(n4599), .A2(n4386), .ZN(n4506) );
  NAND2_X1 U5543 ( .A1(n4785), .A2(n4784), .ZN(n4441) );
  AOI21_X1 U5544 ( .B1(n4787), .B2(n4789), .A(n4404), .ZN(n4784) );
  AND2_X1 U5545 ( .A1(n4988), .A2(n4983), .ZN(n4647) );
  AND2_X1 U5546 ( .A1(n5650), .A2(n5628), .ZN(n5648) );
  AOI21_X1 U5547 ( .B1(n4778), .B2(n4780), .A(n4776), .ZN(n4775) );
  INV_X1 U5548 ( .A(n5623), .ZN(n4776) );
  INV_X1 U5549 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4979) );
  AND2_X1 U5550 ( .A1(n5602), .A2(n5584), .ZN(n5600) );
  OAI21_X1 U5551 ( .B1(n5505), .B2(n4416), .A(n4414), .ZN(n5550) );
  INV_X1 U5552 ( .A(n4417), .ZN(n4416) );
  AOI21_X1 U5553 ( .B1(n4415), .B2(n4417), .A(n4398), .ZN(n4414) );
  NOR2_X1 U5554 ( .A1(n5526), .A2(n4418), .ZN(n4417) );
  INV_X1 U5555 ( .A(SI_20_), .ZN(n5504) );
  INV_X1 U5556 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4975) );
  INV_X1 U5557 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4974) );
  INV_X1 U5558 ( .A(n5046), .ZN(n4962) );
  NAND2_X1 U5559 ( .A1(n5087), .A2(n4410), .ZN(n4409) );
  INV_X1 U5560 ( .A(n4956), .ZN(n4410) );
  OAI21_X1 U5561 ( .B1(n6632), .B2(n4445), .A(n4444), .ZN(n4443) );
  INV_X1 U5562 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n4445) );
  NAND2_X1 U5563 ( .A1(n6632), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U5564 ( .A1(n4443), .A2(SI_7_), .ZN(n4952) );
  OAI21_X1 U5565 ( .B1(n4936), .B2(n4938), .A(n4937), .ZN(n4939) );
  NAND2_X1 U5566 ( .A1(n4936), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U5567 ( .A1(n4936), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4924) );
  AND2_X1 U5568 ( .A1(n8652), .A2(n8543), .ZN(n4670) );
  NAND2_X1 U5569 ( .A1(n4668), .A2(n4358), .ZN(n4667) );
  XNOR2_X1 U5570 ( .A(n8574), .B(n8572), .ZN(n8712) );
  INV_X1 U5571 ( .A(n8726), .ZN(n4671) );
  NAND2_X1 U5572 ( .A1(n5848), .A2(n5847), .ZN(n6270) );
  OAI21_X1 U5573 ( .B1(n7026), .B2(n7261), .A(n4618), .ZN(n7014) );
  NAND2_X1 U5574 ( .A1(n6895), .A2(n7261), .ZN(n4618) );
  NAND2_X1 U5575 ( .A1(n7014), .A2(n7013), .ZN(n7012) );
  XNOR2_X1 U5576 ( .A(n7089), .B(n6910), .ZN(n7088) );
  NAND2_X1 U5577 ( .A1(n4338), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4688) );
  NAND2_X1 U5578 ( .A1(n4406), .A2(n4338), .ZN(n7085) );
  AOI21_X1 U5579 ( .B1(n7164), .B2(n7163), .A(n7165), .ZN(n7455) );
  OR2_X1 U5580 ( .A1(n6073), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U5581 ( .A1(n9899), .A2(n7592), .ZN(n7723) );
  NAND2_X1 U5582 ( .A1(n7774), .A2(n7775), .ZN(n7937) );
  OR2_X1 U5583 ( .A1(n7771), .A2(n4690), .ZN(n4689) );
  NOR2_X1 U5584 ( .A1(n7731), .A2(n7729), .ZN(n4690) );
  NOR2_X1 U5585 ( .A1(n8847), .A2(n8848), .ZN(n8851) );
  NAND2_X1 U5586 ( .A1(n6160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U5587 ( .A1(n6383), .A2(n5849), .ZN(n6467) );
  AOI21_X1 U5588 ( .B1(n4727), .B2(n4725), .A(n4379), .ZN(n4724) );
  INV_X1 U5589 ( .A(n4727), .ZN(n4726) );
  INV_X1 U5590 ( .A(n6467), .ZN(n6468) );
  AND2_X1 U5591 ( .A1(n5813), .A2(n10160), .ZN(n5852) );
  INV_X1 U5592 ( .A(n6207), .ZN(n5808) );
  AOI21_X1 U5593 ( .B1(n4706), .B2(n4708), .A(n4370), .ZN(n4703) );
  INV_X1 U5594 ( .A(n9013), .ZN(n4466) );
  NAND2_X1 U5595 ( .A1(n5804), .A2(n5803), .ZN(n6166) );
  INV_X1 U5596 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5803) );
  INV_X1 U5597 ( .A(n5913), .ZN(n5804) );
  NAND2_X1 U5598 ( .A1(n5802), .A2(n5801), .ZN(n5939) );
  INV_X1 U5599 ( .A(n5937), .ZN(n5802) );
  OR2_X1 U5600 ( .A1(n5939), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U5601 ( .A1(n5800), .A2(n5799), .ZN(n6140) );
  INV_X1 U5602 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5799) );
  INV_X1 U5603 ( .A(n6138), .ZN(n5800) );
  NAND2_X1 U5604 ( .A1(n5798), .A2(n7953), .ZN(n6138) );
  INV_X1 U5605 ( .A(n6122), .ZN(n5798) );
  AND4_X1 U5606 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n8532)
         );
  OR2_X1 U5607 ( .A1(n6103), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U5608 ( .A1(n5797), .A2(n5796), .ZN(n6087) );
  INV_X1 U5609 ( .A(n6059), .ZN(n5797) );
  INV_X1 U5610 ( .A(n6338), .ZN(n4828) );
  AOI21_X1 U5611 ( .B1(n7424), .B2(n6338), .A(n4827), .ZN(n4826) );
  INV_X1 U5612 ( .A(n6339), .ZN(n4827) );
  INV_X1 U5613 ( .A(n4844), .ZN(n4843) );
  NAND2_X1 U5614 ( .A1(n4460), .A2(n4459), .ZN(n7559) );
  AND2_X1 U5615 ( .A1(n8753), .A2(n6077), .ZN(n4459) );
  NAND2_X1 U5616 ( .A1(n4401), .A2(n7427), .ZN(n7560) );
  OR2_X1 U5617 ( .A1(n6029), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U5618 ( .A1(n5795), .A2(n5794), .ZN(n6068) );
  INV_X1 U5619 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5794) );
  INV_X1 U5620 ( .A(n6066), .ZN(n5795) );
  NAND2_X1 U5621 ( .A1(n7284), .A2(n6431), .ZN(n7416) );
  OR2_X1 U5622 ( .A1(n6186), .A2(n9877), .ZN(n5962) );
  NAND2_X1 U5623 ( .A1(n4751), .A2(n6422), .ZN(n7249) );
  INV_X1 U5624 ( .A(n7264), .ZN(n4751) );
  XNOR2_X1 U5625 ( .A(n9926), .B(n8758), .ZN(n7251) );
  NAND2_X1 U5626 ( .A1(n6421), .A2(n6420), .ZN(n7265) );
  NAND2_X1 U5627 ( .A1(n4745), .A2(n4363), .ZN(n8944) );
  NAND2_X1 U5628 ( .A1(n8966), .A2(n6455), .ZN(n4745) );
  AND2_X1 U5629 ( .A1(n6358), .A2(n6359), .ZN(n8995) );
  NAND2_X1 U5630 ( .A1(n6165), .A2(n6164), .ZN(n8700) );
  NAND2_X1 U5631 ( .A1(n4467), .A2(n6352), .ZN(n9038) );
  NOR2_X1 U5632 ( .A1(n4469), .A2(n6147), .ZN(n4468) );
  INV_X1 U5633 ( .A(n6351), .ZN(n4469) );
  AOI21_X1 U5634 ( .B1(n4740), .B2(n4739), .A(n4356), .ZN(n4738) );
  INV_X1 U5635 ( .A(n6444), .ZN(n4739) );
  OR2_X1 U5636 ( .A1(n8100), .A2(n8101), .ZN(n8098) );
  INV_X1 U5637 ( .A(n7390), .ZN(n9934) );
  AND2_X1 U5638 ( .A1(n6826), .A2(n6841), .ZN(n6834) );
  NOR2_X1 U5639 ( .A1(n6821), .A2(n6500), .ZN(n6839) );
  OR2_X1 U5640 ( .A1(n6509), .A2(n5846), .ZN(n6972) );
  NAND2_X1 U5641 ( .A1(n8016), .A2(n7850), .ZN(n9955) );
  AND2_X1 U5642 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  INV_X1 U5643 ( .A(n6295), .ZN(n5841) );
  NAND2_X1 U5644 ( .A1(n4687), .A2(n4362), .ZN(n5783) );
  INV_X1 U5645 ( .A(n4750), .ZN(n4749) );
  INV_X1 U5646 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U5647 ( .A1(n6392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U5648 ( .A1(n6400), .A2(n6393), .ZN(n6395) );
  XNOR2_X1 U5649 ( .A(n6391), .B(n6390), .ZN(n6882) );
  AND2_X1 U5650 ( .A1(n5840), .A2(n6389), .ZN(n6470) );
  NAND2_X1 U5651 ( .A1(n4687), .A2(n4686), .ZN(n6295) );
  XNOR2_X1 U5652 ( .A(n6179), .B(n6178), .ZN(n7045) );
  INV_X1 U5653 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U5654 ( .A1(n6177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6179) );
  NOR2_X1 U5655 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4681) );
  NOR2_X1 U5656 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4680) );
  OR2_X1 U5657 ( .A1(n5897), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6073) );
  AND2_X1 U5658 ( .A1(n9248), .A2(n5572), .ZN(n9199) );
  AND2_X1 U5659 ( .A1(n5666), .A2(n5665), .ZN(n5724) );
  NAND2_X1 U5660 ( .A1(n4715), .A2(n7920), .ZN(n7923) );
  OAI21_X1 U5661 ( .B1(n4916), .B2(n4588), .A(n4587), .ZN(n4589) );
  INV_X1 U5662 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5418) );
  AND2_X1 U5663 ( .A1(n5599), .A2(n5598), .ZN(n9249) );
  OR2_X1 U5664 ( .A1(n5511), .A2(n5510), .ZN(n5535) );
  AOI21_X1 U5665 ( .B1(n4579), .B2(n5500), .A(n4365), .ZN(n4578) );
  NAND2_X1 U5666 ( .A1(n4593), .A2(n4720), .ZN(n7876) );
  NAND2_X1 U5667 ( .A1(n4594), .A2(n4595), .ZN(n4593) );
  NOR2_X1 U5668 ( .A1(n4916), .A2(n4596), .ZN(n4595) );
  NOR2_X1 U5669 ( .A1(n7003), .A2(n4919), .ZN(n5235) );
  NAND2_X1 U5670 ( .A1(n4568), .A2(n4566), .ZN(n5375) );
  OR2_X1 U5671 ( .A1(n4569), .A2(n4567), .ZN(n4566) );
  NOR2_X1 U5672 ( .A1(n5737), .A2(n8463), .ZN(n5744) );
  AND2_X1 U5673 ( .A1(n8459), .A2(n4380), .ZN(n4435) );
  AOI211_X1 U5674 ( .C1(n8456), .C2(n8455), .A(n8464), .B(n8454), .ZN(n8459)
         );
  OR2_X1 U5675 ( .A1(n8392), .A2(n4498), .ZN(n4497) );
  AND2_X1 U5676 ( .A1(n8393), .A2(n4499), .ZN(n4498) );
  NAND2_X1 U5677 ( .A1(n8324), .A2(n4500), .ZN(n4499) );
  INV_X1 U5678 ( .A(n8323), .ZN(n4500) );
  AND2_X1 U5679 ( .A1(n5734), .A2(n5733), .ZN(n8309) );
  AND2_X1 U5680 ( .A1(n5591), .A2(n5590), .ZN(n9221) );
  AND2_X1 U5681 ( .A1(n5474), .A2(n5473), .ZN(n9283) );
  NOR2_X1 U5682 ( .A1(n6743), .A2(n4604), .ZN(n6683) );
  AND2_X1 U5683 ( .A1(n6686), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4604) );
  NOR2_X1 U5684 ( .A1(n6919), .A2(n4609), .ZN(n6921) );
  AND2_X1 U5685 ( .A1(n6920), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U5686 ( .A1(n6921), .A2(n6922), .ZN(n7199) );
  OR2_X1 U5687 ( .A1(n7667), .A2(n7668), .ZN(n4603) );
  OR2_X1 U5688 ( .A1(n7991), .A2(n7990), .ZN(n8068) );
  INV_X1 U5689 ( .A(n9281), .ZN(n9435) );
  NAND2_X1 U5690 ( .A1(n9462), .A2(n4524), .ZN(n9438) );
  INV_X1 U5691 ( .A(n9471), .ZN(n4630) );
  INV_X1 U5692 ( .A(n5683), .ZN(n5681) );
  NAND2_X1 U5693 ( .A1(n9462), .A2(n6598), .ZN(n9463) );
  NAND2_X1 U5694 ( .A1(n4640), .A2(n4637), .ZN(n9521) );
  AND2_X1 U5695 ( .A1(n4644), .A2(n4635), .ZN(n4634) );
  AND2_X1 U5696 ( .A1(n9504), .A2(n9505), .ZN(n4644) );
  NAND2_X1 U5697 ( .A1(n4637), .A2(n4636), .ZN(n4635) );
  NAND2_X1 U5698 ( .A1(n9534), .A2(n6597), .ZN(n9535) );
  NAND2_X1 U5699 ( .A1(n5487), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5511) );
  OR2_X1 U5700 ( .A1(n5419), .A2(n5418), .ZN(n5440) );
  NOR2_X1 U5701 ( .A1(n9706), .A2(n5719), .ZN(n6600) );
  OR2_X1 U5702 ( .A1(n5351), .A2(n9189), .ZN(n5366) );
  NAND2_X1 U5703 ( .A1(n4650), .A2(n4648), .ZN(n7683) );
  INV_X1 U5704 ( .A(n8210), .ZN(n4649) );
  OR2_X1 U5705 ( .A1(n7753), .A2(n9336), .ZN(n6538) );
  OR2_X1 U5706 ( .A1(n5297), .A2(n5093), .ZN(n5095) );
  INV_X1 U5707 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7749) );
  AND2_X1 U5708 ( .A1(n7501), .A2(n4333), .ZN(n7537) );
  NAND2_X1 U5709 ( .A1(n7501), .A2(n4528), .ZN(n7399) );
  INV_X1 U5710 ( .A(n4879), .ZN(n4878) );
  OAI21_X1 U5711 ( .B1(n4881), .B2(n6533), .A(n4378), .ZN(n4879) );
  NAND2_X1 U5712 ( .A1(n7398), .A2(n7397), .ZN(n7396) );
  NAND2_X1 U5713 ( .A1(n7501), .A2(n7442), .ZN(n7441) );
  NOR2_X1 U5714 ( .A1(n6857), .A2(n5178), .ZN(n6946) );
  AND2_X1 U5715 ( .A1(n9850), .A2(n8394), .ZN(n9584) );
  NAND2_X1 U5716 ( .A1(n8315), .A2(n8314), .ZN(n8320) );
  AND2_X1 U5717 ( .A1(n9410), .A2(n9434), .ZN(n9631) );
  AOI21_X1 U5718 ( .B1(n4892), .B2(n4890), .A(n4889), .ZN(n9423) );
  NOR2_X1 U5719 ( .A1(n4895), .A2(n4891), .ZN(n4890) );
  OAI21_X1 U5720 ( .B1(n4893), .B2(n4891), .A(n4376), .ZN(n4889) );
  AND2_X1 U5721 ( .A1(n8359), .A2(n8370), .ZN(n9484) );
  OR2_X1 U5722 ( .A1(n6564), .A2(n9322), .ZN(n6554) );
  INV_X1 U5723 ( .A(n9540), .ZN(n6597) );
  AND2_X1 U5724 ( .A1(n8360), .A2(n8273), .ZN(n9568) );
  AOI21_X1 U5725 ( .B1(n4869), .B2(n4871), .A(n4364), .ZN(n4866) );
  AOI21_X1 U5726 ( .B1(n4906), .B2(n4887), .A(n4371), .ZN(n4886) );
  INV_X1 U5727 ( .A(n9853), .ZN(n9860) );
  NAND2_X1 U5728 ( .A1(n5703), .A2(n9779), .ZN(n7271) );
  AND2_X1 U5729 ( .A1(n7906), .A2(n9706), .ZN(n9845) );
  INV_X1 U5730 ( .A(n8463), .ZN(n9776) );
  XNOR2_X1 U5731 ( .A(n5829), .B(SI_29_), .ZN(n9182) );
  XNOR2_X1 U5732 ( .A(n4441), .B(n5759), .ZN(n5829) );
  XNOR2_X1 U5733 ( .A(n5755), .B(n5754), .ZN(n8205) );
  NAND2_X1 U5734 ( .A1(n4786), .A2(n5677), .ZN(n5755) );
  XNOR2_X1 U5735 ( .A(n5649), .B(n5648), .ZN(n8196) );
  NAND2_X1 U5736 ( .A1(n4425), .A2(n4775), .ZN(n5649) );
  NAND2_X1 U5737 ( .A1(n5601), .A2(n4778), .ZN(n4425) );
  NAND2_X1 U5738 ( .A1(n5008), .A2(n4737), .ZN(n5012) );
  NOR2_X1 U5739 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4737) );
  XNOR2_X1 U5740 ( .A(n5718), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U5741 ( .A1(n5012), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U5742 ( .A1(n4419), .A2(n4420), .ZN(n5527) );
  NAND2_X1 U5743 ( .A1(n5505), .A2(n4421), .ZN(n4419) );
  INV_X1 U5744 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U5745 ( .A1(n4801), .A2(n5408), .ZN(n5429) );
  XNOR2_X1 U5746 ( .A(n5409), .B(n5388), .ZN(n7188) );
  INV_X1 U5747 ( .A(n5380), .ZN(n5381) );
  NAND2_X1 U5748 ( .A1(n4755), .A2(n4756), .ZN(n4972) );
  AOI21_X1 U5749 ( .B1(n4759), .B2(n5069), .A(n4757), .ZN(n4756) );
  INV_X1 U5750 ( .A(n4966), .ZN(n4757) );
  AND2_X1 U5751 ( .A1(n5342), .A2(n4970), .ZN(n4971) );
  OR2_X1 U5752 ( .A1(n5089), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5051) );
  OR2_X1 U5753 ( .A1(n5290), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U5754 ( .A1(n4545), .A2(n4765), .ZN(n5289) );
  AND2_X1 U5755 ( .A1(n4940), .A2(n4941), .ZN(n5203) );
  OR2_X1 U5756 ( .A1(n4939), .A2(SI_4_), .ZN(n4940) );
  NAND2_X1 U5757 ( .A1(n7365), .A2(n7364), .ZN(n7366) );
  INV_X1 U5758 ( .A(n4683), .ZN(n7109) );
  NOR2_X1 U5759 ( .A1(n8622), .A2(n4666), .ZN(n4665) );
  INV_X1 U5760 ( .A(n8552), .ZN(n4666) );
  NAND2_X1 U5761 ( .A1(n8704), .A2(n8552), .ZN(n8623) );
  AND4_X1 U5762 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n7828)
         );
  OAI21_X1 U5763 ( .B1(n7051), .B2(n8564), .A(n7050), .ZN(n7052) );
  NAND2_X1 U5764 ( .A1(n8643), .A2(n8644), .ZN(n4660) );
  NAND2_X1 U5765 ( .A1(n8727), .A2(n8545), .ZN(n8653) );
  AND2_X1 U5766 ( .A1(n7041), .A2(n7040), .ZN(n8729) );
  AND2_X1 U5767 ( .A1(n4331), .A2(n7111), .ZN(n4682) );
  AND2_X1 U5768 ( .A1(n4683), .A2(n4331), .ZN(n7112) );
  NAND2_X1 U5769 ( .A1(n4673), .A2(n4369), .ZN(n4672) );
  NAND2_X1 U5770 ( .A1(n8635), .A2(n4359), .ZN(n8694) );
  NAND2_X1 U5771 ( .A1(n8635), .A2(n8559), .ZN(n8693) );
  NAND2_X1 U5772 ( .A1(n7962), .A2(n4353), .ZN(n8040) );
  AND2_X1 U5773 ( .A1(n7962), .A2(n7961), .ZN(n7965) );
  INV_X1 U5774 ( .A(n8731), .ZN(n8686) );
  INV_X1 U5775 ( .A(n8724), .ZN(n8714) );
  NAND2_X1 U5776 ( .A1(n4671), .A2(n8543), .ZN(n8727) );
  NAND2_X1 U5777 ( .A1(n6829), .A2(n6828), .ZN(n8734) );
  NAND2_X1 U5778 ( .A1(n6327), .A2(n6326), .ZN(n4454) );
  AND2_X1 U5779 ( .A1(n8862), .A2(n4456), .ZN(n4455) );
  AND2_X1 U5780 ( .A1(n4471), .A2(n4470), .ZN(n6387) );
  NOR2_X1 U5781 ( .A1(n6381), .A2(n6382), .ZN(n4471) );
  NAND2_X1 U5782 ( .A1(n6418), .A2(n6383), .ZN(n4470) );
  NAND2_X1 U5783 ( .A1(n6243), .A2(n6242), .ZN(n8934) );
  NAND2_X1 U5784 ( .A1(n6227), .A2(n6226), .ZN(n8923) );
  NAND2_X1 U5785 ( .A1(n5895), .A2(n5894), .ZN(n8935) );
  INV_X1 U5786 ( .A(n8968), .ZN(n8742) );
  INV_X1 U5787 ( .A(n8606), .ZN(n9042) );
  INV_X1 U5788 ( .A(n7828), .ZN(n8752) );
  INV_X1 U5789 ( .A(n7219), .ZN(n8755) );
  INV_X1 U5790 ( .A(n7253), .ZN(n8757) );
  NAND2_X1 U5791 ( .A1(n5974), .A2(n4316), .ZN(n8760) );
  NAND2_X1 U5792 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5965) );
  OR2_X1 U5793 ( .A1(n7158), .A2(n7157), .ZN(n7457) );
  INV_X1 U5794 ( .A(n4537), .ZN(n9906) );
  NAND2_X1 U5795 ( .A1(n4538), .A2(n4328), .ZN(n4537) );
  AND2_X1 U5796 ( .A1(n4529), .A2(n4360), .ZN(n7722) );
  NOR2_X1 U5797 ( .A1(n7722), .A2(n7721), .ZN(n7771) );
  NAND2_X1 U5798 ( .A1(n7727), .A2(n7728), .ZN(n7774) );
  NAND2_X1 U5799 ( .A1(n7776), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U5800 ( .A1(n4692), .A2(n4691), .ZN(n8766) );
  NAND2_X1 U5801 ( .A1(n8120), .A2(n8121), .ZN(n8761) );
  XNOR2_X1 U5802 ( .A(n8797), .B(n8798), .ZN(n8763) );
  AOI21_X1 U5803 ( .B1(n8825), .B2(n9892), .A(n4544), .ZN(n4543) );
  NAND2_X1 U5804 ( .A1(n8828), .A2(n8823), .ZN(n4544) );
  INV_X1 U5805 ( .A(n4700), .ZN(n8831) );
  AND2_X1 U5806 ( .A1(n8820), .A2(n8819), .ZN(n8822) );
  OR2_X1 U5807 ( .A1(n8820), .A2(n8819), .ZN(n4700) );
  NAND2_X1 U5808 ( .A1(n4701), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U5809 ( .A1(n8832), .A2(n4701), .ZN(n4697) );
  INV_X1 U5810 ( .A(n8833), .ZN(n4701) );
  INV_X1 U5811 ( .A(n8875), .ZN(n4627) );
  AOI21_X1 U5812 ( .B1(n8888), .B2(n9046), .A(n8887), .ZN(n9064) );
  NAND2_X1 U5813 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  NAND2_X1 U5814 ( .A1(n9000), .A2(n6453), .ZN(n8982) );
  NAND2_X1 U5815 ( .A1(n4705), .A2(n6448), .ZN(n9022) );
  NAND2_X1 U5816 ( .A1(n9039), .A2(n9040), .ZN(n4705) );
  NAND2_X1 U5817 ( .A1(n7817), .A2(n6342), .ZN(n7893) );
  NAND2_X1 U5818 ( .A1(n4744), .A2(n6434), .ZN(n7554) );
  AOI21_X1 U5819 ( .B1(n4847), .B2(n4845), .A(n4846), .ZN(n4839) );
  INV_X1 U5820 ( .A(n4847), .ZN(n4840) );
  NAND2_X1 U5821 ( .A1(n4848), .A2(n6331), .ZN(n7283) );
  NAND2_X1 U5822 ( .A1(n6330), .A2(n4849), .ZN(n4848) );
  AND2_X1 U5823 ( .A1(n6430), .A2(n6429), .ZN(n4918) );
  NAND2_X1 U5824 ( .A1(n6330), .A2(n6329), .ZN(n7236) );
  INV_X1 U5825 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7389) );
  INV_X1 U5826 ( .A(n9030), .ZN(n9051) );
  NAND2_X1 U5827 ( .A1(n5791), .A2(n4911), .ZN(n5843) );
  AND2_X2 U5828 ( .A1(n6968), .A2(n6519), .ZN(n10005) );
  NAND2_X1 U5829 ( .A1(n6281), .A2(n6614), .ZN(n9112) );
  OR2_X1 U5830 ( .A1(n6004), .A2(n8498), .ZN(n5850) );
  AND2_X1 U5831 ( .A1(n8906), .A2(n8905), .ZN(n9115) );
  INV_X1 U5832 ( .A(n4807), .ZN(n8899) );
  AOI21_X1 U5833 ( .B1(n8911), .B2(n6374), .A(n4810), .ZN(n4807) );
  OAI21_X1 U5834 ( .B1(n6366), .B2(n4829), .A(n4831), .ZN(n8920) );
  NAND2_X1 U5835 ( .A1(n4836), .A2(n6368), .ZN(n8931) );
  NAND2_X1 U5836 ( .A1(n6366), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U5837 ( .A1(n6366), .A2(n6365), .ZN(n8943) );
  NAND2_X1 U5838 ( .A1(n8979), .A2(n6360), .ZN(n8970) );
  NAND2_X1 U5839 ( .A1(n6182), .A2(n6181), .ZN(n9156) );
  INV_X1 U5840 ( .A(n8700), .ZN(n9164) );
  NAND2_X1 U5841 ( .A1(n6350), .A2(n6349), .ZN(n8181) );
  NAND2_X1 U5842 ( .A1(n4814), .A2(n6345), .ZN(n8097) );
  NAND2_X1 U5843 ( .A1(n7976), .A2(n7981), .ZN(n4814) );
  AND2_X1 U5844 ( .A1(n6495), .A2(n6494), .ZN(n9174) );
  NAND2_X1 U5845 ( .A1(n6841), .A2(n6714), .ZN(n10029) );
  INV_X1 U5846 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8024) );
  INV_X1 U5847 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8018) );
  INV_X1 U5848 ( .A(n6470), .ZN(n8016) );
  INV_X1 U5849 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7849) );
  INV_X1 U5850 ( .A(n7044), .ZN(n7850) );
  INV_X1 U5851 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7553) );
  CLKBUF_X1 U5852 ( .A(n7045), .Z(n8862) );
  INV_X1 U5853 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7217) );
  INV_X1 U5854 ( .A(n7946), .ZN(n7938) );
  INV_X1 U5855 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6656) );
  INV_X1 U5856 ( .A(n7598), .ZN(n7589) );
  NOR2_X1 U5857 ( .A1(n6002), .A2(n4851), .ZN(n6035) );
  NAND2_X1 U5858 ( .A1(n5766), .A2(n4853), .ZN(n4851) );
  INV_X1 U5859 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U5860 ( .A1(n7866), .A2(n4570), .ZN(n9186) );
  NAND2_X1 U5861 ( .A1(n7866), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U5862 ( .A1(n9260), .A2(n5501), .ZN(n9209) );
  OAI21_X1 U5863 ( .B1(n4714), .B2(n5500), .A(n4579), .ZN(n9208) );
  INV_X1 U5864 ( .A(n6955), .ZN(n7487) );
  NAND2_X1 U5865 ( .A1(n9239), .A2(n9240), .ZN(n9238) );
  NAND2_X1 U5866 ( .A1(n9228), .A2(n5405), .ZN(n9239) );
  INV_X1 U5867 ( .A(n6564), .ZN(n9499) );
  INV_X1 U5868 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9271) );
  NOR2_X1 U5869 ( .A1(n9197), .A2(n9268), .ZN(n4910) );
  NAND2_X1 U5870 ( .A1(n5742), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9299) );
  AOI21_X1 U5871 ( .B1(n5404), .B2(n9240), .A(n4366), .ZN(n4584) );
  INV_X1 U5872 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9309) );
  INV_X1 U5873 ( .A(n8467), .ZN(n4431) );
  INV_X1 U5874 ( .A(n9254), .ZN(n9321) );
  INV_X1 U5875 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U5876 ( .A1(n5119), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5105) );
  INV_X1 U5877 ( .A(n4608), .ZN(n6678) );
  INV_X1 U5878 ( .A(n4606), .ZN(n6745) );
  NOR2_X1 U5879 ( .A1(n6790), .A2(n6789), .ZN(n6919) );
  NOR2_X1 U5880 ( .A1(n6787), .A2(n4610), .ZN(n6790) );
  AND2_X1 U5881 ( .A1(n6788), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4610) );
  NOR2_X1 U5882 ( .A1(n7335), .A2(n4394), .ZN(n7339) );
  NOR2_X1 U5883 ( .A1(n7339), .A2(n7338), .ZN(n7573) );
  NOR2_X1 U5884 ( .A1(n7573), .A2(n4611), .ZN(n7577) );
  AND2_X1 U5885 ( .A1(n7574), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U5886 ( .A1(n7577), .A2(n7576), .ZN(n7666) );
  INV_X1 U5887 ( .A(n4603), .ZN(n7987) );
  INV_X1 U5888 ( .A(n4601), .ZN(n9359) );
  NAND2_X1 U5889 ( .A1(n9366), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4600) );
  OR2_X1 U5890 ( .A1(n9807), .A2(n8206), .ZN(n9403) );
  AND2_X1 U5891 ( .A1(n6625), .A2(n6624), .ZN(n9804) );
  INV_X1 U5892 ( .A(n9370), .ZN(n9399) );
  NOR2_X1 U5893 ( .A1(n9415), .A2(n9616), .ZN(n9632) );
  NAND2_X1 U5894 ( .A1(n5609), .A2(n5608), .ZN(n9493) );
  NAND2_X1 U5895 ( .A1(n9548), .A2(n8283), .ZN(n9529) );
  NAND2_X1 U5896 ( .A1(n9593), .A2(n8277), .ZN(n9575) );
  NAND2_X1 U5897 ( .A1(n4868), .A2(n4872), .ZN(n9598) );
  NAND2_X1 U5898 ( .A1(n8161), .A2(n4873), .ZN(n4868) );
  NAND2_X1 U5899 ( .A1(n7790), .A2(n6546), .ZN(n7905) );
  NAND2_X1 U5900 ( .A1(n7349), .A2(n4339), .ZN(n7532) );
  AND2_X1 U5901 ( .A1(n7349), .A2(n8236), .ZN(n7533) );
  AND2_X1 U5902 ( .A1(n7497), .A2(n6533), .ZN(n7440) );
  AND2_X1 U5903 ( .A1(n4653), .A2(n8401), .ZN(n6949) );
  NAND2_X1 U5904 ( .A1(n6574), .A2(n4655), .ZN(n4653) );
  NAND2_X1 U5905 ( .A1(n6574), .A2(n6573), .ZN(n6849) );
  OR2_X1 U5906 ( .A1(n9831), .A2(n7275), .ZN(n9834) );
  OR2_X1 U5907 ( .A1(n9831), .A2(n8455), .ZN(n9586) );
  NAND2_X1 U5908 ( .A1(n5125), .A2(n4355), .ZN(n5113) );
  INV_X1 U5909 ( .A(n9834), .ZN(n9590) );
  INV_X1 U5910 ( .A(n9586), .ZN(n9828) );
  AND2_X1 U5911 ( .A1(n6592), .A2(n8398), .ZN(n9850) );
  INV_X1 U5912 ( .A(n9688), .ZN(n9687) );
  INV_X1 U5913 ( .A(n8320), .ZN(n9710) );
  NAND2_X1 U5914 ( .A1(n5656), .A2(n5655), .ZN(n9720) );
  OAI21_X1 U5915 ( .B1(n9496), .B2(n4895), .A(n4893), .ZN(n9445) );
  NAND2_X1 U5916 ( .A1(n4899), .A2(n4896), .ZN(n9461) );
  NOR2_X1 U5917 ( .A1(n4900), .A2(n4901), .ZN(n4896) );
  NAND2_X1 U5918 ( .A1(n9496), .A2(n4902), .ZN(n4899) );
  NAND2_X1 U5919 ( .A1(n4857), .A2(n4861), .ZN(n9533) );
  NAND2_X1 U5920 ( .A1(n9560), .A2(n4862), .ZN(n4857) );
  INV_X1 U5921 ( .A(n9554), .ZN(n9745) );
  AND2_X1 U5922 ( .A1(n4865), .A2(n4347), .ZN(n9544) );
  NAND2_X1 U5923 ( .A1(n9560), .A2(n6551), .ZN(n4865) );
  NAND2_X1 U5924 ( .A1(n4874), .A2(n4875), .ZN(n9608) );
  OR2_X1 U5925 ( .A1(n8161), .A2(n6584), .ZN(n4874) );
  INV_X1 U5926 ( .A(n6548), .ZN(n9774) );
  INV_X1 U5927 ( .A(n9763), .ZN(n9761) );
  AND2_X1 U5928 ( .A1(n9777), .A2(n9776), .ZN(n9841) );
  INV_X1 U5929 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9781) );
  AND2_X1 U5930 ( .A1(n4982), .A2(n4599), .ZN(n4507) );
  INV_X1 U5931 ( .A(n5035), .ZN(n9787) );
  AND2_X1 U5932 ( .A1(n4982), .A2(n4983), .ZN(n4598) );
  INV_X1 U5933 ( .A(n5462), .ZN(n8455) );
  AND2_X1 U5934 ( .A1(n4994), .A2(n5345), .ZN(n7996) );
  NAND2_X1 U5935 ( .A1(n4761), .A2(n4759), .ZN(n5314) );
  NAND2_X1 U5936 ( .A1(n4761), .A2(n4758), .ZN(n5313) );
  NAND2_X1 U5937 ( .A1(n4798), .A2(n4960), .ZN(n5045) );
  NAND2_X1 U5938 ( .A1(n5088), .A2(n5087), .ZN(n4798) );
  NOR2_X1 U5939 ( .A1(n5262), .A2(n4767), .ZN(n4463) );
  NOR2_X1 U5940 ( .A1(n5153), .A2(n4612), .ZN(n9354) );
  NAND2_X1 U5941 ( .A1(n5243), .A2(n4614), .ZN(n4613) );
  NOR2_X2 U5942 ( .A1(n6884), .A2(n6616), .ZN(P2_U3893) );
  OAI21_X1 U5943 ( .B1(n6983), .B2(P2_IR_REG_0__SCAN_IN), .A(n9891), .ZN(n6984) );
  INV_X1 U5944 ( .A(n4529), .ZN(n7719) );
  INV_X1 U5945 ( .A(n4540), .ZN(n8049) );
  NAND2_X1 U5946 ( .A1(n8824), .A2(n4541), .ZN(P2_U3199) );
  INV_X1 U5947 ( .A(n4542), .ZN(n4541) );
  OAI21_X1 U5948 ( .B1(n8831), .B2(n8822), .A(n8821), .ZN(n8824) );
  OAI21_X1 U5949 ( .B1(n8829), .B2(n8877), .A(n4543), .ZN(n4542) );
  NAND2_X1 U5950 ( .A1(n4625), .A2(n4622), .ZN(P2_U3201) );
  NAND2_X1 U5951 ( .A1(n4626), .A2(n9904), .ZN(n4625) );
  INV_X1 U5952 ( .A(n4623), .ZN(n4622) );
  XNOR2_X1 U5953 ( .A(n8876), .B(n4627), .ZN(n4626) );
  NAND2_X1 U5954 ( .A1(n5845), .A2(n6505), .ZN(n6506) );
  INV_X1 U5955 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U5956 ( .A1(n5725), .A2(n9307), .ZN(n5751) );
  NAND2_X1 U5957 ( .A1(n9648), .A2(n9286), .ZN(n4564) );
  NAND2_X1 U5958 ( .A1(n4430), .A2(n4429), .ZN(P1_U3242) );
  OR2_X1 U5959 ( .A1(n8466), .A2(n8465), .ZN(n4429) );
  NAND2_X1 U5960 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  MUX2_X1 U5961 ( .A(n9637), .B(n9716), .S(n9876), .Z(n9638) );
  MUX2_X1 U5962 ( .A(n9717), .B(n9716), .S(n9869), .Z(n9718) );
  AND2_X1 U5963 ( .A1(n4768), .A2(n4771), .ZN(n4327) );
  INV_X1 U5964 ( .A(n6560), .ZN(n6559) );
  OR2_X1 U5965 ( .A1(n7598), .A2(n7582), .ZN(n4328) );
  AND2_X1 U5966 ( .A1(n9594), .A2(n8275), .ZN(n4329) );
  NAND2_X1 U5967 ( .A1(n8751), .A2(n4560), .ZN(n6340) );
  NAND2_X1 U5968 ( .A1(n7108), .A2(n8757), .ZN(n4331) );
  INV_X1 U5969 ( .A(n6293), .ZN(n4687) );
  NAND2_X1 U5970 ( .A1(n4904), .A2(n4982), .ZN(n5003) );
  AND2_X1 U5971 ( .A1(n6598), .A2(n9222), .ZN(n4332) );
  AND2_X1 U5972 ( .A1(n4528), .A2(n4527), .ZN(n4333) );
  INV_X1 U5973 ( .A(n6533), .ZN(n4883) );
  AND2_X1 U5974 ( .A1(n6326), .A2(n8869), .ZN(n4334) );
  INV_X1 U5975 ( .A(n8904), .ZN(n8596) );
  AND2_X1 U5976 ( .A1(n4854), .A2(n5821), .ZN(n4335) );
  AND2_X1 U5977 ( .A1(n4334), .A2(n4456), .ZN(n4336) );
  INV_X1 U5978 ( .A(n4741), .ZN(n4740) );
  NAND2_X1 U5979 ( .A1(n4742), .A2(n6445), .ZN(n4741) );
  INV_X1 U5980 ( .A(n9648), .ZN(n6598) );
  NAND2_X1 U5981 ( .A1(n5630), .A2(n5629), .ZN(n9648) );
  OAI21_X1 U5982 ( .B1(n4401), .B2(n4828), .A(n4826), .ZN(n7704) );
  INV_X1 U5983 ( .A(n8022), .ZN(n4456) );
  OR2_X1 U5984 ( .A1(n8862), .A2(n8022), .ZN(n4337) );
  AND2_X1 U5985 ( .A1(n8341), .A2(n8236), .ZN(n4339) );
  AND2_X1 U5986 ( .A1(n9462), .A2(n4526), .ZN(n4340) );
  AND2_X1 U5987 ( .A1(n6360), .A2(n8969), .ZN(n8983) );
  NAND2_X1 U5988 ( .A1(n8759), .A2(n9920), .ZN(n6421) );
  AND2_X1 U5989 ( .A1(n4457), .A2(n6344), .ZN(n4341) );
  OR2_X1 U5990 ( .A1(n8451), .A2(n7314), .ZN(n4342) );
  AND2_X1 U5991 ( .A1(n4601), .A2(n4600), .ZN(n4343) );
  INV_X1 U5992 ( .A(n6329), .ZN(n4850) );
  AND2_X1 U5993 ( .A1(n9554), .A2(n9325), .ZN(n4344) );
  NAND2_X1 U5994 ( .A1(n6373), .A2(n6372), .ZN(n8911) );
  INV_X1 U5995 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5766) );
  INV_X1 U5996 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4853) );
  INV_X1 U5997 ( .A(n4951), .ZN(n4767) );
  NOR2_X1 U5998 ( .A1(n9986), .A2(n8748), .ZN(n4345) );
  INV_X1 U5999 ( .A(n5069), .ZN(n4762) );
  OR2_X1 U6000 ( .A1(n9122), .A2(n8924), .ZN(n4346) );
  NAND2_X1 U6001 ( .A1(n9563), .A2(n9211), .ZN(n4347) );
  AND2_X1 U6002 ( .A1(n4660), .A2(n8645), .ZN(n4348) );
  OR2_X1 U6003 ( .A1(n4570), .A2(n4571), .ZN(n4349) );
  OR3_X1 U6004 ( .A1(n6388), .A2(n7046), .A3(n4337), .ZN(n4350) );
  AND2_X1 U6005 ( .A1(n4765), .A2(n4413), .ZN(n4351) );
  NOR2_X1 U6006 ( .A1(n9451), .A2(n9452), .ZN(n4352) );
  NAND2_X1 U6007 ( .A1(n4852), .A2(n5766), .ZN(n6019) );
  INV_X1 U6008 ( .A(n8400), .ZN(n4489) );
  AND2_X1 U6009 ( .A1(n7961), .A2(n8037), .ZN(n4353) );
  AND2_X1 U6010 ( .A1(n4640), .A2(n4641), .ZN(n4354) );
  AND2_X1 U6011 ( .A1(n6632), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4355) );
  AND2_X1 U6012 ( .A1(n8537), .A2(n8746), .ZN(n4356) );
  AND2_X1 U6013 ( .A1(n4700), .A2(n4699), .ZN(n4357) );
  NAND2_X1 U6014 ( .A1(n8546), .A2(n9023), .ZN(n4358) );
  AND2_X1 U6015 ( .A1(n8560), .A2(n8559), .ZN(n4359) );
  OR2_X1 U6016 ( .A1(n7718), .A2(n7717), .ZN(n4360) );
  AND2_X1 U6017 ( .A1(n6360), .A2(n4822), .ZN(n4361) );
  AND2_X1 U6018 ( .A1(n5815), .A2(n4749), .ZN(n4362) );
  INV_X1 U6019 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4686) );
  AND2_X1 U6020 ( .A1(n6456), .A2(n6458), .ZN(n4363) );
  INV_X1 U6021 ( .A(n5307), .ZN(n4596) );
  OR2_X1 U6022 ( .A1(n9133), .A2(n8946), .ZN(n6369) );
  INV_X1 U6023 ( .A(n6369), .ZN(n4832) );
  AND2_X1 U6024 ( .A1(n6596), .A2(n8520), .ZN(n4364) );
  INV_X1 U6025 ( .A(n4876), .ZN(n4875) );
  NOR2_X1 U6026 ( .A1(n9774), .A2(n9242), .ZN(n4876) );
  NOR2_X1 U6027 ( .A1(n5523), .A2(n5522), .ZN(n4365) );
  NOR2_X1 U6028 ( .A1(n5428), .A2(n5427), .ZN(n4366) );
  NOR2_X1 U6029 ( .A1(n6597), .A2(n9212), .ZN(n4367) );
  NAND2_X1 U6030 ( .A1(n7136), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U6031 ( .A1(n4576), .A2(n5340), .ZN(n4575) );
  INV_X1 U6032 ( .A(n4575), .ZN(n4572) );
  INV_X1 U6033 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U6034 ( .A1(n4677), .A2(n7837), .ZN(n4369) );
  INV_X1 U6035 ( .A(n8342), .ZN(n7793) );
  AND2_X1 U6036 ( .A1(n8251), .A2(n8414), .ZN(n8342) );
  AND2_X1 U6037 ( .A1(n9100), .A2(n9044), .ZN(n4370) );
  NOR2_X1 U6038 ( .A1(n9702), .A2(n9332), .ZN(n4371) );
  NOR2_X1 U6039 ( .A1(n9540), .A2(n9324), .ZN(n4372) );
  NOR2_X1 U6040 ( .A1(n6596), .A2(n8520), .ZN(n4373) );
  NOR2_X1 U6041 ( .A1(n9618), .A2(n9330), .ZN(n4374) );
  NAND2_X1 U6042 ( .A1(n5869), .A2(n5868), .ZN(n9062) );
  INV_X1 U6043 ( .A(n4638), .ZN(n4637) );
  NAND2_X1 U6044 ( .A1(n4641), .A2(n4639), .ZN(n4638) );
  AND2_X1 U6045 ( .A1(n4797), .A2(n4409), .ZN(n4375) );
  NAND2_X1 U6046 ( .A1(n9446), .A2(n9295), .ZN(n4376) );
  NOR2_X1 U6047 ( .A1(n9062), .A2(n8904), .ZN(n4377) );
  OR2_X1 U6048 ( .A1(n9861), .A2(n9338), .ZN(n4378) );
  AND2_X1 U6049 ( .A1(n9062), .A2(n8904), .ZN(n4379) );
  OR2_X1 U6050 ( .A1(n9168), .A2(n8732), .ZN(n6301) );
  INV_X1 U6051 ( .A(n9594), .ZN(n9597) );
  AND2_X1 U6052 ( .A1(n8276), .A2(n8277), .ZN(n9594) );
  OR2_X1 U6053 ( .A1(n4448), .A2(SI_1_), .ZN(n4447) );
  OR2_X1 U6054 ( .A1(n8457), .A2(n8458), .ZN(n4380) );
  AND2_X1 U6055 ( .A1(n5674), .A2(n9219), .ZN(n4381) );
  AND2_X1 U6056 ( .A1(n4349), .A2(n5373), .ZN(n4382) );
  AND2_X1 U6057 ( .A1(n4651), .A2(n8400), .ZN(n4383) );
  INV_X1 U6058 ( .A(n9414), .ZN(n9714) );
  NAND2_X1 U6059 ( .A1(n8312), .A2(n8311), .ZN(n9414) );
  NOR2_X1 U6060 ( .A1(n5312), .A2(n4760), .ZN(n4759) );
  AND2_X1 U6061 ( .A1(n4688), .A2(n7083), .ZN(n4384) );
  AND2_X1 U6062 ( .A1(n6376), .A2(n4808), .ZN(n4385) );
  INV_X1 U6063 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5013) );
  AND2_X1 U6064 ( .A1(n9133), .A2(n8946), .ZN(n6370) );
  INV_X1 U6065 ( .A(n6370), .ZN(n4830) );
  NOR2_X1 U6066 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4386) );
  AND2_X1 U6067 ( .A1(n9430), .A2(n9429), .ZN(n4387) );
  INV_X1 U6068 ( .A(n4591), .ZN(n4590) );
  NOR2_X1 U6069 ( .A1(n4717), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U6070 ( .A1(n8270), .A2(n8269), .ZN(n4388) );
  AND2_X1 U6071 ( .A1(n6072), .A2(n6070), .ZN(n4389) );
  INV_X1 U6072 ( .A(n4442), .ZN(n5262) );
  OAI21_X1 U6073 ( .B1(n4443), .B2(SI_7_), .A(n4952), .ZN(n4442) );
  NAND2_X1 U6074 ( .A1(n9250), .A2(n5599), .ZN(n9218) );
  AND2_X1 U6075 ( .A1(n4333), .A2(n7542), .ZN(n4390) );
  INV_X1 U6076 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6988) );
  OR2_X1 U6077 ( .A1(n4501), .A2(n8388), .ZN(n4391) );
  INV_X1 U6078 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4721) );
  AND2_X1 U6079 ( .A1(n7365), .A2(n4677), .ZN(n4392) );
  NAND2_X1 U6080 ( .A1(n4867), .A2(n4866), .ZN(n9578) );
  AND2_X1 U6081 ( .A1(n9014), .A2(n6357), .ZN(n8992) );
  AND2_X2 U6082 ( .A1(n6470), .A2(n7044), .ZN(n6508) );
  NAND2_X1 U6083 ( .A1(n4884), .A2(n4886), .ZN(n8001) );
  NAND2_X1 U6084 ( .A1(n8098), .A2(n6444), .ZN(n8143) );
  INV_X1 U6085 ( .A(n8644), .ZN(n4663) );
  INV_X1 U6086 ( .A(n7731), .ZN(n7773) );
  INV_X1 U6087 ( .A(n9520), .ZN(n4639) );
  NAND2_X1 U6088 ( .A1(n5680), .A2(n5679), .ZN(n6560) );
  AND2_X1 U6089 ( .A1(n9610), .A2(n8275), .ZN(n4393) );
  AND2_X1 U6090 ( .A1(n7336), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4394) );
  NOR2_X1 U6091 ( .A1(n4795), .A2(n5379), .ZN(n4395) );
  NOR2_X1 U6092 ( .A1(n9617), .A2(n9618), .ZN(n9599) );
  INV_X1 U6093 ( .A(n9222), .ZN(n9320) );
  AND2_X1 U6094 ( .A1(n5637), .A2(n5636), .ZN(n9222) );
  AND2_X1 U6095 ( .A1(n5342), .A2(n4796), .ZN(n4396) );
  AND4_X1 U6096 ( .A1(n4517), .A2(n4516), .A3(n4515), .A4(n4518), .ZN(n4723)
         );
  NAND2_X1 U6097 ( .A1(n4466), .A2(n6315), .ZN(n9014) );
  INV_X1 U6098 ( .A(n9907), .ZN(n4536) );
  NAND2_X1 U6099 ( .A1(n4574), .A2(n5358), .ZN(n4397) );
  AND2_X1 U6100 ( .A1(n5525), .A2(SI_21_), .ZN(n4398) );
  NAND2_X1 U6101 ( .A1(n4704), .A2(n4703), .ZN(n9006) );
  OR2_X1 U6102 ( .A1(n5407), .A2(SI_16_), .ZN(n4399) );
  AND2_X1 U6103 ( .A1(n4696), .A2(n4695), .ZN(n4400) );
  INV_X1 U6104 ( .A(n7881), .ZN(n4719) );
  OAI21_X1 U6105 ( .B1(n7817), .B2(n4458), .A(n4341), .ZN(n7976) );
  AND2_X1 U6106 ( .A1(n6337), .A2(n6336), .ZN(n4401) );
  INV_X1 U6107 ( .A(n4401), .ZN(n4475) );
  INV_X1 U6108 ( .A(n4779), .ZN(n4778) );
  OAI21_X1 U6109 ( .B1(n5600), .B2(n4780), .A(n5621), .ZN(n4779) );
  OR2_X1 U6110 ( .A1(n8139), .A2(n8156), .ZN(n4402) );
  AND2_X1 U6111 ( .A1(n4537), .A2(n4536), .ZN(n4403) );
  AND2_X1 U6112 ( .A1(n5757), .A2(n5756), .ZN(n4404) );
  AND2_X1 U6113 ( .A1(n6592), .A2(n8455), .ZN(n8458) );
  AND2_X1 U6114 ( .A1(n5745), .A2(n9601), .ZN(n9317) );
  NAND2_X1 U6115 ( .A1(n5056), .A2(n5055), .ZN(n7753) );
  INV_X1 U6116 ( .A(n7753), .ZN(n4527) );
  OR2_X1 U6117 ( .A1(n4384), .A2(n7084), .ZN(n4533) );
  NOR2_X1 U6118 ( .A1(n6406), .A2(n6405), .ZN(n4405) );
  INV_X1 U6119 ( .A(n8401), .ZN(n4654) );
  INV_X1 U6120 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9189) );
  INV_X1 U6121 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4614) );
  INV_X1 U6122 ( .A(n8862), .ZN(n8869) );
  NAND2_X1 U6123 ( .A1(n4507), .A2(n4904), .ZN(n9780) );
  NAND2_X1 U6124 ( .A1(n6296), .A2(n6295), .ZN(n7715) );
  AND2_X1 U6125 ( .A1(n7083), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U6126 ( .A1(n5006), .A2(n5011), .ZN(n8394) );
  INV_X1 U6127 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4408) );
  XNOR2_X1 U6128 ( .A(n8830), .B(n8846), .ZN(n8820) );
  XNOR2_X1 U6129 ( .A(n8845), .B(n8846), .ZN(n8810) );
  AOI211_X2 U6130 ( .C1(n8865), .C2(n8855), .A(n8854), .B(n8853), .ZN(n8856)
         );
  NAND2_X1 U6131 ( .A1(n8761), .A2(n8762), .ZN(n4620) );
  NOR2_X1 U6132 ( .A1(n8810), .A2(n9032), .ZN(n8847) );
  NAND2_X1 U6133 ( .A1(n5601), .A2(n4426), .ZN(n4424) );
  NAND3_X1 U6134 ( .A1(n4434), .A2(n8460), .A3(n4433), .ZN(n4432) );
  NAND3_X1 U6135 ( .A1(n4495), .A2(n4497), .A3(n8395), .ZN(n4433) );
  NAND2_X1 U6136 ( .A1(n4446), .A2(n4923), .ZN(n5149) );
  NAND2_X1 U6137 ( .A1(n4448), .A2(SI_1_), .ZN(n4923) );
  NAND2_X1 U6138 ( .A1(n5109), .A2(n4447), .ZN(n4446) );
  OAI21_X1 U6139 ( .B1(n4936), .B2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .ZN(
        n4451) );
  NAND3_X1 U6140 ( .A1(n4453), .A2(n4452), .A3(n4350), .ZN(P2_U3296) );
  AOI21_X1 U6141 ( .B1(n6327), .B2(n4336), .A(n4405), .ZN(n4452) );
  OAI211_X1 U6142 ( .C1(n7046), .C2(n6388), .A(n4454), .B(n4455), .ZN(n4453)
         );
  NAND2_X1 U6143 ( .A1(n4815), .A2(n7976), .ZN(n4811) );
  INV_X1 U6144 ( .A(n6343), .ZN(n4458) );
  OR2_X1 U6145 ( .A1(n6645), .A2(n6133), .ZN(n4460) );
  NAND2_X1 U6146 ( .A1(n5242), .A2(n4951), .ZN(n4464) );
  NAND2_X1 U6147 ( .A1(n5242), .A2(n4463), .ZN(n5263) );
  NAND2_X1 U6148 ( .A1(n4464), .A2(n5262), .ZN(n5264) );
  NAND2_X1 U6149 ( .A1(n6350), .A2(n4468), .ZN(n4467) );
  NAND3_X1 U6150 ( .A1(n4473), .A2(n4472), .A3(n6371), .ZN(n6373) );
  NAND3_X1 U6151 ( .A1(n4826), .A2(n4477), .A3(n4828), .ZN(n4474) );
  NAND2_X1 U6152 ( .A1(n4383), .A2(n6860), .ZN(n4486) );
  OAI211_X1 U6153 ( .C1(n4488), .C2(n6860), .A(n4651), .B(n4487), .ZN(n6930)
         );
  NAND2_X1 U6154 ( .A1(n4655), .A2(n4489), .ZN(n4487) );
  INV_X1 U6155 ( .A(n4655), .ZN(n4488) );
  NAND2_X1 U6156 ( .A1(n4486), .A2(n4483), .ZN(n8215) );
  INV_X1 U6157 ( .A(n4484), .ZN(n4483) );
  OAI21_X1 U6158 ( .B1(n4655), .B2(n4485), .A(n6929), .ZN(n4484) );
  NAND2_X1 U6159 ( .A1(n4494), .A2(n4490), .ZN(n8258) );
  OAI21_X1 U6160 ( .B1(n4493), .B2(n8416), .A(n4492), .ZN(n4491) );
  NAND3_X1 U6161 ( .A1(n4768), .A2(n4771), .A3(n4496), .ZN(n4495) );
  NOR2_X1 U6162 ( .A1(n8392), .A2(n4391), .ZN(n4496) );
  AOI21_X1 U6163 ( .B1(n4904), .B2(n4505), .A(n5243), .ZN(n5029) );
  AND2_X1 U6164 ( .A1(n4982), .A2(n4506), .ZN(n4505) );
  NAND2_X1 U6165 ( .A1(n4508), .A2(n9612), .ZN(n8279) );
  NAND3_X1 U6166 ( .A1(n4510), .A2(n4388), .A3(n4509), .ZN(n4508) );
  INV_X1 U6167 ( .A(n6570), .ZN(n8325) );
  OAI21_X1 U6168 ( .B1(n6570), .B2(n7313), .A(n7312), .ZN(n9856) );
  OAI21_X1 U6169 ( .B1(n4513), .B2(n4512), .A(n9528), .ZN(n4511) );
  INV_X1 U6170 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4519) );
  NAND3_X1 U6171 ( .A1(n4723), .A2(n4330), .A3(n4990), .ZN(n5389) );
  AND2_X2 U6172 ( .A1(n4520), .A2(n4519), .ZN(n5152) );
  INV_X1 U6173 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4520) );
  NAND3_X1 U6174 ( .A1(n5964), .A2(n6631), .A3(n5125), .ZN(n4521) );
  NAND2_X1 U6175 ( .A1(n4390), .A2(n7501), .ZN(n7689) );
  NAND3_X1 U6176 ( .A1(n4538), .A2(n7584), .A3(n4328), .ZN(n4535) );
  INV_X1 U6177 ( .A(n4538), .ZN(n7583) );
  MUX2_X1 U6178 ( .A(n9185), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6179 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9185), .S(n6614), .Z(n7051) );
  NAND2_X1 U6180 ( .A1(n4764), .A2(n5240), .ZN(n4545) );
  NAND2_X1 U6181 ( .A1(n5218), .A2(n5217), .ZN(n5220) );
  NAND3_X1 U6182 ( .A1(n6150), .A2(n6301), .A3(n8183), .ZN(n4550) );
  NAND2_X1 U6183 ( .A1(n5149), .A2(n5148), .ZN(n5147) );
  NAND3_X1 U6184 ( .A1(n6095), .A2(n7892), .A3(n6308), .ZN(n4557) );
  AND2_X1 U6185 ( .A1(n6080), .A2(n6079), .ZN(n6114) );
  NAND3_X1 U6186 ( .A1(n6309), .A2(n6508), .A3(n6340), .ZN(n4559) );
  NAND4_X1 U6187 ( .A1(n4562), .A2(n4561), .A3(n6257), .A4(n6251), .ZN(n6260)
         );
  AND2_X4 U6188 ( .A1(n4563), .A2(n5035), .ZN(n5165) );
  NAND3_X1 U6189 ( .A1(n9303), .A2(n9302), .A3(n4564), .ZN(P1_U3240) );
  NAND2_X1 U6190 ( .A1(n7866), .A2(n4349), .ZN(n4565) );
  NAND2_X1 U6191 ( .A1(n4565), .A2(n4569), .ZN(n5374) );
  INV_X1 U6192 ( .A(n5373), .ZN(n4567) );
  NAND2_X1 U6193 ( .A1(n7866), .A2(n4382), .ZN(n4568) );
  INV_X1 U6194 ( .A(n5358), .ZN(n4573) );
  INV_X1 U6195 ( .A(n5341), .ZN(n4576) );
  NAND2_X1 U6196 ( .A1(n4714), .A2(n4579), .ZN(n4577) );
  NAND2_X1 U6197 ( .A1(n4577), .A2(n4578), .ZN(n5546) );
  NAND2_X1 U6198 ( .A1(n9229), .A2(n4582), .ZN(n4581) );
  INV_X1 U6199 ( .A(n7294), .ZN(n4594) );
  NAND2_X1 U6200 ( .A1(n4589), .A2(n4586), .ZN(n4715) );
  NAND2_X1 U6201 ( .A1(n7294), .A2(n4591), .ZN(n4586) );
  NOR2_X1 U6202 ( .A1(n7294), .A2(n4916), .ZN(n7476) );
  INV_X1 U6203 ( .A(n9248), .ZN(n4597) );
  NAND2_X1 U6204 ( .A1(n4904), .A2(n4598), .ZN(n4987) );
  OAI21_X1 U6205 ( .B1(n4615), .B2(n5243), .A(n4613), .ZN(n4612) );
  NAND2_X1 U6206 ( .A1(n4616), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n4615) );
  INV_X1 U6207 ( .A(n5152), .ZN(n4616) );
  XNOR2_X1 U6208 ( .A(n4628), .B(n9432), .ZN(n9437) );
  NAND2_X1 U6209 ( .A1(n4629), .A2(n9431), .ZN(n4628) );
  NAND2_X1 U6210 ( .A1(n9454), .A2(n4387), .ZN(n4629) );
  OAI21_X2 U6211 ( .B1(n9548), .B2(n4638), .A(n4634), .ZN(n9506) );
  AOI21_X1 U6212 ( .B1(n4904), .B2(n4646), .A(n4645), .ZN(n4989) );
  NAND2_X1 U6213 ( .A1(n7351), .A2(n4339), .ZN(n4650) );
  AOI21_X1 U6214 ( .B1(n4339), .B2(n7356), .A(n4649), .ZN(n4648) );
  NAND2_X1 U6215 ( .A1(n8568), .A2(n4658), .ZN(n4657) );
  NAND2_X1 U6216 ( .A1(n7856), .A2(n7855), .ZN(n7962) );
  NAND2_X1 U6217 ( .A1(n8040), .A2(n8039), .ZN(n8084) );
  NAND2_X1 U6218 ( .A1(n8704), .A2(n4665), .ZN(n8624) );
  NAND2_X1 U6219 ( .A1(n7223), .A2(n7224), .ZN(n7365) );
  NAND2_X1 U6220 ( .A1(n4674), .A2(n4672), .ZN(n7854) );
  INV_X1 U6221 ( .A(n7836), .ZN(n4673) );
  NAND2_X1 U6222 ( .A1(n7223), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U6223 ( .A1(n8694), .A2(n8562), .ZN(n8613) );
  NAND3_X1 U6224 ( .A1(n5988), .A2(n4679), .A3(n6988), .ZN(n6002) );
  NAND4_X1 U6225 ( .A1(n4681), .A2(n4680), .A3(n6036), .A4(n4853), .ZN(n5897)
         );
  NAND2_X1 U6226 ( .A1(n7072), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U6227 ( .A1(n4683), .A2(n4682), .ZN(n7177) );
  NAND2_X1 U6228 ( .A1(n7072), .A2(n7066), .ZN(n7067) );
  NOR2_X1 U6229 ( .A1(n7068), .A2(n4685), .ZN(n4684) );
  INV_X1 U6230 ( .A(n7066), .ZN(n4685) );
  NAND2_X1 U6231 ( .A1(n8325), .A2(n7305), .ZN(n7304) );
  AOI21_X2 U6232 ( .B1(n6595), .B2(n9609), .A(n6594), .ZN(n8505) );
  NOR2_X2 U6233 ( .A1(n4981), .A2(n4980), .ZN(n4982) );
  NAND2_X1 U6234 ( .A1(n4338), .A2(n7083), .ZN(n6903) );
  INV_X1 U6235 ( .A(n4696), .ZN(n8125) );
  INV_X1 U6236 ( .A(n8126), .ZN(n4695) );
  NAND2_X1 U6237 ( .A1(n6002), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6003) );
  OAI21_X1 U6238 ( .B1(n4698), .B2(n8820), .A(n4697), .ZN(n8860) );
  INV_X1 U6239 ( .A(n8832), .ZN(n4699) );
  NAND2_X2 U6240 ( .A1(n5303), .A2(n5065), .ZN(n5145) );
  NAND2_X2 U6241 ( .A1(n4702), .A2(n5040), .ZN(n5303) );
  NAND2_X1 U6242 ( .A1(n9039), .A2(n4706), .ZN(n4704) );
  OAI21_X1 U6243 ( .B1(n8514), .B2(n8517), .A(n8515), .ZN(n9261) );
  NAND2_X1 U6244 ( .A1(n8514), .A2(n8515), .ZN(n4714) );
  OAI21_X1 U6245 ( .B1(n8913), .B2(n4726), .A(n4724), .ZN(n6469) );
  NAND2_X1 U6246 ( .A1(n8913), .A2(n6465), .ZN(n4732) );
  OAI21_X1 U6247 ( .B1(n8913), .B2(n4730), .A(n4728), .ZN(n4733) );
  INV_X1 U6248 ( .A(n4733), .ZN(n8883) );
  NAND2_X1 U6249 ( .A1(n5008), .A2(n4998), .ZN(n5006) );
  OAI21_X1 U6250 ( .B1(n8100), .B2(n4741), .A(n4738), .ZN(n8182) );
  NAND2_X1 U6251 ( .A1(n4744), .A2(n4743), .ZN(n7557) );
  NAND2_X1 U6252 ( .A1(n9218), .A2(n9219), .ZN(n9291) );
  NAND2_X1 U6253 ( .A1(n4748), .A2(n4746), .ZN(n6409) );
  NAND2_X1 U6254 ( .A1(n9218), .A2(n4381), .ZN(n4748) );
  NAND2_X1 U6255 ( .A1(n9291), .A2(n5647), .ZN(n9292) );
  NOR2_X1 U6256 ( .A1(n6293), .A2(n4750), .ZN(n5836) );
  NAND3_X1 U6257 ( .A1(n7249), .A2(n7250), .A3(n7251), .ZN(n6425) );
  NAND3_X1 U6258 ( .A1(n6422), .A2(n6421), .A3(n6420), .ZN(n7250) );
  NAND2_X4 U6259 ( .A1(n4754), .A2(n4752), .ZN(n4936) );
  INV_X1 U6260 ( .A(n5070), .ZN(n4763) );
  NAND2_X1 U6261 ( .A1(n5070), .A2(n4759), .ZN(n4755) );
  NAND2_X1 U6262 ( .A1(n4769), .A2(n4772), .ZN(n4771) );
  NAND2_X1 U6263 ( .A1(n4773), .A2(n4770), .ZN(n4768) );
  NAND3_X1 U6264 ( .A1(n9714), .A2(n8310), .A3(n4774), .ZN(n4770) );
  NAND3_X1 U6265 ( .A1(n4774), .A2(n8310), .A3(n9414), .ZN(n4769) );
  NAND2_X1 U6266 ( .A1(n5676), .A2(n4787), .ZN(n4785) );
  NAND2_X1 U6267 ( .A1(n5676), .A2(n5675), .ZN(n4786) );
  NAND3_X1 U6268 ( .A1(n8274), .A2(n8432), .A3(n8273), .ZN(n4792) );
  NAND2_X1 U6269 ( .A1(n5343), .A2(n5342), .ZN(n5360) );
  NAND3_X1 U6270 ( .A1(n5385), .A2(n5386), .A3(n4399), .ZN(n4801) );
  NAND2_X1 U6271 ( .A1(n4801), .A2(n4799), .ZN(n5432) );
  NAND2_X1 U6272 ( .A1(n5385), .A2(n5386), .ZN(n5409) );
  NAND2_X4 U6273 ( .A1(n4802), .A2(n9184), .ZN(n6186) );
  NAND2_X1 U6274 ( .A1(n4802), .A2(n5823), .ZN(n5996) );
  INV_X1 U6275 ( .A(n6421), .ZN(n4803) );
  NAND2_X1 U6276 ( .A1(n4804), .A2(n4385), .ZN(n6378) );
  NAND2_X1 U6277 ( .A1(n6373), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U6278 ( .A1(n4811), .A2(n4812), .ZN(n8148) );
  INV_X1 U6279 ( .A(n6368), .ZN(n4835) );
  OAI21_X1 U6280 ( .B1(n4840), .B2(n6330), .A(n4839), .ZN(n7415) );
  NAND2_X1 U6281 ( .A1(n4843), .A2(n4841), .ZN(n6337) );
  NAND2_X1 U6282 ( .A1(n6330), .A2(n4842), .ZN(n4841) );
  INV_X1 U6283 ( .A(n6002), .ZN(n4852) );
  NAND2_X1 U6284 ( .A1(n5841), .A2(n4854), .ZN(n5820) );
  NAND2_X1 U6285 ( .A1(n4335), .A2(n5841), .ZN(n9176) );
  NAND2_X1 U6286 ( .A1(n9560), .A2(n4858), .ZN(n4856) );
  NAND2_X1 U6287 ( .A1(n8161), .A2(n4869), .ZN(n4867) );
  XNOR2_X2 U6288 ( .A(n4989), .B(P1_IR_REG_27__SCAN_IN), .ZN(n9796) );
  NAND2_X1 U6289 ( .A1(n7499), .A2(n4880), .ZN(n4877) );
  NAND2_X1 U6290 ( .A1(n4877), .A2(n4878), .ZN(n7398) );
  INV_X1 U6291 ( .A(n7439), .ZN(n4882) );
  NAND2_X1 U6292 ( .A1(n7791), .A2(n4885), .ZN(n4884) );
  INV_X1 U6293 ( .A(n9496), .ZN(n4892) );
  OAI21_X1 U6294 ( .B1(n9496), .B2(n6555), .A(n6554), .ZN(n9485) );
  NAND2_X1 U6295 ( .A1(n5139), .A2(n5138), .ZN(n6778) );
  NAND2_X1 U6296 ( .A1(n5014), .A2(n5013), .ZN(n5717) );
  OR2_X1 U6297 ( .A1(n5014), .A2(n5013), .ZN(n5015) );
  AND2_X1 U6298 ( .A1(n8464), .A2(n5719), .ZN(n8389) );
  INV_X1 U6299 ( .A(n8464), .ZN(n6592) );
  OR2_X1 U6300 ( .A1(n6769), .A2(n5316), .ZN(n5320) );
  OR2_X1 U6301 ( .A1(n6786), .A2(n5316), .ZN(n4996) );
  NOR2_X2 U6302 ( .A1(n7296), .A2(n7295), .ZN(n7294) );
  XNOR2_X1 U6303 ( .A(n5527), .B(n5507), .ZN(n7806) );
  NAND2_X1 U6304 ( .A1(n7557), .A2(n6435), .ZN(n7706) );
  NOR2_X1 U6305 ( .A1(n7061), .A2(n7049), .ZN(n7053) );
  NAND2_X1 U6306 ( .A1(n5034), .A2(n9787), .ZN(n5442) );
  NOR2_X1 U6307 ( .A1(n5375), .A2(n5377), .ZN(n9306) );
  XNOR2_X1 U6308 ( .A(n5550), .B(n5549), .ZN(n7974) );
  NAND2_X1 U6309 ( .A1(n6524), .A2(n9849), .ZN(n7313) );
  XNOR2_X1 U6310 ( .A(n6526), .B(n6525), .ZN(n6570) );
  NAND2_X1 U6311 ( .A1(n7960), .A2(n7900), .ZN(n7961) );
  NAND2_X1 U6312 ( .A1(n5775), .A2(n5774), .ZN(n6293) );
  INV_X1 U6313 ( .A(n5897), .ZN(n5775) );
  AND2_X1 U6314 ( .A1(n7048), .A2(n8759), .ZN(n7049) );
  AOI21_X2 U6315 ( .B1(n7032), .B2(n7029), .A(n7028), .ZN(n7124) );
  NAND2_X1 U6316 ( .A1(n8589), .A2(n9184), .ZN(n6240) );
  AND2_X1 U6317 ( .A1(n8589), .A2(n9184), .ZN(n5980) );
  NAND2_X1 U6318 ( .A1(n6894), .A2(n6893), .ZN(n9908) );
  OR2_X1 U6319 ( .A1(n9990), .A2(n9955), .ZN(n9163) );
  INV_X1 U6320 ( .A(n9163), .ZN(n6505) );
  INV_X2 U6321 ( .A(n9037), .ZN(n9047) );
  AND2_X1 U6322 ( .A1(n8534), .A2(n8747), .ZN(n4905) );
  OR2_X1 U6323 ( .A1(n6559), .A2(n9699), .ZN(n4907) );
  INV_X1 U6324 ( .A(n8718), .ZN(n8914) );
  NAND2_X1 U6325 ( .A1(n8700), .A2(n9024), .ZN(n4908) );
  AND2_X1 U6326 ( .A1(n5689), .A2(n5688), .ZN(n9420) );
  INV_X1 U6327 ( .A(n9420), .ZN(n6558) );
  OR2_X1 U6328 ( .A1(n6559), .A2(n9773), .ZN(n4909) );
  OR2_X1 U6329 ( .A1(n6004), .A2(n10044), .ZN(n4911) );
  NAND2_X1 U6330 ( .A1(n5128), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4912) );
  AND2_X1 U6331 ( .A1(n4985), .A2(n4984), .ZN(n4913) );
  XNOR2_X1 U6332 ( .A(n5135), .B(n5136), .ZN(n6770) );
  INV_X1 U6333 ( .A(n9684), .ZN(n6596) );
  AND3_X1 U6334 ( .A1(n5446), .A2(n5445), .A3(n5444), .ZN(n8520) );
  NAND2_X1 U6335 ( .A1(n9047), .A2(n7235), .ZN(n9055) );
  INV_X1 U6336 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4925) );
  INV_X1 U6337 ( .A(n7813), .ZN(n6545) );
  AND2_X1 U6338 ( .A1(n5305), .A2(n5304), .ZN(n4916) );
  NOR2_X1 U6339 ( .A1(n5724), .A2(n9288), .ZN(n4917) );
  XOR2_X1 U6340 ( .A(n5233), .B(n5640), .Z(n4919) );
  NOR2_X1 U6341 ( .A1(n7854), .A2(n7853), .ZN(n7960) );
  INV_X2 U6342 ( .A(n9831), .ZN(n9624) );
  NOR2_X1 U6343 ( .A1(n6441), .A2(n7977), .ZN(n4920) );
  INV_X1 U6344 ( .A(n7699), .ZN(n6542) );
  OAI21_X1 U6345 ( .B1(n6374), .B2(n5846), .A(n6253), .ZN(n6255) );
  INV_X1 U6346 ( .A(n6260), .ZN(n6261) );
  OAI21_X1 U6347 ( .B1(n5846), .B2(n6376), .A(n6261), .ZN(n6263) );
  NOR2_X1 U6348 ( .A1(n6467), .A2(n6264), .ZN(n6265) );
  NAND2_X1 U6349 ( .A1(n6382), .A2(n5846), .ZN(n5847) );
  NAND2_X1 U6350 ( .A1(n6298), .A2(n6508), .ZN(n5848) );
  NAND2_X1 U6351 ( .A1(n6271), .A2(n6383), .ZN(n6298) );
  INV_X1 U6352 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5771) );
  INV_X1 U6353 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4984) );
  OR2_X1 U6354 ( .A1(n7238), .A2(n7060), .ZN(n6430) );
  INV_X1 U6355 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U6356 ( .A1(n6899), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9884) );
  INV_X1 U6357 ( .A(n7581), .ZN(n7582) );
  INV_X1 U6358 ( .A(n9908), .ZN(n8821) );
  INV_X1 U6359 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5801) );
  INV_X1 U6360 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5796) );
  NOR2_X1 U6361 ( .A1(n4345), .A2(n4920), .ZN(n6442) );
  OR2_X1 U6362 ( .A1(n7474), .A2(n5306), .ZN(n5307) );
  AND2_X1 U6363 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5193) );
  OR3_X1 U6364 ( .A1(n5610), .A2(n9256), .A3(n9224), .ZN(n5631) );
  INV_X1 U6365 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5439) );
  INV_X1 U6366 ( .A(SI_27_), .ZN(n10185) );
  INV_X1 U6367 ( .A(SI_23_), .ZN(n5552) );
  INV_X1 U6368 ( .A(SI_19_), .ZN(n5458) );
  INV_X1 U6369 ( .A(SI_17_), .ZN(n5411) );
  INV_X1 U6370 ( .A(n7362), .ZN(n7363) );
  AND2_X1 U6371 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  OR2_X1 U6372 ( .A1(n5860), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5862) );
  AND2_X1 U6373 ( .A1(n7453), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7454) );
  OR2_X1 U6374 ( .A1(n6209), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5889) );
  INV_X1 U6375 ( .A(n6183), .ZN(n5806) );
  OR2_X1 U6376 ( .A1(n6140), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5937) );
  AND2_X1 U6377 ( .A1(n6482), .A2(n6715), .ZN(n6967) );
  OR3_X1 U6378 ( .A1(n6497), .A2(n7044), .A3(n7715), .ZN(n6832) );
  INV_X1 U6379 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5816) );
  INV_X1 U6380 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6161) );
  INV_X1 U6381 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5093) );
  INV_X1 U6382 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6383 ( .A1(n6999), .A2(n5235), .ZN(n6990) );
  NAND2_X1 U6384 ( .A1(n4322), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5108) );
  INV_X1 U6385 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6733) );
  INV_X1 U6386 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U6387 ( .A1(n8205), .A2(n8313), .ZN(n5680) );
  NAND2_X1 U6388 ( .A1(n9599), .A2(n6596), .ZN(n9583) );
  AOI21_X1 U6389 ( .B1(n9318), .B2(n8164), .A(n8001), .ZN(n6547) );
  OR2_X1 U6390 ( .A1(n7889), .A2(n9335), .ZN(n6540) );
  OR2_X1 U6391 ( .A1(n5316), .A2(n6640), .ZN(n5177) );
  OR2_X1 U6392 ( .A1(n5316), .A2(n6642), .ZN(n5155) );
  AND2_X1 U6393 ( .A1(n5578), .A2(n5555), .ZN(n5576) );
  NAND2_X1 U6394 ( .A1(n5412), .A2(n5411), .ZN(n5431) );
  NAND2_X1 U6395 ( .A1(n8754), .A2(n7363), .ZN(n7364) );
  NAND2_X1 U6396 ( .A1(n8576), .A2(n8914), .ZN(n8577) );
  NAND2_X1 U6397 ( .A1(n7964), .A2(n8749), .ZN(n8039) );
  INV_X1 U6398 ( .A(n9024), .ZN(n8997) );
  OR2_X1 U6399 ( .A1(n6194), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U6400 ( .A1(n5808), .A2(n5807), .ZN(n6209) );
  OR2_X1 U6401 ( .A1(n6166), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6183) );
  OR2_X1 U6402 ( .A1(n6831), .A2(n7040), .ZN(n8731) );
  INV_X1 U6403 ( .A(n5862), .ZN(n8512) );
  NAND2_X1 U6404 ( .A1(n5852), .A2(n5814), .ZN(n5860) );
  NAND2_X1 U6405 ( .A1(n5806), .A2(n5805), .ZN(n6194) );
  NOR2_X1 U6406 ( .A1(n9971), .A2(n7044), .ZN(n6840) );
  AND3_X1 U6407 ( .A1(n6510), .A2(n6841), .A3(n6818), .ZN(n6511) );
  OR2_X1 U6408 ( .A1(n7040), .A2(n5846), .ZN(n9012) );
  INV_X1 U6409 ( .A(n9046), .ZN(n9007) );
  OR2_X1 U6410 ( .A1(n6499), .A2(n6470), .ZN(n9971) );
  NAND2_X1 U6411 ( .A1(n6096), .A2(n5919), .ZN(n6118) );
  NAND2_X1 U6412 ( .A1(n5075), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5324) );
  INV_X1 U6413 ( .A(n9409), .ZN(n9244) );
  OR2_X1 U6414 ( .A1(n5324), .A2(n5032), .ZN(n5351) );
  INV_X1 U6415 ( .A(n8451), .ZN(n5738) );
  AND3_X1 U6416 ( .A1(n6764), .A2(n6763), .A3(n6762), .ZN(n8382) );
  INV_X1 U6417 ( .A(n9599), .ZN(n9615) );
  INV_X1 U6418 ( .A(n8339), .ZN(n7909) );
  AND2_X1 U6419 ( .A1(n8221), .A2(n8227), .ZN(n7439) );
  NAND2_X1 U6420 ( .A1(n8389), .A2(n8206), .ZN(n9281) );
  OR2_X1 U6421 ( .A1(n9777), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U6422 ( .A1(n5392), .A2(n5391), .ZN(n6548) );
  INV_X1 U6423 ( .A(n7688), .ZN(n7800) );
  INV_X1 U6424 ( .A(n8335), .ZN(n7356) );
  XNOR2_X1 U6425 ( .A(n9344), .B(n9835), .ZN(n6859) );
  AND2_X1 U6426 ( .A1(n6599), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7272) );
  AND2_X1 U6427 ( .A1(n5623), .A2(n5607), .ZN(n5621) );
  NAND2_X1 U6428 ( .A1(n6842), .A2(n9030), .ZN(n8657) );
  AND4_X1 U6429 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n8606)
         );
  NOR2_X1 U6430 ( .A1(n8784), .A2(n8783), .ZN(n8786) );
  AND2_X1 U6431 ( .A1(P2_U3893), .A2(n6403), .ZN(n9892) );
  NAND2_X1 U6432 ( .A1(n6841), .A2(n6840), .ZN(n9030) );
  INV_X1 U6433 ( .A(n9099), .ZN(n9105) );
  AND2_X1 U6434 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  NOR2_X1 U6435 ( .A1(n4832), .A2(n6370), .ZN(n8932) );
  INV_X1 U6436 ( .A(n8983), .ZN(n8978) );
  AND2_X1 U6437 ( .A1(n7822), .A2(n9971), .ZN(n9982) );
  INV_X1 U6438 ( .A(n9955), .ZN(n9987) );
  INV_X1 U6439 ( .A(n9982), .ZN(n9949) );
  OR2_X1 U6440 ( .A1(n6714), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6495) );
  XNOR2_X1 U6441 ( .A(n6402), .B(n6401), .ZN(n6480) );
  AND2_X1 U6442 ( .A1(n6099), .A2(n6118), .ZN(n7946) );
  INV_X1 U6443 ( .A(n9301), .ZN(n9311) );
  INV_X1 U6444 ( .A(n8382), .ZN(n9410) );
  AND2_X1 U6445 ( .A1(n5541), .A2(n5540), .ZN(n9212) );
  AND2_X1 U6446 ( .A1(n9381), .A2(n9380), .ZN(n9396) );
  INV_X1 U6447 ( .A(n9626), .ZN(n9838) );
  NOR2_X1 U6448 ( .A1(n9874), .A2(n9845), .ZN(n9688) );
  INV_X1 U6449 ( .A(n9773), .ZN(n9721) );
  INV_X1 U6450 ( .A(n9845), .ZN(n9858) );
  AND2_X1 U6451 ( .A1(n5362), .A2(n5348), .ZN(n7997) );
  AND2_X1 U6452 ( .A1(n5054), .A2(n5071), .ZN(n7336) );
  CLKBUF_X1 U6453 ( .A(n9790), .Z(n9786) );
  INV_X1 U6454 ( .A(n6717), .ZN(n6616) );
  AND2_X1 U6455 ( .A1(n6838), .A2(n6837), .ZN(n8724) );
  INV_X1 U6456 ( .A(n8657), .ZN(n8738) );
  NAND2_X1 U6457 ( .A1(n5867), .A2(n5866), .ZN(n8904) );
  INV_X1 U6458 ( .A(n9009), .ZN(n9044) );
  INV_X1 U6459 ( .A(n8532), .ZN(n8747) );
  OR2_X1 U6460 ( .A1(P2_U3150), .A2(n6885), .ZN(n9896) );
  AND2_X1 U6461 ( .A1(n6970), .A2(n9030), .ZN(n9037) );
  NAND2_X1 U6462 ( .A1(n5845), .A2(n9105), .ZN(n6522) );
  NAND2_X1 U6463 ( .A1(n10005), .A2(n9949), .ZN(n9108) );
  INV_X1 U6464 ( .A(n10005), .ZN(n10003) );
  INV_X1 U6465 ( .A(n6457), .ZN(n9145) );
  OR2_X1 U6466 ( .A1(n9990), .A2(n9982), .ZN(n9171) );
  AND2_X1 U6467 ( .A1(n6503), .A2(n6502), .ZN(n9990) );
  INV_X1 U6468 ( .A(n10029), .ZN(n6767) );
  AND2_X1 U6469 ( .A1(n6882), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6717) );
  XNOR2_X1 U6470 ( .A(n6397), .B(n6396), .ZN(n8178) );
  INV_X1 U6471 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10037) );
  INV_X1 U6472 ( .A(n6415), .ZN(n6416) );
  AOI21_X1 U6473 ( .B1(n6409), .B2(n5751), .A(n5750), .ZN(n5752) );
  INV_X1 U6474 ( .A(n9493), .ZN(n9731) );
  INV_X1 U6475 ( .A(n9307), .ZN(n9288) );
  INV_X1 U6476 ( .A(n9212), .ZN(n9324) );
  AND3_X1 U6477 ( .A1(n5400), .A2(n5399), .A3(n5398), .ZN(n9242) );
  OR2_X1 U6478 ( .A1(n9807), .A2(n8203), .ZN(n9370) );
  OR2_X1 U6479 ( .A1(n9807), .A2(n8461), .ZN(n9387) );
  OR2_X1 U6480 ( .A1(n9831), .A2(n7315), .ZN(n9626) );
  AND2_X1 U6481 ( .A1(n7273), .A2(n9601), .ZN(n9831) );
  NAND2_X1 U6482 ( .A1(n9876), .A2(n9860), .ZN(n9699) );
  OR2_X2 U6483 ( .A1(n6609), .A2(n7271), .ZN(n9874) );
  INV_X1 U6484 ( .A(n9618), .ZN(n9769) );
  AND3_X1 U6485 ( .A1(n9866), .A2(n9865), .A3(n9864), .ZN(n9875) );
  OR2_X1 U6486 ( .A1(n6609), .A2(n6608), .ZN(n9867) );
  INV_X2 U6487 ( .A(n9867), .ZN(n9869) );
  INV_X1 U6488 ( .A(n9841), .ZN(n9842) );
  INV_X1 U6489 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5123) );
  OAI21_X1 U6490 ( .B1(n4936), .B2(n4925), .A(n4924), .ZN(n4926) );
  NAND2_X1 U6491 ( .A1(n4926), .A2(SI_2_), .ZN(n4930) );
  INV_X1 U6492 ( .A(n4926), .ZN(n4928) );
  INV_X1 U6493 ( .A(SI_2_), .ZN(n4927) );
  NAND2_X1 U6494 ( .A1(n4928), .A2(n4927), .ZN(n4929) );
  AND2_X1 U6495 ( .A1(n4930), .A2(n4929), .ZN(n5148) );
  NAND2_X1 U6496 ( .A1(n5147), .A2(n4930), .ZN(n5171) );
  MUX2_X1 U6497 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4936), .Z(n4931) );
  NAND2_X1 U6498 ( .A1(n4931), .A2(SI_3_), .ZN(n4935) );
  INV_X1 U6499 ( .A(n4931), .ZN(n4933) );
  INV_X1 U6500 ( .A(SI_3_), .ZN(n4932) );
  NAND2_X1 U6501 ( .A1(n4933), .A2(n4932), .ZN(n4934) );
  AND2_X1 U6502 ( .A1(n4935), .A2(n4934), .ZN(n5170) );
  NAND2_X1 U6503 ( .A1(n5171), .A2(n5170), .ZN(n5173) );
  NAND2_X1 U6504 ( .A1(n5173), .A2(n4935), .ZN(n5204) );
  NAND2_X1 U6505 ( .A1(n4939), .A2(SI_4_), .ZN(n4941) );
  NAND2_X1 U6506 ( .A1(n5204), .A2(n5203), .ZN(n5206) );
  NAND2_X1 U6507 ( .A1(n5206), .A2(n4941), .ZN(n5218) );
  MUX2_X1 U6508 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4936), .Z(n4942) );
  NAND2_X1 U6509 ( .A1(n4942), .A2(SI_5_), .ZN(n4946) );
  INV_X1 U6510 ( .A(n4942), .ZN(n4944) );
  INV_X1 U6511 ( .A(SI_5_), .ZN(n4943) );
  NAND2_X1 U6512 ( .A1(n4944), .A2(n4943), .ZN(n4945) );
  AND2_X1 U6513 ( .A1(n4946), .A2(n4945), .ZN(n5217) );
  MUX2_X1 U6514 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4936), .Z(n4947) );
  NAND2_X1 U6515 ( .A1(n4947), .A2(SI_6_), .ZN(n4951) );
  INV_X1 U6516 ( .A(n4947), .ZN(n4949) );
  INV_X1 U6517 ( .A(SI_6_), .ZN(n4948) );
  NAND2_X1 U6518 ( .A1(n4949), .A2(n4948), .ZN(n4950) );
  AND2_X1 U6519 ( .A1(n4951), .A2(n4950), .ZN(n5239) );
  MUX2_X1 U6520 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6631), .Z(n4953) );
  XNOR2_X1 U6521 ( .A(n4953), .B(SI_8_), .ZN(n5288) );
  INV_X1 U6522 ( .A(n4953), .ZN(n4955) );
  INV_X1 U6523 ( .A(SI_8_), .ZN(n4954) );
  NAND2_X1 U6524 ( .A1(n4955), .A2(n4954), .ZN(n4956) );
  INV_X1 U6525 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4957) );
  MUX2_X1 U6526 ( .A(n6656), .B(n4957), .S(n6631), .Z(n4959) );
  XNOR2_X1 U6527 ( .A(n4959), .B(SI_9_), .ZN(n5087) );
  INV_X1 U6528 ( .A(SI_9_), .ZN(n4958) );
  NAND2_X1 U6529 ( .A1(n4959), .A2(n4958), .ZN(n4960) );
  MUX2_X1 U6530 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6631), .Z(n4961) );
  NAND2_X1 U6531 ( .A1(n4961), .A2(SI_10_), .ZN(n4963) );
  OAI21_X1 U6532 ( .B1(n4961), .B2(SI_10_), .A(n4963), .ZN(n5046) );
  NAND2_X1 U6533 ( .A1(n5048), .A2(n4963), .ZN(n5070) );
  MUX2_X1 U6534 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6631), .Z(n4964) );
  XNOR2_X1 U6535 ( .A(n4964), .B(SI_11_), .ZN(n5069) );
  MUX2_X1 U6536 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6631), .Z(n4965) );
  NAND2_X1 U6537 ( .A1(n4965), .A2(SI_12_), .ZN(n4966) );
  OAI21_X1 U6538 ( .B1(n4965), .B2(SI_12_), .A(n4966), .ZN(n5312) );
  MUX2_X1 U6539 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6631), .Z(n4967) );
  INV_X1 U6540 ( .A(n4967), .ZN(n4969) );
  INV_X1 U6541 ( .A(SI_13_), .ZN(n4968) );
  NAND2_X1 U6542 ( .A1(n4969), .A2(n4968), .ZN(n4970) );
  OR2_X1 U6543 ( .A1(n4972), .A2(n4971), .ZN(n4973) );
  NAND2_X1 U6544 ( .A1(n5343), .A2(n4973), .ZN(n6786) );
  INV_X1 U6545 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4976) );
  NOR2_X1 U6546 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4978) );
  NAND4_X1 U6547 ( .A1(n4978), .A2(n5013), .A3(n4721), .A4(n5018), .ZN(n4981)
         );
  NAND4_X1 U6548 ( .A1(n4999), .A2(n4998), .A3(n5020), .A4(n4979), .ZN(n4980)
         );
  INV_X1 U6549 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4983) );
  XNOR2_X1 U6550 ( .A(n5025), .B(n4986), .ZN(n5727) );
  NAND2_X1 U6551 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n4988) );
  NAND2_X1 U6552 ( .A1(n5199), .A2(n4723), .ZN(n5317) );
  NOR2_X1 U6553 ( .A1(n5317), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n4993) );
  OR2_X1 U6554 ( .A1(n4993), .A2(n5243), .ZN(n4991) );
  MUX2_X1 U6555 ( .A(n4991), .B(P1_IR_REG_31__SCAN_IN), .S(n4992), .Z(n4994)
         );
  NAND2_X1 U6556 ( .A1(n4993), .A2(n4992), .ZN(n5345) );
  AOI22_X1 U6557 ( .A1(n4326), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4319), .B2(
        n7996), .ZN(n4995) );
  NAND2_X1 U6558 ( .A1(n5013), .A2(n4999), .ZN(n5000) );
  NAND2_X1 U6559 ( .A1(n5003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5004) );
  AND2_X1 U6560 ( .A1(n8197), .A2(n8175), .ZN(n5005) );
  INV_X1 U6561 ( .A(n5008), .ZN(n5009) );
  NAND2_X1 U6562 ( .A1(n5009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5010) );
  MUX2_X1 U6563 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5010), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5011) );
  INV_X1 U6564 ( .A(n5016), .ZN(n5017) );
  NAND2_X1 U6565 ( .A1(n5415), .A2(n5018), .ZN(n5019) );
  NAND2_X1 U6566 ( .A1(n5019), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6567 ( .A1(n5434), .A2(n5433), .ZN(n5436) );
  XNOR2_X2 U6568 ( .A(n5021), .B(n5020), .ZN(n5462) );
  INV_X1 U6569 ( .A(n6562), .ZN(n5023) );
  INV_X1 U6570 ( .A(n5128), .ZN(n5040) );
  INV_X2 U6571 ( .A(n5303), .ZN(n5376) );
  NAND2_X1 U6572 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5024) );
  NAND2_X1 U6573 ( .A1(n5025), .A2(n5024), .ZN(n5026) );
  XNOR2_X2 U6574 ( .A(n5026), .B(n9781), .ZN(n5034) );
  INV_X1 U6575 ( .A(n5029), .ZN(n5028) );
  NAND2_X1 U6576 ( .A1(n5028), .A2(n5027), .ZN(n5031) );
  NAND2_X1 U6577 ( .A1(n5029), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U6578 ( .A1(n5225), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5272) );
  NOR2_X1 U6579 ( .A1(n5272), .A2(n6733), .ZN(n5271) );
  NAND2_X1 U6580 ( .A1(n5271), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6581 ( .A1(n5324), .A2(n5032), .ZN(n5033) );
  AND2_X1 U6582 ( .A1(n5351), .A2(n5033), .ZN(n7873) );
  NAND2_X1 U6583 ( .A1(n5140), .A2(n7873), .ZN(n5039) );
  NAND2_X1 U6584 ( .A1(n4323), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6585 ( .A1(n4322), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6586 ( .A1(n5165), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5036) );
  NAND4_X1 U6587 ( .A1(n5039), .A2(n5038), .A3(n5037), .A4(n5036), .ZN(n9333)
         );
  AOI22_X1 U6588 ( .A1(n7813), .A2(n5695), .B1(n5376), .B2(n9333), .ZN(n5340)
         );
  NOR2_X1 U6589 ( .A1(n6562), .A2(n7314), .ZN(n5041) );
  NAND2_X1 U6590 ( .A1(n7813), .A2(n5657), .ZN(n5043) );
  NAND2_X1 U6591 ( .A1(n9333), .A2(n5695), .ZN(n5042) );
  NAND2_X1 U6592 ( .A1(n5043), .A2(n5042), .ZN(n5044) );
  XNOR2_X1 U6593 ( .A(n5044), .B(n5619), .ZN(n5341) );
  NAND2_X1 U6594 ( .A1(n5045), .A2(n5046), .ZN(n5047) );
  NAND2_X1 U6595 ( .A1(n5048), .A2(n5047), .ZN(n6660) );
  OR2_X1 U6596 ( .A1(n6660), .A2(n5316), .ZN(n5056) );
  INV_X1 U6597 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U6598 ( .A1(n5199), .A2(n5049), .ZN(n5221) );
  NOR2_X1 U6599 ( .A1(n5221), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5244) );
  NOR2_X1 U6600 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5050) );
  NAND2_X1 U6601 ( .A1(n5244), .A2(n5050), .ZN(n5290) );
  NAND2_X1 U6602 ( .A1(n5051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5053) );
  INV_X1 U6603 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5052) );
  OR2_X1 U6604 ( .A1(n5053), .A2(n5052), .ZN(n5054) );
  NAND2_X1 U6605 ( .A1(n5053), .A2(n5052), .ZN(n5071) );
  AOI22_X1 U6606 ( .A1(n4326), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4320), .B2(
        n7336), .ZN(n5055) );
  NAND2_X1 U6607 ( .A1(n7753), .A2(n5657), .ZN(n5064) );
  INV_X1 U6608 ( .A(n5057), .ZN(n5077) );
  NAND2_X1 U6609 ( .A1(n5095), .A2(n7749), .ZN(n5058) );
  AND2_X1 U6610 ( .A1(n5077), .A2(n5058), .ZN(n7752) );
  NAND2_X1 U6611 ( .A1(n5140), .A2(n7752), .ZN(n5062) );
  NAND2_X1 U6612 ( .A1(n4323), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6613 ( .A1(n4324), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6614 ( .A1(n5165), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5059) );
  NAND4_X1 U6615 ( .A1(n5062), .A2(n5061), .A3(n5060), .A4(n5059), .ZN(n9336)
         );
  NAND2_X1 U6616 ( .A1(n9336), .A2(n5281), .ZN(n5063) );
  NAND2_X1 U6617 ( .A1(n5064), .A2(n5063), .ZN(n5066) );
  XNOR2_X1 U6618 ( .A(n5066), .B(n5640), .ZN(n7748) );
  NAND2_X1 U6619 ( .A1(n7753), .A2(n5695), .ZN(n5068) );
  NAND2_X1 U6620 ( .A1(n9336), .A2(n5376), .ZN(n5067) );
  NAND2_X1 U6621 ( .A1(n5068), .A2(n5067), .ZN(n5308) );
  XNOR2_X1 U6622 ( .A(n5070), .B(n5069), .ZN(n6720) );
  NAND2_X1 U6623 ( .A1(n6720), .A2(n8313), .ZN(n5074) );
  NAND2_X1 U6624 ( .A1(n5071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5072) );
  XNOR2_X1 U6625 ( .A(n5072), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7574) );
  AOI22_X1 U6626 ( .A1(n4326), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7574), .B2(
        n4320), .ZN(n5073) );
  NAND2_X1 U6627 ( .A1(n7889), .A2(n5657), .ZN(n5084) );
  INV_X1 U6628 ( .A(n5075), .ZN(n5322) );
  INV_X1 U6629 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6630 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  AND2_X1 U6631 ( .A1(n5322), .A2(n5078), .ZN(n7884) );
  NAND2_X1 U6632 ( .A1(n5140), .A2(n7884), .ZN(n5082) );
  NAND2_X1 U6633 ( .A1(n4323), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6634 ( .A1(n4324), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6635 ( .A1(n5165), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5079) );
  NAND4_X1 U6636 ( .A1(n5082), .A2(n5081), .A3(n5080), .A4(n5079), .ZN(n9335)
         );
  NAND2_X1 U6637 ( .A1(n9335), .A2(n5695), .ZN(n5083) );
  NAND2_X1 U6638 ( .A1(n5084), .A2(n5083), .ZN(n5085) );
  INV_X2 U6639 ( .A(n5640), .ZN(n5693) );
  XNOR2_X1 U6640 ( .A(n5085), .B(n5693), .ZN(n5310) );
  AND2_X1 U6641 ( .A1(n5376), .A2(n9335), .ZN(n5086) );
  AOI21_X1 U6642 ( .B1(n7889), .B2(n5695), .A(n5086), .ZN(n5309) );
  NOR2_X1 U6643 ( .A1(n5310), .A2(n5309), .ZN(n7881) );
  XNOR2_X1 U6644 ( .A(n5088), .B(n5087), .ZN(n6654) );
  NAND2_X1 U6645 ( .A1(n6654), .A2(n8313), .ZN(n5092) );
  NAND2_X1 U6646 ( .A1(n5089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6647 ( .A(n5090), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7200) );
  AOI22_X1 U6648 ( .A1(n4326), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4319), .B2(
        n7200), .ZN(n5091) );
  NAND2_X1 U6649 ( .A1(n7524), .A2(n5657), .ZN(n5101) );
  NAND2_X1 U6650 ( .A1(n5297), .A2(n5093), .ZN(n5094) );
  AND2_X1 U6651 ( .A1(n5095), .A2(n5094), .ZN(n7481) );
  NAND2_X1 U6652 ( .A1(n5140), .A2(n7481), .ZN(n5099) );
  NAND2_X1 U6653 ( .A1(n4323), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6654 ( .A1(n5165), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6655 ( .A1(n4322), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5096) );
  NAND4_X1 U6656 ( .A1(n5099), .A2(n5098), .A3(n5097), .A4(n5096), .ZN(n9337)
         );
  NAND2_X1 U6657 ( .A1(n9337), .A2(n5695), .ZN(n5100) );
  NAND2_X1 U6658 ( .A1(n5101), .A2(n5100), .ZN(n5102) );
  XNOR2_X1 U6659 ( .A(n5102), .B(n5619), .ZN(n7474) );
  NAND2_X1 U6660 ( .A1(n7524), .A2(n5695), .ZN(n5104) );
  NAND2_X1 U6661 ( .A1(n9337), .A2(n5376), .ZN(n5103) );
  NAND2_X1 U6662 ( .A1(n5104), .A2(n5103), .ZN(n5306) );
  INV_X1 U6663 ( .A(n5306), .ZN(n7473) );
  NAND2_X1 U6664 ( .A1(n5140), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6665 ( .A1(n5165), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6666 ( .A1(n6526), .A2(n5122), .ZN(n5115) );
  XNOR2_X1 U6667 ( .A(n5110), .B(n5109), .ZN(n5964) );
  INV_X1 U6668 ( .A(n5964), .ZN(n6643) );
  NAND2_X1 U6669 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9798), .ZN(n5111) );
  XNOR2_X1 U6670 ( .A(n5111), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U6671 ( .A1(n4318), .A2(n6666), .ZN(n5112) );
  NAND2_X1 U6672 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  AOI22_X1 U6673 ( .A1(n6526), .A2(n5376), .B1(n5122), .B2(n7321), .ZN(n5136)
         );
  NAND2_X1 U6674 ( .A1(n4324), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6675 ( .A1(n5140), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U6676 ( .A1(n5165), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U6677 ( .A1(n5119), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U6678 ( .A1(n6524), .A2(n5122), .ZN(n5127) );
  NAND2_X1 U6679 ( .A1(n6631), .A2(SI_0_), .ZN(n5124) );
  XNOR2_X1 U6680 ( .A(n5124), .B(n5123), .ZN(n9794) );
  MUX2_X1 U6681 ( .A(n4519), .B(n9794), .S(n5125), .Z(n7317) );
  INV_X1 U6682 ( .A(n7317), .ZN(n9849) );
  NAND2_X1 U6683 ( .A1(n5145), .A2(n9849), .ZN(n5126) );
  NAND2_X1 U6684 ( .A1(n6524), .A2(n5376), .ZN(n5132) );
  NAND2_X1 U6685 ( .A1(n5128), .A2(n9798), .ZN(n5129) );
  OAI21_X1 U6686 ( .B1(n5690), .B2(n7317), .A(n5129), .ZN(n5130) );
  INV_X1 U6687 ( .A(n5130), .ZN(n5131) );
  NAND2_X1 U6688 ( .A1(n5132), .A2(n5131), .ZN(n6750) );
  NAND2_X1 U6689 ( .A1(n6751), .A2(n6750), .ZN(n6749) );
  NAND2_X1 U6690 ( .A1(n5133), .A2(n5693), .ZN(n5134) );
  NAND2_X1 U6691 ( .A1(n6770), .A2(n6771), .ZN(n5139) );
  INV_X1 U6692 ( .A(n5135), .ZN(n5137) );
  NAND2_X1 U6693 ( .A1(n5137), .A2(n5136), .ZN(n5138) );
  NAND2_X1 U6694 ( .A1(n5140), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6695 ( .A1(n4324), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6696 ( .A1(n5165), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6697 ( .A1(n9344), .A2(n5281), .ZN(n5158) );
  NAND2_X1 U6698 ( .A1(n5146), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5156) );
  OR2_X1 U6699 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  NAND2_X1 U6700 ( .A1(n5147), .A2(n5150), .ZN(n6642) );
  NAND2_X1 U6701 ( .A1(n4318), .A2(n9354), .ZN(n5154) );
  NAND2_X1 U6702 ( .A1(n5145), .A2(n6963), .ZN(n5157) );
  NAND2_X1 U6703 ( .A1(n5158), .A2(n5157), .ZN(n5159) );
  XNOR2_X1 U6704 ( .A(n5159), .B(n5693), .ZN(n5164) );
  NAND2_X1 U6705 ( .A1(n9344), .A2(n5376), .ZN(n5161) );
  NAND2_X1 U6706 ( .A1(n6963), .A2(n5281), .ZN(n5160) );
  NAND2_X1 U6707 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  XNOR2_X1 U6708 ( .A(n5164), .B(n5162), .ZN(n6777) );
  NAND2_X1 U6709 ( .A1(n6778), .A2(n6777), .ZN(n6803) );
  INV_X1 U6710 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6711 ( .A1(n5164), .A2(n5163), .ZN(n6802) );
  INV_X1 U6712 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7376) );
  NAND2_X1 U6713 ( .A1(n5140), .A2(n7376), .ZN(n5169) );
  NAND2_X1 U6714 ( .A1(n4323), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6715 ( .A1(n5165), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6716 ( .A1(n4324), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6717 ( .A1(n9343), .A2(n5281), .ZN(n5180) );
  OR2_X1 U6718 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  NAND2_X1 U6719 ( .A1(n5173), .A2(n5172), .ZN(n6640) );
  NAND2_X1 U6720 ( .A1(n4326), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5176) );
  OR2_X1 U6721 ( .A1(n5153), .A2(n5243), .ZN(n5174) );
  XNOR2_X1 U6722 ( .A(n5174), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U6723 ( .A1(n4319), .A2(n6685), .ZN(n5175) );
  AND3_X2 U6724 ( .A1(n5177), .A2(n5176), .A3(n5175), .ZN(n7379) );
  NAND2_X1 U6725 ( .A1(n5145), .A2(n5178), .ZN(n5179) );
  NAND2_X1 U6726 ( .A1(n5180), .A2(n5179), .ZN(n5181) );
  XNOR2_X1 U6727 ( .A(n5181), .B(n5693), .ZN(n5187) );
  NAND2_X1 U6728 ( .A1(n9343), .A2(n5376), .ZN(n5183) );
  NAND2_X1 U6729 ( .A1(n5178), .A2(n5281), .ZN(n5182) );
  NAND2_X1 U6730 ( .A1(n5183), .A2(n5182), .ZN(n5186) );
  INV_X1 U6731 ( .A(n5186), .ZN(n5184) );
  NAND2_X1 U6732 ( .A1(n5187), .A2(n5184), .ZN(n5188) );
  AND2_X1 U6733 ( .A1(n6802), .A2(n5188), .ZN(n5185) );
  NAND2_X1 U6734 ( .A1(n6803), .A2(n5185), .ZN(n5191) );
  XNOR2_X1 U6735 ( .A(n5187), .B(n5186), .ZN(n6805) );
  INV_X1 U6736 ( .A(n6805), .ZN(n5189) );
  NAND2_X1 U6737 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  NAND2_X1 U6738 ( .A1(n5191), .A2(n5190), .ZN(n6999) );
  INV_X1 U6739 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6740 ( .A1(n7376), .A2(n5192), .ZN(n5194) );
  INV_X1 U6741 ( .A(n5193), .ZN(n5226) );
  AND2_X1 U6742 ( .A1(n5194), .A2(n5226), .ZN(n7327) );
  NAND2_X1 U6743 ( .A1(n5140), .A2(n7327), .ZN(n5198) );
  NAND2_X1 U6744 ( .A1(n4323), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6745 ( .A1(n4324), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6746 ( .A1(n5165), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6747 ( .A1(n9342), .A2(n5281), .ZN(n5210) );
  NOR2_X1 U6748 ( .A1(n5199), .A2(n5243), .ZN(n5200) );
  MUX2_X1 U6749 ( .A(n5243), .B(n5200), .S(P1_IR_REG_4__SCAN_IN), .Z(n5202) );
  INV_X1 U6750 ( .A(n5221), .ZN(n5201) );
  NOR2_X1 U6751 ( .A1(n5202), .A2(n5201), .ZN(n6686) );
  AOI22_X1 U6752 ( .A1(n4326), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n4320), .B2(
        n6686), .ZN(n5208) );
  OR2_X1 U6753 ( .A1(n5204), .A2(n5203), .ZN(n5205) );
  NAND2_X1 U6754 ( .A1(n5206), .A2(n5205), .ZN(n6635) );
  OR2_X1 U6755 ( .A1(n6635), .A2(n5316), .ZN(n5207) );
  INV_X1 U6756 ( .A(n7326), .ZN(n7004) );
  NAND2_X1 U6757 ( .A1(n5145), .A2(n7004), .ZN(n5209) );
  NAND2_X1 U6758 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  XNOR2_X1 U6759 ( .A(n5211), .B(n5619), .ZN(n5214) );
  NAND2_X1 U6760 ( .A1(n9342), .A2(n5376), .ZN(n5212) );
  OAI21_X1 U6761 ( .B1(n7326), .B2(n5690), .A(n5212), .ZN(n5213) );
  NAND2_X1 U6762 ( .A1(n5214), .A2(n5213), .ZN(n5236) );
  OR2_X1 U6763 ( .A1(n5214), .A2(n5213), .ZN(n5215) );
  NAND2_X1 U6764 ( .A1(n5236), .A2(n5215), .ZN(n7003) );
  INV_X1 U6765 ( .A(n7003), .ZN(n5216) );
  NAND2_X1 U6766 ( .A1(n6999), .A2(n5216), .ZN(n7000) );
  INV_X1 U6767 ( .A(n5145), .ZN(n5496) );
  OR2_X1 U6768 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  NAND2_X1 U6769 ( .A1(n5220), .A2(n5219), .ZN(n6649) );
  OR2_X1 U6770 ( .A1(n6649), .A2(n5316), .ZN(n5224) );
  NAND2_X1 U6771 ( .A1(n5221), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5222) );
  XNOR2_X1 U6772 ( .A(n5222), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6698) );
  AOI22_X1 U6773 ( .A1(n4326), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n4320), .B2(
        n6698), .ZN(n5223) );
  INV_X1 U6774 ( .A(n5225), .ZN(n5248) );
  INV_X1 U6775 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U6776 ( .A1(n5226), .A2(n6693), .ZN(n5227) );
  AND2_X1 U6777 ( .A1(n5248), .A2(n5227), .ZN(n7486) );
  NAND2_X1 U6778 ( .A1(n5140), .A2(n7486), .ZN(n5231) );
  NAND2_X1 U6779 ( .A1(n4323), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6780 ( .A1(n4324), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6781 ( .A1(n5165), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5228) );
  NAND4_X1 U6782 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n9341)
         );
  NAND2_X1 U6783 ( .A1(n9341), .A2(n5281), .ZN(n5232) );
  OAI21_X1 U6784 ( .B1(n5496), .B2(n6955), .A(n5232), .ZN(n5233) );
  AND2_X1 U6785 ( .A1(n4919), .A2(n5236), .ZN(n5234) );
  NAND2_X1 U6786 ( .A1(n7000), .A2(n5234), .ZN(n6992) );
  OR2_X1 U6787 ( .A1(n4919), .A2(n5236), .ZN(n6989) );
  AOI22_X1 U6788 ( .A1(n7487), .A2(n5695), .B1(n5376), .B2(n9341), .ZN(n6993)
         );
  AND2_X1 U6789 ( .A1(n6989), .A2(n6993), .ZN(n5237) );
  NAND2_X1 U6790 ( .A1(n6990), .A2(n5237), .ZN(n5238) );
  NAND2_X1 U6791 ( .A1(n6992), .A2(n5238), .ZN(n7032) );
  OR2_X1 U6792 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6793 ( .A1(n5242), .A2(n5241), .ZN(n6647) );
  OR2_X1 U6794 ( .A1(n6647), .A2(n5316), .ZN(n5246) );
  OR2_X1 U6795 ( .A1(n5244), .A2(n5243), .ZN(n5266) );
  XNOR2_X1 U6796 ( .A(n5266), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6727) );
  AOI22_X1 U6797 ( .A1(n4326), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n4320), .B2(
        n6727), .ZN(n5245) );
  NAND2_X1 U6798 ( .A1(n5246), .A2(n5245), .ZN(n9818) );
  NAND2_X1 U6799 ( .A1(n9818), .A2(n5145), .ZN(n5255) );
  INV_X1 U6800 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6801 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  AND2_X1 U6802 ( .A1(n5272), .A2(n5249), .ZN(n9820) );
  NAND2_X1 U6803 ( .A1(n5140), .A2(n9820), .ZN(n5253) );
  NAND2_X1 U6804 ( .A1(n4323), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6805 ( .A1(n5165), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6806 ( .A1(n4324), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5250) );
  NAND4_X1 U6807 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n9340)
         );
  NAND2_X1 U6808 ( .A1(n9340), .A2(n5281), .ZN(n5254) );
  NAND2_X1 U6809 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  XNOR2_X1 U6810 ( .A(n5256), .B(n5693), .ZN(n5261) );
  INV_X1 U6811 ( .A(n5261), .ZN(n5259) );
  AND2_X1 U6812 ( .A1(n5376), .A2(n9340), .ZN(n5257) );
  AOI21_X1 U6813 ( .B1(n9818), .B2(n5695), .A(n5257), .ZN(n5260) );
  INV_X1 U6814 ( .A(n5260), .ZN(n5258) );
  NAND2_X1 U6815 ( .A1(n5259), .A2(n5258), .ZN(n7029) );
  AND2_X1 U6816 ( .A1(n5261), .A2(n5260), .ZN(n7028) );
  NAND2_X1 U6817 ( .A1(n5264), .A2(n5263), .ZN(n6645) );
  OR2_X1 U6818 ( .A1(n6645), .A2(n5316), .ZN(n5270) );
  INV_X1 U6819 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6820 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  NAND2_X1 U6821 ( .A1(n5267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5268) );
  XNOR2_X1 U6822 ( .A(n5268), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U6823 ( .A1(n4326), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4319), .B2(
        n6788), .ZN(n5269) );
  NAND2_X1 U6824 ( .A1(n5270), .A2(n5269), .ZN(n7514) );
  NAND2_X1 U6825 ( .A1(n7514), .A2(n5145), .ZN(n5279) );
  INV_X1 U6826 ( .A(n5271), .ZN(n5295) );
  NAND2_X1 U6827 ( .A1(n5272), .A2(n6733), .ZN(n5273) );
  AND2_X1 U6828 ( .A1(n5295), .A2(n5273), .ZN(n9808) );
  NAND2_X1 U6829 ( .A1(n5140), .A2(n9808), .ZN(n5277) );
  NAND2_X1 U6830 ( .A1(n4323), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6831 ( .A1(n4322), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6832 ( .A1(n5165), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5274) );
  NAND4_X1 U6833 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(n9339)
         );
  NAND2_X1 U6834 ( .A1(n9339), .A2(n5281), .ZN(n5278) );
  NAND2_X1 U6835 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  XNOR2_X1 U6836 ( .A(n5280), .B(n5619), .ZN(n5287) );
  INV_X1 U6837 ( .A(n5287), .ZN(n5285) );
  NAND2_X1 U6838 ( .A1(n7514), .A2(n5281), .ZN(n5283) );
  NAND2_X1 U6839 ( .A1(n9339), .A2(n5376), .ZN(n5282) );
  NAND2_X1 U6840 ( .A1(n5283), .A2(n5282), .ZN(n5286) );
  INV_X1 U6841 ( .A(n5286), .ZN(n5284) );
  NAND2_X1 U6842 ( .A1(n5285), .A2(n5284), .ZN(n7120) );
  AND2_X1 U6843 ( .A1(n5287), .A2(n5286), .ZN(n7121) );
  AOI21_X2 U6844 ( .B1(n7124), .B2(n7120), .A(n7121), .ZN(n5305) );
  XNOR2_X1 U6845 ( .A(n5289), .B(n5288), .ZN(n6650) );
  NAND2_X1 U6846 ( .A1(n6650), .A2(n8313), .ZN(n5293) );
  NAND2_X1 U6847 ( .A1(n5290), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5291) );
  XNOR2_X1 U6848 ( .A(n5291), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6920) );
  AOI22_X1 U6849 ( .A1(n4326), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4319), .B2(
        n6920), .ZN(n5292) );
  NAND2_X1 U6850 ( .A1(n5293), .A2(n5292), .ZN(n9861) );
  INV_X1 U6851 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6852 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  AND2_X1 U6853 ( .A1(n5297), .A2(n5296), .ZN(n7443) );
  NAND2_X1 U6854 ( .A1(n5140), .A2(n7443), .ZN(n5301) );
  NAND2_X1 U6855 ( .A1(n4323), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6856 ( .A1(n5165), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6857 ( .A1(n4324), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5298) );
  NAND4_X1 U6858 ( .A1(n5301), .A2(n5300), .A3(n5299), .A4(n5298), .ZN(n9338)
         );
  AOI22_X1 U6859 ( .A1(n9861), .A2(n5145), .B1(n5695), .B2(n9338), .ZN(n5302)
         );
  XNOR2_X1 U6860 ( .A(n5302), .B(n5640), .ZN(n5304) );
  XNOR2_X1 U6861 ( .A(n5305), .B(n5304), .ZN(n7296) );
  INV_X1 U6862 ( .A(n9861), .ZN(n7442) );
  INV_X1 U6863 ( .A(n9338), .ZN(n7125) );
  OAI22_X1 U6864 ( .A1(n7442), .A2(n5690), .B1(n7125), .B2(n5697), .ZN(n7295)
         );
  INV_X1 U6865 ( .A(n7748), .ZN(n7877) );
  INV_X1 U6866 ( .A(n5308), .ZN(n7879) );
  NAND2_X1 U6867 ( .A1(n7877), .A2(n7879), .ZN(n5311) );
  NAND2_X1 U6868 ( .A1(n5310), .A2(n5309), .ZN(n7919) );
  OAI21_X1 U6869 ( .B1(n7881), .B2(n5311), .A(n7919), .ZN(n5338) );
  NAND2_X1 U6870 ( .A1(n5313), .A2(n5312), .ZN(n5315) );
  NAND2_X1 U6871 ( .A1(n5315), .A2(n5314), .ZN(n6769) );
  NAND2_X1 U6872 ( .A1(n5317), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6873 ( .A(n5318), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7669) );
  AOI22_X1 U6874 ( .A1(n4326), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4320), .B2(
        n7669), .ZN(n5319) );
  NAND2_X1 U6875 ( .A1(n7699), .A2(n5657), .ZN(n5330) );
  INV_X1 U6876 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6877 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  AND2_X1 U6878 ( .A1(n5324), .A2(n5323), .ZN(n7929) );
  NAND2_X1 U6879 ( .A1(n5140), .A2(n7929), .ZN(n5328) );
  NAND2_X1 U6880 ( .A1(n4323), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6881 ( .A1(n5165), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6882 ( .A1(n4324), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5325) );
  NAND4_X1 U6883 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n9334)
         );
  NAND2_X1 U6884 ( .A1(n9334), .A2(n5695), .ZN(n5329) );
  NAND2_X1 U6885 ( .A1(n5330), .A2(n5329), .ZN(n5331) );
  XNOR2_X1 U6886 ( .A(n5331), .B(n5693), .ZN(n5333) );
  AND2_X1 U6887 ( .A1(n5376), .A2(n9334), .ZN(n5332) );
  AOI21_X1 U6888 ( .B1(n7699), .B2(n5695), .A(n5332), .ZN(n5334) );
  NAND2_X1 U6889 ( .A1(n5333), .A2(n5334), .ZN(n5339) );
  INV_X1 U6890 ( .A(n5333), .ZN(n5336) );
  INV_X1 U6891 ( .A(n5334), .ZN(n5335) );
  NAND2_X1 U6892 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  AND2_X1 U6893 ( .A1(n5339), .A2(n5337), .ZN(n7920) );
  XNOR2_X1 U6894 ( .A(n5341), .B(n5340), .ZN(n7868) );
  MUX2_X1 U6895 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6631), .Z(n5359) );
  XNOR2_X1 U6896 ( .A(n5359), .B(SI_14_), .ZN(n5344) );
  XNOR2_X1 U6897 ( .A(n5360), .B(n5344), .ZN(n6816) );
  NAND2_X1 U6898 ( .A1(n6816), .A2(n8313), .ZN(n5350) );
  NAND2_X1 U6899 ( .A1(n5345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6900 ( .A1(n5347), .A2(n5346), .ZN(n5362) );
  OR2_X1 U6901 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  AOI22_X1 U6902 ( .A1(n4326), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4320), .B2(
        n7997), .ZN(n5349) );
  NAND2_X1 U6903 ( .A1(n5351), .A2(n9189), .ZN(n5352) );
  AND2_X1 U6904 ( .A1(n5366), .A2(n5352), .ZN(n9194) );
  NAND2_X1 U6905 ( .A1(n5140), .A2(n9194), .ZN(n5356) );
  NAND2_X1 U6906 ( .A1(n4323), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6907 ( .A1(n4324), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6908 ( .A1(n5165), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5353) );
  NAND4_X1 U6909 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n9332)
         );
  AOI22_X1 U6910 ( .A1(n9702), .A2(n5657), .B1(n5695), .B2(n9332), .ZN(n5357)
         );
  XNOR2_X1 U6911 ( .A(n5357), .B(n5640), .ZN(n5358) );
  AOI22_X1 U6912 ( .A1(n9702), .A2(n5695), .B1(n5376), .B2(n9332), .ZN(n9187)
         );
  MUX2_X1 U6913 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6631), .Z(n5382) );
  XNOR2_X1 U6914 ( .A(n5382), .B(SI_15_), .ZN(n5361) );
  XNOR2_X1 U6915 ( .A(n5381), .B(n5361), .ZN(n7038) );
  NAND2_X1 U6916 ( .A1(n7038), .A2(n8313), .ZN(n5365) );
  NAND2_X1 U6917 ( .A1(n5362), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5363) );
  XNOR2_X1 U6918 ( .A(n5363), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8481) );
  AOI22_X1 U6919 ( .A1(n4326), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4319), .B2(
        n8481), .ZN(n5364) );
  INV_X1 U6920 ( .A(n5394), .ZN(n5396) );
  NAND2_X1 U6921 ( .A1(n5366), .A2(n9309), .ZN(n5367) );
  AND2_X1 U6922 ( .A1(n5396), .A2(n5367), .ZN(n9314) );
  NAND2_X1 U6923 ( .A1(n5140), .A2(n9314), .ZN(n5371) );
  NAND2_X1 U6924 ( .A1(n4323), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6925 ( .A1(n4322), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6926 ( .A1(n5165), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5368) );
  NAND4_X1 U6927 ( .A1(n5371), .A2(n5370), .A3(n5369), .A4(n5368), .ZN(n9331)
         );
  INV_X1 U6928 ( .A(n9331), .ZN(n8164) );
  OAI22_X1 U6929 ( .A1(n9318), .A2(n5496), .B1(n8164), .B2(n5690), .ZN(n5372)
         );
  XNOR2_X1 U6930 ( .A(n5372), .B(n5619), .ZN(n5373) );
  NOR2_X1 U6931 ( .A1(n5374), .A2(n5373), .ZN(n5377) );
  AOI22_X1 U6932 ( .A1(n8012), .A2(n5695), .B1(n5376), .B2(n9331), .ZN(n9305)
         );
  NAND2_X1 U6933 ( .A1(n9306), .A2(n9305), .ZN(n9304) );
  INV_X1 U6934 ( .A(n5377), .ZN(n5378) );
  NAND2_X1 U6935 ( .A1(n9304), .A2(n5378), .ZN(n9229) );
  INV_X1 U6936 ( .A(SI_15_), .ZN(n5379) );
  NAND2_X1 U6937 ( .A1(n5380), .A2(n5379), .ZN(n5386) );
  INV_X1 U6938 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U6939 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  MUX2_X1 U6940 ( .A(n7217), .B(n5387), .S(n4936), .Z(n5406) );
  XNOR2_X1 U6941 ( .A(n5406), .B(SI_16_), .ZN(n5388) );
  NAND2_X1 U6942 ( .A1(n7188), .A2(n8313), .ZN(n5392) );
  NAND2_X1 U6943 ( .A1(n5389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5390) );
  XNOR2_X1 U6944 ( .A(n5390), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9366) );
  AOI22_X1 U6945 ( .A1(n4326), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4319), .B2(
        n9366), .ZN(n5391) );
  INV_X1 U6946 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9697) );
  INV_X1 U6947 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9771) );
  OAI22_X1 U6948 ( .A1(n5515), .A2(n9697), .B1(n8318), .B2(n9771), .ZN(n5393)
         );
  INV_X1 U6949 ( .A(n5393), .ZN(n5400) );
  NAND2_X1 U6950 ( .A1(n5394), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5419) );
  INV_X1 U6951 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6952 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  AND2_X1 U6953 ( .A1(n5419), .A2(n5397), .ZN(n9232) );
  NAND2_X1 U6954 ( .A1(n9232), .A2(n5140), .ZN(n5399) );
  NAND2_X1 U6955 ( .A1(n4323), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5398) );
  OAI22_X1 U6956 ( .A1(n9774), .A2(n5496), .B1(n9242), .B2(n5690), .ZN(n5401)
         );
  XNOR2_X1 U6957 ( .A(n5401), .B(n5640), .ZN(n5403) );
  OAI22_X1 U6958 ( .A1(n9774), .A2(n5690), .B1(n9242), .B2(n5697), .ZN(n5402)
         );
  NOR2_X1 U6959 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  AOI21_X1 U6960 ( .B1(n5403), .B2(n5402), .A(n5404), .ZN(n9230) );
  INV_X1 U6961 ( .A(n5404), .ZN(n5405) );
  NAND2_X1 U6962 ( .A1(n5407), .A2(SI_16_), .ZN(n5408) );
  MUX2_X1 U6963 ( .A(n10037), .B(n5410), .S(n6631), .Z(n5412) );
  INV_X1 U6964 ( .A(n5412), .ZN(n5413) );
  NAND2_X1 U6965 ( .A1(n5413), .A2(SI_17_), .ZN(n5414) );
  NAND2_X1 U6966 ( .A1(n5431), .A2(n5414), .ZN(n5430) );
  XNOR2_X1 U6967 ( .A(n5429), .B(n5430), .ZN(n7232) );
  NAND2_X1 U6968 ( .A1(n7232), .A2(n8313), .ZN(n5417) );
  XNOR2_X1 U6969 ( .A(n5415), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9375) );
  AOI22_X1 U6970 ( .A1(n4326), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4320), .B2(
        n9375), .ZN(n5416) );
  NAND2_X1 U6971 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  AND2_X1 U6972 ( .A1(n5440), .A2(n5420), .ZN(n9619) );
  NAND2_X1 U6973 ( .A1(n9619), .A2(n5140), .ZN(n5423) );
  AOI22_X1 U6974 ( .A1(n4322), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n5165), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6975 ( .A1(n4323), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5421) );
  OAI22_X1 U6976 ( .A1(n9769), .A2(n5690), .B1(n9282), .B2(n5697), .ZN(n5427)
         );
  NAND2_X1 U6977 ( .A1(n9618), .A2(n5657), .ZN(n5425) );
  OR2_X1 U6978 ( .A1(n9282), .A2(n5690), .ZN(n5424) );
  NAND2_X1 U6979 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  XNOR2_X1 U6980 ( .A(n5426), .B(n5619), .ZN(n5428) );
  XOR2_X1 U6981 ( .A(n5427), .B(n5428), .Z(n9240) );
  NAND2_X1 U6982 ( .A1(n5432), .A2(n5431), .ZN(n5453) );
  MUX2_X1 U6983 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6631), .Z(n5455) );
  XNOR2_X1 U6984 ( .A(n5455), .B(n10197), .ZN(n5454) );
  XNOR2_X1 U6985 ( .A(n5453), .B(n5454), .ZN(n7372) );
  NAND2_X1 U6986 ( .A1(n7372), .A2(n8313), .ZN(n5438) );
  OR2_X1 U6987 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  AND2_X1 U6988 ( .A1(n5436), .A2(n5435), .ZN(n9386) );
  AOI22_X1 U6989 ( .A1(n4326), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4319), .B2(
        n9386), .ZN(n5437) );
  NAND2_X1 U6990 ( .A1(n9684), .A2(n5657), .ZN(n5448) );
  INV_X1 U6991 ( .A(n5465), .ZN(n5467) );
  NAND2_X1 U6992 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  NAND2_X1 U6993 ( .A1(n5467), .A2(n5441), .ZN(n9602) );
  OR2_X1 U6994 ( .A1(n9602), .A2(n5728), .ZN(n5446) );
  INV_X1 U6995 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9685) );
  INV_X1 U6996 ( .A(n5165), .ZN(n8318) );
  INV_X1 U6997 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10202) );
  OAI22_X1 U6998 ( .A1(n5515), .A2(n9685), .B1(n8318), .B2(n10202), .ZN(n5443)
         );
  INV_X1 U6999 ( .A(n5443), .ZN(n5445) );
  NAND2_X1 U7000 ( .A1(n4323), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5444) );
  INV_X1 U7001 ( .A(n8520), .ZN(n9329) );
  NAND2_X1 U7002 ( .A1(n9329), .A2(n5695), .ZN(n5447) );
  NAND2_X1 U7003 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  XNOR2_X1 U7004 ( .A(n5449), .B(n5693), .ZN(n5452) );
  NOR2_X1 U7005 ( .A1(n8520), .A2(n5697), .ZN(n5450) );
  AOI21_X1 U7006 ( .B1(n9684), .B2(n5695), .A(n5450), .ZN(n5451) );
  AND2_X1 U7007 ( .A1(n5452), .A2(n5451), .ZN(n9276) );
  OR2_X1 U7008 ( .A1(n5452), .A2(n5451), .ZN(n9277) );
  NAND2_X1 U7009 ( .A1(n5455), .A2(SI_18_), .ZN(n5456) );
  MUX2_X1 U7010 ( .A(n7553), .B(n5457), .S(n4936), .Z(n5459) );
  INV_X1 U7011 ( .A(n5459), .ZN(n5460) );
  NAND2_X1 U7012 ( .A1(n5460), .A2(SI_19_), .ZN(n5461) );
  NAND2_X1 U7013 ( .A1(n5481), .A2(n5461), .ZN(n5482) );
  XNOR2_X1 U7014 ( .A(n5483), .B(n5482), .ZN(n7527) );
  NAND2_X1 U7015 ( .A1(n7527), .A2(n8313), .ZN(n5464) );
  AOI22_X1 U7016 ( .A1(n4326), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8455), .B2(
        n4320), .ZN(n5463) );
  NAND2_X1 U7017 ( .A1(n9589), .A2(n5657), .ZN(n5476) );
  INV_X1 U7018 ( .A(n5487), .ZN(n5489) );
  INV_X1 U7019 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7020 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  AND2_X1 U7021 ( .A1(n5489), .A2(n5468), .ZN(n8519) );
  NAND2_X1 U7022 ( .A1(n8519), .A2(n5140), .ZN(n5474) );
  INV_X1 U7023 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U7024 ( .A1(n4324), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7025 ( .A1(n5165), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5470) );
  OAI211_X1 U7026 ( .C1(n5731), .C2(n9582), .A(n5471), .B(n5470), .ZN(n5472)
         );
  INV_X1 U7027 ( .A(n5472), .ZN(n5473) );
  INV_X1 U7028 ( .A(n9283), .ZN(n9328) );
  NAND2_X1 U7029 ( .A1(n9328), .A2(n5695), .ZN(n5475) );
  NAND2_X1 U7030 ( .A1(n5476), .A2(n5475), .ZN(n5477) );
  XNOR2_X1 U7031 ( .A(n5477), .B(n5693), .ZN(n5480) );
  NOR2_X1 U7032 ( .A1(n9283), .A2(n5697), .ZN(n5478) );
  AOI21_X1 U7033 ( .B1(n9589), .B2(n5695), .A(n5478), .ZN(n5479) );
  NOR2_X1 U7034 ( .A1(n5480), .A2(n5479), .ZN(n8517) );
  NAND2_X1 U7035 ( .A1(n5480), .A2(n5479), .ZN(n8515) );
  MUX2_X1 U7036 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6631), .Z(n5502) );
  XNOR2_X1 U7037 ( .A(n5502), .B(n5504), .ZN(n5484) );
  XNOR2_X1 U7038 ( .A(n5505), .B(n5484), .ZN(n7702) );
  NAND2_X1 U7039 ( .A1(n7702), .A2(n8313), .ZN(n5486) );
  NAND2_X1 U7040 ( .A1(n4326), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5485) );
  INV_X1 U7041 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7042 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  NAND2_X1 U7043 ( .A1(n5511), .A2(n5490), .ZN(n9564) );
  OR2_X1 U7044 ( .A1(n9564), .A2(n5728), .ZN(n5495) );
  INV_X1 U7045 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U7046 ( .A1(n4324), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7047 ( .A1(n5165), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5491) );
  OAI211_X1 U7048 ( .C1(n5731), .C2(n9565), .A(n5492), .B(n5491), .ZN(n5493)
         );
  INV_X1 U7049 ( .A(n5493), .ZN(n5494) );
  OAI22_X1 U7050 ( .A1(n9563), .A2(n5496), .B1(n9211), .B2(n5690), .ZN(n5497)
         );
  XNOR2_X1 U7051 ( .A(n5497), .B(n5640), .ZN(n5499) );
  OAI22_X1 U7052 ( .A1(n9563), .A2(n5690), .B1(n9211), .B2(n5697), .ZN(n5498)
         );
  NOR2_X1 U7053 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AOI21_X1 U7054 ( .B1(n5499), .B2(n5498), .A(n5500), .ZN(n9262) );
  INV_X1 U7055 ( .A(n5500), .ZN(n5501) );
  INV_X1 U7056 ( .A(n5502), .ZN(n5503) );
  INV_X1 U7057 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n5506) );
  MUX2_X1 U7058 ( .A(n7849), .B(n5506), .S(n6631), .Z(n5524) );
  XNOR2_X1 U7059 ( .A(n5524), .B(SI_21_), .ZN(n5507) );
  NAND2_X1 U7060 ( .A1(n7806), .A2(n8313), .ZN(n5509) );
  NAND2_X1 U7061 ( .A1(n4326), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5508) );
  INV_X1 U7062 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7063 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  AND2_X1 U7064 ( .A1(n5535), .A2(n5512), .ZN(n9553) );
  NAND2_X1 U7065 ( .A1(n9553), .A2(n5140), .ZN(n5518) );
  INV_X1 U7066 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U7067 ( .A1(n4323), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7068 ( .A1(n5165), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5513) );
  OAI211_X1 U7069 ( .C1(n5515), .C2(n10171), .A(n5514), .B(n5513), .ZN(n5516)
         );
  INV_X1 U7070 ( .A(n5516), .ZN(n5517) );
  OAI22_X1 U7071 ( .A1(n9745), .A2(n5690), .B1(n9269), .B2(n5697), .ZN(n5522)
         );
  NAND2_X1 U7072 ( .A1(n9554), .A2(n5657), .ZN(n5520) );
  OR2_X1 U7073 ( .A1(n9269), .A2(n5690), .ZN(n5519) );
  NAND2_X1 U7074 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  XNOR2_X1 U7075 ( .A(n5521), .B(n5619), .ZN(n5523) );
  XOR2_X1 U7076 ( .A(n5522), .B(n5523), .Z(n9210) );
  INV_X1 U7077 ( .A(n5546), .ZN(n5544) );
  NOR2_X1 U7078 ( .A1(n5525), .A2(SI_21_), .ZN(n5526) );
  MUX2_X1 U7079 ( .A(n8018), .B(n5528), .S(n4936), .Z(n5530) );
  INV_X1 U7080 ( .A(SI_22_), .ZN(n5529) );
  NAND2_X1 U7081 ( .A1(n5530), .A2(n5529), .ZN(n5548) );
  INV_X1 U7082 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7083 ( .A1(n5531), .A2(SI_22_), .ZN(n5532) );
  NAND2_X1 U7084 ( .A1(n5548), .A2(n5532), .ZN(n5549) );
  NAND2_X1 U7085 ( .A1(n7974), .A2(n8313), .ZN(n5534) );
  NAND2_X1 U7086 ( .A1(n4326), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5533) );
  INV_X1 U7087 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U7088 ( .A1(n5535), .A2(n9271), .ZN(n5536) );
  NAND2_X1 U7089 ( .A1(n5559), .A2(n5536), .ZN(n9538) );
  OR2_X1 U7090 ( .A1(n9538), .A2(n5728), .ZN(n5541) );
  INV_X1 U7091 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U7092 ( .A1(n4322), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7093 ( .A1(n5165), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5537) );
  OAI211_X1 U7094 ( .C1(n5731), .C2(n9537), .A(n5538), .B(n5537), .ZN(n5539)
         );
  INV_X1 U7095 ( .A(n5539), .ZN(n5540) );
  AOI22_X1 U7096 ( .A1(n9540), .A2(n5657), .B1(n5695), .B2(n9324), .ZN(n5542)
         );
  XNOR2_X1 U7097 ( .A(n5542), .B(n5640), .ZN(n5545) );
  INV_X1 U7098 ( .A(n5545), .ZN(n5543) );
  NAND2_X1 U7099 ( .A1(n5544), .A2(n5543), .ZN(n5547) );
  NAND2_X1 U7100 ( .A1(n5546), .A2(n5545), .ZN(n9198) );
  OAI22_X1 U7101 ( .A1(n6597), .A2(n5690), .B1(n9212), .B2(n5697), .ZN(n9268)
         );
  INV_X1 U7102 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5551) );
  MUX2_X1 U7103 ( .A(n8024), .B(n5551), .S(n4936), .Z(n5553) );
  NAND2_X1 U7104 ( .A1(n5553), .A2(n5552), .ZN(n5578) );
  INV_X1 U7105 ( .A(n5553), .ZN(n5554) );
  NAND2_X1 U7106 ( .A1(n5554), .A2(SI_23_), .ZN(n5555) );
  XNOR2_X1 U7107 ( .A(n5577), .B(n5576), .ZN(n5886) );
  NAND2_X1 U7108 ( .A1(n5886), .A2(n8313), .ZN(n5557) );
  NAND2_X1 U7109 ( .A1(n4326), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7110 ( .A1(n6589), .A2(n5657), .ZN(n5567) );
  INV_X1 U7111 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U7112 ( .A1(n5559), .A2(n9204), .ZN(n5560) );
  NAND2_X1 U7113 ( .A1(n5610), .A2(n5560), .ZN(n9524) );
  OR2_X1 U7114 ( .A1(n9524), .A2(n5728), .ZN(n5565) );
  INV_X1 U7115 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9517) );
  NAND2_X1 U7116 ( .A1(n4324), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7117 ( .A1(n5165), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5561) );
  OAI211_X1 U7118 ( .C1(n5731), .C2(n9517), .A(n5562), .B(n5561), .ZN(n5563)
         );
  INV_X1 U7119 ( .A(n5563), .ZN(n5564) );
  OR2_X1 U7120 ( .A1(n9270), .A2(n5690), .ZN(n5566) );
  NAND2_X1 U7121 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  XNOR2_X1 U7122 ( .A(n5568), .B(n5693), .ZN(n5571) );
  NOR2_X1 U7123 ( .A1(n9270), .A2(n5697), .ZN(n5569) );
  AOI21_X1 U7124 ( .B1(n6589), .B2(n5695), .A(n5569), .ZN(n5570) );
  NAND2_X1 U7125 ( .A1(n5571), .A2(n5570), .ZN(n9248) );
  OR2_X1 U7126 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  INV_X1 U7127 ( .A(n9199), .ZN(n5573) );
  OR2_X1 U7128 ( .A1(n9268), .A2(n5573), .ZN(n5574) );
  NAND2_X1 U7129 ( .A1(n5577), .A2(n5576), .ZN(n5579) );
  NAND2_X1 U7130 ( .A1(n5579), .A2(n5578), .ZN(n5601) );
  INV_X1 U7131 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8094) );
  INV_X1 U7132 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5580) );
  MUX2_X1 U7133 ( .A(n8094), .B(n5580), .S(n6631), .Z(n5582) );
  INV_X1 U7134 ( .A(SI_24_), .ZN(n5581) );
  NAND2_X1 U7135 ( .A1(n5582), .A2(n5581), .ZN(n5602) );
  INV_X1 U7136 ( .A(n5582), .ZN(n5583) );
  NAND2_X1 U7137 ( .A1(n5583), .A2(SI_24_), .ZN(n5584) );
  XNOR2_X1 U7138 ( .A(n5601), .B(n5600), .ZN(n8081) );
  NAND2_X1 U7139 ( .A1(n8081), .A2(n8313), .ZN(n5586) );
  NAND2_X1 U7140 ( .A1(n4326), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7141 ( .A1(n6564), .A2(n5657), .ZN(n5593) );
  XNOR2_X1 U7142 ( .A(n5610), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U7143 ( .A1(n9255), .A2(n5140), .ZN(n5591) );
  INV_X1 U7144 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U7145 ( .A1(n5165), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7146 ( .A1(n4322), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5587) );
  OAI211_X1 U7147 ( .C1(n5731), .C2(n9500), .A(n5588), .B(n5587), .ZN(n5589)
         );
  INV_X1 U7148 ( .A(n5589), .ZN(n5590) );
  OR2_X1 U7149 ( .A1(n9221), .A2(n5690), .ZN(n5592) );
  NAND2_X1 U7150 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  XNOR2_X1 U7151 ( .A(n5594), .B(n5693), .ZN(n5597) );
  NOR2_X1 U7152 ( .A1(n9221), .A2(n5697), .ZN(n5595) );
  AOI21_X1 U7153 ( .B1(n6564), .B2(n5695), .A(n5595), .ZN(n5596) );
  NAND2_X1 U7154 ( .A1(n5597), .A2(n5596), .ZN(n5599) );
  OR2_X1 U7155 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  INV_X1 U7156 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8177) );
  INV_X1 U7157 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5603) );
  MUX2_X1 U7158 ( .A(n8177), .B(n5603), .S(n6631), .Z(n5605) );
  INV_X1 U7159 ( .A(SI_25_), .ZN(n5604) );
  NAND2_X1 U7160 ( .A1(n5605), .A2(n5604), .ZN(n5623) );
  INV_X1 U7161 ( .A(n5605), .ZN(n5606) );
  NAND2_X1 U7162 ( .A1(n5606), .A2(SI_25_), .ZN(n5607) );
  XNOR2_X1 U7163 ( .A(n5622), .B(n5621), .ZN(n8174) );
  NAND2_X1 U7164 ( .A1(n8174), .A2(n8313), .ZN(n5609) );
  NAND2_X1 U7165 ( .A1(n4326), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5608) );
  INV_X1 U7166 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9256) );
  INV_X1 U7167 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9224) );
  OAI21_X1 U7168 ( .B1(n5610), .B2(n9256), .A(n9224), .ZN(n5611) );
  AND2_X1 U7169 ( .A1(n5611), .A2(n5631), .ZN(n9223) );
  NAND2_X1 U7170 ( .A1(n9223), .A2(n5140), .ZN(n5616) );
  INV_X1 U7171 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U7172 ( .A1(n4322), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7173 ( .A1(n5165), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5612) );
  OAI211_X1 U7174 ( .C1(n5731), .C2(n9487), .A(n5613), .B(n5612), .ZN(n5614)
         );
  INV_X1 U7175 ( .A(n5614), .ZN(n5615) );
  OAI22_X1 U7176 ( .A1(n9731), .A2(n5690), .B1(n9254), .B2(n5697), .ZN(n5644)
         );
  NAND2_X1 U7177 ( .A1(n9493), .A2(n5657), .ZN(n5618) );
  NAND2_X1 U7178 ( .A1(n9321), .A2(n5695), .ZN(n5617) );
  NAND2_X1 U7179 ( .A1(n5618), .A2(n5617), .ZN(n5620) );
  XNOR2_X1 U7180 ( .A(n5620), .B(n5619), .ZN(n5643) );
  XOR2_X1 U7181 ( .A(n5644), .B(n5643), .Z(n9219) );
  INV_X1 U7182 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8201) );
  INV_X1 U7183 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5624) );
  MUX2_X1 U7184 ( .A(n8201), .B(n5624), .S(n6631), .Z(n5626) );
  INV_X1 U7185 ( .A(SI_26_), .ZN(n5625) );
  NAND2_X1 U7186 ( .A1(n5626), .A2(n5625), .ZN(n5650) );
  INV_X1 U7187 ( .A(n5626), .ZN(n5627) );
  NAND2_X1 U7188 ( .A1(n5627), .A2(SI_26_), .ZN(n5628) );
  NAND2_X1 U7189 ( .A1(n8196), .A2(n8313), .ZN(n5630) );
  NAND2_X1 U7190 ( .A1(n4326), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7191 ( .A1(n9648), .A2(n5657), .ZN(n5639) );
  INV_X1 U7192 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U7193 ( .A1(n5631), .A2(n9298), .ZN(n5632) );
  NAND2_X1 U7194 ( .A1(n5681), .A2(n5632), .ZN(n9466) );
  OR2_X1 U7195 ( .A1(n9466), .A2(n5728), .ZN(n5637) );
  INV_X1 U7196 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U7197 ( .A1(n4322), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7198 ( .A1(n5165), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5633) );
  OAI211_X1 U7199 ( .C1(n5731), .C2(n9465), .A(n5634), .B(n5633), .ZN(n5635)
         );
  INV_X1 U7200 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U7201 ( .A1(n9320), .A2(n5695), .ZN(n5638) );
  NAND2_X1 U7202 ( .A1(n5639), .A2(n5638), .ZN(n5641) );
  XNOR2_X1 U7203 ( .A(n5641), .B(n5640), .ZN(n5669) );
  NOR2_X1 U7204 ( .A1(n9222), .A2(n5697), .ZN(n5642) );
  AOI21_X1 U7205 ( .B1(n9648), .B2(n5695), .A(n5642), .ZN(n5670) );
  XNOR2_X1 U7206 ( .A(n5669), .B(n5670), .ZN(n9293) );
  INV_X1 U7207 ( .A(n5643), .ZN(n5646) );
  INV_X1 U7208 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U7209 ( .A1(n5646), .A2(n5645), .ZN(n9290) );
  INV_X1 U7210 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8498) );
  INV_X1 U7211 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5651) );
  MUX2_X1 U7212 ( .A(n8498), .B(n5651), .S(n4936), .Z(n5652) );
  NAND2_X1 U7213 ( .A1(n5652), .A2(n10185), .ZN(n5677) );
  INV_X1 U7214 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7215 ( .A1(n5653), .A2(SI_27_), .ZN(n5654) );
  NAND2_X1 U7216 ( .A1(n8202), .A2(n8313), .ZN(n5656) );
  NAND2_X1 U7217 ( .A1(n4326), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7218 ( .A1(n9720), .A2(n5657), .ZN(n5662) );
  XNOR2_X1 U7219 ( .A(n5681), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n6411) );
  INV_X1 U7220 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U7221 ( .A1(n5165), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7222 ( .A1(n4324), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5658) );
  OAI211_X1 U7223 ( .C1(n5731), .C2(n9447), .A(n5659), .B(n5658), .ZN(n5660)
         );
  AOI21_X1 U7224 ( .B1(n6411), .B2(n5140), .A(n5660), .ZN(n9295) );
  OR2_X1 U7225 ( .A1(n9295), .A2(n5690), .ZN(n5661) );
  NAND2_X1 U7226 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  XNOR2_X1 U7227 ( .A(n5663), .B(n5693), .ZN(n5666) );
  INV_X1 U7228 ( .A(n5666), .ZN(n5668) );
  NOR2_X1 U7229 ( .A1(n9295), .A2(n5697), .ZN(n5664) );
  AOI21_X1 U7230 ( .B1(n9720), .B2(n5695), .A(n5664), .ZN(n5665) );
  INV_X1 U7231 ( .A(n5665), .ZN(n5667) );
  AOI21_X1 U7232 ( .B1(n5668), .B2(n5667), .A(n5724), .ZN(n6407) );
  INV_X1 U7233 ( .A(n6407), .ZN(n5673) );
  INV_X1 U7234 ( .A(n5669), .ZN(n5671) );
  OR2_X1 U7235 ( .A1(n5671), .A2(n5670), .ZN(n6408) );
  INV_X1 U7236 ( .A(n6408), .ZN(n5672) );
  NOR2_X1 U7237 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  INV_X1 U7238 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8585) );
  INV_X1 U7239 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5678) );
  MUX2_X1 U7240 ( .A(n8585), .B(n5678), .S(n6631), .Z(n5757) );
  XNOR2_X1 U7241 ( .A(n5757), .B(SI_28_), .ZN(n5754) );
  NAND2_X1 U7242 ( .A1(n4326), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7243 ( .A1(n6560), .A2(n5657), .ZN(n5692) );
  INV_X1 U7244 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6412) );
  INV_X1 U7245 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5743) );
  OAI21_X1 U7246 ( .B1(n5681), .B2(n6412), .A(n5743), .ZN(n5684) );
  AND2_X1 U7247 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n5682) );
  NAND2_X1 U7248 ( .A1(n5683), .A2(n5682), .ZN(n9426) );
  NAND2_X1 U7249 ( .A1(n5684), .A2(n9426), .ZN(n8501) );
  OR2_X1 U7250 ( .A1(n8501), .A2(n5728), .ZN(n5689) );
  INV_X1 U7251 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U7252 ( .A1(n5165), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7253 ( .A1(n4322), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5685) );
  OAI211_X1 U7254 ( .C1(n5731), .C2(n8500), .A(n5686), .B(n5685), .ZN(n5687)
         );
  INV_X1 U7255 ( .A(n5687), .ZN(n5688) );
  OR2_X1 U7256 ( .A1(n9420), .A2(n5690), .ZN(n5691) );
  NAND2_X1 U7257 ( .A1(n5692), .A2(n5691), .ZN(n5694) );
  XNOR2_X1 U7258 ( .A(n5694), .B(n5693), .ZN(n5699) );
  NAND2_X1 U7259 ( .A1(n6560), .A2(n5695), .ZN(n5696) );
  OAI21_X1 U7260 ( .B1(n9420), .B2(n5697), .A(n5696), .ZN(n5698) );
  XNOR2_X1 U7261 ( .A(n5699), .B(n5698), .ZN(n5725) );
  INV_X1 U7262 ( .A(n5725), .ZN(n5722) );
  INV_X1 U7263 ( .A(P1_B_REG_SCAN_IN), .ZN(n9407) );
  MUX2_X1 U7264 ( .A(n5701), .B(P1_B_REG_SCAN_IN), .S(n5700), .Z(n5702) );
  OR2_X1 U7265 ( .A1(n5700), .A2(n8197), .ZN(n9779) );
  NOR4_X1 U7266 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5707) );
  NOR4_X1 U7267 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5706) );
  NOR4_X1 U7268 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5705) );
  NOR4_X1 U7269 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5704) );
  AND4_X1 U7270 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n5704), .ZN(n5713)
         );
  NOR2_X1 U7271 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n5711) );
  NOR4_X1 U7272 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5710) );
  NOR4_X1 U7273 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5709) );
  NOR4_X1 U7274 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5708) );
  AND4_X1 U7275 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .ZN(n5712)
         );
  NAND2_X1 U7276 ( .A1(n5713), .A2(n5712), .ZN(n6601) );
  INV_X1 U7277 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5714) );
  NOR2_X1 U7278 ( .A1(n6601), .A2(n5714), .ZN(n5715) );
  OR2_X1 U7279 ( .A1(n9777), .A2(n5715), .ZN(n7270) );
  OR2_X1 U7280 ( .A1(n8197), .A2(n8175), .ZN(n9778) );
  NAND2_X1 U7281 ( .A1(n7270), .A2(n9778), .ZN(n5716) );
  OR2_X1 U7282 ( .A1(n7271), .A2(n5716), .ZN(n5737) );
  NAND2_X1 U7283 ( .A1(n5717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5718) );
  INV_X1 U7284 ( .A(n8389), .ZN(n5720) );
  INV_X1 U7285 ( .A(n5719), .ZN(n8398) );
  NAND2_X1 U7286 ( .A1(n5738), .A2(n9850), .ZN(n9853) );
  AND2_X1 U7287 ( .A1(n5720), .A2(n9853), .ZN(n5721) );
  NAND2_X1 U7288 ( .A1(n5722), .A2(n4917), .ZN(n5723) );
  NAND3_X1 U7289 ( .A1(n5725), .A2(n9307), .A3(n5724), .ZN(n5749) );
  INV_X1 U7290 ( .A(n5744), .ZN(n5726) );
  NOR2_X2 U7291 ( .A1(n5726), .A2(n5738), .ZN(n9301) );
  INV_X1 U7292 ( .A(n5727), .ZN(n8206) );
  OR2_X1 U7293 ( .A1(n9295), .A2(n9281), .ZN(n5736) );
  OR2_X1 U7294 ( .A1(n9426), .A2(n5728), .ZN(n5734) );
  INV_X1 U7295 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U7296 ( .A1(n4324), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U7297 ( .A1(n5165), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5729) );
  OAI211_X1 U7298 ( .C1(n5731), .C2(n9425), .A(n5730), .B(n5729), .ZN(n5732)
         );
  INV_X1 U7299 ( .A(n5732), .ZN(n5733) );
  INV_X1 U7300 ( .A(n8309), .ZN(n9319) );
  NAND2_X1 U7301 ( .A1(n8389), .A2(n5727), .ZN(n9409) );
  NAND2_X1 U7302 ( .A1(n9319), .A2(n9244), .ZN(n5735) );
  NAND2_X1 U7303 ( .A1(n5736), .A2(n5735), .ZN(n6594) );
  INV_X1 U7304 ( .A(n9850), .ZN(n6561) );
  NOR2_X1 U7305 ( .A1(n6561), .A2(n8394), .ZN(n7274) );
  OAI21_X1 U7306 ( .B1(n7274), .B2(n9853), .A(n5737), .ZN(n5741) );
  NOR2_X1 U7307 ( .A1(n5128), .A2(n6618), .ZN(n5740) );
  NAND2_X1 U7308 ( .A1(n8389), .A2(n5738), .ZN(n5739) );
  AND2_X1 U7309 ( .A1(n5740), .A2(n5739), .ZN(n6599) );
  NAND2_X1 U7310 ( .A1(n5741), .A2(n6599), .ZN(n5742) );
  OAI22_X1 U7311 ( .A1(n8501), .A2(n9299), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5743), .ZN(n5747) );
  NAND2_X1 U7312 ( .A1(n5744), .A2(n7274), .ZN(n5745) );
  NAND2_X1 U7313 ( .A1(n8458), .A2(n8394), .ZN(n9706) );
  NOR2_X1 U7314 ( .A1(n6559), .A2(n9317), .ZN(n5746) );
  AOI211_X1 U7315 ( .C1(n9301), .C2(n6594), .A(n5747), .B(n5746), .ZN(n5748)
         );
  NAND2_X1 U7316 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U7317 ( .A1(n5753), .A2(n5752), .ZN(P1_U3220) );
  INV_X1 U7318 ( .A(SI_28_), .ZN(n5756) );
  INV_X1 U7319 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9183) );
  INV_X1 U7320 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5758) );
  MUX2_X1 U7321 ( .A(n9183), .B(n5758), .S(n6631), .Z(n5759) );
  INV_X1 U7322 ( .A(SI_29_), .ZN(n5760) );
  INV_X1 U7323 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10044) );
  INV_X1 U7324 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n5761) );
  MUX2_X1 U7325 ( .A(n10044), .B(n5761), .S(n6631), .Z(n5763) );
  INV_X1 U7326 ( .A(SI_30_), .ZN(n5762) );
  NAND2_X1 U7327 ( .A1(n5763), .A2(n5762), .ZN(n6273) );
  INV_X1 U7328 ( .A(n5763), .ZN(n5764) );
  NAND2_X1 U7329 ( .A1(n5764), .A2(SI_30_), .ZN(n5765) );
  NAND2_X1 U7330 ( .A1(n6273), .A2(n5765), .ZN(n6274) );
  NOR2_X1 U7331 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5772) );
  NAND4_X1 U7332 ( .A1(n5772), .A2(n5899), .A3(n10173), .A4(n5771), .ZN(n5773)
         );
  NAND2_X1 U7333 ( .A1(n6393), .A2(n6396), .ZN(n6398) );
  INV_X1 U7334 ( .A(n6398), .ZN(n5778) );
  NOR2_X1 U7335 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5777) );
  XNOR2_X2 U7336 ( .A(n5781), .B(n5816), .ZN(n6403) );
  NAND3_X1 U7337 ( .A1(n6392), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n5790) );
  XNOR2_X1 U7338 ( .A(n9177), .B(P2_IR_REG_27__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7339 ( .A1(n6401), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5784) );
  NOR2_X1 U7340 ( .A1(n6398), .A2(n5784), .ZN(n5785) );
  NAND2_X2 U7341 ( .A1(n6403), .A2(n6404), .ZN(n5966) );
  NAND2_X1 U7342 ( .A1(n8588), .A2(n6229), .ZN(n5791) );
  NAND2_X2 U7343 ( .A1(n5966), .A2(n6631), .ZN(n6004) );
  INV_X1 U7344 ( .A(n5843), .ZN(n6380) );
  NAND2_X1 U7345 ( .A1(n10068), .A2(n7389), .ZN(n6027) );
  INV_X1 U7346 ( .A(n6027), .ZN(n5793) );
  NAND2_X1 U7347 ( .A1(n5793), .A2(n5792), .ZN(n6029) );
  INV_X1 U7348 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5805) );
  INV_X1 U7349 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5807) );
  INV_X1 U7350 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5809) );
  INV_X1 U7351 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5811) );
  INV_X1 U7352 ( .A(n6234), .ZN(n5813) );
  INV_X1 U7353 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10160) );
  INV_X1 U7354 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5814) );
  XNOR2_X2 U7355 ( .A(n5819), .B(n5818), .ZN(n8589) );
  XNOR2_X2 U7356 ( .A(n5822), .B(n5821), .ZN(n9184) );
  NAND2_X1 U7357 ( .A1(n8512), .A2(n6235), .ZN(n6288) );
  INV_X1 U7358 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7359 ( .A1(n6282), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7360 ( .A1(n8589), .A2(n5823), .ZN(n5982) );
  NAND2_X1 U7361 ( .A1(n6237), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5824) );
  OAI211_X1 U7362 ( .C1(n5826), .C2(n6186), .A(n5825), .B(n5824), .ZN(n5827)
         );
  INV_X1 U7363 ( .A(n5827), .ZN(n5828) );
  NAND2_X1 U7364 ( .A1(n6288), .A2(n5828), .ZN(n8740) );
  NAND2_X1 U7365 ( .A1(n6380), .A2(n8740), .ZN(n6271) );
  NAND2_X1 U7366 ( .A1(n9182), .A2(n6229), .ZN(n5831) );
  OR2_X1 U7367 ( .A1(n6004), .A2(n9183), .ZN(n5830) );
  NAND2_X1 U7368 ( .A1(n5831), .A2(n5830), .ZN(n5845) );
  INV_X1 U7369 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U7370 ( .A1(n6237), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7371 ( .A1(n6282), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5832) );
  OAI211_X1 U7372 ( .C1(n6186), .C2(n8527), .A(n5833), .B(n5832), .ZN(n5834)
         );
  INV_X1 U7373 ( .A(n5834), .ZN(n5835) );
  INV_X1 U7374 ( .A(n5836), .ZN(n5837) );
  NAND2_X1 U7375 ( .A1(n5837), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5838) );
  MUX2_X1 U7376 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5838), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5840) );
  NAND2_X1 U7377 ( .A1(n6295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5842) );
  INV_X1 U7378 ( .A(n8740), .ZN(n5844) );
  NAND2_X1 U7379 ( .A1(n5843), .A2(n5844), .ZN(n6272) );
  NAND2_X1 U7380 ( .A1(n5845), .A2(n8741), .ZN(n5849) );
  NAND2_X1 U7381 ( .A1(n6272), .A2(n5849), .ZN(n6382) );
  NAND2_X1 U7382 ( .A1(n8202), .A2(n6229), .ZN(n5851) );
  INV_X1 U7383 ( .A(n5852), .ZN(n5853) );
  NAND2_X1 U7384 ( .A1(n5853), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7385 ( .A1(n5860), .A2(n5854), .ZN(n8908) );
  NAND2_X1 U7386 ( .A1(n8908), .A2(n6235), .ZN(n5859) );
  INV_X1 U7387 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U7388 ( .A1(n6282), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7389 ( .A1(n6237), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5855) );
  OAI211_X1 U7390 ( .C1(n8907), .C2(n6186), .A(n5856), .B(n5855), .ZN(n5857)
         );
  INV_X1 U7391 ( .A(n5857), .ZN(n5858) );
  NAND2_X1 U7392 ( .A1(n5860), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7393 ( .A1(n5862), .A2(n5861), .ZN(n8889) );
  NAND2_X1 U7394 ( .A1(n8889), .A2(n6235), .ZN(n5867) );
  INV_X1 U7395 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U7396 ( .A1(n6237), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7397 ( .A1(n6282), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5863) );
  OAI211_X1 U7398 ( .C1(n8890), .C2(n6186), .A(n5864), .B(n5863), .ZN(n5865)
         );
  INV_X1 U7399 ( .A(n5865), .ZN(n5866) );
  NAND2_X1 U7400 ( .A1(n6376), .A2(n8904), .ZN(n5870) );
  NAND2_X1 U7401 ( .A1(n8205), .A2(n6229), .ZN(n5869) );
  OR2_X1 U7402 ( .A1(n6004), .A2(n8585), .ZN(n5868) );
  INV_X1 U7403 ( .A(n9062), .ZN(n6466) );
  MUX2_X1 U7404 ( .A(n5870), .B(n6466), .S(n5846), .Z(n6258) );
  NAND2_X1 U7405 ( .A1(n8196), .A2(n6229), .ZN(n5872) );
  OR2_X1 U7406 ( .A1(n6004), .A2(n8201), .ZN(n5871) );
  NAND2_X1 U7407 ( .A1(n8917), .A2(n6235), .ZN(n5877) );
  INV_X1 U7408 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U7409 ( .A1(n6237), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7410 ( .A1(n6282), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5873) );
  OAI211_X1 U7411 ( .C1(n8916), .C2(n6186), .A(n5874), .B(n5873), .ZN(n5875)
         );
  INV_X1 U7412 ( .A(n5875), .ZN(n5876) );
  NAND2_X2 U7413 ( .A1(n5877), .A2(n5876), .ZN(n8924) );
  NAND2_X1 U7414 ( .A1(n7974), .A2(n6229), .ZN(n5879) );
  OR2_X1 U7415 ( .A1(n6004), .A2(n8018), .ZN(n5878) );
  XNOR2_X1 U7416 ( .A(n6209), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U7417 ( .A1(n8961), .A2(n6235), .ZN(n5885) );
  INV_X1 U7418 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7419 ( .A1(n6237), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7420 ( .A1(n6282), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5880) );
  OAI211_X1 U7421 ( .C1(n5882), .C2(n6186), .A(n5881), .B(n5880), .ZN(n5883)
         );
  INV_X1 U7422 ( .A(n5883), .ZN(n5884) );
  NAND2_X1 U7423 ( .A1(n5886), .A2(n6229), .ZN(n5888) );
  OR2_X1 U7424 ( .A1(n6004), .A2(n8024), .ZN(n5887) );
  NAND2_X1 U7425 ( .A1(n5889), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7426 ( .A1(n6220), .A2(n5890), .ZN(n8949) );
  NAND2_X1 U7427 ( .A1(n8949), .A2(n6235), .ZN(n5895) );
  INV_X1 U7428 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U7429 ( .A1(n6282), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7430 ( .A1(n6237), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5891) );
  OAI211_X1 U7431 ( .C1(n8948), .C2(n6186), .A(n5892), .B(n5891), .ZN(n5893)
         );
  INV_X1 U7432 ( .A(n5893), .ZN(n5894) );
  NAND2_X1 U7433 ( .A1(n8950), .A2(n8958), .ZN(n6368) );
  NAND2_X1 U7434 ( .A1(n6457), .A2(n8968), .ZN(n6364) );
  AND2_X1 U7435 ( .A1(n6368), .A2(n6364), .ZN(n5896) );
  MUX2_X1 U7436 ( .A(n6365), .B(n5896), .S(n5846), .Z(n6217) );
  NAND2_X1 U7437 ( .A1(n7232), .A2(n6229), .ZN(n5902) );
  NAND2_X1 U7438 ( .A1(n5908), .A2(n5899), .ZN(n6158) );
  NAND2_X1 U7439 ( .A1(n6158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U7440 ( .A(n5900), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8846) );
  AOI22_X1 U7441 ( .A1(n6180), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6880), .B2(
        n8846), .ZN(n5901) );
  NAND2_X1 U7442 ( .A1(n6282), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5907) );
  INV_X1 U7443 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8819) );
  OR2_X1 U7444 ( .A1(n6185), .A2(n8819), .ZN(n5906) );
  NAND2_X1 U7445 ( .A1(n5913), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5903) );
  AND2_X1 U7446 ( .A1(n6166), .A2(n5903), .ZN(n9031) );
  OR2_X1 U7447 ( .A1(n6141), .A2(n9031), .ZN(n5905) );
  INV_X1 U7448 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9032) );
  OR2_X1 U7449 ( .A1(n6186), .A2(n9032), .ZN(n5904) );
  OR2_X1 U7450 ( .A1(n9100), .A2(n9009), .ZN(n6172) );
  NAND2_X1 U7451 ( .A1(n9100), .A2(n9009), .ZN(n6355) );
  NAND2_X1 U7452 ( .A1(n6172), .A2(n6355), .ZN(n6449) );
  NAND2_X1 U7453 ( .A1(n7188), .A2(n6229), .ZN(n5911) );
  OR2_X1 U7454 ( .A1(n5908), .A2(n9177), .ZN(n5909) );
  XNOR2_X1 U7455 ( .A(n5909), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8806) );
  AOI22_X1 U7456 ( .A1(n6180), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6880), .B2(
        n8806), .ZN(n5910) );
  NAND2_X1 U7457 ( .A1(n6282), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5917) );
  INV_X1 U7458 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9104) );
  OR2_X1 U7459 ( .A1(n5982), .A2(n9104), .ZN(n5916) );
  NAND2_X1 U7460 ( .A1(n5939), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5912) );
  AND2_X1 U7461 ( .A1(n5913), .A2(n5912), .ZN(n9049) );
  OR2_X1 U7462 ( .A1(n6141), .A2(n9049), .ZN(n5915) );
  INV_X1 U7463 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9048) );
  OR2_X1 U7464 ( .A1(n6186), .A2(n9048), .ZN(n5914) );
  INV_X1 U7465 ( .A(n6301), .ZN(n6353) );
  NAND2_X1 U7466 ( .A1(n7038), .A2(n6229), .ZN(n5927) );
  NOR2_X1 U7467 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5918) );
  INV_X1 U7468 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7469 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6134) );
  INV_X1 U7470 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7471 ( .A1(n6134), .A2(n5921), .ZN(n5922) );
  NAND2_X1 U7472 ( .A1(n5922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5928) );
  INV_X1 U7473 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7474 ( .A1(n5928), .A2(n5923), .ZN(n5924) );
  NAND2_X1 U7475 ( .A1(n5924), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5925) );
  XNOR2_X1 U7476 ( .A(n5925), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8798) );
  AOI22_X1 U7477 ( .A1(n8798), .A2(n6880), .B1(n6180), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7478 ( .A1(n6816), .A2(n6229), .ZN(n5930) );
  XNOR2_X1 U7479 ( .A(n5928), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8139) );
  AOI22_X1 U7480 ( .A1(n6180), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6880), .B2(
        n8139), .ZN(n5929) );
  NAND2_X1 U7481 ( .A1(n6282), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5936) );
  INV_X1 U7482 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8156) );
  OR2_X1 U7483 ( .A1(n5982), .A2(n8156), .ZN(n5935) );
  NAND2_X1 U7484 ( .A1(n6140), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5931) );
  AND2_X1 U7485 ( .A1(n5937), .A2(n5931), .ZN(n8607) );
  OR2_X1 U7486 ( .A1(n6141), .A2(n8607), .ZN(n5934) );
  INV_X1 U7487 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5932) );
  OR2_X1 U7488 ( .A1(n6186), .A2(n5932), .ZN(n5933) );
  NAND4_X1 U7489 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n8746)
         );
  INV_X1 U7490 ( .A(n8746), .ZN(n8539) );
  NAND3_X1 U7491 ( .A1(n8537), .A2(n8539), .A3(n5846), .ZN(n5944) );
  NAND2_X1 U7492 ( .A1(n6282), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5943) );
  INV_X1 U7493 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8767) );
  OR2_X1 U7494 ( .A1(n6185), .A2(n8767), .ZN(n5942) );
  NAND2_X1 U7495 ( .A1(n5937), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5938) );
  AND2_X1 U7496 ( .A1(n5939), .A2(n5938), .ZN(n8192) );
  OR2_X1 U7497 ( .A1(n6141), .A2(n8192), .ZN(n5941) );
  INV_X1 U7498 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8191) );
  OR2_X1 U7499 ( .A1(n6186), .A2(n8191), .ZN(n5940) );
  NAND2_X1 U7500 ( .A1(n8606), .A2(n5846), .ZN(n5945) );
  NAND2_X1 U7501 ( .A1(n5944), .A2(n5945), .ZN(n5947) );
  NOR2_X1 U7502 ( .A1(n5945), .A2(n8746), .ZN(n5946) );
  AOI22_X1 U7503 ( .A1(n8542), .A2(n5947), .B1(n5946), .B2(n8537), .ZN(n6156)
         );
  NAND2_X1 U7504 ( .A1(n6237), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5953) );
  INV_X1 U7505 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5948) );
  OR2_X1 U7506 ( .A1(n6240), .A2(n5948), .ZN(n5952) );
  NAND2_X1 U7507 ( .A1(n6029), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5949) );
  AND2_X1 U7508 ( .A1(n6066), .A2(n5949), .ZN(n7225) );
  OR2_X1 U7509 ( .A1(n6141), .A2(n7225), .ZN(n5951) );
  INV_X1 U7510 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7419) );
  OR2_X1 U7511 ( .A1(n6186), .A2(n7419), .ZN(n5950) );
  OR2_X1 U7512 ( .A1(n6647), .A2(n6133), .ZN(n5958) );
  NAND2_X1 U7513 ( .A1(n5897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5954) );
  MUX2_X1 U7514 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5954), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5955) );
  NAND2_X1 U7515 ( .A1(n5955), .A2(n6073), .ZN(n7453) );
  OR2_X1 U7516 ( .A1(n6614), .A2(n7453), .ZN(n5957) );
  INV_X1 U7517 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6646) );
  OR2_X1 U7518 ( .A1(n6004), .A2(n6646), .ZN(n5956) );
  INV_X1 U7519 ( .A(n9951), .ZN(n7421) );
  NAND2_X1 U7520 ( .A1(n7429), .A2(n7421), .ZN(n6336) );
  INV_X1 U7521 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7522 ( .A1(n5982), .A2(n5959), .ZN(n5963) );
  INV_X1 U7523 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U7524 ( .A1(n5980), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5961) );
  INV_X1 U7525 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9888) );
  OR2_X1 U7526 ( .A1(n5996), .A2(n9888), .ZN(n5960) );
  AND4_X2 U7527 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n7254)
         );
  OR2_X1 U7528 ( .A1(n6004), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5968) );
  OR2_X1 U7529 ( .A1(n6133), .A2(n5964), .ZN(n5969) );
  OR2_X1 U7530 ( .A1(n5966), .A2(n6897), .ZN(n5967) );
  NAND3_X1 U7531 ( .A1(n5968), .A2(n5969), .A3(n5967), .ZN(n9920) );
  INV_X1 U7532 ( .A(n6186), .ZN(n6236) );
  NAND2_X1 U7533 ( .A1(n6236), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5974) );
  INV_X1 U7534 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5970) );
  INV_X1 U7535 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10057) );
  OR2_X1 U7536 ( .A1(n5982), .A2(n10057), .ZN(n5972) );
  INV_X1 U7537 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6845) );
  OR2_X1 U7538 ( .A1(n5996), .A2(n6845), .ZN(n5971) );
  NAND2_X1 U7539 ( .A1(n6632), .A2(SI_0_), .ZN(n5975) );
  XNOR2_X1 U7540 ( .A(n5975), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9185) );
  INV_X1 U7541 ( .A(n7051), .ZN(n6980) );
  NAND2_X1 U7542 ( .A1(n8760), .A2(n6980), .ZN(n6302) );
  NAND2_X1 U7543 ( .A1(n6302), .A2(n6508), .ZN(n5994) );
  NAND2_X1 U7544 ( .A1(n6302), .A2(n7044), .ZN(n5976) );
  NAND2_X1 U7545 ( .A1(n7050), .A2(n5976), .ZN(n5977) );
  NAND2_X1 U7546 ( .A1(n5977), .A2(n6421), .ZN(n5978) );
  NAND2_X1 U7547 ( .A1(n5978), .A2(n6420), .ZN(n5979) );
  MUX2_X1 U7548 ( .A(n5979), .B(n6420), .S(n6508), .Z(n5993) );
  NAND2_X1 U7549 ( .A1(n6282), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5986) );
  INV_X1 U7550 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5981) );
  OR2_X1 U7551 ( .A1(n5982), .A2(n5981), .ZN(n5985) );
  INV_X1 U7552 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7079) );
  OR2_X1 U7553 ( .A1(n5996), .A2(n7079), .ZN(n5984) );
  INV_X1 U7554 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7261) );
  OR2_X1 U7555 ( .A1(n6186), .A2(n7261), .ZN(n5983) );
  OR2_X1 U7556 ( .A1(n6004), .A2(n4925), .ZN(n5992) );
  OR2_X1 U7557 ( .A1(n6133), .A2(n6642), .ZN(n5991) );
  OR2_X1 U7558 ( .A1(n6614), .A2(n7026), .ZN(n5990) );
  OAI211_X1 U7559 ( .C1(n7265), .C2(n5994), .A(n5993), .B(n4321), .ZN(n6012)
         );
  NAND2_X1 U7560 ( .A1(n6282), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6001) );
  INV_X1 U7561 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5995) );
  OR2_X1 U7562 ( .A1(n6141), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5999) );
  INV_X1 U7563 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5997) );
  OR2_X1 U7564 ( .A1(n6186), .A2(n5997), .ZN(n5998) );
  XNOR2_X1 U7565 ( .A(n6003), .B(n5766), .ZN(n7098) );
  INV_X1 U7566 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6633) );
  OR2_X1 U7567 ( .A1(n6004), .A2(n6633), .ZN(n6006) );
  OR2_X1 U7568 ( .A1(n6133), .A2(n6640), .ZN(n6005) );
  OAI211_X1 U7569 ( .C1(n6614), .C2(n7098), .A(n6006), .B(n6005), .ZN(n7390)
         );
  NAND2_X1 U7570 ( .A1(n8757), .A2(n9934), .ZN(n6304) );
  NAND2_X1 U7571 ( .A1(n8758), .A2(n9926), .ZN(n6007) );
  NAND2_X1 U7572 ( .A1(n6304), .A2(n6007), .ZN(n6009) );
  NAND2_X1 U7573 ( .A1(n7253), .A2(n7390), .ZN(n6329) );
  INV_X1 U7574 ( .A(n8758), .ZN(n6423) );
  INV_X1 U7575 ( .A(n9926), .ZN(n7258) );
  NAND2_X1 U7576 ( .A1(n6423), .A2(n7258), .ZN(n6328) );
  NAND2_X1 U7577 ( .A1(n6329), .A2(n6328), .ZN(n6008) );
  MUX2_X1 U7578 ( .A(n6009), .B(n6008), .S(n5846), .Z(n6010) );
  INV_X1 U7579 ( .A(n6010), .ZN(n6011) );
  NAND2_X1 U7580 ( .A1(n6012), .A2(n6011), .ZN(n6025) );
  NAND2_X1 U7581 ( .A1(n6282), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6018) );
  INV_X1 U7582 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7583 ( .A1(n5982), .A2(n6013), .ZN(n6017) );
  NAND2_X1 U7584 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6014) );
  AND2_X1 U7585 ( .A1(n6027), .A2(n6014), .ZN(n7241) );
  OR2_X1 U7586 ( .A1(n5996), .A2(n7241), .ZN(n6016) );
  INV_X1 U7587 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7240) );
  OR2_X1 U7588 ( .A1(n6186), .A2(n7240), .ZN(n6015) );
  NAND2_X1 U7589 ( .A1(n6019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6020) );
  XNOR2_X1 U7590 ( .A(n6020), .B(n4853), .ZN(n7136) );
  OR2_X1 U7591 ( .A1(n6004), .A2(n4938), .ZN(n6022) );
  OR2_X1 U7592 ( .A1(n6133), .A2(n6635), .ZN(n6021) );
  OAI211_X1 U7593 ( .C1(n6614), .C2(n7136), .A(n6022), .B(n6021), .ZN(n7243)
         );
  NAND2_X1 U7594 ( .A1(n8756), .A2(n9940), .ZN(n6331) );
  INV_X1 U7595 ( .A(n6331), .ZN(n6023) );
  NOR2_X1 U7596 ( .A1(n8756), .A2(n9940), .ZN(n6332) );
  OR2_X1 U7597 ( .A1(n6023), .A2(n6332), .ZN(n7237) );
  INV_X1 U7598 ( .A(n7237), .ZN(n6024) );
  NAND2_X1 U7599 ( .A1(n6025), .A2(n6024), .ZN(n6046) );
  NAND2_X1 U7600 ( .A1(n6236), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6034) );
  INV_X1 U7601 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6026) );
  OR2_X1 U7602 ( .A1(n6185), .A2(n6026), .ZN(n6033) );
  NAND2_X1 U7603 ( .A1(n6027), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6028) );
  AND2_X1 U7604 ( .A1(n6029), .A2(n6028), .ZN(n7181) );
  OR2_X1 U7605 ( .A1(n6141), .A2(n7181), .ZN(n6032) );
  INV_X1 U7606 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6030) );
  OR2_X1 U7607 ( .A1(n6240), .A2(n6030), .ZN(n6031) );
  OR2_X1 U7608 ( .A1(n6035), .A2(n9177), .ZN(n6037) );
  XNOR2_X1 U7609 ( .A(n6037), .B(n6036), .ZN(n7155) );
  OR2_X1 U7610 ( .A1(n6133), .A2(n6649), .ZN(n6039) );
  INV_X1 U7611 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6648) );
  OR2_X1 U7612 ( .A1(n6004), .A2(n6648), .ZN(n6038) );
  OAI211_X1 U7613 ( .C1(n6614), .C2(n7155), .A(n6039), .B(n6038), .ZN(n7289)
         );
  INV_X1 U7614 ( .A(n7289), .ZN(n9946) );
  NAND2_X1 U7615 ( .A1(n8755), .A2(n9946), .ZN(n6333) );
  OAI211_X1 U7616 ( .C1(n6046), .C2(n4850), .A(n6333), .B(n6331), .ZN(n6042)
         );
  NAND2_X1 U7617 ( .A1(n7219), .A2(n7289), .ZN(n6334) );
  AND2_X1 U7618 ( .A1(n6336), .A2(n6334), .ZN(n6041) );
  NAND2_X1 U7619 ( .A1(n8754), .A2(n9951), .ZN(n6306) );
  INV_X1 U7620 ( .A(n6306), .ZN(n6040) );
  AOI21_X1 U7621 ( .B1(n6042), .B2(n6041), .A(n6040), .ZN(n6043) );
  MUX2_X1 U7622 ( .A(n6336), .B(n6043), .S(n6508), .Z(n6080) );
  INV_X1 U7623 ( .A(n6304), .ZN(n6045) );
  INV_X1 U7624 ( .A(n6332), .ZN(n6044) );
  OAI211_X1 U7625 ( .C1(n6046), .C2(n6045), .A(n6334), .B(n6044), .ZN(n6047)
         );
  NAND4_X1 U7626 ( .A1(n6047), .A2(n5846), .A3(n6333), .A4(n6306), .ZN(n6078)
         );
  NAND2_X1 U7627 ( .A1(n6650), .A2(n6229), .ZN(n6050) );
  NAND2_X1 U7628 ( .A1(n6075), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6048) );
  AOI22_X1 U7629 ( .A1(n6180), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6880), .B2(
        n9903), .ZN(n6049) );
  NAND2_X1 U7630 ( .A1(n6050), .A2(n6049), .ZN(n9964) );
  NAND2_X1 U7631 ( .A1(n6282), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6055) );
  INV_X1 U7632 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7594) );
  OR2_X1 U7633 ( .A1(n6185), .A2(n7594), .ZN(n6054) );
  NAND2_X1 U7634 ( .A1(n6068), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6051) );
  AND2_X1 U7635 ( .A1(n6059), .A2(n6051), .ZN(n7762) );
  OR2_X1 U7636 ( .A1(n6141), .A2(n7762), .ZN(n6053) );
  INV_X1 U7637 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7595) );
  OR2_X1 U7638 ( .A1(n6186), .A2(n7595), .ZN(n6052) );
  NAND2_X1 U7639 ( .A1(n9964), .A2(n7828), .ZN(n6339) );
  NAND2_X1 U7640 ( .A1(n6654), .A2(n6229), .ZN(n6058) );
  OR2_X1 U7641 ( .A1(n6056), .A2(n9177), .ZN(n6082) );
  XNOR2_X1 U7642 ( .A(n6082), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7718) );
  AOI22_X1 U7643 ( .A1(n6180), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6880), .B2(
        n7718), .ZN(n6057) );
  NAND2_X1 U7644 ( .A1(n6282), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6064) );
  INV_X1 U7645 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7601) );
  OR2_X1 U7646 ( .A1(n6185), .A2(n7601), .ZN(n6063) );
  NAND2_X1 U7647 ( .A1(n6059), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6060) );
  AND2_X1 U7648 ( .A1(n6087), .A2(n6060), .ZN(n7841) );
  OR2_X1 U7649 ( .A1(n6141), .A2(n7841), .ZN(n6062) );
  INV_X1 U7650 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7710) );
  OR2_X1 U7651 ( .A1(n6186), .A2(n7710), .ZN(n6061) );
  NAND4_X1 U7652 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n8751)
         );
  INV_X1 U7653 ( .A(n8751), .ZN(n7555) );
  OR2_X1 U7654 ( .A1(n9964), .A2(n7828), .ZN(n6309) );
  NAND2_X1 U7655 ( .A1(n9969), .A2(n7555), .ZN(n6308) );
  AND2_X1 U7656 ( .A1(n6065), .A2(n6308), .ZN(n6110) );
  INV_X1 U7657 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7460) );
  OR2_X1 U7658 ( .A1(n6186), .A2(n7460), .ZN(n6072) );
  NAND2_X1 U7659 ( .A1(n6066), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6067) );
  AND2_X1 U7660 ( .A1(n6068), .A2(n6067), .ZN(n7434) );
  OR2_X1 U7661 ( .A1(n6141), .A2(n7434), .ZN(n6071) );
  INV_X1 U7662 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6069) );
  OR2_X1 U7663 ( .A1(n6240), .A2(n6069), .ZN(n6070) );
  NAND2_X1 U7664 ( .A1(n6073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6074) );
  MUX2_X1 U7665 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6074), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6076) );
  AOI22_X1 U7666 ( .A1(n6180), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6880), .B2(
        n7598), .ZN(n6077) );
  NAND2_X1 U7667 ( .A1(n7758), .A2(n7436), .ZN(n6093) );
  NAND2_X1 U7668 ( .A1(n6093), .A2(n7559), .ZN(n7424) );
  INV_X1 U7669 ( .A(n7424), .ZN(n7427) );
  AND3_X1 U7670 ( .A1(n6078), .A2(n6110), .A3(n7427), .ZN(n6079) );
  OR2_X1 U7671 ( .A1(n6660), .A2(n6133), .ZN(n6086) );
  INV_X1 U7672 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7673 ( .A1(n6082), .A2(n6081), .ZN(n6083) );
  NAND2_X1 U7674 ( .A1(n6083), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7675 ( .A(n6084), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7731) );
  AOI22_X1 U7676 ( .A1(n6180), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6880), .B2(
        n7731), .ZN(n6085) );
  NAND2_X1 U7677 ( .A1(n6282), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6092) );
  INV_X1 U7678 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7729) );
  OR2_X1 U7679 ( .A1(n6185), .A2(n7729), .ZN(n6091) );
  INV_X1 U7680 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7730) );
  OR2_X1 U7681 ( .A1(n6186), .A2(n7730), .ZN(n6090) );
  NAND2_X1 U7682 ( .A1(n6087), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6088) );
  AND2_X1 U7683 ( .A1(n6103), .A2(n6088), .ZN(n7858) );
  OR2_X1 U7684 ( .A1(n6141), .A2(n7858), .ZN(n6089) );
  NAND4_X1 U7685 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n8750)
         );
  NAND2_X1 U7686 ( .A1(n9975), .A2(n7900), .ZN(n7892) );
  NAND2_X1 U7687 ( .A1(n6339), .A2(n6093), .ZN(n6094) );
  NAND2_X1 U7688 ( .A1(n6110), .A2(n6094), .ZN(n6095) );
  OR2_X1 U7689 ( .A1(n9975), .A2(n7900), .ZN(n6342) );
  NAND2_X1 U7690 ( .A1(n6720), .A2(n6229), .ZN(n6101) );
  NOR2_X1 U7691 ( .A1(n6096), .A2(n9177), .ZN(n6097) );
  MUX2_X1 U7692 ( .A(n9177), .B(n6097), .S(P2_IR_REG_11__SCAN_IN), .Z(n6098)
         );
  INV_X1 U7693 ( .A(n6098), .ZN(n6099) );
  AOI22_X1 U7694 ( .A1(n6180), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6880), .B2(
        n7946), .ZN(n6100) );
  NAND2_X1 U7695 ( .A1(n6101), .A2(n6100), .ZN(n9980) );
  NAND2_X1 U7696 ( .A1(n6282), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6108) );
  INV_X1 U7697 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6102) );
  OR2_X1 U7698 ( .A1(n5982), .A2(n6102), .ZN(n6107) );
  INV_X1 U7699 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7901) );
  OR2_X1 U7700 ( .A1(n6186), .A2(n7901), .ZN(n6106) );
  NAND2_X1 U7701 ( .A1(n6103), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6104) );
  AND2_X1 U7702 ( .A1(n6122), .A2(n6104), .ZN(n7966) );
  OR2_X1 U7703 ( .A1(n6141), .A2(n7966), .ZN(n6105) );
  NAND4_X1 U7704 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n8749)
         );
  INV_X1 U7705 ( .A(n8749), .ZN(n8038) );
  OR2_X1 U7706 ( .A1(n9980), .A2(n8038), .ZN(n6344) );
  NAND2_X1 U7707 ( .A1(n9980), .A2(n8038), .ZN(n6112) );
  NAND2_X1 U7708 ( .A1(n6109), .A2(n6112), .ZN(n6117) );
  INV_X1 U7709 ( .A(n6110), .ZN(n6111) );
  AND2_X1 U7710 ( .A1(n6309), .A2(n7559), .ZN(n6338) );
  OAI211_X1 U7711 ( .C1(n6111), .C2(n6338), .A(n6342), .B(n6340), .ZN(n6113)
         );
  AND2_X1 U7712 ( .A1(n6112), .A2(n7892), .ZN(n6343) );
  OAI21_X1 U7713 ( .B1(n6114), .B2(n6113), .A(n6343), .ZN(n6115) );
  NAND2_X1 U7714 ( .A1(n6115), .A2(n6344), .ZN(n6116) );
  MUX2_X1 U7715 ( .A(n6117), .B(n6116), .S(n5846), .Z(n6128) );
  OR2_X1 U7716 ( .A1(n6769), .A2(n6133), .ZN(n6121) );
  NAND2_X1 U7717 ( .A1(n6118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6119) );
  XNOR2_X1 U7718 ( .A(n6119), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8053) );
  AOI22_X1 U7719 ( .A1(n6180), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6880), .B2(
        n8053), .ZN(n6120) );
  NAND2_X1 U7720 ( .A1(n6282), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6127) );
  INV_X1 U7721 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7947) );
  OR2_X1 U7722 ( .A1(n6185), .A2(n7947), .ZN(n6126) );
  NAND2_X1 U7723 ( .A1(n6122), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6123) );
  AND2_X1 U7724 ( .A1(n6138), .A2(n6123), .ZN(n8045) );
  OR2_X1 U7725 ( .A1(n6141), .A2(n8045), .ZN(n6125) );
  INV_X1 U7726 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7948) );
  OR2_X1 U7727 ( .A1(n6186), .A2(n7948), .ZN(n6124) );
  NAND4_X1 U7728 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n8748)
         );
  XNOR2_X1 U7729 ( .A(n9986), .B(n8748), .ZN(n7981) );
  NAND2_X1 U7730 ( .A1(n6128), .A2(n7981), .ZN(n6132) );
  OR2_X1 U7731 ( .A1(n9986), .A2(n6508), .ZN(n6130) );
  NAND2_X1 U7732 ( .A1(n9986), .A2(n6508), .ZN(n6129) );
  INV_X1 U7733 ( .A(n8748), .ZN(n8035) );
  MUX2_X1 U7734 ( .A(n6130), .B(n6129), .S(n8035), .Z(n6131) );
  NAND2_X1 U7735 ( .A1(n6132), .A2(n6131), .ZN(n6146) );
  OR2_X1 U7736 ( .A1(n6786), .A2(n6133), .ZN(n6136) );
  XNOR2_X1 U7737 ( .A(n6134), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8124) );
  AOI22_X1 U7738 ( .A1(n6180), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6880), .B2(
        n8124), .ZN(n6135) );
  NAND2_X1 U7739 ( .A1(n6282), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6145) );
  INV_X1 U7740 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8107) );
  OR2_X1 U7741 ( .A1(n6185), .A2(n8107), .ZN(n6144) );
  INV_X1 U7742 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6137) );
  OR2_X1 U7743 ( .A1(n6186), .A2(n6137), .ZN(n6143) );
  NAND2_X1 U7744 ( .A1(n6138), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6139) );
  AND2_X1 U7745 ( .A1(n6140), .A2(n6139), .ZN(n8112) );
  OR2_X1 U7746 ( .A1(n6141), .A2(n8112), .ZN(n6142) );
  NAND2_X1 U7747 ( .A1(n8111), .A2(n8532), .ZN(n6346) );
  OR2_X1 U7748 ( .A1(n8542), .A2(n8606), .ZN(n6352) );
  NAND2_X1 U7749 ( .A1(n8542), .A2(n8606), .ZN(n6351) );
  NAND2_X1 U7750 ( .A1(n6352), .A2(n6351), .ZN(n8180) );
  INV_X1 U7751 ( .A(n8180), .ZN(n8183) );
  INV_X1 U7752 ( .A(n8537), .ZN(n8612) );
  AND2_X1 U7753 ( .A1(n8612), .A2(n8746), .ZN(n6348) );
  NAND2_X1 U7754 ( .A1(n8537), .A2(n8539), .ZN(n6349) );
  INV_X1 U7755 ( .A(n6349), .ZN(n6147) );
  NAND3_X1 U7756 ( .A1(n8111), .A2(n8532), .A3(n6508), .ZN(n6148) );
  OAI21_X1 U7757 ( .B1(n6347), .B2(n6508), .A(n6148), .ZN(n6149) );
  NOR2_X1 U7758 ( .A1(n8147), .A2(n6149), .ZN(n6150) );
  INV_X1 U7759 ( .A(n8542), .ZN(n8739) );
  NAND2_X1 U7760 ( .A1(n6348), .A2(n6508), .ZN(n6151) );
  OR2_X1 U7761 ( .A1(n8606), .A2(n5846), .ZN(n6152) );
  NAND2_X1 U7762 ( .A1(n6151), .A2(n6152), .ZN(n6154) );
  INV_X1 U7763 ( .A(n6152), .ZN(n6153) );
  AOI22_X1 U7764 ( .A1(n8739), .A2(n6154), .B1(n6348), .B2(n6153), .ZN(n6155)
         );
  NAND2_X1 U7765 ( .A1(n9168), .A2(n8732), .ZN(n6354) );
  NAND2_X1 U7766 ( .A1(n9027), .A2(n6157), .ZN(n6174) );
  NOR2_X1 U7767 ( .A1(n6174), .A2(n6353), .ZN(n6176) );
  INV_X1 U7768 ( .A(n6354), .ZN(n6173) );
  NAND2_X1 U7769 ( .A1(n7372), .A2(n6229), .ZN(n6165) );
  INV_X1 U7770 ( .A(n6158), .ZN(n6159) );
  NAND2_X1 U7771 ( .A1(n6159), .A2(n10173), .ZN(n6160) );
  NAND2_X1 U7772 ( .A1(n6162), .A2(n6161), .ZN(n6177) );
  OR2_X1 U7773 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  AND2_X1 U7774 ( .A1(n6177), .A2(n6163), .ZN(n8865) );
  AOI22_X1 U7775 ( .A1(n6180), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6880), .B2(
        n8865), .ZN(n6164) );
  NAND2_X1 U7776 ( .A1(n6166), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7777 ( .A1(n6183), .A2(n6167), .ZN(n9017) );
  NAND2_X1 U7778 ( .A1(n6235), .A2(n9017), .ZN(n6171) );
  INV_X1 U7779 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9161) );
  OR2_X1 U7780 ( .A1(n6240), .A2(n9161), .ZN(n6170) );
  INV_X1 U7781 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9097) );
  OR2_X1 U7782 ( .A1(n6185), .A2(n9097), .ZN(n6169) );
  OR2_X1 U7783 ( .A1(n6186), .A2(n10034), .ZN(n6168) );
  NAND4_X1 U7784 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(n9024)
         );
  OAI211_X1 U7785 ( .C1(n6174), .C2(n6173), .A(n6357), .B(n6172), .ZN(n6175)
         );
  MUX2_X1 U7786 ( .A(n6176), .B(n6175), .S(n5846), .Z(n6201) );
  NAND2_X1 U7787 ( .A1(n7527), .A2(n6229), .ZN(n6182) );
  AOI22_X1 U7788 ( .A1(n6180), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8869), .B2(
        n6880), .ZN(n6181) );
  NAND2_X1 U7789 ( .A1(n6183), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7790 ( .A1(n6194), .A2(n6184), .ZN(n9003) );
  NAND2_X1 U7791 ( .A1(n9003), .A2(n6235), .ZN(n6191) );
  INV_X1 U7792 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9092) );
  OR2_X1 U7793 ( .A1(n6185), .A2(n9092), .ZN(n6188) );
  INV_X1 U7794 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9002) );
  OR2_X1 U7795 ( .A1(n6186), .A2(n9002), .ZN(n6187) );
  AND2_X1 U7796 ( .A1(n6188), .A2(n6187), .ZN(n6190) );
  NAND2_X1 U7797 ( .A1(n6282), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7798 ( .A1(n9156), .A2(n9011), .ZN(n6359) );
  NAND2_X1 U7799 ( .A1(n8700), .A2(n8997), .ZN(n6300) );
  NAND3_X1 U7800 ( .A1(n6201), .A2(n6359), .A3(n6300), .ZN(n6199) );
  NAND2_X1 U7801 ( .A1(n7702), .A2(n6229), .ZN(n6193) );
  INV_X1 U7802 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7714) );
  OR2_X1 U7803 ( .A1(n6004), .A2(n7714), .ZN(n6192) );
  NAND2_X1 U7804 ( .A1(n6194), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7805 ( .A1(n6207), .A2(n6195), .ZN(n8986) );
  NAND2_X1 U7806 ( .A1(n8986), .A2(n6235), .ZN(n6198) );
  AOI22_X1 U7807 ( .A1(n6282), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n6237), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7808 ( .A1(n6236), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6196) );
  NAND3_X1 U7809 ( .A1(n6199), .A2(n6358), .A3(n6360), .ZN(n6204) );
  NAND2_X1 U7810 ( .A1(n6300), .A2(n6355), .ZN(n6200) );
  OAI211_X1 U7811 ( .C1(n6201), .C2(n6200), .A(n6358), .B(n6357), .ZN(n6202)
         );
  NAND2_X1 U7812 ( .A1(n6202), .A2(n6359), .ZN(n6203) );
  NAND2_X1 U7813 ( .A1(n9089), .A2(n8998), .ZN(n8969) );
  INV_X1 U7814 ( .A(n8969), .ZN(n6215) );
  NAND2_X1 U7815 ( .A1(n7806), .A2(n6229), .ZN(n6206) );
  OR2_X1 U7816 ( .A1(n6004), .A2(n7849), .ZN(n6205) );
  NAND2_X1 U7817 ( .A1(n6207), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7818 ( .A1(n6209), .A2(n6208), .ZN(n8973) );
  NAND2_X1 U7819 ( .A1(n8973), .A2(n6235), .ZN(n6212) );
  AOI22_X1 U7820 ( .A1(n6282), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n6237), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7821 ( .A1(n6236), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7822 ( .A1(n9085), .A2(n8985), .ZN(n6299) );
  AND2_X1 U7823 ( .A1(n6299), .A2(n8969), .ZN(n6361) );
  AND2_X1 U7824 ( .A1(n6362), .A2(n6360), .ZN(n6213) );
  MUX2_X1 U7825 ( .A(n6361), .B(n6213), .S(n6508), .Z(n6214) );
  NAND2_X1 U7826 ( .A1(n6365), .A2(n6364), .ZN(n8960) );
  INV_X1 U7827 ( .A(n8960), .ZN(n8955) );
  MUX2_X1 U7828 ( .A(n6362), .B(n6299), .S(n6508), .Z(n6216) );
  NAND2_X1 U7829 ( .A1(n8081), .A2(n6229), .ZN(n6219) );
  OR2_X1 U7830 ( .A1(n6004), .A2(n8094), .ZN(n6218) );
  NAND2_X1 U7831 ( .A1(n6220), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7832 ( .A1(n6232), .A2(n6221), .ZN(n8940) );
  NAND2_X1 U7833 ( .A1(n8940), .A2(n6235), .ZN(n6227) );
  INV_X1 U7834 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7835 ( .A1(n6282), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7836 ( .A1(n6237), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6222) );
  OAI211_X1 U7837 ( .C1(n6224), .C2(n6186), .A(n6223), .B(n6222), .ZN(n6225)
         );
  INV_X1 U7838 ( .A(n6225), .ZN(n6226) );
  INV_X1 U7839 ( .A(n8950), .ZN(n9138) );
  INV_X1 U7840 ( .A(n6367), .ZN(n6228) );
  NAND3_X1 U7841 ( .A1(n6247), .A2(n6369), .A3(n6228), .ZN(n6245) );
  NOR2_X1 U7842 ( .A1(n6370), .A2(n6508), .ZN(n6244) );
  NAND2_X1 U7843 ( .A1(n8174), .A2(n6229), .ZN(n6231) );
  OR2_X1 U7844 ( .A1(n6004), .A2(n8177), .ZN(n6230) );
  NAND2_X1 U7845 ( .A1(n6232), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7846 ( .A1(n6234), .A2(n6233), .ZN(n8928) );
  NAND2_X1 U7847 ( .A1(n8928), .A2(n6235), .ZN(n6243) );
  INV_X1 U7848 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U7849 ( .A1(n6236), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7850 ( .A1(n6237), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6238) );
  OAI211_X1 U7851 ( .C1(n6240), .C2(n10187), .A(n6239), .B(n6238), .ZN(n6241)
         );
  INV_X1 U7852 ( .A(n6241), .ZN(n6242) );
  OR2_X1 U7853 ( .A1(n9127), .A2(n8934), .ZN(n6463) );
  NAND2_X1 U7854 ( .A1(n9127), .A2(n8934), .ZN(n6462) );
  NAND2_X1 U7855 ( .A1(n6463), .A2(n6462), .ZN(n8922) );
  NAND4_X1 U7856 ( .A1(n6374), .A2(n6245), .A3(n6244), .A4(n8922), .ZN(n6246)
         );
  OAI211_X1 U7857 ( .C1(n6247), .C2(n6367), .A(n4830), .B(n6368), .ZN(n6249)
         );
  AND2_X1 U7858 ( .A1(n6369), .A2(n6508), .ZN(n6248) );
  NAND4_X1 U7859 ( .A1(n6249), .A2(n6248), .A3(n6375), .A4(n8922), .ZN(n6250)
         );
  OR3_X1 U7860 ( .A1(n9116), .A2(n6508), .A3(n8718), .ZN(n6251) );
  NAND2_X1 U7861 ( .A1(n9127), .A2(n8717), .ZN(n6371) );
  NAND2_X1 U7862 ( .A1(n6371), .A2(n6508), .ZN(n6252) );
  NAND2_X1 U7863 ( .A1(n6374), .A2(n6252), .ZN(n6253) );
  OR2_X1 U7864 ( .A1(n9127), .A2(n8717), .ZN(n6372) );
  NAND3_X1 U7865 ( .A1(n6375), .A2(n5846), .A3(n6372), .ZN(n6254) );
  OAI211_X1 U7866 ( .C1(n6375), .C2(n5846), .A(n6255), .B(n6254), .ZN(n6256)
         );
  NOR3_X1 U7867 ( .A1(n6467), .A2(n6258), .A3(n6260), .ZN(n6259) );
  INV_X1 U7868 ( .A(n6259), .ZN(n6268) );
  MUX2_X1 U7869 ( .A(n8596), .B(n6466), .S(n5846), .Z(n6262) );
  NAND2_X1 U7870 ( .A1(n6263), .A2(n6262), .ZN(n6266) );
  MUX2_X1 U7871 ( .A(n8904), .B(n9062), .S(n6508), .Z(n6264) );
  NAND2_X1 U7872 ( .A1(n6266), .A2(n6265), .ZN(n6267) );
  NAND2_X1 U7873 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  INV_X1 U7874 ( .A(n6271), .ZN(n6384) );
  AOI21_X1 U7875 ( .B1(n6508), .B2(n6272), .A(n6384), .ZN(n6290) );
  NAND2_X1 U7876 ( .A1(n6291), .A2(n5846), .ZN(n6289) );
  INV_X1 U7877 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6277) );
  INV_X1 U7878 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6276) );
  MUX2_X1 U7879 ( .A(n6277), .B(n6276), .S(n4936), .Z(n6278) );
  XNOR2_X1 U7880 ( .A(n6278), .B(SI_31_), .ZN(n6279) );
  MUX2_X1 U7881 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9175), .S(n6632), .Z(n6281) );
  INV_X1 U7882 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7883 ( .A1(n6282), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6284) );
  INV_X1 U7884 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10069) );
  OR2_X1 U7885 ( .A1(n5982), .A2(n10069), .ZN(n6283) );
  OAI211_X1 U7886 ( .C1(n6285), .C2(n6186), .A(n6284), .B(n6283), .ZN(n6286)
         );
  INV_X1 U7887 ( .A(n6286), .ZN(n6287) );
  NAND2_X1 U7888 ( .A1(n6288), .A2(n6287), .ZN(n8510) );
  OR2_X1 U7889 ( .A1(n9112), .A2(n8510), .ZN(n6322) );
  OAI211_X1 U7890 ( .C1(n6291), .C2(n6290), .A(n6289), .B(n6322), .ZN(n6292)
         );
  NAND2_X1 U7891 ( .A1(n9112), .A2(n8510), .ZN(n6386) );
  NAND2_X1 U7892 ( .A1(n6292), .A2(n6386), .ZN(n6297) );
  NAND2_X1 U7893 ( .A1(n6293), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6294) );
  MUX2_X1 U7894 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6294), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6296) );
  NAND2_X1 U7895 ( .A1(n6297), .A2(n7715), .ZN(n6327) );
  INV_X1 U7896 ( .A(n6382), .ZN(n6321) );
  INV_X1 U7897 ( .A(n6298), .ZN(n6320) );
  NAND2_X1 U7898 ( .A1(n6375), .A2(n6374), .ZN(n8912) );
  NAND2_X1 U7899 ( .A1(n6362), .A2(n6299), .ZN(n8971) );
  NAND2_X1 U7900 ( .A1(n6357), .A2(n6300), .ZN(n9016) );
  INV_X1 U7901 ( .A(n9016), .ZN(n6315) );
  NAND2_X1 U7902 ( .A1(n6301), .A2(n6354), .ZN(n9040) );
  INV_X1 U7903 ( .A(n6302), .ZN(n6303) );
  INV_X1 U7904 ( .A(n7050), .ZN(n7263) );
  NOR2_X1 U7905 ( .A1(n6303), .A2(n7263), .ZN(n6971) );
  NAND2_X1 U7906 ( .A1(n6329), .A2(n6304), .ZN(n7385) );
  INV_X1 U7907 ( .A(n7385), .ZN(n7387) );
  NAND2_X1 U7908 ( .A1(n6971), .A2(n7387), .ZN(n6305) );
  AND2_X1 U7909 ( .A1(n6334), .A2(n6333), .ZN(n7282) );
  INV_X1 U7910 ( .A(n7282), .ZN(n7285) );
  NOR4_X1 U7911 ( .A1(n6305), .A2(n7265), .A3(n7285), .A4(n7237), .ZN(n6307)
         );
  NAND4_X1 U7912 ( .A1(n6307), .A2(n7417), .A3(n7427), .A4(n4321), .ZN(n6311)
         );
  XNOR2_X1 U7913 ( .A(n9975), .B(n7900), .ZN(n7818) );
  NAND2_X1 U7914 ( .A1(n6340), .A2(n6308), .ZN(n7705) );
  INV_X1 U7915 ( .A(n7561), .ZN(n6310) );
  NOR4_X1 U7916 ( .A1(n6311), .A2(n7818), .A3(n7705), .A4(n6310), .ZN(n6312)
         );
  OR2_X1 U7917 ( .A1(n9980), .A2(n8749), .ZN(n6440) );
  NAND2_X1 U7918 ( .A1(n9980), .A2(n8749), .ZN(n7979) );
  NAND2_X1 U7919 ( .A1(n6440), .A2(n7979), .ZN(n7963) );
  NAND4_X1 U7920 ( .A1(n8101), .A2(n6312), .A3(n7981), .A4(n7963), .ZN(n6313)
         );
  NOR4_X1 U7921 ( .A1(n8180), .A2(n9040), .A3(n6313), .A4(n8147), .ZN(n6314)
         );
  NAND4_X1 U7922 ( .A1(n8995), .A2(n9027), .A3(n6315), .A4(n6314), .ZN(n6316)
         );
  NOR4_X1 U7923 ( .A1(n8960), .A2(n8971), .A3(n8978), .A4(n6316), .ZN(n6317)
         );
  NAND4_X1 U7924 ( .A1(n4914), .A2(n8922), .A3(n8932), .A4(n6317), .ZN(n6318)
         );
  NOR4_X1 U7925 ( .A1(n8895), .A2(n8900), .A3(n8912), .A4(n6318), .ZN(n6319)
         );
  NAND4_X1 U7926 ( .A1(n6386), .A2(n6321), .A3(n6320), .A4(n6319), .ZN(n6324)
         );
  INV_X1 U7927 ( .A(n6322), .ZN(n6323) );
  AOI21_X1 U7928 ( .B1(n7850), .B2(n6324), .A(n6323), .ZN(n6325) );
  NAND2_X1 U7929 ( .A1(n6325), .A2(n7234), .ZN(n6326) );
  NAND2_X1 U7930 ( .A1(n7248), .A2(n4321), .ZN(n7246) );
  NAND2_X1 U7931 ( .A1(n7246), .A2(n6328), .ZN(n7388) );
  NAND2_X1 U7932 ( .A1(n7388), .A2(n7387), .ZN(n6330) );
  INV_X1 U7933 ( .A(n6333), .ZN(n6335) );
  INV_X1 U7934 ( .A(n6341), .ZN(n7817) );
  OR2_X1 U7935 ( .A1(n9986), .A2(n8035), .ZN(n6345) );
  AOI21_X1 U7936 ( .B1(n9038), .B2(n6354), .A(n6353), .ZN(n9026) );
  NAND2_X1 U7937 ( .A1(n9026), .A2(n9027), .ZN(n6356) );
  NAND2_X1 U7938 ( .A1(n6356), .A2(n6355), .ZN(n9013) );
  NAND2_X1 U7939 ( .A1(n6363), .A2(n6362), .ZN(n8959) );
  NAND2_X1 U7940 ( .A1(n6378), .A2(n6377), .ZN(n8894) );
  NAND2_X1 U7941 ( .A1(n9062), .A2(n8596), .ZN(n6379) );
  INV_X1 U7942 ( .A(n9112), .ZN(n6385) );
  NOR2_X1 U7943 ( .A1(n6385), .A2(n6380), .ZN(n6381) );
  AOI22_X1 U7944 ( .A1(n6387), .A2(n6386), .B1(n6385), .B2(n6384), .ZN(n6388)
         );
  INV_X1 U7945 ( .A(n7715), .ZN(n7234) );
  NAND2_X1 U7946 ( .A1(n6389), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6391) );
  OR2_X1 U7947 ( .A1(n6882), .A2(P2_U3151), .ZN(n8022) );
  OR2_X1 U7948 ( .A1(n6400), .A2(n6393), .ZN(n6394) );
  NAND2_X1 U7949 ( .A1(n6398), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U7950 ( .A1(n6400), .A2(n6399), .ZN(n6402) );
  INV_X1 U7951 ( .A(n6841), .ZN(n9173) );
  INV_X1 U7952 ( .A(n6403), .ZN(n6879) );
  INV_X1 U7953 ( .A(n6404), .ZN(n6869) );
  INV_X2 U7954 ( .A(n6869), .ZN(n8811) );
  NAND2_X1 U7955 ( .A1(n6879), .A2(n8811), .ZN(n6892) );
  NAND2_X1 U7956 ( .A1(n8862), .A2(n7715), .ZN(n6509) );
  NOR3_X1 U7957 ( .A1(n9173), .A2(n6892), .A3(n6972), .ZN(n6406) );
  OAI21_X1 U7958 ( .B1(n8022), .B2(n6470), .A(P2_B_REG_SCAN_IN), .ZN(n6405) );
  AOI21_X1 U7959 ( .B1(n9292), .B2(n6408), .A(n6407), .ZN(n6410) );
  OAI21_X1 U7960 ( .B1(n6410), .B2(n6409), .A(n9307), .ZN(n6417) );
  INV_X1 U7961 ( .A(n9720), .ZN(n9446) );
  OAI22_X1 U7962 ( .A1(n9420), .A2(n9409), .B1(n9222), .B2(n9281), .ZN(n9455)
         );
  INV_X1 U7963 ( .A(n6411), .ZN(n9448) );
  OAI22_X1 U7964 ( .A1(n9448), .A2(n9299), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6412), .ZN(n6413) );
  AOI21_X1 U7965 ( .B1(n9455), .B2(n9301), .A(n6413), .ZN(n6414) );
  OAI21_X1 U7966 ( .B1(n9446), .B2(n9317), .A(n6414), .ZN(n6415) );
  NAND2_X1 U7967 ( .A1(n6417), .A2(n6416), .ZN(P1_U3214) );
  INV_X1 U7968 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U7969 ( .A1(n8869), .A2(n7715), .ZN(n6499) );
  INV_X1 U7970 ( .A(n9971), .ZN(n6478) );
  INV_X1 U7971 ( .A(n6476), .ZN(n6477) );
  NAND2_X1 U7972 ( .A1(n8862), .A2(n6470), .ZN(n6512) );
  NAND2_X1 U7973 ( .A1(n6509), .A2(n6512), .ZN(n6419) );
  NAND3_X1 U7974 ( .A1(n6972), .A2(n9955), .A3(n6419), .ZN(n7822) );
  NAND2_X1 U7975 ( .A1(n7254), .A2(n9920), .ZN(n6422) );
  NAND2_X1 U7976 ( .A1(n8760), .A2(n7051), .ZN(n7264) );
  NAND2_X1 U7977 ( .A1(n6423), .A2(n9926), .ZN(n6424) );
  NAND2_X1 U7978 ( .A1(n6425), .A2(n6424), .ZN(n7384) );
  NAND2_X1 U7979 ( .A1(n7384), .A2(n7385), .ZN(n6427) );
  NAND2_X1 U7980 ( .A1(n7253), .A2(n9934), .ZN(n6426) );
  NAND2_X1 U7981 ( .A1(n6427), .A2(n6426), .ZN(n7238) );
  NAND2_X1 U7982 ( .A1(n7238), .A2(n7060), .ZN(n6428) );
  NAND2_X1 U7983 ( .A1(n6428), .A2(n7243), .ZN(n6429) );
  NAND2_X1 U7984 ( .A1(n7219), .A2(n9946), .ZN(n6431) );
  NAND2_X1 U7985 ( .A1(n7416), .A2(n7429), .ZN(n6432) );
  NAND2_X1 U7986 ( .A1(n6433), .A2(n6432), .ZN(n7428) );
  NAND2_X1 U7987 ( .A1(n7758), .A2(n9956), .ZN(n6434) );
  NAND2_X1 U7988 ( .A1(n9964), .A2(n8752), .ZN(n6435) );
  OR2_X1 U7989 ( .A1(n9969), .A2(n8751), .ZN(n6436) );
  NAND2_X1 U7990 ( .A1(n7706), .A2(n6436), .ZN(n6438) );
  NAND2_X1 U7991 ( .A1(n9969), .A2(n8751), .ZN(n6437) );
  AND2_X1 U7992 ( .A1(n9975), .A2(n8750), .ZN(n7895) );
  NAND2_X1 U7993 ( .A1(n9986), .A2(n8748), .ZN(n6439) );
  NAND2_X1 U7994 ( .A1(n6439), .A2(n7979), .ZN(n6441) );
  OR2_X1 U7995 ( .A1(n7895), .A2(n6441), .ZN(n6443) );
  OR2_X1 U7996 ( .A1(n9975), .A2(n8750), .ZN(n7897) );
  AND2_X1 U7997 ( .A1(n7897), .A2(n6440), .ZN(n7977) );
  NAND2_X1 U7998 ( .A1(n8111), .A2(n8747), .ZN(n6444) );
  OR2_X1 U7999 ( .A1(n8537), .A2(n8746), .ZN(n6445) );
  NAND2_X1 U8000 ( .A1(n8182), .A2(n8180), .ZN(n6447) );
  NAND2_X1 U8001 ( .A1(n8542), .A2(n9042), .ZN(n6446) );
  NAND2_X1 U8002 ( .A1(n6447), .A2(n6446), .ZN(n9039) );
  NAND2_X1 U8003 ( .A1(n9168), .A2(n9023), .ZN(n6448) );
  INV_X1 U8004 ( .A(n9006), .ZN(n6450) );
  INV_X1 U8005 ( .A(n8995), .ZN(n6451) );
  OR2_X1 U8006 ( .A1(n8700), .A2(n9024), .ZN(n8993) );
  AND2_X1 U8007 ( .A1(n6451), .A2(n8993), .ZN(n6452) );
  INV_X1 U8008 ( .A(n9011), .ZN(n8745) );
  NAND2_X1 U8009 ( .A1(n9156), .A2(n8745), .ZN(n6453) );
  INV_X1 U8010 ( .A(n8998), .ZN(n8744) );
  OR2_X1 U8011 ( .A1(n9089), .A2(n8744), .ZN(n6454) );
  NAND2_X1 U8012 ( .A1(n8980), .A2(n6454), .ZN(n8966) );
  AND2_X1 U8013 ( .A1(n8971), .A2(n8960), .ZN(n6455) );
  INV_X1 U8014 ( .A(n8985), .ZN(n8743) );
  OR2_X1 U8015 ( .A1(n9085), .A2(n8743), .ZN(n8953) );
  OR2_X1 U8016 ( .A1(n6457), .A2(n8742), .ZN(n6458) );
  NOR2_X1 U8017 ( .A1(n8950), .A2(n8935), .ZN(n6460) );
  NAND2_X1 U8018 ( .A1(n8950), .A2(n8935), .ZN(n6459) );
  AND2_X1 U8019 ( .A1(n9133), .A2(n8923), .ZN(n6461) );
  OAI22_X1 U8020 ( .A1(n8933), .A2(n6461), .B1(n8923), .B2(n9133), .ZN(n8921)
         );
  NAND2_X1 U8021 ( .A1(n8921), .A2(n6462), .ZN(n6464) );
  NAND2_X1 U8022 ( .A1(n6464), .A2(n6463), .ZN(n8913) );
  NAND2_X1 U8023 ( .A1(n9122), .A2(n8924), .ZN(n6465) );
  XNOR2_X1 U8024 ( .A(n6469), .B(n6468), .ZN(n6471) );
  NAND2_X1 U8025 ( .A1(n8869), .A2(n6470), .ZN(n6497) );
  NAND2_X1 U8026 ( .A1(n6471), .A2(n9046), .ZN(n6475) );
  NAND2_X1 U8027 ( .A1(n6403), .A2(n6869), .ZN(n6472) );
  NAND2_X1 U8028 ( .A1(n6892), .A2(n6472), .ZN(n7040) );
  AND2_X1 U8029 ( .A1(n6614), .A2(P2_B_REG_SCAN_IN), .ZN(n6473) );
  NOR2_X1 U8030 ( .A1(n9012), .A2(n6473), .ZN(n8509) );
  AOI22_X1 U8031 ( .A1(n9041), .A2(n8904), .B1(n8740), .B2(n8509), .ZN(n6474)
         );
  AOI21_X1 U8032 ( .B1(n6478), .B2(n6477), .A(n8525), .ZN(n6520) );
  XNOR2_X1 U8033 ( .A(n8095), .B(P2_B_REG_SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8034 ( .A1(n8178), .A2(n6479), .ZN(n6481) );
  OR2_X1 U8035 ( .A1(n6714), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U8036 ( .A1(n8200), .A2(n8095), .ZN(n6715) );
  NOR2_X1 U8037 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n6486) );
  NOR4_X1 U8038 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6485) );
  NOR4_X1 U8039 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6484) );
  NOR4_X1 U8040 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6483) );
  NAND4_X1 U8041 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n6492)
         );
  NOR4_X1 U8042 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6490) );
  NOR4_X1 U8043 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6489) );
  NOR4_X1 U8044 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6488) );
  NOR4_X1 U8045 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6487) );
  NAND4_X1 U8046 ( .A1(n6490), .A2(n6489), .A3(n6488), .A4(n6487), .ZN(n6491)
         );
  NOR2_X1 U8047 ( .A1(n6492), .A2(n6491), .ZN(n6493) );
  INV_X1 U8048 ( .A(n6510), .ZN(n6820) );
  NOR2_X1 U8049 ( .A1(n6967), .A2(n6820), .ZN(n6496) );
  NAND2_X1 U8050 ( .A1(n8178), .A2(n8200), .ZN(n6494) );
  INV_X1 U8051 ( .A(n9174), .ZN(n6516) );
  NOR2_X1 U8052 ( .A1(n6508), .A2(n9987), .ZN(n6498) );
  NAND2_X1 U8053 ( .A1(n6832), .A2(n6498), .ZN(n6835) );
  NAND2_X1 U8054 ( .A1(n6499), .A2(n9987), .ZN(n8937) );
  NAND2_X1 U8055 ( .A1(n6835), .A2(n8937), .ZN(n6819) );
  NAND2_X1 U8056 ( .A1(n6834), .A2(n6819), .ZN(n6503) );
  NAND2_X1 U8057 ( .A1(n6510), .A2(n6841), .ZN(n6500) );
  NAND2_X1 U8058 ( .A1(n6972), .A2(n6832), .ZN(n6501) );
  NAND2_X1 U8059 ( .A1(n6839), .A2(n6501), .ZN(n6502) );
  MUX2_X1 U8060 ( .A(n6504), .B(n6520), .S(n9988), .Z(n6507) );
  NAND2_X1 U8061 ( .A1(n6507), .A2(n6506), .ZN(P2_U3456) );
  INV_X1 U8062 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U8063 ( .A1(n6509), .A2(n6508), .ZN(n6818) );
  INV_X1 U8064 ( .A(n6967), .ZN(n6514) );
  OR2_X1 U8065 ( .A1(n6512), .A2(n7715), .ZN(n6513) );
  AND2_X1 U8066 ( .A1(n6513), .A2(n5846), .ZN(n6966) );
  OAI21_X1 U8067 ( .B1(n6514), .B2(n6840), .A(n6966), .ZN(n6518) );
  INV_X1 U8068 ( .A(n6966), .ZN(n6515) );
  NAND2_X1 U8069 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  MUX2_X1 U8070 ( .A(n6521), .B(n6520), .S(n10005), .Z(n6523) );
  NAND2_X1 U8071 ( .A1(n10005), .A2(n9987), .ZN(n9099) );
  NAND2_X1 U8072 ( .A1(n6523), .A2(n6522), .ZN(P2_U3488) );
  INV_X1 U8073 ( .A(n9589), .ZN(n9754) );
  NAND2_X1 U8074 ( .A1(n7313), .A2(n6570), .ZN(n7312) );
  INV_X1 U8075 ( .A(n6526), .ZN(n6780) );
  NAND2_X1 U8076 ( .A1(n6780), .A2(n6525), .ZN(n6527) );
  NAND2_X1 U8077 ( .A1(n7312), .A2(n6527), .ZN(n6856) );
  NAND2_X1 U8078 ( .A1(n6856), .A2(n6859), .ZN(n6855) );
  INV_X1 U8079 ( .A(n9344), .ZN(n6572) );
  NAND2_X1 U8080 ( .A1(n6572), .A2(n9835), .ZN(n6528) );
  NAND2_X1 U8081 ( .A1(n6855), .A2(n6528), .ZN(n6847) );
  XNOR2_X1 U8082 ( .A(n9343), .B(n5178), .ZN(n8327) );
  INV_X1 U8083 ( .A(n8327), .ZN(n6848) );
  NAND2_X1 U8084 ( .A1(n6847), .A2(n6848), .ZN(n6846) );
  INV_X1 U8085 ( .A(n9343), .ZN(n6779) );
  NAND2_X1 U8086 ( .A1(n6779), .A2(n7379), .ZN(n6529) );
  NAND2_X1 U8087 ( .A1(n6846), .A2(n6529), .ZN(n6945) );
  XNOR2_X1 U8088 ( .A(n9342), .B(n7326), .ZN(n8331) );
  NAND2_X1 U8089 ( .A1(n6945), .A2(n8331), .ZN(n6944) );
  INV_X1 U8090 ( .A(n9342), .ZN(n6576) );
  NAND2_X1 U8091 ( .A1(n6576), .A2(n7326), .ZN(n6530) );
  NAND2_X1 U8092 ( .A1(n6944), .A2(n6530), .ZN(n6941) );
  INV_X1 U8093 ( .A(n9341), .ZN(n7034) );
  NAND2_X1 U8094 ( .A1(n7034), .A2(n7487), .ZN(n8216) );
  NAND2_X1 U8095 ( .A1(n6955), .A2(n9341), .ZN(n8404) );
  NAND2_X1 U8096 ( .A1(n8216), .A2(n8404), .ZN(n8330) );
  NAND2_X1 U8097 ( .A1(n6941), .A2(n8330), .ZN(n6940) );
  NAND2_X1 U8098 ( .A1(n7034), .A2(n6955), .ZN(n6531) );
  NAND2_X1 U8099 ( .A1(n6940), .A2(n6531), .ZN(n7206) );
  INV_X1 U8100 ( .A(n9340), .ZN(n7126) );
  OR2_X1 U8101 ( .A1(n9818), .A2(n7126), .ZN(n8218) );
  NAND2_X1 U8102 ( .A1(n9818), .A2(n7126), .ZN(n8332) );
  NAND2_X1 U8103 ( .A1(n8218), .A2(n8332), .ZN(n7208) );
  NAND2_X1 U8104 ( .A1(n7206), .A2(n7208), .ZN(n7205) );
  OR2_X1 U8105 ( .A1(n9818), .A2(n9340), .ZN(n6532) );
  NAND2_X1 U8106 ( .A1(n7205), .A2(n6532), .ZN(n7499) );
  INV_X1 U8107 ( .A(n9339), .ZN(n7033) );
  OR2_X1 U8108 ( .A1(n7514), .A2(n7033), .ZN(n8220) );
  NAND2_X1 U8109 ( .A1(n7514), .A2(n7033), .ZN(n8333) );
  INV_X1 U8110 ( .A(n8223), .ZN(n7498) );
  OR2_X1 U8111 ( .A1(n7514), .A2(n9339), .ZN(n6533) );
  OR2_X1 U8112 ( .A1(n9861), .A2(n7125), .ZN(n8221) );
  NAND2_X1 U8113 ( .A1(n9861), .A2(n7125), .ZN(n8227) );
  INV_X1 U8114 ( .A(n9337), .ZN(n6534) );
  OR2_X1 U8115 ( .A1(n7524), .A2(n6534), .ZN(n8244) );
  NAND2_X1 U8116 ( .A1(n7524), .A2(n6534), .ZN(n8235) );
  NAND2_X1 U8117 ( .A1(n8244), .A2(n8235), .ZN(n7397) );
  NAND2_X1 U8118 ( .A1(n7396), .A2(n6535), .ZN(n7357) );
  INV_X1 U8119 ( .A(n9336), .ZN(n6536) );
  NOR2_X1 U8120 ( .A1(n7753), .A2(n6536), .ZN(n8211) );
  INV_X1 U8121 ( .A(n8211), .ZN(n6537) );
  AND2_X1 U8122 ( .A1(n7753), .A2(n6536), .ZN(n8243) );
  INV_X1 U8123 ( .A(n8243), .ZN(n8236) );
  NAND2_X1 U8124 ( .A1(n7357), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U8125 ( .A1(n7355), .A2(n6538), .ZN(n7531) );
  INV_X1 U8126 ( .A(n9335), .ZN(n6539) );
  OR2_X1 U8127 ( .A1(n7889), .A2(n6539), .ZN(n8210) );
  AND2_X1 U8128 ( .A1(n7889), .A2(n6539), .ZN(n8246) );
  INV_X1 U8129 ( .A(n8246), .ZN(n8237) );
  INV_X1 U8130 ( .A(n8341), .ZN(n7530) );
  NAND2_X1 U8131 ( .A1(n7531), .A2(n7530), .ZN(n7529) );
  NAND2_X1 U8132 ( .A1(n7529), .A2(n6540), .ZN(n7682) );
  INV_X1 U8133 ( .A(n9334), .ZN(n6541) );
  NAND2_X1 U8134 ( .A1(n7699), .A2(n6541), .ZN(n8249) );
  NAND2_X1 U8135 ( .A1(n8247), .A2(n8249), .ZN(n8338) );
  NAND2_X1 U8136 ( .A1(n7682), .A2(n8338), .ZN(n7681) );
  NAND2_X1 U8137 ( .A1(n6542), .A2(n6541), .ZN(n6543) );
  NAND2_X1 U8138 ( .A1(n7681), .A2(n6543), .ZN(n7791) );
  INV_X1 U8139 ( .A(n9333), .ZN(n6544) );
  OR2_X1 U8140 ( .A1(n7813), .A2(n6544), .ZN(n8251) );
  NAND2_X1 U8141 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  INV_X1 U8142 ( .A(n9702), .ZN(n9191) );
  INV_X1 U8143 ( .A(n9332), .ZN(n8253) );
  NAND2_X1 U8144 ( .A1(n8267), .A2(n8424), .ZN(n8344) );
  INV_X1 U8145 ( .A(n8344), .ZN(n6584) );
  NOR2_X1 U8146 ( .A1(n9769), .A2(n9282), .ZN(n6549) );
  INV_X1 U8147 ( .A(n9282), .ZN(n9330) );
  INV_X1 U8148 ( .A(n9211), .ZN(n9327) );
  NAND2_X1 U8149 ( .A1(n9673), .A2(n9327), .ZN(n6551) );
  NAND2_X1 U8150 ( .A1(n9745), .A2(n9269), .ZN(n6552) );
  INV_X1 U8151 ( .A(n9269), .ZN(n9325) );
  INV_X1 U8152 ( .A(n9270), .ZN(n9323) );
  NOR2_X1 U8153 ( .A1(n6589), .A2(n9323), .ZN(n6553) );
  INV_X1 U8154 ( .A(n6589), .ZN(n9518) );
  NOR2_X1 U8155 ( .A1(n9499), .A2(n9221), .ZN(n6555) );
  INV_X1 U8156 ( .A(n9221), .ZN(n9322) );
  NOR2_X1 U8157 ( .A1(n9493), .A2(n9321), .ZN(n6556) );
  NOR2_X1 U8158 ( .A1(n6598), .A2(n9222), .ZN(n6557) );
  NAND2_X1 U8159 ( .A1(n9720), .A2(n9295), .ZN(n8303) );
  NAND2_X1 U8160 ( .A1(n9429), .A2(n8303), .ZN(n9451) );
  NAND2_X1 U8161 ( .A1(n6560), .A2(n9420), .ZN(n9431) );
  NAND2_X1 U8162 ( .A1(n8353), .A2(n9431), .ZN(n9428) );
  XNOR2_X1 U8163 ( .A(n9423), .B(n9428), .ZN(n8508) );
  NAND2_X1 U8164 ( .A1(n6562), .A2(n7314), .ZN(n8462) );
  NAND2_X1 U8165 ( .A1(n8462), .A2(n6561), .ZN(n7277) );
  NOR2_X1 U8166 ( .A1(n6562), .A2(n8451), .ZN(n6563) );
  OR2_X1 U8167 ( .A1(n7277), .A2(n6563), .ZN(n7906) );
  NAND2_X1 U8168 ( .A1(n9493), .A2(n9254), .ZN(n8370) );
  NAND2_X1 U8169 ( .A1(n6564), .A2(n9221), .ZN(n8366) );
  NAND2_X1 U8170 ( .A1(n6589), .A2(n9270), .ZN(n9505) );
  OR2_X1 U8171 ( .A1(n9618), .A2(n9282), .ZN(n8275) );
  NAND2_X1 U8172 ( .A1(n9618), .A2(n9282), .ZN(n8271) );
  OR2_X1 U8173 ( .A1(n8012), .A2(n8164), .ZN(n8209) );
  NAND2_X1 U8174 ( .A1(n8012), .A2(n8164), .ZN(n8265) );
  NAND2_X1 U8175 ( .A1(n8209), .A2(n8265), .ZN(n8345) );
  INV_X1 U8176 ( .A(n8345), .ZN(n8002) );
  AND2_X1 U8177 ( .A1(n8244), .A2(n8221), .ZN(n8231) );
  INV_X1 U8178 ( .A(n8231), .ZN(n6567) );
  INV_X1 U8179 ( .A(n8220), .ZN(n6565) );
  INV_X1 U8180 ( .A(n8218), .ZN(n8212) );
  OR3_X1 U8181 ( .A1(n6567), .A2(n6565), .A3(n8212), .ZN(n8408) );
  AND2_X1 U8182 ( .A1(n8235), .A2(n8227), .ZN(n8232) );
  INV_X1 U8183 ( .A(n8232), .ZN(n8337) );
  INV_X1 U8184 ( .A(n8333), .ZN(n6566) );
  OR2_X1 U8185 ( .A1(n8337), .A2(n6566), .ZN(n6569) );
  NAND2_X1 U8186 ( .A1(n6567), .A2(n8235), .ZN(n6568) );
  NAND2_X1 U8187 ( .A1(n6569), .A2(n6568), .ZN(n8409) );
  NAND2_X1 U8188 ( .A1(n8408), .A2(n8409), .ZN(n6579) );
  NOR2_X1 U8189 ( .A1(n6524), .A2(n7317), .ZN(n7305) );
  NAND2_X1 U8190 ( .A1(n6780), .A2(n7321), .ZN(n6571) );
  NAND2_X1 U8191 ( .A1(n7304), .A2(n6571), .ZN(n6860) );
  NAND2_X1 U8192 ( .A1(n9344), .A2(n9835), .ZN(n8400) );
  NAND2_X1 U8193 ( .A1(n6572), .A2(n6963), .ZN(n6573) );
  NOR2_X1 U8194 ( .A1(n9343), .A2(n7379), .ZN(n6575) );
  NAND2_X1 U8195 ( .A1(n9343), .A2(n7379), .ZN(n8401) );
  NAND2_X1 U8196 ( .A1(n9342), .A2(n7326), .ZN(n8403) );
  NAND2_X1 U8197 ( .A1(n6576), .A2(n7004), .ZN(n6929) );
  AND2_X1 U8198 ( .A1(n8216), .A2(n6929), .ZN(n6577) );
  NAND2_X1 U8199 ( .A1(n6930), .A2(n6577), .ZN(n6933) );
  NAND2_X1 U8200 ( .A1(n6933), .A2(n8404), .ZN(n8213) );
  NAND3_X1 U8201 ( .A1(n8407), .A2(n8232), .A3(n8333), .ZN(n6578) );
  NAND2_X1 U8202 ( .A1(n6579), .A2(n6578), .ZN(n7351) );
  INV_X1 U8203 ( .A(n8338), .ZN(n7684) );
  INV_X1 U8204 ( .A(n8247), .ZN(n6580) );
  NOR2_X1 U8205 ( .A1(n7793), .A2(n6580), .ZN(n6581) );
  NAND2_X1 U8206 ( .A1(n7792), .A2(n6581), .ZN(n6582) );
  NAND2_X1 U8207 ( .A1(n6582), .A2(n8414), .ZN(n7908) );
  XNOR2_X1 U8208 ( .A(n9702), .B(n9332), .ZN(n8339) );
  OR2_X1 U8209 ( .A1(n9702), .A2(n8253), .ZN(n8252) );
  NAND3_X1 U8210 ( .A1(n8002), .A2(n8003), .A3(n8252), .ZN(n6583) );
  NAND2_X1 U8211 ( .A1(n6584), .A2(n8162), .ZN(n6585) );
  NAND2_X1 U8212 ( .A1(n6585), .A2(n8267), .ZN(n9611) );
  NAND2_X1 U8213 ( .A1(n9612), .A2(n9611), .ZN(n9610) );
  OR2_X1 U8214 ( .A1(n9684), .A2(n8520), .ZN(n8276) );
  NAND2_X1 U8215 ( .A1(n9684), .A2(n8520), .ZN(n8277) );
  OR2_X1 U8216 ( .A1(n9589), .A2(n9283), .ZN(n8281) );
  NAND2_X1 U8217 ( .A1(n9589), .A2(n9283), .ZN(n8432) );
  NAND2_X1 U8218 ( .A1(n6586), .A2(n8432), .ZN(n8362) );
  INV_X1 U8219 ( .A(n8362), .ZN(n9569) );
  NAND2_X1 U8220 ( .A1(n9673), .A2(n9211), .ZN(n8273) );
  NAND2_X1 U8221 ( .A1(n9569), .A2(n9568), .ZN(n6587) );
  NAND2_X1 U8222 ( .A1(n6587), .A2(n8360), .ZN(n9546) );
  NAND2_X1 U8223 ( .A1(n9554), .A2(n9269), .ZN(n8283) );
  NAND2_X1 U8224 ( .A1(n8436), .A2(n8283), .ZN(n9545) );
  XNOR2_X1 U8225 ( .A(n9540), .B(n9324), .ZN(n9528) );
  NAND2_X1 U8226 ( .A1(n9540), .A2(n9212), .ZN(n8289) );
  INV_X1 U8227 ( .A(n8289), .ZN(n6588) );
  OR2_X1 U8228 ( .A1(n6589), .A2(n9270), .ZN(n8292) );
  NAND2_X1 U8229 ( .A1(n8292), .A2(n9505), .ZN(n9520) );
  NAND3_X1 U8230 ( .A1(n9484), .A2(n9479), .A3(n9506), .ZN(n6590) );
  NAND2_X1 U8231 ( .A1(n6590), .A2(n8370), .ZN(n9469) );
  OR2_X1 U8232 ( .A1(n9648), .A2(n9222), .ZN(n8373) );
  NAND2_X1 U8233 ( .A1(n9648), .A2(n9222), .ZN(n8375) );
  INV_X1 U8234 ( .A(n8375), .ZN(n9452) );
  NAND2_X1 U8235 ( .A1(n9454), .A2(n9429), .ZN(n6591) );
  XNOR2_X1 U8236 ( .A(n6591), .B(n9428), .ZN(n6595) );
  NOR2_X1 U8237 ( .A1(n6592), .A2(n5462), .ZN(n8323) );
  INV_X1 U8238 ( .A(n8394), .ZN(n8395) );
  NAND2_X1 U8239 ( .A1(n8395), .A2(n5719), .ZN(n8454) );
  INV_X1 U8240 ( .A(n8454), .ZN(n6593) );
  NAND2_X1 U8241 ( .A1(n6525), .A2(n7317), .ZN(n7316) );
  OR2_X1 U8242 ( .A1(n7316), .A2(n6963), .ZN(n6857) );
  NAND2_X1 U8243 ( .A1(n6946), .A2(n7326), .ZN(n6938) );
  INV_X1 U8244 ( .A(n7514), .ZN(n9810) );
  AND2_X2 U8245 ( .A1(n7500), .A2(n9810), .ZN(n7501) );
  INV_X1 U8246 ( .A(n7889), .ZN(n7542) );
  NOR2_X1 U8247 ( .A1(n9702), .A2(n7914), .ZN(n8009) );
  NAND2_X1 U8248 ( .A1(n9318), .A2(n8009), .ZN(n8168) );
  NOR2_X1 U8249 ( .A1(n9589), .A2(n9583), .ZN(n9561) );
  NAND2_X1 U8250 ( .A1(n9563), .A2(n9561), .ZN(n9551) );
  NOR2_X2 U8251 ( .A1(n9489), .A2(n9493), .ZN(n9462) );
  OAI211_X1 U8252 ( .C1(n6559), .C2(n4340), .A(n9584), .B(n9438), .ZN(n8502)
         );
  OAI211_X1 U8253 ( .C1(n8508), .C2(n9845), .A(n8505), .B(n8502), .ZN(n6610)
         );
  INV_X1 U8254 ( .A(n6600), .ZN(n6605) );
  OAI21_X1 U8255 ( .B1(n9777), .B2(P1_D_REG_1__SCAN_IN), .A(n9778), .ZN(n6604)
         );
  INV_X1 U8256 ( .A(n6601), .ZN(n6602) );
  OR2_X1 U8257 ( .A1(n9777), .A2(n6602), .ZN(n6603) );
  NAND4_X1 U8258 ( .A1(n7272), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n6609)
         );
  MUX2_X1 U8259 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n6610), .S(n9876), .Z(n6606)
         );
  INV_X1 U8260 ( .A(n6606), .ZN(n6607) );
  NAND2_X1 U8261 ( .A1(n6607), .A2(n4907), .ZN(P1_U3550) );
  INV_X1 U8262 ( .A(n7271), .ZN(n6608) );
  MUX2_X1 U8263 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n6610), .S(n9869), .Z(n6611)
         );
  INV_X1 U8264 ( .A(n6611), .ZN(n6612) );
  NAND2_X1 U8265 ( .A1(n6612), .A2(n4909), .ZN(P1_U3518) );
  INV_X1 U8266 ( .A(n6618), .ZN(n6617) );
  NAND2_X1 U8267 ( .A1(n6884), .A2(n5846), .ZN(n6613) );
  NAND2_X1 U8268 ( .A1(n6613), .A2(n6882), .ZN(n6878) );
  NAND2_X1 U8269 ( .A1(n6878), .A2(n6614), .ZN(n6615) );
  NAND2_X1 U8270 ( .A1(n6615), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U8271 ( .A1(n9798), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6620) );
  INV_X1 U8272 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9872) );
  MUX2_X1 U8273 ( .A(n9872), .B(P1_REG1_REG_1__SCAN_IN), .S(n6666), .Z(n6619)
         );
  NOR2_X1 U8274 ( .A1(n6619), .A2(n6620), .ZN(n6665) );
  AOI21_X1 U8275 ( .B1(n6617), .B2(n8389), .A(n4319), .ZN(n6623) );
  NAND2_X1 U8276 ( .A1(n6618), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8467) );
  NAND2_X1 U8277 ( .A1(n8463), .A2(n8467), .ZN(n6624) );
  NAND2_X1 U8278 ( .A1(n6623), .A2(n6624), .ZN(n9807) );
  INV_X1 U8279 ( .A(n9796), .ZN(n8203) );
  AOI211_X1 U8280 ( .C1(n6620), .C2(n6619), .A(n6665), .B(n9370), .ZN(n6629)
         );
  NAND2_X1 U8281 ( .A1(n9798), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6753) );
  XNOR2_X1 U8282 ( .A(n6666), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6621) );
  NOR2_X1 U8283 ( .A1(n6621), .A2(n6753), .ZN(n6662) );
  NAND2_X1 U8284 ( .A1(n8206), .A2(n8203), .ZN(n8461) );
  AOI211_X1 U8285 ( .C1(n6753), .C2(n6621), .A(n6662), .B(n9387), .ZN(n6628)
         );
  INV_X1 U8286 ( .A(n6666), .ZN(n6622) );
  NOR2_X1 U8287 ( .A1(n9403), .A2(n6622), .ZN(n6627) );
  INV_X1 U8288 ( .A(n6623), .ZN(n6625) );
  INV_X1 U8289 ( .A(n9804), .ZN(n8496) );
  INV_X1 U8290 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7617) );
  INV_X1 U8291 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7311) );
  OAI22_X1 U8292 ( .A1(n8496), .A2(n7617), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7311), .ZN(n6626) );
  OR4_X1 U8293 ( .A1(n6629), .A2(n6628), .A3(n6627), .A4(n6626), .ZN(P1_U3244)
         );
  NOR2_X1 U8294 ( .A1(n6631), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9790) );
  AOI22_X1 U8295 ( .A1(n9790), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n6666), .ZN(n6630) );
  OAI21_X1 U8296 ( .B1(n6643), .B2(n9792), .A(n6630), .ZN(P1_U3354) );
  AND2_X1 U8297 ( .A1(n6631), .A2(P2_U3151), .ZN(n9180) );
  INV_X2 U8298 ( .A(n9180), .ZN(n8590) );
  AND2_X1 U8299 ( .A1(n6632), .A2(P2_U3151), .ZN(n8021) );
  INV_X2 U8300 ( .A(n8021), .ZN(n8587) );
  OAI222_X1 U8301 ( .A1(n8590), .A2(n6633), .B1(n7098), .B2(P2_U3151), .C1(
        n8587), .C2(n6640), .ZN(P2_U3292) );
  OAI222_X1 U8302 ( .A1(n8590), .A2(n4925), .B1(n7026), .B2(P2_U3151), .C1(
        n8587), .C2(n6642), .ZN(P2_U3293) );
  OAI222_X1 U8303 ( .A1(n8590), .A2(n4938), .B1(n7136), .B2(P2_U3151), .C1(
        n8587), .C2(n6635), .ZN(P2_U3291) );
  AOI22_X1 U8304 ( .A1(n6686), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n9786), .ZN(n6634) );
  OAI21_X1 U8305 ( .B1(n6635), .B2(n9792), .A(n6634), .ZN(P1_U3351) );
  AOI22_X1 U8306 ( .A1(n6788), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9786), .ZN(n6636) );
  OAI21_X1 U8307 ( .B1(n6645), .B2(n9792), .A(n6636), .ZN(P1_U3348) );
  AOI22_X1 U8308 ( .A1(n6727), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9786), .ZN(n6637) );
  OAI21_X1 U8309 ( .B1(n6647), .B2(n9792), .A(n6637), .ZN(P1_U3349) );
  AOI22_X1 U8310 ( .A1(n6698), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9786), .ZN(n6638) );
  OAI21_X1 U8311 ( .B1(n6649), .B2(n9792), .A(n6638), .ZN(P1_U3350) );
  AOI22_X1 U8312 ( .A1(n6685), .A2(P1_STATE_REG_SCAN_IN), .B1(n9786), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6639) );
  OAI21_X1 U8313 ( .B1(n6640), .B2(n9792), .A(n6639), .ZN(P1_U3352) );
  AOI22_X1 U8314 ( .A1(n9354), .A2(P1_STATE_REG_SCAN_IN), .B1(n9786), .B2(
        P2_DATAO_REG_2__SCAN_IN), .ZN(n6641) );
  OAI21_X1 U8315 ( .B1(n6642), .B2(n9792), .A(n6641), .ZN(P1_U3353) );
  INV_X1 U8316 ( .A(n6897), .ZN(n6871) );
  OAI222_X1 U8317 ( .A1(n8587), .A2(n6643), .B1(n8590), .B2(n4921), .C1(
        P2_U3151), .C2(n6871), .ZN(P2_U3294) );
  INV_X1 U8318 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6644) );
  OAI222_X1 U8319 ( .A1(n8587), .A2(n6645), .B1(n7589), .B2(P2_U3151), .C1(
        n6644), .C2(n8590), .ZN(P2_U3288) );
  OAI222_X1 U8320 ( .A1(n8587), .A2(n6647), .B1(n7453), .B2(P2_U3151), .C1(
        n6646), .C2(n8590), .ZN(P2_U3289) );
  OAI222_X1 U8321 ( .A1(n8587), .A2(n6649), .B1(n7155), .B2(P2_U3151), .C1(
        n6648), .C2(n8590), .ZN(P2_U3290) );
  NOR2_X1 U8322 ( .A1(n9804), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8323 ( .A(n6650), .ZN(n6652) );
  AOI22_X1 U8324 ( .A1(n6920), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9786), .ZN(n6651) );
  OAI21_X1 U8325 ( .B1(n6652), .B2(n9792), .A(n6651), .ZN(P1_U3347) );
  INV_X1 U8326 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6653) );
  INV_X1 U8327 ( .A(n9903), .ZN(n7586) );
  OAI222_X1 U8328 ( .A1(n8590), .A2(n6653), .B1(n8587), .B2(n6652), .C1(
        P2_U3151), .C2(n7586), .ZN(P2_U3287) );
  INV_X1 U8329 ( .A(n6654), .ZN(n6657) );
  AOI22_X1 U8330 ( .A1(n7200), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9786), .ZN(n6655) );
  OAI21_X1 U8331 ( .B1(n6657), .B2(n9792), .A(n6655), .ZN(P1_U3346) );
  INV_X1 U8332 ( .A(n7718), .ZN(n7724) );
  OAI222_X1 U8333 ( .A1(n8587), .A2(n6657), .B1(n7724), .B2(P2_U3151), .C1(
        n6656), .C2(n8590), .ZN(P2_U3286) );
  AOI22_X1 U8334 ( .A1(n7336), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9790), .ZN(n6658) );
  OAI21_X1 U8335 ( .B1(n6660), .B2(n9792), .A(n6658), .ZN(P1_U3345) );
  INV_X1 U8336 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6659) );
  OAI222_X1 U8337 ( .A1(n8587), .A2(n6660), .B1(n7773), .B2(P2_U3151), .C1(
        n6659), .C2(n8590), .ZN(P2_U3285) );
  INV_X1 U8338 ( .A(P1_U3973), .ZN(n9326) );
  NAND2_X1 U8339 ( .A1(n9326), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6661) );
  OAI21_X1 U8340 ( .B1(n9242), .B2(n9326), .A(n6661), .ZN(P1_U3570) );
  INV_X1 U8341 ( .A(n6685), .ZN(n6677) );
  AOI21_X1 U8342 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6666), .A(n6662), .ZN(
        n9347) );
  XNOR2_X1 U8343 ( .A(n9354), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9346) );
  NOR2_X1 U8344 ( .A1(n9347), .A2(n9346), .ZN(n9345) );
  AOI21_X1 U8345 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n9354), .A(n9345), .ZN(
        n6664) );
  XNOR2_X1 U8346 ( .A(n6685), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6663) );
  AOI211_X1 U8347 ( .C1(n6664), .C2(n6663), .A(n6678), .B(n9387), .ZN(n6673)
         );
  AOI21_X1 U8348 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n6666), .A(n6665), .ZN(
        n9351) );
  INV_X1 U8349 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6667) );
  MUX2_X1 U8350 ( .A(n6667), .B(P1_REG1_REG_2__SCAN_IN), .S(n9354), .Z(n9350)
         );
  OR2_X1 U8351 ( .A1(n9351), .A2(n9350), .ZN(n9348) );
  NAND2_X1 U8352 ( .A1(n9354), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6670) );
  INV_X1 U8353 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6668) );
  MUX2_X1 U8354 ( .A(n6668), .B(P1_REG1_REG_3__SCAN_IN), .S(n6685), .Z(n6669)
         );
  AOI21_X1 U8355 ( .B1(n9348), .B2(n6670), .A(n6669), .ZN(n6684) );
  AND3_X1 U8356 ( .A1(n9348), .A2(n6670), .A3(n6669), .ZN(n6671) );
  NOR3_X1 U8357 ( .A1(n9370), .A2(n6684), .A3(n6671), .ZN(n6672) );
  NOR2_X1 U8358 ( .A1(n6673), .A2(n6672), .ZN(n6676) );
  AND2_X1 U8359 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6674) );
  AOI21_X1 U8360 ( .B1(n9804), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6674), .ZN(
        n6675) );
  OAI211_X1 U8361 ( .C1(n6677), .C2(n9403), .A(n6676), .B(n6675), .ZN(P1_U3246) );
  INV_X1 U8362 ( .A(n6698), .ZN(n6701) );
  INV_X1 U8363 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6679) );
  MUX2_X1 U8364 ( .A(n6679), .B(P1_REG2_REG_4__SCAN_IN), .S(n6686), .Z(n6744)
         );
  INV_X1 U8365 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6680) );
  MUX2_X1 U8366 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6680), .S(n6698), .Z(n6681)
         );
  INV_X1 U8367 ( .A(n6681), .ZN(n6682) );
  NOR2_X1 U8368 ( .A1(n6683), .A2(n6682), .ZN(n6697) );
  AOI211_X1 U8369 ( .C1(n6683), .C2(n6682), .A(n9387), .B(n6697), .ZN(n6692)
         );
  AOI21_X1 U8370 ( .B1(n6685), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6684), .ZN(
        n6739) );
  INV_X1 U8371 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6687) );
  MUX2_X1 U8372 ( .A(n6687), .B(P1_REG1_REG_4__SCAN_IN), .S(n6686), .Z(n6740)
         );
  INV_X1 U8373 ( .A(n6686), .ZN(n6742) );
  OAI22_X1 U8374 ( .A1(n6739), .A2(n6740), .B1(n6687), .B2(n6742), .ZN(n6688)
         );
  INV_X1 U8375 ( .A(n6688), .ZN(n6690) );
  INV_X1 U8376 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10038) );
  MUX2_X1 U8377 ( .A(n10038), .B(P1_REG1_REG_5__SCAN_IN), .S(n6698), .Z(n6689)
         );
  NOR2_X1 U8378 ( .A1(n6690), .A2(n6689), .ZN(n6705) );
  AOI211_X1 U8379 ( .C1(n6690), .C2(n6689), .A(n6705), .B(n9370), .ZN(n6691)
         );
  NOR2_X1 U8380 ( .A1(n6692), .A2(n6691), .ZN(n6696) );
  NOR2_X1 U8381 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6693), .ZN(n6694) );
  AOI21_X1 U8382 ( .B1(n9804), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6694), .ZN(
        n6695) );
  OAI211_X1 U8383 ( .C1(n6701), .C2(n9403), .A(n6696), .B(n6695), .ZN(P1_U3248) );
  INV_X1 U8384 ( .A(n6727), .ZN(n6713) );
  AOI21_X1 U8385 ( .B1(n6698), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6697), .ZN(
        n6700) );
  XNOR2_X1 U8386 ( .A(n6727), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6699) );
  NOR2_X1 U8387 ( .A1(n6701), .A2(n10038), .ZN(n6704) );
  INV_X1 U8388 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6702) );
  MUX2_X1 U8389 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6702), .S(n6727), .Z(n6703)
         );
  OAI21_X1 U8390 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6730) );
  INV_X1 U8391 ( .A(n6730), .ZN(n6707) );
  NOR3_X1 U8392 ( .A1(n6705), .A2(n6704), .A3(n6703), .ZN(n6706) );
  NOR3_X1 U8393 ( .A1(n6707), .A2(n6706), .A3(n9370), .ZN(n6708) );
  NOR2_X1 U8394 ( .A1(n6709), .A2(n6708), .ZN(n6712) );
  AND2_X1 U8395 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6710) );
  AOI21_X1 U8396 ( .B1(n9804), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6710), .ZN(
        n6711) );
  OAI211_X1 U8397 ( .C1(n6713), .C2(n9403), .A(n6712), .B(n6711), .ZN(P1_U3249) );
  INV_X1 U8398 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6718) );
  INV_X1 U8399 ( .A(n6715), .ZN(n6716) );
  AOI22_X1 U8400 ( .A1(n10029), .A2(n6718), .B1(n6717), .B2(n6716), .ZN(
        P2_U3376) );
  NAND2_X1 U8401 ( .A1(n6526), .A2(P1_U3973), .ZN(n6719) );
  OAI21_X1 U8402 ( .B1(P1_U3973), .B2(n4921), .A(n6719), .ZN(P1_U3555) );
  INV_X1 U8403 ( .A(n6720), .ZN(n6759) );
  AOI22_X1 U8404 ( .A1(n7574), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9790), .ZN(n6721) );
  OAI21_X1 U8405 ( .B1(n6759), .B2(n9792), .A(n6721), .ZN(P1_U3344) );
  AND2_X1 U8406 ( .A1(n10029), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8407 ( .A1(n10029), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8408 ( .A1(n10029), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8409 ( .A1(n10029), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8410 ( .A1(n10029), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8411 ( .A1(n10029), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8412 ( .A1(n10029), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8413 ( .A1(n10029), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8414 ( .A1(n10029), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8415 ( .A1(n10029), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8416 ( .A1(n10029), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8417 ( .A1(n10029), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8418 ( .A1(n10029), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8419 ( .A1(n10029), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8420 ( .A1(n10029), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8421 ( .A1(n10029), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8422 ( .A1(n10029), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8423 ( .A1(n10029), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8424 ( .A1(n10029), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8425 ( .A1(n10029), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8426 ( .A1(n10029), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8427 ( .A1(n10029), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8428 ( .A1(n10029), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8429 ( .A1(n10029), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  INV_X1 U8430 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6723) );
  MUX2_X1 U8431 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6723), .S(n6788), .Z(n6724)
         );
  INV_X1 U8432 ( .A(n6724), .ZN(n6725) );
  NOR2_X1 U8433 ( .A1(n6726), .A2(n6725), .ZN(n6787) );
  AOI211_X1 U8434 ( .C1(n6726), .C2(n6725), .A(n9387), .B(n6787), .ZN(n6738)
         );
  INV_X1 U8435 ( .A(n6788), .ZN(n6792) );
  NAND2_X1 U8436 ( .A1(n6727), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6729) );
  INV_X1 U8437 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6791) );
  MUX2_X1 U8438 ( .A(n6791), .B(P1_REG1_REG_7__SCAN_IN), .S(n6788), .Z(n6728)
         );
  AOI21_X1 U8439 ( .B1(n6730), .B2(n6729), .A(n6728), .ZN(n6795) );
  INV_X1 U8440 ( .A(n6795), .ZN(n6732) );
  NAND3_X1 U8441 ( .A1(n6730), .A2(n6729), .A3(n6728), .ZN(n6731) );
  NAND3_X1 U8442 ( .A1(n6732), .A2(n9399), .A3(n6731), .ZN(n6736) );
  NOR2_X1 U8443 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6733), .ZN(n6734) );
  AOI21_X1 U8444 ( .B1(n9804), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6734), .ZN(
        n6735) );
  OAI211_X1 U8445 ( .C1(n9403), .C2(n6792), .A(n6736), .B(n6735), .ZN(n6737)
         );
  OR2_X1 U8446 ( .A1(n6738), .A2(n6737), .ZN(P1_U3250) );
  XOR2_X1 U8447 ( .A(n6740), .B(n6739), .Z(n6748) );
  NAND2_X1 U8448 ( .A1(n9804), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6741) );
  NAND2_X1 U8449 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7005) );
  OAI211_X1 U8450 ( .C1(n9403), .C2(n6742), .A(n6741), .B(n7005), .ZN(n6747)
         );
  AOI211_X1 U8451 ( .C1(n6745), .C2(n6744), .A(n6743), .B(n9387), .ZN(n6746)
         );
  AOI211_X1 U8452 ( .C1(n9399), .C2(n6748), .A(n6747), .B(n6746), .ZN(n6758)
         );
  OAI21_X1 U8453 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(n6811) );
  NAND3_X1 U8454 ( .A1(n6811), .A2(n9796), .A3(n8206), .ZN(n6757) );
  OR2_X1 U8455 ( .A1(n9796), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U8456 ( .A1(n8206), .A2(n6752), .ZN(n9797) );
  NAND2_X1 U8457 ( .A1(n9797), .A2(n4519), .ZN(n9801) );
  INV_X1 U8458 ( .A(n8461), .ZN(n6755) );
  INV_X1 U8459 ( .A(n6753), .ZN(n6754) );
  NAND2_X1 U8460 ( .A1(n6755), .A2(n6754), .ZN(n6756) );
  NAND4_X1 U8461 ( .A1(n6757), .A2(P1_U3973), .A3(n9801), .A4(n6756), .ZN(
        n9356) );
  NAND2_X1 U8462 ( .A1(n6758), .A2(n9356), .ZN(P1_U3247) );
  INV_X1 U8463 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6760) );
  OAI222_X1 U8464 ( .A1(n8590), .A2(n6760), .B1(n8587), .B2(n6759), .C1(
        P2_U3151), .C2(n7938), .ZN(P2_U3284) );
  AOI22_X1 U8465 ( .A1(n7669), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9790), .ZN(n6761) );
  OAI21_X1 U8466 ( .B1(n6769), .B2(n9792), .A(n6761), .ZN(P1_U3343) );
  NAND2_X1 U8467 ( .A1(n4323), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U8468 ( .A1(n4322), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6763) );
  NAND2_X1 U8469 ( .A1(n5165), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6762) );
  NAND2_X1 U8470 ( .A1(n9410), .A2(P1_U3973), .ZN(n6765) );
  OAI21_X1 U8471 ( .B1(P1_U3973), .B2(n6277), .A(n6765), .ZN(P1_U3585) );
  INV_X1 U8472 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10157) );
  NOR2_X1 U8473 ( .A1(n6767), .A2(n10157), .ZN(P2_U3253) );
  INV_X1 U8474 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10161) );
  NOR2_X1 U8475 ( .A1(n6767), .A2(n10161), .ZN(P2_U3236) );
  INV_X1 U8476 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10158) );
  NOR2_X1 U8477 ( .A1(n6767), .A2(n10158), .ZN(P2_U3243) );
  INV_X1 U8478 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10188) );
  NOR2_X1 U8479 ( .A1(n6767), .A2(n10188), .ZN(P2_U3262) );
  INV_X1 U8480 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6766) );
  NOR2_X1 U8481 ( .A1(n6767), .A2(n6766), .ZN(P2_U3234) );
  INV_X1 U8482 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6768) );
  OAI222_X1 U8483 ( .A1(n8587), .A2(n6769), .B1(n8050), .B2(P2_U3151), .C1(
        n6768), .C2(n8590), .ZN(P2_U3283) );
  XOR2_X1 U8484 ( .A(n6771), .B(n6770), .Z(n6776) );
  INV_X1 U8485 ( .A(n9317), .ZN(n9286) );
  NAND2_X1 U8486 ( .A1(n6524), .A2(n9435), .ZN(n6773) );
  NAND2_X1 U8487 ( .A1(n9344), .A2(n9244), .ZN(n6772) );
  NAND2_X1 U8488 ( .A1(n6773), .A2(n6772), .ZN(n7307) );
  AOI22_X1 U8489 ( .A1(n9286), .A2(n7321), .B1(n9301), .B2(n7307), .ZN(n6775)
         );
  NAND2_X1 U8490 ( .A1(n9299), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6810) );
  NAND2_X1 U8491 ( .A1(n6810), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6774) );
  OAI211_X1 U8492 ( .C1(n6776), .C2(n9288), .A(n6775), .B(n6774), .ZN(P1_U3222) );
  XOR2_X1 U8493 ( .A(n6778), .B(n6777), .Z(n6783) );
  OAI22_X1 U8494 ( .A1(n6780), .A2(n9281), .B1(n6779), .B2(n9409), .ZN(n6861)
         );
  AOI22_X1 U8495 ( .A1(n9286), .A2(n6963), .B1(n9301), .B2(n6861), .ZN(n6782)
         );
  NAND2_X1 U8496 ( .A1(n6810), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6781) );
  OAI211_X1 U8497 ( .C1(n6783), .C2(n9288), .A(n6782), .B(n6781), .ZN(P1_U3237) );
  AOI22_X1 U8498 ( .A1(n7996), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9790), .ZN(n6784) );
  OAI21_X1 U8499 ( .B1(n6786), .B2(n9792), .A(n6784), .ZN(P1_U3342) );
  INV_X1 U8500 ( .A(n8124), .ZN(n8129) );
  INV_X1 U8501 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6785) );
  OAI222_X1 U8502 ( .A1(n8587), .A2(n6786), .B1(n8129), .B2(P2_U3151), .C1(
        n6785), .C2(n8590), .ZN(P2_U3282) );
  XNOR2_X1 U8503 ( .A(n6920), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6789) );
  AOI211_X1 U8504 ( .C1(n6790), .C2(n6789), .A(n9387), .B(n6919), .ZN(n6801)
         );
  INV_X1 U8505 ( .A(n6920), .ZN(n6914) );
  NOR2_X1 U8506 ( .A1(n6792), .A2(n6791), .ZN(n6794) );
  INV_X1 U8507 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6915) );
  MUX2_X1 U8508 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6915), .S(n6920), .Z(n6793)
         );
  OAI21_X1 U8509 ( .B1(n6795), .B2(n6794), .A(n6793), .ZN(n6913) );
  OR3_X1 U8510 ( .A1(n6795), .A2(n6794), .A3(n6793), .ZN(n6796) );
  NAND3_X1 U8511 ( .A1(n6913), .A2(n9399), .A3(n6796), .ZN(n6799) );
  AND2_X1 U8512 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6797) );
  AOI21_X1 U8513 ( .B1(n9804), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6797), .ZN(
        n6798) );
  OAI211_X1 U8514 ( .C1(n9403), .C2(n6914), .A(n6799), .B(n6798), .ZN(n6800)
         );
  OR2_X1 U8515 ( .A1(n6801), .A2(n6800), .ZN(P1_U3251) );
  NAND2_X1 U8516 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  XOR2_X1 U8517 ( .A(n6805), .B(n6804), .Z(n6809) );
  AOI22_X1 U8518 ( .A1(n9435), .A2(n9344), .B1(n9342), .B2(n9244), .ZN(n6850)
         );
  INV_X1 U8519 ( .A(n6850), .ZN(n6806) );
  AOI22_X1 U8520 ( .A1(n9286), .A2(n5178), .B1(n9301), .B2(n6806), .ZN(n6808)
         );
  MUX2_X1 U8521 ( .A(n9299), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6807) );
  OAI211_X1 U8522 ( .C1(n6809), .C2(n9288), .A(n6808), .B(n6807), .ZN(P1_U3218) );
  INV_X1 U8523 ( .A(n6810), .ZN(n6815) );
  INV_X1 U8524 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U8525 ( .A1(n6526), .A2(n9244), .ZN(n9843) );
  OAI22_X1 U8526 ( .A1(n9311), .A2(n9843), .B1(n9288), .B2(n6811), .ZN(n6812)
         );
  AOI21_X1 U8527 ( .B1(n9849), .B2(n9286), .A(n6812), .ZN(n6813) );
  OAI21_X1 U8528 ( .B1(n6815), .B2(n6814), .A(n6813), .ZN(P1_U3232) );
  INV_X1 U8529 ( .A(n6816), .ZN(n6867) );
  AOI22_X1 U8530 ( .A1(n7997), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9790), .ZN(n6817) );
  OAI21_X1 U8531 ( .B1(n6867), .B2(n9792), .A(n6817), .ZN(P1_U3341) );
  AND2_X1 U8532 ( .A1(n6884), .A2(n6818), .ZN(n6823) );
  OAI21_X1 U8533 ( .B1(n6821), .B2(n6820), .A(n6819), .ZN(n6822) );
  OAI211_X1 U8534 ( .C1(n6826), .C2(n6832), .A(n6823), .B(n6822), .ZN(n6824)
         );
  NAND2_X1 U8535 ( .A1(n6824), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6829) );
  INV_X1 U8536 ( .A(n6972), .ZN(n6830) );
  NAND2_X1 U8537 ( .A1(n6841), .A2(n6830), .ZN(n6825) );
  OAI21_X1 U8538 ( .B1(n6826), .B2(n6825), .A(n8022), .ZN(n6827) );
  INV_X1 U8539 ( .A(n6827), .ZN(n6828) );
  NOR2_X1 U8540 ( .A1(n8734), .A2(P2_U3151), .ZN(n7080) );
  AND2_X1 U8541 ( .A1(n6834), .A2(n6830), .ZN(n7041) );
  INV_X1 U8542 ( .A(n7041), .ZN(n6831) );
  INV_X1 U8543 ( .A(n6832), .ZN(n6833) );
  NAND2_X1 U8544 ( .A1(n6834), .A2(n6833), .ZN(n6838) );
  INV_X1 U8545 ( .A(n6835), .ZN(n6836) );
  NAND2_X1 U8546 ( .A1(n6839), .A2(n6836), .ZN(n6837) );
  NAND2_X1 U8547 ( .A1(n6839), .A2(n9987), .ZN(n6842) );
  OAI22_X1 U8548 ( .A1(n6971), .A2(n8724), .B1(n8738), .B2(n6980), .ZN(n6843)
         );
  AOI21_X1 U8549 ( .B1(n8686), .B2(n8759), .A(n6843), .ZN(n6844) );
  OAI21_X1 U8550 ( .B1(n7080), .B2(n6845), .A(n6844), .ZN(P2_U3172) );
  OAI21_X1 U8551 ( .B1(n6847), .B2(n6848), .A(n6846), .ZN(n7381) );
  AOI211_X1 U8552 ( .C1(n5178), .C2(n6857), .A(n9616), .B(n6946), .ZN(n7375)
         );
  XNOR2_X1 U8553 ( .A(n6849), .B(n6848), .ZN(n6851) );
  OAI21_X1 U8554 ( .B1(n6851), .B2(n9846), .A(n6850), .ZN(n7374) );
  AOI211_X1 U8555 ( .C1(n9858), .C2(n7381), .A(n7375), .B(n7374), .ZN(n6960)
         );
  INV_X1 U8556 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6852) );
  OAI22_X1 U8557 ( .A1(n9773), .A2(n7379), .B1(n9869), .B2(n6852), .ZN(n6853)
         );
  INV_X1 U8558 ( .A(n6853), .ZN(n6854) );
  OAI21_X1 U8559 ( .B1(n6960), .B2(n9867), .A(n6854), .ZN(P1_U3462) );
  OAI21_X1 U8560 ( .B1(n6856), .B2(n6859), .A(n6855), .ZN(n9837) );
  INV_X1 U8561 ( .A(n6857), .ZN(n6858) );
  AOI211_X1 U8562 ( .C1(n6963), .C2(n7316), .A(n9616), .B(n6858), .ZN(n9829)
         );
  INV_X1 U8563 ( .A(n6859), .ZN(n8326) );
  XNOR2_X1 U8564 ( .A(n6860), .B(n8326), .ZN(n6862) );
  AOI21_X1 U8565 ( .B1(n6862), .B2(n9609), .A(n6861), .ZN(n9840) );
  INV_X1 U8566 ( .A(n9840), .ZN(n6863) );
  AOI211_X1 U8567 ( .C1(n9858), .C2(n9837), .A(n9829), .B(n6863), .ZN(n6965)
         );
  INV_X1 U8568 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6864) );
  OAI22_X1 U8569 ( .A1(n9773), .A2(n9835), .B1(n9869), .B2(n6864), .ZN(n6865)
         );
  INV_X1 U8570 ( .A(n6865), .ZN(n6866) );
  OAI21_X1 U8571 ( .B1(n6965), .B2(n9867), .A(n6866), .ZN(P1_U3459) );
  INV_X1 U8572 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6868) );
  INV_X1 U8573 ( .A(n8139), .ZN(n8769) );
  OAI222_X1 U8574 ( .A1(n8590), .A2(n6868), .B1(n8587), .B2(n6867), .C1(
        P2_U3151), .C2(n8769), .ZN(P2_U3281) );
  MUX2_X1 U8575 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8811), .Z(n7099) );
  XNOR2_X1 U8576 ( .A(n7099), .B(n7098), .ZN(n6877) );
  MUX2_X1 U8577 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6404), .Z(n6872) );
  XNOR2_X1 U8578 ( .A(n6872), .B(n6897), .ZN(n9890) );
  INV_X1 U8579 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6870) );
  MUX2_X1 U8580 ( .A(n6870), .B(n10057), .S(n8811), .Z(n6983) );
  AOI22_X1 U8581 ( .A1(n9890), .A2(n9891), .B1(n6872), .B2(n6871), .ZN(n7010)
         );
  MUX2_X1 U8582 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8811), .Z(n6873) );
  XNOR2_X1 U8583 ( .A(n6873), .B(n7026), .ZN(n7011) );
  INV_X1 U8584 ( .A(n7026), .ZN(n6875) );
  INV_X1 U8585 ( .A(n6873), .ZN(n6874) );
  OAI22_X1 U8586 ( .A1(n7010), .A2(n7011), .B1(n6875), .B2(n6874), .ZN(n6876)
         );
  NOR2_X1 U8587 ( .A1(n6876), .A2(n6877), .ZN(n7101) );
  AOI21_X1 U8588 ( .B1(n6877), .B2(n6876), .A(n7101), .ZN(n6912) );
  INV_X1 U8589 ( .A(n9892), .ZN(n9913) );
  INV_X1 U8590 ( .A(n7098), .ZN(n6910) );
  AND2_X1 U8591 ( .A1(n6878), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6894) );
  INV_X1 U8592 ( .A(n6894), .ZN(n6982) );
  MUX2_X1 U8593 ( .A(n6982), .B(n8841), .S(n6879), .Z(n6881) );
  INV_X1 U8594 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6908) );
  INV_X1 U8595 ( .A(n6882), .ZN(n6883) );
  NOR2_X1 U8596 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  NOR2_X1 U8597 ( .A1(n6403), .A2(n8811), .ZN(n6886) );
  NAND2_X1 U8598 ( .A1(n6894), .A2(n6886), .ZN(n8877) );
  INV_X1 U8599 ( .A(n8877), .ZN(n9904) );
  NAND2_X1 U8600 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n6988), .ZN(n6887) );
  NAND2_X1 U8601 ( .A1(n6897), .A2(n6887), .ZN(n6888) );
  NAND2_X1 U8602 ( .A1(n5987), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U8603 ( .A1(n6888), .A2(n6889), .ZN(n9878) );
  OR2_X1 U8604 ( .A1(n9878), .A2(n9877), .ZN(n9880) );
  NAND2_X1 U8605 ( .A1(n9880), .A2(n6889), .ZN(n7013) );
  NAND2_X1 U8606 ( .A1(n7026), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6890) );
  XNOR2_X1 U8607 ( .A(n7088), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n6891) );
  NOR2_X1 U8608 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7389), .ZN(n7057) );
  AOI21_X1 U8609 ( .B1(n9904), .B2(n6891), .A(n7057), .ZN(n6907) );
  INV_X1 U8610 ( .A(n6892), .ZN(n6893) );
  MUX2_X1 U8611 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5981), .S(n6895), .Z(n7018)
         );
  NAND2_X1 U8612 ( .A1(n6988), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8613 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8614 ( .A1(n5987), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6900) );
  INV_X1 U8615 ( .A(n9882), .ZN(n6899) );
  NAND2_X1 U8616 ( .A1(n9884), .A2(n6900), .ZN(n7017) );
  NAND2_X1 U8617 ( .A1(n7018), .A2(n7017), .ZN(n7016) );
  NAND2_X1 U8618 ( .A1(n7026), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U8619 ( .A1(n7016), .A2(n6901), .ZN(n6902) );
  NAND2_X1 U8620 ( .A1(n6902), .A2(n7098), .ZN(n7083) );
  NAND2_X1 U8621 ( .A1(n6903), .A2(n5995), .ZN(n6904) );
  NAND2_X1 U8622 ( .A1(n7085), .A2(n6904), .ZN(n6905) );
  NAND2_X1 U8623 ( .A1(n8821), .A2(n6905), .ZN(n6906) );
  OAI211_X1 U8624 ( .C1(n6908), .C2(n9896), .A(n6907), .B(n6906), .ZN(n6909)
         );
  AOI21_X1 U8625 ( .B1(n6910), .B2(n9902), .A(n6909), .ZN(n6911) );
  OAI21_X1 U8626 ( .B1(n6912), .B2(n9913), .A(n6911), .ZN(P2_U3185) );
  OAI21_X1 U8627 ( .B1(n6915), .B2(n6914), .A(n6913), .ZN(n6917) );
  INV_X1 U8628 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10047) );
  INV_X1 U8629 ( .A(n7200), .ZN(n6924) );
  AOI22_X1 U8630 ( .A1(n7200), .A2(n10047), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6924), .ZN(n6916) );
  NOR2_X1 U8631 ( .A1(n6916), .A2(n6917), .ZN(n7190) );
  AOI21_X1 U8632 ( .B1(n6917), .B2(n6916), .A(n7190), .ZN(n6928) );
  NOR2_X1 U8633 ( .A1(n7200), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6918) );
  AOI21_X1 U8634 ( .B1(n7200), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6918), .ZN(
        n6922) );
  OAI21_X1 U8635 ( .B1(n6922), .B2(n6921), .A(n7199), .ZN(n6923) );
  INV_X1 U8636 ( .A(n9387), .ZN(n8490) );
  NAND2_X1 U8637 ( .A1(n6923), .A2(n8490), .ZN(n6927) );
  AND2_X1 U8638 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7480) );
  NOR2_X1 U8639 ( .A1(n9403), .A2(n6924), .ZN(n6925) );
  AOI211_X1 U8640 ( .C1(n9804), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7480), .B(
        n6925), .ZN(n6926) );
  OAI211_X1 U8641 ( .C1(n6928), .C2(n9370), .A(n6927), .B(n6926), .ZN(P1_U3252) );
  INV_X1 U8642 ( .A(n8404), .ZN(n6932) );
  NAND2_X1 U8643 ( .A1(n8215), .A2(n8330), .ZN(n6931) );
  OAI211_X1 U8644 ( .C1(n6933), .C2(n6932), .A(n6931), .B(n9609), .ZN(n6937)
         );
  NAND2_X1 U8645 ( .A1(n9342), .A2(n9435), .ZN(n6935) );
  NAND2_X1 U8646 ( .A1(n9340), .A2(n9244), .ZN(n6934) );
  NAND2_X1 U8647 ( .A1(n6935), .A2(n6934), .ZN(n6995) );
  INV_X1 U8648 ( .A(n6995), .ZN(n6936) );
  NAND2_X1 U8649 ( .A1(n6937), .A2(n6936), .ZN(n7490) );
  INV_X1 U8650 ( .A(n6938), .ZN(n6947) );
  OAI211_X1 U8651 ( .C1(n6947), .C2(n6955), .A(n9584), .B(n7207), .ZN(n7489)
         );
  INV_X1 U8652 ( .A(n7489), .ZN(n6939) );
  NOR2_X1 U8653 ( .A1(n7490), .A2(n6939), .ZN(n6958) );
  OAI21_X1 U8654 ( .B1(n6941), .B2(n8330), .A(n6940), .ZN(n7493) );
  OAI22_X1 U8655 ( .A1(n9699), .A2(n6955), .B1(n9876), .B2(n10038), .ZN(n6942)
         );
  AOI21_X1 U8656 ( .B1(n7493), .B2(n9688), .A(n6942), .ZN(n6943) );
  OAI21_X1 U8657 ( .B1(n6958), .B2(n9874), .A(n6943), .ZN(P1_U3527) );
  OAI21_X1 U8658 ( .B1(n6945), .B2(n8331), .A(n6944), .ZN(n7324) );
  INV_X1 U8659 ( .A(n6946), .ZN(n6948) );
  AOI211_X1 U8660 ( .C1(n7004), .C2(n6948), .A(n9616), .B(n6947), .ZN(n7331)
         );
  XNOR2_X1 U8661 ( .A(n6949), .B(n8331), .ZN(n6950) );
  AOI22_X1 U8662 ( .A1(n9435), .A2(n9343), .B1(n9341), .B2(n9244), .ZN(n7007)
         );
  OAI21_X1 U8663 ( .B1(n6950), .B2(n9846), .A(n7007), .ZN(n7325) );
  AOI211_X1 U8664 ( .C1(n9858), .C2(n7324), .A(n7331), .B(n7325), .ZN(n6962)
         );
  INV_X1 U8665 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6951) );
  OAI22_X1 U8666 ( .A1(n9773), .A2(n7326), .B1(n9869), .B2(n6951), .ZN(n6952)
         );
  INV_X1 U8667 ( .A(n6952), .ZN(n6953) );
  OAI21_X1 U8668 ( .B1(n6962), .B2(n9867), .A(n6953), .ZN(P1_U3465) );
  INV_X1 U8669 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6954) );
  OAI22_X1 U8670 ( .A1(n9773), .A2(n6955), .B1(n9869), .B2(n6954), .ZN(n6956)
         );
  AOI21_X1 U8671 ( .B1(n7493), .B2(n9763), .A(n6956), .ZN(n6957) );
  OAI21_X1 U8672 ( .B1(n6958), .B2(n9867), .A(n6957), .ZN(P1_U3468) );
  AOI22_X1 U8673 ( .A1(n9640), .A2(n5178), .B1(n9874), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6959) );
  OAI21_X1 U8674 ( .B1(n6960), .B2(n9874), .A(n6959), .ZN(P1_U3525) );
  AOI22_X1 U8675 ( .A1(n9640), .A2(n7004), .B1(n9874), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6961) );
  OAI21_X1 U8676 ( .B1(n6962), .B2(n9874), .A(n6961), .ZN(P1_U3526) );
  AOI22_X1 U8677 ( .A1(n9640), .A2(n6963), .B1(n9874), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6964) );
  OAI21_X1 U8678 ( .B1(n6965), .B2(n9874), .A(n6964), .ZN(P1_U3524) );
  MUX2_X1 U8679 ( .A(n6967), .B(n9174), .S(n6966), .Z(n6969) );
  NAND2_X1 U8680 ( .A1(n6969), .A2(n6968), .ZN(n6970) );
  INV_X1 U8681 ( .A(n4315), .ZN(n9028) );
  INV_X1 U8682 ( .A(n6971), .ZN(n6977) );
  NAND3_X1 U8683 ( .A1(n6977), .A2(n6972), .A3(n9955), .ZN(n6973) );
  NAND2_X1 U8684 ( .A1(n8759), .A2(n9043), .ZN(n6978) );
  AOI21_X1 U8685 ( .B1(n6973), .B2(n6978), .A(n9037), .ZN(n6974) );
  AOI21_X1 U8686 ( .B1(n9037), .B2(P2_REG2_REG_0__SCAN_IN), .A(n6974), .ZN(
        n6976) );
  NAND2_X1 U8687 ( .A1(n9051), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6975) );
  OAI211_X1 U8688 ( .C1(n9028), .C2(n6980), .A(n6976), .B(n6975), .ZN(P2_U3233) );
  OAI21_X1 U8689 ( .B1(n9046), .B2(n9949), .A(n6977), .ZN(n6979) );
  OAI211_X1 U8690 ( .C1(n9955), .C2(n6980), .A(n6979), .B(n6978), .ZN(n9109)
         );
  NAND2_X1 U8691 ( .A1(n9109), .A2(n9988), .ZN(n6981) );
  OAI21_X1 U8692 ( .B1(n5970), .B2(n9988), .A(n6981), .ZN(P2_U3390) );
  OAI21_X1 U8693 ( .B1(n6982), .B2(n6403), .A(n9913), .ZN(n6985) );
  AOI22_X1 U8694 ( .A1(n6985), .A2(n6984), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6987) );
  INV_X1 U8695 ( .A(n9896), .ZN(n9898) );
  NAND2_X1 U8696 ( .A1(n9898), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n6986) );
  OAI211_X1 U8697 ( .C1(n8840), .C2(n6988), .A(n6987), .B(n6986), .ZN(P2_U3182) );
  AND2_X1 U8698 ( .A1(n6990), .A2(n6989), .ZN(n6991) );
  NAND2_X1 U8699 ( .A1(n6992), .A2(n6991), .ZN(n6994) );
  XNOR2_X1 U8700 ( .A(n6994), .B(n6993), .ZN(n6998) );
  AOI22_X1 U8701 ( .A1(n9301), .A2(n6995), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n6997) );
  INV_X1 U8702 ( .A(n9299), .ZN(n9313) );
  AOI22_X1 U8703 ( .A1(n9286), .A2(n7487), .B1(n7486), .B2(n9313), .ZN(n6996)
         );
  OAI211_X1 U8704 ( .C1(n6998), .C2(n9288), .A(n6997), .B(n6996), .ZN(P1_U3227) );
  INV_X1 U8705 ( .A(n6999), .ZN(n7002) );
  INV_X1 U8706 ( .A(n7000), .ZN(n7001) );
  AOI211_X1 U8707 ( .C1(n7003), .C2(n7002), .A(n9288), .B(n7001), .ZN(n7009)
         );
  AOI22_X1 U8708 ( .A1(n9286), .A2(n7004), .B1(n9313), .B2(n7327), .ZN(n7006)
         );
  OAI211_X1 U8709 ( .C1(n7007), .C2(n9311), .A(n7006), .B(n7005), .ZN(n7008)
         );
  OR2_X1 U8710 ( .A1(n7009), .A2(n7008), .ZN(P1_U3230) );
  XOR2_X1 U8711 ( .A(n7011), .B(n7010), .Z(n7024) );
  INV_X1 U8712 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7022) );
  OAI21_X1 U8713 ( .B1(n7014), .B2(n7013), .A(n7012), .ZN(n7015) );
  AOI22_X1 U8714 ( .A1(n9904), .A2(n7015), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n7021) );
  OAI21_X1 U8715 ( .B1(n7018), .B2(n7017), .A(n7016), .ZN(n7019) );
  NAND2_X1 U8716 ( .A1(n8821), .A2(n7019), .ZN(n7020) );
  OAI211_X1 U8717 ( .C1(n7022), .C2(n9896), .A(n7021), .B(n7020), .ZN(n7023)
         );
  AOI21_X1 U8718 ( .B1(n9892), .B2(n7024), .A(n7023), .ZN(n7025) );
  OAI21_X1 U8719 ( .B1(n7026), .B2(n8840), .A(n7025), .ZN(P2_U3184) );
  NAND2_X1 U8720 ( .A1(n9326), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7027) );
  OAI21_X1 U8721 ( .B1(n9295), .B2(n9326), .A(n7027), .ZN(P1_U3581) );
  INV_X1 U8722 ( .A(n7028), .ZN(n7030) );
  NAND2_X1 U8723 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  XNOR2_X1 U8724 ( .A(n7032), .B(n7031), .ZN(n7037) );
  OAI22_X1 U8725 ( .A1(n7034), .A2(n9281), .B1(n7033), .B2(n9409), .ZN(n7209)
         );
  AOI22_X1 U8726 ( .A1(n9301), .A2(n7209), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7036) );
  AOI22_X1 U8727 ( .A1(n9286), .A2(n9818), .B1(n9313), .B2(n9820), .ZN(n7035)
         );
  OAI211_X1 U8728 ( .C1(n7037), .C2(n9288), .A(n7036), .B(n7035), .ZN(P1_U3239) );
  INV_X1 U8729 ( .A(n7038), .ZN(n7081) );
  AOI22_X1 U8730 ( .A1(n8481), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9790), .ZN(n7039) );
  OAI21_X1 U8731 ( .B1(n7081), .B2(n9792), .A(n7039), .ZN(P1_U3340) );
  INV_X1 U8732 ( .A(n8729), .ZN(n8716) );
  OAI22_X1 U8733 ( .A1(n8716), .A2(n7042), .B1(n8738), .B2(n9920), .ZN(n7043)
         );
  AOI21_X1 U8734 ( .B1(n8686), .B2(n8758), .A(n7043), .ZN(n7056) );
  NAND2_X4 U8735 ( .A1(n7047), .A2(n7046), .ZN(n7064) );
  XNOR2_X1 U8736 ( .A(n7267), .B(n7064), .ZN(n7048) );
  NOR2_X1 U8737 ( .A1(n8759), .A2(n7048), .ZN(n7061) );
  NAND2_X1 U8738 ( .A1(n7053), .A2(n7052), .ZN(n7063) );
  OAI21_X1 U8739 ( .B1(n7053), .B2(n7052), .A(n7063), .ZN(n7054) );
  NAND2_X1 U8740 ( .A1(n7054), .A2(n8714), .ZN(n7055) );
  OAI211_X1 U8741 ( .C1(n7080), .C2(n9888), .A(n7056), .B(n7055), .ZN(P2_U3162) );
  NAND2_X1 U8742 ( .A1(n8729), .A2(n8758), .ZN(n7059) );
  AOI21_X1 U8743 ( .B1(n8657), .B2(n7390), .A(n7057), .ZN(n7058) );
  OAI211_X1 U8744 ( .C1(n7060), .C2(n8731), .A(n7059), .B(n7058), .ZN(n7070)
         );
  XNOR2_X1 U8745 ( .A(n9934), .B(n7064), .ZN(n7107) );
  XNOR2_X1 U8746 ( .A(n7107), .B(n7253), .ZN(n7068) );
  INV_X1 U8747 ( .A(n7061), .ZN(n7062) );
  NAND2_X1 U8748 ( .A1(n7063), .A2(n7062), .ZN(n7073) );
  XNOR2_X1 U8749 ( .A(n9926), .B(n7064), .ZN(n7065) );
  XNOR2_X1 U8750 ( .A(n7065), .B(n8758), .ZN(n7074) );
  NAND2_X1 U8751 ( .A1(n7073), .A2(n7074), .ZN(n7072) );
  NAND2_X1 U8752 ( .A1(n7065), .A2(n6423), .ZN(n7066) );
  AOI211_X1 U8753 ( .C1(n7068), .C2(n7067), .A(n8724), .B(n7109), .ZN(n7069)
         );
  AOI211_X1 U8754 ( .C1(n7389), .C2(n8734), .A(n7070), .B(n7069), .ZN(n7071)
         );
  INV_X1 U8755 ( .A(n7071), .ZN(P2_U3158) );
  OAI21_X1 U8756 ( .B1(n7074), .B2(n7073), .A(n7072), .ZN(n7075) );
  NAND2_X1 U8757 ( .A1(n7075), .A2(n8714), .ZN(n7078) );
  OAI22_X1 U8758 ( .A1(n8716), .A2(n7254), .B1(n9926), .B2(n8738), .ZN(n7076)
         );
  AOI21_X1 U8759 ( .B1(n8686), .B2(n8757), .A(n7076), .ZN(n7077) );
  OAI211_X1 U8760 ( .C1(n7080), .C2(n7079), .A(n7078), .B(n7077), .ZN(P2_U3177) );
  INV_X1 U8761 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7082) );
  INV_X1 U8762 ( .A(n8798), .ZN(n8787) );
  OAI222_X1 U8763 ( .A1(n8590), .A2(n7082), .B1(n8587), .B2(n7081), .C1(
        P2_U3151), .C2(n8787), .ZN(P2_U3280) );
  INV_X1 U8764 ( .A(n7136), .ZN(n7135) );
  XNOR2_X1 U8765 ( .A(n7136), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7084) );
  NAND3_X1 U8766 ( .A1(n7085), .A2(n7084), .A3(n7083), .ZN(n7086) );
  NAND2_X1 U8767 ( .A1(n4533), .A2(n7086), .ZN(n7087) );
  NOR2_X1 U8768 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10068), .ZN(n7113) );
  AOI21_X1 U8769 ( .B1(n8821), .B2(n7087), .A(n7113), .ZN(n7097) );
  NAND2_X1 U8770 ( .A1(n9898), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7096) );
  MUX2_X1 U8771 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7240), .S(n7136), .Z(n7093)
         );
  NAND2_X1 U8772 ( .A1(n7088), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7091) );
  NAND2_X1 U8773 ( .A1(n7089), .A2(n7098), .ZN(n7090) );
  NAND2_X1 U8774 ( .A1(n7091), .A2(n7090), .ZN(n7092) );
  NAND2_X1 U8775 ( .A1(n7092), .A2(n7093), .ZN(n7134) );
  OAI21_X1 U8776 ( .B1(n7093), .B2(n7092), .A(n7134), .ZN(n7094) );
  NAND2_X1 U8777 ( .A1(n9904), .A2(n7094), .ZN(n7095) );
  NAND3_X1 U8778 ( .A1(n7097), .A2(n7096), .A3(n7095), .ZN(n7105) );
  MUX2_X1 U8779 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8811), .Z(n7133) );
  XNOR2_X1 U8780 ( .A(n7133), .B(n7136), .ZN(n7103) );
  NOR2_X1 U8781 ( .A1(n7099), .A2(n7098), .ZN(n7100) );
  OR2_X1 U8782 ( .A1(n7101), .A2(n7100), .ZN(n7102) );
  NOR3_X1 U8783 ( .A1(n7101), .A2(n7100), .A3(n7103), .ZN(n7132) );
  AOI211_X1 U8784 ( .C1(n7103), .C2(n7102), .A(n9913), .B(n7132), .ZN(n7104)
         );
  AOI211_X1 U8785 ( .C1(n9902), .C2(n7135), .A(n7105), .B(n7104), .ZN(n7106)
         );
  INV_X1 U8786 ( .A(n7106), .ZN(P2_U3186) );
  INV_X1 U8787 ( .A(n7107), .ZN(n7108) );
  XNOR2_X1 U8788 ( .A(n7243), .B(n7064), .ZN(n7110) );
  NOR2_X1 U8789 ( .A1(n8756), .A2(n7110), .ZN(n7176) );
  AOI21_X1 U8790 ( .B1(n8756), .B2(n7110), .A(n7176), .ZN(n7111) );
  OAI21_X1 U8791 ( .B1(n7112), .B2(n7111), .A(n7177), .ZN(n7118) );
  INV_X1 U8792 ( .A(n8734), .ZN(n8664) );
  NOR2_X1 U8793 ( .A1(n8664), .A2(n7241), .ZN(n7117) );
  NAND2_X1 U8794 ( .A1(n8729), .A2(n8757), .ZN(n7115) );
  AOI21_X1 U8795 ( .B1(n8657), .B2(n7243), .A(n7113), .ZN(n7114) );
  OAI211_X1 U8796 ( .C1(n7219), .C2(n8731), .A(n7115), .B(n7114), .ZN(n7116)
         );
  AOI211_X1 U8797 ( .C1(n7118), .C2(n8714), .A(n7117), .B(n7116), .ZN(n7119)
         );
  INV_X1 U8798 ( .A(n7119), .ZN(P2_U3170) );
  INV_X1 U8799 ( .A(n7120), .ZN(n7122) );
  NOR2_X1 U8800 ( .A1(n7122), .A2(n7121), .ZN(n7123) );
  XNOR2_X1 U8801 ( .A(n7124), .B(n7123), .ZN(n7131) );
  INV_X1 U8802 ( .A(n9808), .ZN(n7128) );
  OAI22_X1 U8803 ( .A1(n7126), .A2(n9281), .B1(n7125), .B2(n9409), .ZN(n7507)
         );
  AOI22_X1 U8804 ( .A1(n9301), .A2(n7507), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7127) );
  OAI21_X1 U8805 ( .B1(n7128), .B2(n9299), .A(n7127), .ZN(n7129) );
  AOI21_X1 U8806 ( .B1(n7514), .B2(n9286), .A(n7129), .ZN(n7130) );
  OAI21_X1 U8807 ( .B1(n7131), .B2(n9288), .A(n7130), .ZN(P1_U3213) );
  AOI21_X1 U8808 ( .B1(n7133), .B2(n7136), .A(n7132), .ZN(n7149) );
  MUX2_X1 U8809 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8811), .Z(n7145) );
  XNOR2_X1 U8810 ( .A(n7145), .B(n7155), .ZN(n7148) );
  XNOR2_X1 U8811 ( .A(n7149), .B(n7148), .ZN(n7144) );
  INV_X1 U8812 ( .A(n7155), .ZN(n7147) );
  XNOR2_X1 U8813 ( .A(n7154), .B(n7147), .ZN(n7156) );
  XNOR2_X1 U8814 ( .A(n7156), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7142) );
  NAND2_X1 U8815 ( .A1(n7137), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7164) );
  OAI21_X1 U8816 ( .B1(n7137), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7164), .ZN(
        n7138) );
  AND2_X1 U8817 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7182) );
  AOI21_X1 U8818 ( .B1(n7138), .B2(n8821), .A(n7182), .ZN(n7140) );
  NAND2_X1 U8819 ( .A1(n9898), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7139) );
  OAI211_X1 U8820 ( .C1(n8840), .C2(n7155), .A(n7140), .B(n7139), .ZN(n7141)
         );
  AOI21_X1 U8821 ( .B1(n9904), .B2(n7142), .A(n7141), .ZN(n7143) );
  OAI21_X1 U8822 ( .B1(n7144), .B2(n9913), .A(n7143), .ZN(P2_U3187) );
  INV_X1 U8823 ( .A(n7145), .ZN(n7146) );
  OAI22_X1 U8824 ( .A1(n7149), .A2(n7148), .B1(n7147), .B2(n7146), .ZN(n7153)
         );
  INV_X1 U8825 ( .A(n7453), .ZN(n7458) );
  INV_X1 U8826 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7162) );
  MUX2_X1 U8827 ( .A(n7419), .B(n7162), .S(n8811), .Z(n7151) );
  AND2_X1 U8828 ( .A1(n7151), .A2(n7458), .ZN(n7462) );
  INV_X1 U8829 ( .A(n7462), .ZN(n7150) );
  OAI21_X1 U8830 ( .B1(n7458), .B2(n7151), .A(n7150), .ZN(n7152) );
  NOR2_X1 U8831 ( .A1(n7152), .A2(n7153), .ZN(n7461) );
  AOI21_X1 U8832 ( .B1(n7153), .B2(n7152), .A(n7461), .ZN(n7175) );
  AOI22_X1 U8833 ( .A1(n7156), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n7155), .B2(
        n7154), .ZN(n7158) );
  INV_X1 U8834 ( .A(n7158), .ZN(n7160) );
  MUX2_X1 U8835 ( .A(n7419), .B(P2_REG2_REG_6__SCAN_IN), .S(n7453), .Z(n7157)
         );
  INV_X1 U8836 ( .A(n7157), .ZN(n7159) );
  OAI21_X1 U8837 ( .B1(n7160), .B2(n7159), .A(n7457), .ZN(n7173) );
  INV_X1 U8838 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7161) );
  NOR2_X1 U8839 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7161), .ZN(n7226) );
  AOI21_X1 U8840 ( .B1(n9898), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7226), .ZN(
        n7171) );
  INV_X1 U8841 ( .A(n7167), .ZN(n7163) );
  MUX2_X1 U8842 ( .A(n7162), .B(P2_REG1_REG_6__SCAN_IN), .S(n7453), .Z(n7165)
         );
  INV_X1 U8843 ( .A(n7164), .ZN(n7168) );
  INV_X1 U8844 ( .A(n7165), .ZN(n7166) );
  NOR3_X1 U8845 ( .A1(n7168), .A2(n7167), .A3(n7166), .ZN(n7169) );
  OAI21_X1 U8846 ( .B1(n7455), .B2(n7169), .A(n8821), .ZN(n7170) );
  OAI211_X1 U8847 ( .C1(n8840), .C2(n7453), .A(n7171), .B(n7170), .ZN(n7172)
         );
  AOI21_X1 U8848 ( .B1(n9904), .B2(n7173), .A(n7172), .ZN(n7174) );
  OAI21_X1 U8849 ( .B1(n7175), .B2(n9913), .A(n7174), .ZN(P2_U3188) );
  INV_X1 U8850 ( .A(n7176), .ZN(n7179) );
  XNOR2_X1 U8851 ( .A(n7289), .B(n8564), .ZN(n7220) );
  XNOR2_X1 U8852 ( .A(n7219), .B(n7220), .ZN(n7178) );
  AOI21_X1 U8853 ( .B1(n7177), .B2(n7179), .A(n7178), .ZN(n7222) );
  AND3_X1 U8854 ( .A1(n7177), .A2(n7179), .A3(n7178), .ZN(n7180) );
  OAI21_X1 U8855 ( .B1(n7222), .B2(n7180), .A(n8714), .ZN(n7187) );
  INV_X1 U8856 ( .A(n7181), .ZN(n7288) );
  NAND2_X1 U8857 ( .A1(n8729), .A2(n8756), .ZN(n7184) );
  AOI21_X1 U8858 ( .B1(n8657), .B2(n7289), .A(n7182), .ZN(n7183) );
  OAI211_X1 U8859 ( .C1(n7429), .C2(n8731), .A(n7184), .B(n7183), .ZN(n7185)
         );
  AOI21_X1 U8860 ( .B1(n7288), .B2(n8734), .A(n7185), .ZN(n7186) );
  NAND2_X1 U8861 ( .A1(n7187), .A2(n7186), .ZN(P2_U3167) );
  INV_X1 U8862 ( .A(n7188), .ZN(n7218) );
  AOI22_X1 U8863 ( .A1(n9366), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9786), .ZN(n7189) );
  OAI21_X1 U8864 ( .B1(n7218), .B2(n9792), .A(n7189), .ZN(P1_U3339) );
  INV_X1 U8865 ( .A(n7336), .ZN(n7341) );
  NOR2_X1 U8866 ( .A1(n7200), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7191) );
  NOR2_X1 U8867 ( .A1(n7191), .A2(n7190), .ZN(n7194) );
  INV_X1 U8868 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7192) );
  MUX2_X1 U8869 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7192), .S(n7336), .Z(n7193)
         );
  NAND2_X1 U8870 ( .A1(n7193), .A2(n7194), .ZN(n7340) );
  OAI211_X1 U8871 ( .C1(n7194), .C2(n7193), .A(n7340), .B(n9399), .ZN(n7197)
         );
  AND2_X1 U8872 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7195) );
  AOI21_X1 U8873 ( .B1(n9804), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7195), .ZN(
        n7196) );
  OAI211_X1 U8874 ( .C1(n9403), .C2(n7341), .A(n7197), .B(n7196), .ZN(n7204)
         );
  INV_X1 U8875 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7198) );
  AOI22_X1 U8876 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7341), .B1(n7336), .B2(
        n7198), .ZN(n7202) );
  OAI21_X1 U8877 ( .B1(n7200), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7199), .ZN(
        n7201) );
  NOR2_X1 U8878 ( .A1(n7202), .A2(n7201), .ZN(n7335) );
  AOI211_X1 U8879 ( .C1(n7202), .C2(n7201), .A(n7335), .B(n9387), .ZN(n7203)
         );
  OR2_X1 U8880 ( .A1(n7204), .A2(n7203), .ZN(P1_U3253) );
  OAI21_X1 U8881 ( .B1(n7206), .B2(n7208), .A(n7205), .ZN(n9825) );
  AOI211_X1 U8882 ( .C1(n9818), .C2(n7207), .A(n9616), .B(n7500), .ZN(n9819)
         );
  XNOR2_X1 U8883 ( .A(n8213), .B(n7208), .ZN(n7210) );
  AOI21_X1 U8884 ( .B1(n7210), .B2(n9609), .A(n7209), .ZN(n9827) );
  INV_X1 U8885 ( .A(n9827), .ZN(n7211) );
  AOI211_X1 U8886 ( .C1(n9858), .C2(n9825), .A(n9819), .B(n7211), .ZN(n7216)
         );
  INV_X1 U8887 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7212) );
  NOR2_X1 U8888 ( .A1(n9869), .A2(n7212), .ZN(n7213) );
  AOI21_X1 U8889 ( .B1(n9721), .B2(n9818), .A(n7213), .ZN(n7214) );
  OAI21_X1 U8890 ( .B1(n7216), .B2(n9867), .A(n7214), .ZN(P1_U3471) );
  AOI22_X1 U8891 ( .A1(n9640), .A2(n9818), .B1(n9874), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7215) );
  OAI21_X1 U8892 ( .B1(n7216), .B2(n9874), .A(n7215), .ZN(P1_U3528) );
  INV_X1 U8893 ( .A(n8806), .ZN(n8818) );
  OAI222_X1 U8894 ( .A1(n8587), .A2(n7218), .B1(n8818), .B2(P2_U3151), .C1(
        n7217), .C2(n8590), .ZN(P2_U3279) );
  NOR2_X1 U8895 ( .A1(n7222), .A2(n7221), .ZN(n7223) );
  XNOR2_X1 U8896 ( .A(n9951), .B(n7064), .ZN(n7362) );
  XNOR2_X1 U8897 ( .A(n8754), .B(n7362), .ZN(n7224) );
  OAI211_X1 U8898 ( .C1(n7223), .C2(n7224), .A(n7365), .B(n8714), .ZN(n7231)
         );
  INV_X1 U8899 ( .A(n7225), .ZN(n7420) );
  NAND2_X1 U8900 ( .A1(n8729), .A2(n8755), .ZN(n7228) );
  AOI21_X1 U8901 ( .B1(n8657), .B2(n7421), .A(n7226), .ZN(n7227) );
  OAI211_X1 U8902 ( .C1(n7758), .C2(n8731), .A(n7228), .B(n7227), .ZN(n7229)
         );
  AOI21_X1 U8903 ( .B1(n7420), .B2(n8734), .A(n7229), .ZN(n7230) );
  NAND2_X1 U8904 ( .A1(n7231), .A2(n7230), .ZN(P2_U3179) );
  INV_X1 U8905 ( .A(n7232), .ZN(n7293) );
  AOI22_X1 U8906 ( .A1(n9375), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9786), .ZN(n7233) );
  OAI21_X1 U8907 ( .B1(n7293), .B2(n9792), .A(n7233), .ZN(P1_U3338) );
  OR3_X1 U8908 ( .A1(n8862), .A2(n7234), .A3(n7850), .ZN(n7426) );
  NAND2_X1 U8909 ( .A1(n7822), .A2(n7426), .ZN(n7235) );
  XNOR2_X1 U8910 ( .A(n7236), .B(n7237), .ZN(n9938) );
  XNOR2_X1 U8911 ( .A(n7238), .B(n7237), .ZN(n7239) );
  AOI222_X1 U8912 ( .A1(n9046), .A2(n7239), .B1(n8755), .B2(n9043), .C1(n8757), 
        .C2(n9041), .ZN(n9939) );
  MUX2_X1 U8913 ( .A(n7240), .B(n9939), .S(n9047), .Z(n7245) );
  INV_X1 U8914 ( .A(n7241), .ZN(n7242) );
  AOI22_X1 U8915 ( .A1(n4315), .A2(n7243), .B1(n9051), .B2(n7242), .ZN(n7244)
         );
  OAI211_X1 U8916 ( .C1(n9055), .C2(n9938), .A(n7245), .B(n7244), .ZN(P2_U3229) );
  OAI21_X1 U8917 ( .B1(n7248), .B2(n4321), .A(n7246), .ZN(n9930) );
  INV_X1 U8918 ( .A(n9930), .ZN(n9927) );
  AND2_X1 U8919 ( .A1(n7250), .A2(n7249), .ZN(n7252) );
  XNOR2_X1 U8920 ( .A(n7252), .B(n7251), .ZN(n7256) );
  OAI22_X1 U8921 ( .A1(n7254), .A2(n9010), .B1(n7253), .B2(n9012), .ZN(n7255)
         );
  AOI21_X1 U8922 ( .B1(n7256), .B2(n9046), .A(n7255), .ZN(n9925) );
  INV_X1 U8923 ( .A(n8937), .ZN(n7257) );
  AOI22_X1 U8924 ( .A1(n7258), .A2(n7257), .B1(n9051), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7259) );
  AND2_X1 U8925 ( .A1(n9925), .A2(n7259), .ZN(n7260) );
  MUX2_X1 U8926 ( .A(n7261), .B(n7260), .S(n9047), .Z(n7262) );
  OAI21_X1 U8927 ( .B1(n9927), .B2(n9055), .A(n7262), .ZN(P2_U3231) );
  XNOR2_X1 U8928 ( .A(n7265), .B(n7263), .ZN(n9921) );
  XNOR2_X1 U8929 ( .A(n7265), .B(n7264), .ZN(n7266) );
  AOI222_X1 U8930 ( .A1(n9046), .A2(n7266), .B1(n8760), .B2(n9041), .C1(n8758), 
        .C2(n9043), .ZN(n9919) );
  MUX2_X1 U8931 ( .A(n9877), .B(n9919), .S(n9047), .Z(n7269) );
  AOI22_X1 U8932 ( .A1(n4315), .A2(n7267), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9051), .ZN(n7268) );
  OAI211_X1 U8933 ( .C1(n9921), .C2(n9055), .A(n7269), .B(n7268), .ZN(P2_U3232) );
  NAND4_X1 U8934 ( .A1(n7272), .A2(n7271), .A3(n7270), .A4(n9778), .ZN(n7273)
         );
  INV_X1 U8935 ( .A(n7274), .ZN(n7275) );
  AOI21_X1 U8936 ( .B1(n9828), .B2(n9850), .A(n9590), .ZN(n7281) );
  INV_X1 U8937 ( .A(n7305), .ZN(n7276) );
  NAND2_X1 U8938 ( .A1(n6524), .A2(n7317), .ZN(n8399) );
  AND2_X1 U8939 ( .A1(n7276), .A2(n8399), .ZN(n9844) );
  OAI21_X1 U8940 ( .B1(n9844), .B2(n7277), .A(n9843), .ZN(n7278) );
  INV_X1 U8941 ( .A(n9601), .ZN(n9830) );
  AOI22_X1 U8942 ( .A1(n7278), .A2(n9624), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9830), .ZN(n7280) );
  NAND2_X1 U8943 ( .A1(n9620), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7279) );
  OAI211_X1 U8944 ( .C1(n7281), .C2(n7317), .A(n7280), .B(n7279), .ZN(P1_U3293) );
  XNOR2_X1 U8945 ( .A(n7283), .B(n7282), .ZN(n9944) );
  INV_X1 U8946 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7287) );
  OAI21_X1 U8947 ( .B1(n4918), .B2(n7285), .A(n7284), .ZN(n7286) );
  AOI222_X1 U8948 ( .A1(n9046), .A2(n7286), .B1(n8754), .B2(n9043), .C1(n8756), 
        .C2(n9041), .ZN(n9945) );
  MUX2_X1 U8949 ( .A(n7287), .B(n9945), .S(n9047), .Z(n7291) );
  AOI22_X1 U8950 ( .A1(n4315), .A2(n7289), .B1(n9051), .B2(n7288), .ZN(n7290)
         );
  OAI211_X1 U8951 ( .C1(n9944), .C2(n9055), .A(n7291), .B(n7290), .ZN(P2_U3228) );
  INV_X1 U8952 ( .A(n8846), .ZN(n7292) );
  OAI222_X1 U8953 ( .A1(n8590), .A2(n10037), .B1(n8587), .B2(n7293), .C1(
        P2_U3151), .C2(n7292), .ZN(P2_U3278) );
  AOI21_X1 U8954 ( .B1(n7296), .B2(n7295), .A(n7294), .ZN(n7303) );
  INV_X1 U8955 ( .A(n7443), .ZN(n7300) );
  NAND2_X1 U8956 ( .A1(n9337), .A2(n9244), .ZN(n7298) );
  NAND2_X1 U8957 ( .A1(n9339), .A2(n9435), .ZN(n7297) );
  NAND2_X1 U8958 ( .A1(n7298), .A2(n7297), .ZN(n7447) );
  AOI22_X1 U8959 ( .A1(n9301), .A2(n7447), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7299) );
  OAI21_X1 U8960 ( .B1(n7300), .B2(n9299), .A(n7299), .ZN(n7301) );
  AOI21_X1 U8961 ( .B1(n9861), .B2(n9286), .A(n7301), .ZN(n7302) );
  OAI21_X1 U8962 ( .B1(n7303), .B2(n9288), .A(n7302), .ZN(P1_U3221) );
  OAI21_X1 U8963 ( .B1(n7305), .B2(n8325), .A(n7304), .ZN(n7306) );
  NAND2_X1 U8964 ( .A1(n7306), .A2(n9609), .ZN(n7309) );
  INV_X1 U8965 ( .A(n7307), .ZN(n7308) );
  NAND2_X1 U8966 ( .A1(n7309), .A2(n7308), .ZN(n9854) );
  INV_X1 U8967 ( .A(n9854), .ZN(n7323) );
  NAND2_X1 U8968 ( .A1(n9620), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7310) );
  OAI21_X1 U8969 ( .B1(n7311), .B2(n9601), .A(n7310), .ZN(n7320) );
  INV_X1 U8970 ( .A(n9856), .ZN(n7318) );
  NAND2_X1 U8971 ( .A1(n7314), .A2(n8455), .ZN(n7913) );
  AND2_X1 U8972 ( .A1(n7906), .A2(n7913), .ZN(n7315) );
  OAI211_X1 U8973 ( .C1(n6525), .C2(n7317), .A(n9584), .B(n7316), .ZN(n9852)
         );
  OAI22_X1 U8974 ( .A1(n7318), .A2(n9626), .B1(n9586), .B2(n9852), .ZN(n7319)
         );
  AOI211_X1 U8975 ( .C1(n9590), .C2(n7321), .A(n7320), .B(n7319), .ZN(n7322)
         );
  OAI21_X1 U8976 ( .B1(n9831), .B2(n7323), .A(n7322), .ZN(P1_U3292) );
  INV_X1 U8977 ( .A(n7324), .ZN(n7334) );
  NAND2_X1 U8978 ( .A1(n7325), .A2(n9624), .ZN(n7333) );
  NOR2_X1 U8979 ( .A1(n9834), .A2(n7326), .ZN(n7330) );
  INV_X1 U8980 ( .A(n7327), .ZN(n7328) );
  OAI22_X1 U8981 ( .A1(n9624), .A2(n6679), .B1(n7328), .B2(n9601), .ZN(n7329)
         );
  AOI211_X1 U8982 ( .C1(n7331), .C2(n9828), .A(n7330), .B(n7329), .ZN(n7332)
         );
  OAI211_X1 U8983 ( .C1(n7334), .C2(n9626), .A(n7333), .B(n7332), .ZN(P1_U3289) );
  INV_X1 U8984 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7337) );
  INV_X1 U8985 ( .A(n7574), .ZN(n7568) );
  AOI22_X1 U8986 ( .A1(n7574), .A2(n7337), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7568), .ZN(n7338) );
  AOI211_X1 U8987 ( .C1(n7339), .C2(n7338), .A(n7573), .B(n9387), .ZN(n7348)
         );
  XNOR2_X1 U8988 ( .A(n7568), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7343) );
  OAI21_X1 U8989 ( .B1(n7341), .B2(n7192), .A(n7340), .ZN(n7342) );
  NAND2_X1 U8990 ( .A1(n7343), .A2(n7342), .ZN(n7566) );
  OAI211_X1 U8991 ( .C1(n7343), .C2(n7342), .A(n9399), .B(n7566), .ZN(n7346)
         );
  NAND2_X1 U8992 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7886) );
  INV_X1 U8993 ( .A(n7886), .ZN(n7344) );
  AOI21_X1 U8994 ( .B1(n9804), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7344), .ZN(
        n7345) );
  OAI211_X1 U8995 ( .C1(n9403), .C2(n7568), .A(n7346), .B(n7345), .ZN(n7347)
         );
  OR2_X1 U8996 ( .A1(n7348), .A2(n7347), .ZN(P1_U3254) );
  INV_X1 U8997 ( .A(n7349), .ZN(n7350) );
  AOI21_X1 U8998 ( .B1(n7351), .B2(n7356), .A(n7350), .ZN(n7354) );
  NAND2_X1 U8999 ( .A1(n9335), .A2(n9244), .ZN(n7353) );
  NAND2_X1 U9000 ( .A1(n9337), .A2(n9435), .ZN(n7352) );
  AND2_X1 U9001 ( .A1(n7353), .A2(n7352), .ZN(n7750) );
  OAI21_X1 U9002 ( .B1(n7354), .B2(n9846), .A(n7750), .ZN(n7407) );
  AOI21_X1 U9003 ( .B1(n7752), .B2(n9830), .A(n7407), .ZN(n7361) );
  OAI21_X1 U9004 ( .B1(n7357), .B2(n7356), .A(n7355), .ZN(n7409) );
  NAND2_X1 U9005 ( .A1(n7409), .A2(n9838), .ZN(n7360) );
  AOI211_X1 U9006 ( .C1(n7753), .C2(n7399), .A(n9616), .B(n7537), .ZN(n7408)
         );
  OAI22_X1 U9007 ( .A1(n4527), .A2(n9834), .B1(n9624), .B2(n7198), .ZN(n7358)
         );
  AOI21_X1 U9008 ( .B1(n7408), .B2(n9828), .A(n7358), .ZN(n7359) );
  OAI211_X1 U9009 ( .C1(n9831), .C2(n7361), .A(n7360), .B(n7359), .ZN(P1_U3283) );
  XNOR2_X1 U9010 ( .A(n7436), .B(n7064), .ZN(n7757) );
  XNOR2_X1 U9011 ( .A(n7757), .B(n8753), .ZN(n7367) );
  AOI21_X1 U9012 ( .B1(n7367), .B2(n7366), .A(n4392), .ZN(n7371) );
  AOI22_X1 U9013 ( .A1(n8686), .A2(n8752), .B1(n7436), .B2(n8657), .ZN(n7370)
         );
  AND2_X1 U9014 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7467) );
  NOR2_X1 U9015 ( .A1(n8664), .A2(n7434), .ZN(n7368) );
  AOI211_X1 U9016 ( .C1(n8729), .C2(n8754), .A(n7467), .B(n7368), .ZN(n7369)
         );
  OAI211_X1 U9017 ( .C1(n7371), .C2(n8724), .A(n7370), .B(n7369), .ZN(P2_U3153) );
  INV_X1 U9018 ( .A(n7372), .ZN(n7495) );
  AOI22_X1 U9019 ( .A1(n9386), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9786), .ZN(n7373) );
  OAI21_X1 U9020 ( .B1(n7495), .B2(n9792), .A(n7373), .ZN(P1_U3337) );
  INV_X1 U9021 ( .A(n7374), .ZN(n7383) );
  NAND2_X1 U9022 ( .A1(n7375), .A2(n9828), .ZN(n7378) );
  AOI22_X1 U9023 ( .A1(n9831), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9830), .B2(
        n7376), .ZN(n7377) );
  OAI211_X1 U9024 ( .C1(n7379), .C2(n9834), .A(n7378), .B(n7377), .ZN(n7380)
         );
  AOI21_X1 U9025 ( .B1(n9838), .B2(n7381), .A(n7380), .ZN(n7382) );
  OAI21_X1 U9026 ( .B1(n9831), .B2(n7383), .A(n7382), .ZN(P1_U3290) );
  XNOR2_X1 U9027 ( .A(n7385), .B(n7384), .ZN(n7386) );
  AOI222_X1 U9028 ( .A1(n9046), .A2(n7386), .B1(n8756), .B2(n9043), .C1(n8758), 
        .C2(n9041), .ZN(n9933) );
  XNOR2_X1 U9029 ( .A(n7388), .B(n7387), .ZN(n9936) );
  INV_X1 U9030 ( .A(n9055), .ZN(n9035) );
  AOI22_X1 U9031 ( .A1(n4315), .A2(n7390), .B1(n9051), .B2(n7389), .ZN(n7391)
         );
  OAI21_X1 U9032 ( .B1(n5997), .B2(n9047), .A(n7391), .ZN(n7392) );
  AOI21_X1 U9033 ( .B1(n9936), .B2(n9035), .A(n7392), .ZN(n7393) );
  OAI21_X1 U9034 ( .B1(n9933), .B2(n9037), .A(n7393), .ZN(P2_U3230) );
  NOR2_X1 U9035 ( .A1(n8407), .A2(n8212), .ZN(n7504) );
  NAND2_X1 U9036 ( .A1(n7504), .A2(n8223), .ZN(n7503) );
  NAND2_X1 U9037 ( .A1(n7503), .A2(n8333), .ZN(n7446) );
  OR2_X1 U9038 ( .A1(n7446), .A2(n4882), .ZN(n7448) );
  NAND2_X1 U9039 ( .A1(n7448), .A2(n8221), .ZN(n7394) );
  XOR2_X1 U9040 ( .A(n7397), .B(n7394), .Z(n7395) );
  NAND2_X1 U9041 ( .A1(n9338), .A2(n9435), .ZN(n7478) );
  OAI21_X1 U9042 ( .B1(n7395), .B2(n9846), .A(n7478), .ZN(n7517) );
  INV_X1 U9043 ( .A(n7517), .ZN(n7406) );
  OAI21_X1 U9044 ( .B1(n7398), .B2(n7397), .A(n7396), .ZN(n7519) );
  INV_X1 U9045 ( .A(n7524), .ZN(n7521) );
  INV_X1 U9046 ( .A(n7441), .ZN(n7400) );
  OAI211_X1 U9047 ( .C1(n7400), .C2(n7521), .A(n9584), .B(n7399), .ZN(n7401)
         );
  NAND2_X1 U9048 ( .A1(n9336), .A2(n9244), .ZN(n7477) );
  NAND2_X1 U9049 ( .A1(n7401), .A2(n7477), .ZN(n7518) );
  NAND2_X1 U9050 ( .A1(n7518), .A2(n9828), .ZN(n7403) );
  AOI22_X1 U9051 ( .A1(n9620), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7481), .B2(
        n9830), .ZN(n7402) );
  OAI211_X1 U9052 ( .C1(n7521), .C2(n9834), .A(n7403), .B(n7402), .ZN(n7404)
         );
  AOI21_X1 U9053 ( .B1(n7519), .B2(n9838), .A(n7404), .ZN(n7405) );
  OAI21_X1 U9054 ( .B1(n7406), .B2(n9620), .A(n7405), .ZN(P1_U3284) );
  AOI211_X1 U9055 ( .C1(n7409), .C2(n9858), .A(n7408), .B(n7407), .ZN(n7414)
         );
  INV_X1 U9056 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7410) );
  NOR2_X1 U9057 ( .A1(n9869), .A2(n7410), .ZN(n7411) );
  AOI21_X1 U9058 ( .B1(n7753), .B2(n9721), .A(n7411), .ZN(n7412) );
  OAI21_X1 U9059 ( .B1(n7414), .B2(n9867), .A(n7412), .ZN(P1_U3483) );
  AOI22_X1 U9060 ( .A1(n7753), .A2(n9640), .B1(n9874), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7413) );
  OAI21_X1 U9061 ( .B1(n7414), .B2(n9874), .A(n7413), .ZN(P1_U3532) );
  XOR2_X1 U9062 ( .A(n7415), .B(n7417), .Z(n9952) );
  XOR2_X1 U9063 ( .A(n7417), .B(n7416), .Z(n7418) );
  AOI222_X1 U9064 ( .A1(n9046), .A2(n7418), .B1(n8755), .B2(n9041), .C1(n8753), 
        .C2(n9043), .ZN(n9950) );
  MUX2_X1 U9065 ( .A(n7419), .B(n9950), .S(n9047), .Z(n7423) );
  AOI22_X1 U9066 ( .A1(n4315), .A2(n7421), .B1(n9051), .B2(n7420), .ZN(n7422)
         );
  OAI211_X1 U9067 ( .C1(n9055), .C2(n9952), .A(n7423), .B(n7422), .ZN(P2_U3227) );
  NAND2_X1 U9068 ( .A1(n4475), .A2(n7424), .ZN(n7425) );
  AND2_X1 U9069 ( .A1(n7560), .A2(n7425), .ZN(n7431) );
  INV_X1 U9070 ( .A(n7431), .ZN(n9957) );
  OR2_X1 U9071 ( .A1(n9037), .A2(n7426), .ZN(n8531) );
  XNOR2_X1 U9072 ( .A(n7428), .B(n7427), .ZN(n7433) );
  INV_X1 U9073 ( .A(n7822), .ZN(n9931) );
  OAI22_X1 U9074 ( .A1(n7429), .A2(n9010), .B1(n7828), .B2(n9012), .ZN(n7430)
         );
  AOI21_X1 U9075 ( .B1(n7431), .B2(n9931), .A(n7430), .ZN(n7432) );
  OAI21_X1 U9076 ( .B1(n9007), .B2(n7433), .A(n7432), .ZN(n9959) );
  NAND2_X1 U9077 ( .A1(n9959), .A2(n9047), .ZN(n7438) );
  OAI22_X1 U9078 ( .A1(n9047), .A2(n7460), .B1(n7434), .B2(n9030), .ZN(n7435)
         );
  AOI21_X1 U9079 ( .B1(n4315), .B2(n7436), .A(n7435), .ZN(n7437) );
  OAI211_X1 U9080 ( .C1(n9957), .C2(n8531), .A(n7438), .B(n7437), .ZN(P2_U3226) );
  XNOR2_X1 U9081 ( .A(n7440), .B(n7439), .ZN(n9859) );
  OAI211_X1 U9082 ( .C1(n7501), .C2(n7442), .A(n9584), .B(n7441), .ZN(n9863)
         );
  AOI22_X1 U9083 ( .A1(n9620), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7443), .B2(
        n9830), .ZN(n7445) );
  NAND2_X1 U9084 ( .A1(n9861), .A2(n9590), .ZN(n7444) );
  OAI211_X1 U9085 ( .C1(n9863), .C2(n9586), .A(n7445), .B(n7444), .ZN(n7451)
         );
  AOI21_X1 U9086 ( .B1(n7446), .B2(n4882), .A(n9846), .ZN(n7449) );
  AOI21_X1 U9087 ( .B1(n7449), .B2(n7448), .A(n7447), .ZN(n9865) );
  NOR2_X1 U9088 ( .A1(n9865), .A2(n9831), .ZN(n7450) );
  AOI211_X1 U9089 ( .C1(n9838), .C2(n9859), .A(n7451), .B(n7450), .ZN(n7452)
         );
  INV_X1 U9090 ( .A(n7452), .ZN(P1_U3285) );
  INV_X1 U9091 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9997) );
  AOI21_X1 U9092 ( .B1(n7456), .B2(n9997), .A(n7583), .ZN(n7472) );
  OAI21_X1 U9093 ( .B1(n7458), .B2(n7419), .A(n7457), .ZN(n7588) );
  XNOR2_X1 U9094 ( .A(n7588), .B(n7598), .ZN(n7459) );
  NAND2_X1 U9095 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(n7459), .ZN(n7590) );
  OAI21_X1 U9096 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7459), .A(n7590), .ZN(
        n7470) );
  MUX2_X1 U9097 ( .A(n7460), .B(n9997), .S(n8811), .Z(n7599) );
  XNOR2_X1 U9098 ( .A(n7599), .B(n7598), .ZN(n7464) );
  NOR2_X1 U9099 ( .A1(n7462), .A2(n7461), .ZN(n7463) );
  NOR2_X1 U9100 ( .A1(n7463), .A2(n7464), .ZN(n7597) );
  AOI21_X1 U9101 ( .B1(n7464), .B2(n7463), .A(n7597), .ZN(n7465) );
  NOR2_X1 U9102 ( .A1(n9913), .A2(n7465), .ZN(n7466) );
  AOI211_X1 U9103 ( .C1(n9898), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7467), .B(
        n7466), .ZN(n7468) );
  OAI21_X1 U9104 ( .B1(n7589), .B2(n8840), .A(n7468), .ZN(n7469) );
  AOI21_X1 U9105 ( .B1(n9904), .B2(n7470), .A(n7469), .ZN(n7471) );
  OAI21_X1 U9106 ( .B1(n7472), .B2(n9908), .A(n7471), .ZN(P2_U3189) );
  XNOR2_X1 U9107 ( .A(n7474), .B(n7473), .ZN(n7475) );
  XNOR2_X1 U9108 ( .A(n7476), .B(n7475), .ZN(n7484) );
  AOI21_X1 U9109 ( .B1(n7478), .B2(n7477), .A(n9311), .ZN(n7479) );
  AOI211_X1 U9110 ( .C1(n9313), .C2(n7481), .A(n7480), .B(n7479), .ZN(n7483)
         );
  NAND2_X1 U9111 ( .A1(n7524), .A2(n9286), .ZN(n7482) );
  OAI211_X1 U9112 ( .C1(n7484), .C2(n9288), .A(n7483), .B(n7482), .ZN(P1_U3231) );
  NAND2_X1 U9113 ( .A1(n8510), .A2(P2_U3893), .ZN(n7485) );
  OAI21_X1 U9114 ( .B1(P2_U3893), .B2(n6276), .A(n7485), .ZN(P2_U3522) );
  AOI22_X1 U9115 ( .A1(n9590), .A2(n7487), .B1(n7486), .B2(n9830), .ZN(n7488)
         );
  OAI21_X1 U9116 ( .B1(n7489), .B2(n9586), .A(n7488), .ZN(n7492) );
  MUX2_X1 U9117 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7490), .S(n9624), .Z(n7491)
         );
  AOI211_X1 U9118 ( .C1(n9838), .C2(n7493), .A(n7492), .B(n7491), .ZN(n7494)
         );
  INV_X1 U9119 ( .A(n7494), .ZN(P1_U3288) );
  INV_X1 U9120 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7496) );
  INV_X1 U9121 ( .A(n8865), .ZN(n8849) );
  OAI222_X1 U9122 ( .A1(n8590), .A2(n7496), .B1(n8849), .B2(P2_U3151), .C1(
        n8587), .C2(n7495), .ZN(P2_U3277) );
  INV_X1 U9123 ( .A(n9706), .ZN(n7510) );
  OAI21_X1 U9124 ( .B1(n7499), .B2(n7498), .A(n7497), .ZN(n9814) );
  INV_X1 U9125 ( .A(n7500), .ZN(n7502) );
  AOI211_X1 U9126 ( .C1(n7514), .C2(n7502), .A(n9616), .B(n7501), .ZN(n9812)
         );
  OAI21_X1 U9127 ( .B1(n8223), .B2(n7504), .A(n7503), .ZN(n7508) );
  INV_X1 U9128 ( .A(n9814), .ZN(n7505) );
  NOR2_X1 U9129 ( .A1(n7505), .A2(n7906), .ZN(n7506) );
  AOI211_X1 U9130 ( .C1(n9609), .C2(n7508), .A(n7507), .B(n7506), .ZN(n9817)
         );
  INV_X1 U9131 ( .A(n9817), .ZN(n7509) );
  AOI211_X1 U9132 ( .C1(n7510), .C2(n9814), .A(n9812), .B(n7509), .ZN(n7516)
         );
  INV_X1 U9133 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7511) );
  OAI22_X1 U9134 ( .A1(n9773), .A2(n9810), .B1(n9869), .B2(n7511), .ZN(n7512)
         );
  INV_X1 U9135 ( .A(n7512), .ZN(n7513) );
  OAI21_X1 U9136 ( .B1(n7516), .B2(n9867), .A(n7513), .ZN(P1_U3474) );
  AOI22_X1 U9137 ( .A1(n9640), .A2(n7514), .B1(n9874), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7515) );
  OAI21_X1 U9138 ( .B1(n7516), .B2(n9874), .A(n7515), .ZN(P1_U3529) );
  AOI211_X1 U9139 ( .C1(n9858), .C2(n7519), .A(n7518), .B(n7517), .ZN(n7526)
         );
  INV_X1 U9140 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7520) );
  OAI22_X1 U9141 ( .A1(n7521), .A2(n9773), .B1(n9869), .B2(n7520), .ZN(n7522)
         );
  INV_X1 U9142 ( .A(n7522), .ZN(n7523) );
  OAI21_X1 U9143 ( .B1(n7526), .B2(n9867), .A(n7523), .ZN(P1_U3480) );
  AOI22_X1 U9144 ( .A1(n7524), .A2(n9640), .B1(n9874), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7525) );
  OAI21_X1 U9145 ( .B1(n7526), .B2(n9874), .A(n7525), .ZN(P1_U3531) );
  INV_X1 U9146 ( .A(n7527), .ZN(n7552) );
  AOI22_X1 U9147 ( .A1(n8455), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n9786), .ZN(n7528) );
  OAI21_X1 U9148 ( .B1(n7552), .B2(n9792), .A(n7528), .ZN(P1_U3336) );
  OAI21_X1 U9149 ( .B1(n7531), .B2(n7530), .A(n7529), .ZN(n7548) );
  INV_X1 U9150 ( .A(n7548), .ZN(n7545) );
  OAI211_X1 U9151 ( .C1(n7533), .C2(n8341), .A(n7532), .B(n9609), .ZN(n7536)
         );
  NAND2_X1 U9152 ( .A1(n9336), .A2(n9435), .ZN(n7535) );
  NAND2_X1 U9153 ( .A1(n9334), .A2(n9244), .ZN(n7534) );
  AND2_X1 U9154 ( .A1(n7535), .A2(n7534), .ZN(n7887) );
  NAND2_X1 U9155 ( .A1(n7536), .A2(n7887), .ZN(n7546) );
  INV_X1 U9156 ( .A(n7537), .ZN(n7539) );
  INV_X1 U9157 ( .A(n7689), .ZN(n7538) );
  AOI211_X1 U9158 ( .C1(n7889), .C2(n7539), .A(n9616), .B(n7538), .ZN(n7547)
         );
  NAND2_X1 U9159 ( .A1(n7547), .A2(n9828), .ZN(n7541) );
  AOI22_X1 U9160 ( .A1(n9620), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7884), .B2(
        n9830), .ZN(n7540) );
  OAI211_X1 U9161 ( .C1(n7542), .C2(n9834), .A(n7541), .B(n7540), .ZN(n7543)
         );
  AOI21_X1 U9162 ( .B1(n9624), .B2(n7546), .A(n7543), .ZN(n7544) );
  OAI21_X1 U9163 ( .B1(n7545), .B2(n9626), .A(n7544), .ZN(P1_U3282) );
  AOI211_X1 U9164 ( .C1(n7548), .C2(n9858), .A(n7547), .B(n7546), .ZN(n7551)
         );
  AOI22_X1 U9165 ( .A1(n7889), .A2(n9721), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n9867), .ZN(n7549) );
  OAI21_X1 U9166 ( .B1(n7551), .B2(n9867), .A(n7549), .ZN(P1_U3486) );
  AOI22_X1 U9167 ( .A1(n7889), .A2(n9640), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n9874), .ZN(n7550) );
  OAI21_X1 U9168 ( .B1(n7551), .B2(n9874), .A(n7550), .ZN(P1_U3533) );
  OAI222_X1 U9169 ( .A1(n8590), .A2(n7553), .B1(n8587), .B2(n7552), .C1(
        P2_U3151), .C2(n8862), .ZN(P2_U3276) );
  AOI21_X1 U9170 ( .B1(n7554), .B2(n7561), .A(n9007), .ZN(n7558) );
  OAI22_X1 U9171 ( .A1(n7555), .A2(n9012), .B1(n7758), .B2(n9010), .ZN(n7556)
         );
  AOI21_X1 U9172 ( .B1(n7558), .B2(n7557), .A(n7556), .ZN(n9961) );
  OAI22_X1 U9173 ( .A1(n9047), .A2(n7595), .B1(n7762), .B2(n9030), .ZN(n7564)
         );
  NAND2_X1 U9174 ( .A1(n7560), .A2(n7559), .ZN(n7562) );
  XNOR2_X1 U9175 ( .A(n7562), .B(n7561), .ZN(n9960) );
  NOR2_X1 U9176 ( .A1(n9960), .A2(n9055), .ZN(n7563) );
  AOI211_X1 U9177 ( .C1(n4315), .C2(n9964), .A(n7564), .B(n7563), .ZN(n7565)
         );
  OAI21_X1 U9178 ( .B1(n9037), .B2(n9961), .A(n7565), .ZN(P2_U3225) );
  INV_X1 U9179 ( .A(n9403), .ZN(n9367) );
  INV_X1 U9180 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7567) );
  OAI21_X1 U9181 ( .B1(n7568), .B2(n7567), .A(n7566), .ZN(n7570) );
  XNOR2_X1 U9182 ( .A(n7669), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7569) );
  NOR2_X1 U9183 ( .A1(n7570), .A2(n7569), .ZN(n7670) );
  AOI21_X1 U9184 ( .B1(n7570), .B2(n7569), .A(n7670), .ZN(n7572) );
  AND2_X1 U9185 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7928) );
  AOI21_X1 U9186 ( .B1(n9804), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7928), .ZN(
        n7571) );
  OAI21_X1 U9187 ( .B1(n7572), .B2(n9370), .A(n7571), .ZN(n7579) );
  NOR2_X1 U9188 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7669), .ZN(n7575) );
  AOI21_X1 U9189 ( .B1(n7669), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7575), .ZN(
        n7576) );
  AOI221_X1 U9190 ( .B1(n7577), .B2(n7666), .C1(n7576), .C2(n7666), .A(n9387), 
        .ZN(n7578) );
  AOI211_X1 U9191 ( .C1(n9367), .C2(n7669), .A(n7579), .B(n7578), .ZN(n7580)
         );
  INV_X1 U9192 ( .A(n7580), .ZN(P1_U3255) );
  XNOR2_X1 U9193 ( .A(n9903), .B(n7594), .ZN(n9907) );
  NAND2_X1 U9194 ( .A1(n7586), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7584) );
  XNOR2_X1 U9195 ( .A(n7718), .B(n7717), .ZN(n7585) );
  AOI21_X1 U9196 ( .B1(n7601), .B2(n7585), .A(n7719), .ZN(n7615) );
  NAND2_X1 U9197 ( .A1(n7586), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7592) );
  MUX2_X1 U9198 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7595), .S(n9903), .Z(n7587)
         );
  INV_X1 U9199 ( .A(n7587), .ZN(n9900) );
  NAND2_X1 U9200 ( .A1(n7589), .A2(n7588), .ZN(n7591) );
  NAND2_X1 U9201 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n7593), .ZN(n7725) );
  OAI21_X1 U9202 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7593), .A(n7725), .ZN(
        n7613) );
  NOR2_X1 U9203 ( .A1(n8840), .A2(n7724), .ZN(n7612) );
  INV_X1 U9204 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7633) );
  MUX2_X1 U9205 ( .A(n7595), .B(n7594), .S(n8811), .Z(n7596) );
  NAND2_X1 U9206 ( .A1(n7596), .A2(n9903), .ZN(n7600) );
  OAI21_X1 U9207 ( .B1(n7596), .B2(n9903), .A(n7600), .ZN(n9911) );
  AOI21_X1 U9208 ( .B1(n7599), .B2(n7598), .A(n7597), .ZN(n9912) );
  NOR2_X1 U9209 ( .A1(n9911), .A2(n9912), .ZN(n9910) );
  INV_X1 U9210 ( .A(n7600), .ZN(n7606) );
  MUX2_X1 U9211 ( .A(n7710), .B(n7601), .S(n8811), .Z(n7602) );
  NAND2_X1 U9212 ( .A1(n7602), .A2(n7718), .ZN(n7736) );
  INV_X1 U9213 ( .A(n7602), .ZN(n7603) );
  NAND2_X1 U9214 ( .A1(n7603), .A2(n7724), .ZN(n7604) );
  AND2_X1 U9215 ( .A1(n7736), .A2(n7604), .ZN(n7605) );
  OAI21_X1 U9216 ( .B1(n9910), .B2(n7606), .A(n7605), .ZN(n7737) );
  INV_X1 U9217 ( .A(n7737), .ZN(n7608) );
  NOR3_X1 U9218 ( .A1(n9910), .A2(n7606), .A3(n7605), .ZN(n7607) );
  OAI21_X1 U9219 ( .B1(n7608), .B2(n7607), .A(n9892), .ZN(n7610) );
  AND2_X1 U9220 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7840) );
  INV_X1 U9221 ( .A(n7840), .ZN(n7609) );
  OAI211_X1 U9222 ( .C1(n7633), .C2(n9896), .A(n7610), .B(n7609), .ZN(n7611)
         );
  AOI211_X1 U9223 ( .C1(n7613), .C2(n9904), .A(n7612), .B(n7611), .ZN(n7614)
         );
  OAI21_X1 U9224 ( .B1(n7615), .B2(n9908), .A(n7614), .ZN(P2_U3191) );
  NOR2_X1 U9225 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7660) );
  NOR2_X1 U9226 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7657) );
  NOR2_X1 U9227 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7654) );
  NOR2_X1 U9228 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7651) );
  NOR2_X1 U9229 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7648) );
  NOR2_X1 U9230 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7646) );
  NOR2_X1 U9231 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7642) );
  NOR2_X1 U9232 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7639) );
  NOR2_X1 U9233 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7636) );
  NOR2_X1 U9234 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7632) );
  NOR2_X1 U9235 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7630) );
  NOR2_X1 U9236 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7628) );
  NOR2_X1 U9237 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7626) );
  NOR2_X1 U9238 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7624) );
  NAND2_X1 U9239 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7622) );
  XOR2_X1 U9240 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10233) );
  NAND2_X1 U9241 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7620) );
  AOI21_X1 U9242 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10006) );
  NAND2_X1 U9243 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7616) );
  NOR2_X1 U9244 ( .A1(n7617), .A2(n7616), .ZN(n10007) );
  NOR2_X1 U9245 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10007), .ZN(n7618) );
  NOR2_X1 U9246 ( .A1(n10006), .A2(n7618), .ZN(n10231) );
  XOR2_X1 U9247 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10230) );
  NAND2_X1 U9248 ( .A1(n10231), .A2(n10230), .ZN(n7619) );
  NAND2_X1 U9249 ( .A1(n7620), .A2(n7619), .ZN(n10232) );
  NAND2_X1 U9250 ( .A1(n10233), .A2(n10232), .ZN(n7621) );
  NAND2_X1 U9251 ( .A1(n7622), .A2(n7621), .ZN(n10235) );
  XNOR2_X1 U9252 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10234) );
  NOR2_X1 U9253 ( .A1(n10235), .A2(n10234), .ZN(n7623) );
  NOR2_X1 U9254 ( .A1(n7624), .A2(n7623), .ZN(n10223) );
  XNOR2_X1 U9255 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10222) );
  NOR2_X1 U9256 ( .A1(n10223), .A2(n10222), .ZN(n7625) );
  NOR2_X1 U9257 ( .A1(n7626), .A2(n7625), .ZN(n10221) );
  XNOR2_X1 U9258 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10220) );
  NOR2_X1 U9259 ( .A1(n10221), .A2(n10220), .ZN(n7627) );
  NOR2_X1 U9260 ( .A1(n7628), .A2(n7627), .ZN(n10227) );
  XNOR2_X1 U9261 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10226) );
  NOR2_X1 U9262 ( .A1(n10227), .A2(n10226), .ZN(n7629) );
  NOR2_X1 U9263 ( .A1(n7630), .A2(n7629), .ZN(n10229) );
  XNOR2_X1 U9264 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10228) );
  NOR2_X1 U9265 ( .A1(n10229), .A2(n10228), .ZN(n7631) );
  NOR2_X1 U9266 ( .A1(n7632), .A2(n7631), .ZN(n10225) );
  INV_X1 U9267 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7634) );
  AOI22_X1 U9268 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7634), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7633), .ZN(n10224) );
  NOR2_X1 U9269 ( .A1(n10225), .A2(n10224), .ZN(n7635) );
  NOR2_X1 U9270 ( .A1(n7636), .A2(n7635), .ZN(n10028) );
  INV_X1 U9271 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7637) );
  INV_X1 U9272 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7742) );
  AOI22_X1 U9273 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7637), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7742), .ZN(n10027) );
  NOR2_X1 U9274 ( .A1(n10028), .A2(n10027), .ZN(n7638) );
  NOR2_X1 U9275 ( .A1(n7639), .A2(n7638), .ZN(n10026) );
  INV_X1 U9276 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7640) );
  INV_X1 U9277 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7782) );
  AOI22_X1 U9278 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n7640), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7782), .ZN(n10025) );
  NOR2_X1 U9279 ( .A1(n10026), .A2(n10025), .ZN(n7641) );
  NOR2_X1 U9280 ( .A1(n7642), .A2(n7641), .ZN(n10024) );
  INV_X1 U9281 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7644) );
  INV_X1 U9282 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7643) );
  AOI22_X1 U9283 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7644), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7643), .ZN(n10023) );
  NOR2_X1 U9284 ( .A1(n10024), .A2(n10023), .ZN(n7645) );
  NOR2_X1 U9285 ( .A1(n7646), .A2(n7645), .ZN(n10022) );
  XNOR2_X1 U9286 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10021) );
  NOR2_X1 U9287 ( .A1(n10022), .A2(n10021), .ZN(n7647) );
  NOR2_X1 U9288 ( .A1(n7648), .A2(n7647), .ZN(n10020) );
  INV_X1 U9289 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7649) );
  INV_X1 U9290 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8137) );
  AOI22_X1 U9291 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n7649), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n8137), .ZN(n10019) );
  NOR2_X1 U9292 ( .A1(n10020), .A2(n10019), .ZN(n7650) );
  NOR2_X1 U9293 ( .A1(n7651), .A2(n7650), .ZN(n10018) );
  INV_X1 U9294 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7652) );
  INV_X1 U9295 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8765) );
  AOI22_X1 U9296 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7652), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8765), .ZN(n10017) );
  NOR2_X1 U9297 ( .A1(n10018), .A2(n10017), .ZN(n7653) );
  NOR2_X1 U9298 ( .A1(n7654), .A2(n7653), .ZN(n10016) );
  INV_X1 U9299 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7655) );
  INV_X1 U9300 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8796) );
  AOI22_X1 U9301 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7655), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8796), .ZN(n10015) );
  NOR2_X1 U9302 ( .A1(n10016), .A2(n10015), .ZN(n7656) );
  NOR2_X1 U9303 ( .A1(n7657), .A2(n7656), .ZN(n10014) );
  INV_X1 U9304 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7658) );
  INV_X1 U9305 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8826) );
  AOI22_X1 U9306 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7658), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n8826), .ZN(n10013) );
  NOR2_X1 U9307 ( .A1(n10014), .A2(n10013), .ZN(n7659) );
  NOR2_X1 U9308 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  NOR2_X1 U9309 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7661), .ZN(n10009) );
  AND2_X1 U9310 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7661), .ZN(n10010) );
  NOR2_X1 U9311 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10010), .ZN(n7662) );
  NOR2_X1 U9312 ( .A1(n10009), .A2(n7662), .ZN(n7664) );
  XNOR2_X1 U9313 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7663) );
  XNOR2_X1 U9314 ( .A(n7664), .B(n7663), .ZN(ADD_1068_U4) );
  INV_X1 U9315 ( .A(n7996), .ZN(n7678) );
  INV_X1 U9316 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7665) );
  AOI22_X1 U9317 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7678), .B1(n7996), .B2(
        n7665), .ZN(n7668) );
  OAI21_X1 U9318 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7669), .A(n7666), .ZN(
        n7667) );
  AOI211_X1 U9319 ( .C1(n7668), .C2(n7667), .A(n7987), .B(n9387), .ZN(n7680)
         );
  INV_X1 U9320 ( .A(n7669), .ZN(n7672) );
  INV_X1 U9321 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7671) );
  AOI21_X1 U9322 ( .B1(n7672), .B2(n7671), .A(n7670), .ZN(n7674) );
  XNOR2_X1 U9323 ( .A(n7678), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U9324 ( .A1(n7673), .A2(n7674), .ZN(n7994) );
  OAI211_X1 U9325 ( .C1(n7674), .C2(n7673), .A(n9399), .B(n7994), .ZN(n7677)
         );
  NAND2_X1 U9326 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n7870) );
  INV_X1 U9327 ( .A(n7870), .ZN(n7675) );
  AOI21_X1 U9328 ( .B1(n9804), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7675), .ZN(
        n7676) );
  OAI211_X1 U9329 ( .C1(n9403), .C2(n7678), .A(n7677), .B(n7676), .ZN(n7679)
         );
  OR2_X1 U9330 ( .A1(n7680), .A2(n7679), .ZN(P1_U3256) );
  OAI21_X1 U9331 ( .B1(n7682), .B2(n8338), .A(n7681), .ZN(n7697) );
  INV_X1 U9332 ( .A(n7697), .ZN(n7694) );
  OAI211_X1 U9333 ( .C1(n7684), .C2(n7683), .A(n7792), .B(n9609), .ZN(n7687)
         );
  NAND2_X1 U9334 ( .A1(n9335), .A2(n9435), .ZN(n7686) );
  NAND2_X1 U9335 ( .A1(n9333), .A2(n9244), .ZN(n7685) );
  AND2_X1 U9336 ( .A1(n7686), .A2(n7685), .ZN(n7926) );
  NAND2_X1 U9337 ( .A1(n7687), .A2(n7926), .ZN(n7695) );
  AOI211_X1 U9338 ( .C1(n7699), .C2(n7689), .A(n9616), .B(n7688), .ZN(n7696)
         );
  NAND2_X1 U9339 ( .A1(n7696), .A2(n9828), .ZN(n7691) );
  AOI22_X1 U9340 ( .A1(n9620), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7929), .B2(
        n9830), .ZN(n7690) );
  OAI211_X1 U9341 ( .C1(n6542), .C2(n9834), .A(n7691), .B(n7690), .ZN(n7692)
         );
  AOI21_X1 U9342 ( .B1(n9624), .B2(n7695), .A(n7692), .ZN(n7693) );
  OAI21_X1 U9343 ( .B1(n7694), .B2(n9626), .A(n7693), .ZN(P1_U3281) );
  AOI211_X1 U9344 ( .C1(n7697), .C2(n9858), .A(n7696), .B(n7695), .ZN(n7701)
         );
  AOI22_X1 U9345 ( .A1(n7699), .A2(n9640), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n9874), .ZN(n7698) );
  OAI21_X1 U9346 ( .B1(n7701), .B2(n9874), .A(n7698), .ZN(P1_U3534) );
  AOI22_X1 U9347 ( .A1(n7699), .A2(n9721), .B1(P1_REG0_REG_12__SCAN_IN), .B2(
        n9867), .ZN(n7700) );
  OAI21_X1 U9348 ( .B1(n7701), .B2(n9867), .A(n7700), .ZN(P1_U3489) );
  INV_X1 U9349 ( .A(n7702), .ZN(n7716) );
  AOI22_X1 U9350 ( .A1(n8395), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n9786), .ZN(n7703) );
  OAI21_X1 U9351 ( .B1(n7716), .B2(n9792), .A(n7703), .ZN(P1_U3335) );
  XNOR2_X1 U9352 ( .A(n7704), .B(n7705), .ZN(n9966) );
  XOR2_X1 U9353 ( .A(n7706), .B(n7705), .Z(n7707) );
  NAND2_X1 U9354 ( .A1(n7707), .A2(n9046), .ZN(n7709) );
  AOI22_X1 U9355 ( .A1(n8752), .A2(n9041), .B1(n9043), .B2(n8750), .ZN(n7708)
         );
  OAI211_X1 U9356 ( .C1(n7822), .C2(n9966), .A(n7709), .B(n7708), .ZN(n9967)
         );
  NAND2_X1 U9357 ( .A1(n9967), .A2(n9047), .ZN(n7713) );
  OAI22_X1 U9358 ( .A1(n9047), .A2(n7710), .B1(n7841), .B2(n9030), .ZN(n7711)
         );
  AOI21_X1 U9359 ( .B1(n4315), .B2(n9969), .A(n7711), .ZN(n7712) );
  OAI211_X1 U9360 ( .C1(n9966), .C2(n8531), .A(n7713), .B(n7712), .ZN(P2_U3224) );
  OAI222_X1 U9361 ( .A1(n8587), .A2(n7716), .B1(n7715), .B2(P2_U3151), .C1(
        n7714), .C2(n8590), .ZN(P2_U3275) );
  NAND2_X1 U9362 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7773), .ZN(n7720) );
  OAI21_X1 U9363 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7773), .A(n7720), .ZN(
        n7721) );
  AOI21_X1 U9364 ( .B1(n7722), .B2(n7721), .A(n7771), .ZN(n7747) );
  AOI22_X1 U9365 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7773), .B1(n7731), .B2(
        n7730), .ZN(n7728) );
  NAND2_X1 U9366 ( .A1(n7724), .A2(n7723), .ZN(n7726) );
  NAND2_X1 U9367 ( .A1(n7726), .A2(n7725), .ZN(n7727) );
  OAI21_X1 U9368 ( .B1(n7728), .B2(n7727), .A(n7774), .ZN(n7745) );
  NOR2_X1 U9369 ( .A1(n8840), .A2(n7773), .ZN(n7744) );
  MUX2_X1 U9370 ( .A(n7730), .B(n7729), .S(n8811), .Z(n7732) );
  NAND2_X1 U9371 ( .A1(n7732), .A2(n7731), .ZN(n7777) );
  INV_X1 U9372 ( .A(n7732), .ZN(n7733) );
  NAND2_X1 U9373 ( .A1(n7733), .A2(n7773), .ZN(n7734) );
  NAND2_X1 U9374 ( .A1(n7777), .A2(n7734), .ZN(n7735) );
  AOI21_X1 U9375 ( .B1(n7737), .B2(n7736), .A(n7735), .ZN(n7779) );
  AND3_X1 U9376 ( .A1(n7737), .A2(n7736), .A3(n7735), .ZN(n7738) );
  OAI21_X1 U9377 ( .B1(n7779), .B2(n7738), .A(n9892), .ZN(n7741) );
  INV_X1 U9378 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7739) );
  NOR2_X1 U9379 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7739), .ZN(n7859) );
  INV_X1 U9380 ( .A(n7859), .ZN(n7740) );
  OAI211_X1 U9381 ( .C1(n7742), .C2(n9896), .A(n7741), .B(n7740), .ZN(n7743)
         );
  AOI211_X1 U9382 ( .C1(n7745), .C2(n9904), .A(n7744), .B(n7743), .ZN(n7746)
         );
  OAI21_X1 U9383 ( .B1(n7747), .B2(n9908), .A(n7746), .ZN(P2_U3192) );
  XNOR2_X1 U9384 ( .A(n7876), .B(n7748), .ZN(n7880) );
  XNOR2_X1 U9385 ( .A(n7880), .B(n7879), .ZN(n7756) );
  OAI22_X1 U9386 ( .A1(n9311), .A2(n7750), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7749), .ZN(n7751) );
  AOI21_X1 U9387 ( .B1(n7752), .B2(n9313), .A(n7751), .ZN(n7755) );
  NAND2_X1 U9388 ( .A1(n7753), .A2(n9286), .ZN(n7754) );
  OAI211_X1 U9389 ( .C1(n7756), .C2(n9288), .A(n7755), .B(n7754), .ZN(P1_U3217) );
  XNOR2_X1 U9390 ( .A(n9964), .B(n7064), .ZN(n7831) );
  INV_X1 U9391 ( .A(n7757), .ZN(n7759) );
  AND2_X1 U9392 ( .A1(n7759), .A2(n7758), .ZN(n7829) );
  NOR2_X1 U9393 ( .A1(n4392), .A2(n7829), .ZN(n7827) );
  XOR2_X1 U9394 ( .A(n7831), .B(n7827), .Z(n7760) );
  NAND2_X1 U9395 ( .A1(n7760), .A2(n7828), .ZN(n7826) );
  OAI21_X1 U9396 ( .B1(n7760), .B2(n7828), .A(n7826), .ZN(n7769) );
  INV_X1 U9397 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7761) );
  NOR2_X1 U9398 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7761), .ZN(n9897) );
  AOI21_X1 U9399 ( .B1(n8686), .B2(n8751), .A(n9897), .ZN(n7767) );
  NAND2_X1 U9400 ( .A1(n8657), .A2(n9964), .ZN(n7766) );
  INV_X1 U9401 ( .A(n7762), .ZN(n7763) );
  NAND2_X1 U9402 ( .A1(n8734), .A2(n7763), .ZN(n7765) );
  NAND2_X1 U9403 ( .A1(n8729), .A2(n8753), .ZN(n7764) );
  NAND4_X1 U9404 ( .A1(n7767), .A2(n7766), .A3(n7765), .A4(n7764), .ZN(n7768)
         );
  AOI21_X1 U9405 ( .B1(n7769), .B2(n8714), .A(n7768), .ZN(n7770) );
  INV_X1 U9406 ( .A(n7770), .ZN(P2_U3161) );
  AOI21_X1 U9407 ( .B1(n6102), .B2(n7772), .A(n7933), .ZN(n7789) );
  NAND2_X1 U9408 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7773), .ZN(n7775) );
  XNOR2_X1 U9409 ( .A(n7937), .B(n7946), .ZN(n7776) );
  OAI21_X1 U9410 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7776), .A(n7939), .ZN(
        n7787) );
  INV_X1 U9411 ( .A(n7777), .ZN(n7778) );
  NOR2_X1 U9412 ( .A1(n7779), .A2(n7778), .ZN(n7781) );
  MUX2_X1 U9413 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8811), .Z(n7943) );
  XNOR2_X1 U9414 ( .A(n7943), .B(n7938), .ZN(n7780) );
  NOR2_X1 U9415 ( .A1(n7781), .A2(n7780), .ZN(n7944) );
  AOI21_X1 U9416 ( .B1(n7781), .B2(n7780), .A(n7944), .ZN(n7785) );
  INV_X1 U9417 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U9418 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10196), .ZN(n7967) );
  NOR2_X1 U9419 ( .A1(n9896), .A2(n7782), .ZN(n7783) );
  AOI211_X1 U9420 ( .C1(n9902), .C2(n7946), .A(n7967), .B(n7783), .ZN(n7784)
         );
  OAI21_X1 U9421 ( .B1(n7785), .B2(n9913), .A(n7784), .ZN(n7786) );
  AOI21_X1 U9422 ( .B1(n7787), .B2(n9904), .A(n7786), .ZN(n7788) );
  OAI21_X1 U9423 ( .B1(n7789), .B2(n9908), .A(n7788), .ZN(P2_U3193) );
  OAI21_X1 U9424 ( .B1(n7791), .B2(n7793), .A(n7790), .ZN(n7812) );
  INV_X1 U9425 ( .A(n7812), .ZN(n7805) );
  NAND2_X1 U9426 ( .A1(n7792), .A2(n8247), .ZN(n7794) );
  XNOR2_X1 U9427 ( .A(n7794), .B(n7793), .ZN(n7795) );
  NAND2_X1 U9428 ( .A1(n7795), .A2(n9609), .ZN(n7798) );
  NAND2_X1 U9429 ( .A1(n9332), .A2(n9244), .ZN(n7797) );
  NAND2_X1 U9430 ( .A1(n9334), .A2(n9435), .ZN(n7796) );
  AND2_X1 U9431 ( .A1(n7797), .A2(n7796), .ZN(n7871) );
  NAND2_X1 U9432 ( .A1(n7798), .A2(n7871), .ZN(n7809) );
  INV_X1 U9433 ( .A(n7914), .ZN(n7799) );
  AOI211_X1 U9434 ( .C1(n7813), .C2(n7800), .A(n9616), .B(n7799), .ZN(n7808)
         );
  NAND2_X1 U9435 ( .A1(n7808), .A2(n9828), .ZN(n7802) );
  AOI22_X1 U9436 ( .A1(n9620), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7873), .B2(
        n9830), .ZN(n7801) );
  OAI211_X1 U9437 ( .C1(n6545), .C2(n9834), .A(n7802), .B(n7801), .ZN(n7803)
         );
  AOI21_X1 U9438 ( .B1(n9624), .B2(n7809), .A(n7803), .ZN(n7804) );
  OAI21_X1 U9439 ( .B1(n7805), .B2(n9626), .A(n7804), .ZN(P1_U3280) );
  INV_X1 U9440 ( .A(n7806), .ZN(n7851) );
  AOI22_X1 U9441 ( .A1(n5719), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n9786), .ZN(n7807) );
  OAI21_X1 U9442 ( .B1(n7851), .B2(n9792), .A(n7807), .ZN(P1_U3334) );
  NOR2_X1 U9443 ( .A1(n7809), .A2(n7808), .ZN(n7816) );
  NAND2_X1 U9444 ( .A1(n7812), .A2(n9688), .ZN(n7811) );
  AOI22_X1 U9445 ( .A1(n7813), .A2(n9640), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n9874), .ZN(n7810) );
  OAI211_X1 U9446 ( .C1(n7816), .C2(n9874), .A(n7811), .B(n7810), .ZN(P1_U3535) );
  NAND2_X1 U9447 ( .A1(n7812), .A2(n9763), .ZN(n7815) );
  AOI22_X1 U9448 ( .A1(n7813), .A2(n9721), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n9867), .ZN(n7814) );
  OAI211_X1 U9449 ( .C1(n7816), .C2(n9867), .A(n7815), .B(n7814), .ZN(P1_U3492) );
  XNOR2_X1 U9450 ( .A(n7817), .B(n7818), .ZN(n9972) );
  XOR2_X1 U9451 ( .A(n7818), .B(n7896), .Z(n7819) );
  NAND2_X1 U9452 ( .A1(n7819), .A2(n9046), .ZN(n7821) );
  AOI22_X1 U9453 ( .A1(n9043), .A2(n8749), .B1(n8751), .B2(n9041), .ZN(n7820)
         );
  OAI211_X1 U9454 ( .C1(n7822), .C2(n9972), .A(n7821), .B(n7820), .ZN(n9973)
         );
  NAND2_X1 U9455 ( .A1(n9973), .A2(n9047), .ZN(n7825) );
  OAI22_X1 U9456 ( .A1(n9047), .A2(n7730), .B1(n7858), .B2(n9030), .ZN(n7823)
         );
  AOI21_X1 U9457 ( .B1(n4315), .B2(n9975), .A(n7823), .ZN(n7824) );
  OAI211_X1 U9458 ( .C1(n9972), .C2(n8531), .A(n7825), .B(n7824), .ZN(P2_U3223) );
  OAI21_X1 U9459 ( .B1(n7827), .B2(n7831), .A(n7826), .ZN(n7839) );
  XNOR2_X1 U9460 ( .A(n9969), .B(n7064), .ZN(n7852) );
  XNOR2_X1 U9461 ( .A(n7852), .B(n8751), .ZN(n7838) );
  NAND2_X1 U9462 ( .A1(n7831), .A2(n8752), .ZN(n7837) );
  NOR2_X1 U9463 ( .A1(n7829), .A2(n7828), .ZN(n7832) );
  INV_X1 U9464 ( .A(n7829), .ZN(n7830) );
  OAI22_X1 U9465 ( .A1(n7832), .A2(n7831), .B1(n8752), .B2(n7830), .ZN(n7833)
         );
  INV_X1 U9466 ( .A(n7833), .ZN(n7835) );
  INV_X1 U9467 ( .A(n7838), .ZN(n7834) );
  NAND2_X1 U9468 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  AOI211_X1 U9469 ( .C1(n7839), .C2(n7838), .A(n8724), .B(n7854), .ZN(n7848)
         );
  AOI21_X1 U9470 ( .B1(n8729), .B2(n8752), .A(n7840), .ZN(n7846) );
  NAND2_X1 U9471 ( .A1(n9969), .A2(n8657), .ZN(n7845) );
  INV_X1 U9472 ( .A(n7841), .ZN(n7842) );
  NAND2_X1 U9473 ( .A1(n8734), .A2(n7842), .ZN(n7844) );
  NAND2_X1 U9474 ( .A1(n8686), .A2(n8750), .ZN(n7843) );
  NAND4_X1 U9475 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n7843), .ZN(n7847)
         );
  OR2_X1 U9476 ( .A1(n7848), .A2(n7847), .ZN(P2_U3171) );
  OAI222_X1 U9477 ( .A1(n8587), .A2(n7851), .B1(n7850), .B2(P2_U3151), .C1(
        n7849), .C2(n8590), .ZN(P2_U3274) );
  INV_X1 U9478 ( .A(n9975), .ZN(n7865) );
  AND2_X1 U9479 ( .A1(n7852), .A2(n8751), .ZN(n7853) );
  XNOR2_X1 U9480 ( .A(n7960), .B(n8750), .ZN(n7856) );
  XOR2_X1 U9481 ( .A(n7064), .B(n9975), .Z(n7855) );
  OAI21_X1 U9482 ( .B1(n7856), .B2(n7855), .A(n7962), .ZN(n7857) );
  NAND2_X1 U9483 ( .A1(n7857), .A2(n8714), .ZN(n7864) );
  INV_X1 U9484 ( .A(n7858), .ZN(n7862) );
  AOI21_X1 U9485 ( .B1(n8729), .B2(n8751), .A(n7859), .ZN(n7860) );
  OAI21_X1 U9486 ( .B1(n8038), .B2(n8731), .A(n7860), .ZN(n7861) );
  AOI21_X1 U9487 ( .B1(n7862), .B2(n8734), .A(n7861), .ZN(n7863) );
  OAI211_X1 U9488 ( .C1(n7865), .C2(n8738), .A(n7864), .B(n7863), .ZN(P2_U3157) );
  OAI21_X1 U9489 ( .B1(n7868), .B2(n7867), .A(n7866), .ZN(n7869) );
  NAND2_X1 U9490 ( .A1(n7869), .A2(n9307), .ZN(n7875) );
  OAI21_X1 U9491 ( .B1(n9311), .B2(n7871), .A(n7870), .ZN(n7872) );
  AOI21_X1 U9492 ( .B1(n7873), .B2(n9313), .A(n7872), .ZN(n7874) );
  OAI211_X1 U9493 ( .C1(n6545), .C2(n9317), .A(n7875), .B(n7874), .ZN(P1_U3234) );
  INV_X1 U9494 ( .A(n7876), .ZN(n7878) );
  OAI22_X1 U9495 ( .A1(n7880), .A2(n7879), .B1(n7878), .B2(n7877), .ZN(n7883)
         );
  NAND2_X1 U9496 ( .A1(n4719), .A2(n7919), .ZN(n7882) );
  NOR2_X1 U9497 ( .A1(n7883), .A2(n7882), .ZN(n7922) );
  AOI21_X1 U9498 ( .B1(n7883), .B2(n7882), .A(n7922), .ZN(n7891) );
  NAND2_X1 U9499 ( .A1(n9313), .A2(n7884), .ZN(n7885) );
  OAI211_X1 U9500 ( .C1(n9311), .C2(n7887), .A(n7886), .B(n7885), .ZN(n7888)
         );
  AOI21_X1 U9501 ( .B1(n7889), .B2(n9286), .A(n7888), .ZN(n7890) );
  OAI21_X1 U9502 ( .B1(n7891), .B2(n9288), .A(n7890), .ZN(P1_U3236) );
  NAND2_X1 U9503 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  XOR2_X1 U9504 ( .A(n7963), .B(n7894), .Z(n9977) );
  OR2_X1 U9505 ( .A1(n7896), .A2(n7895), .ZN(n7978) );
  NAND2_X1 U9506 ( .A1(n7978), .A2(n7897), .ZN(n7898) );
  XNOR2_X1 U9507 ( .A(n7898), .B(n7963), .ZN(n7899) );
  OAI222_X1 U9508 ( .A1(n9010), .A2(n7900), .B1(n9012), .B2(n8035), .C1(n7899), 
        .C2(n9007), .ZN(n9978) );
  NAND2_X1 U9509 ( .A1(n9978), .A2(n9047), .ZN(n7904) );
  OAI22_X1 U9510 ( .A1(n9047), .A2(n7901), .B1(n7966), .B2(n9030), .ZN(n7902)
         );
  AOI21_X1 U9511 ( .B1(n9980), .B2(n4315), .A(n7902), .ZN(n7903) );
  OAI211_X1 U9512 ( .C1(n9977), .C2(n9055), .A(n7904), .B(n7903), .ZN(P2_U3222) );
  XNOR2_X1 U9513 ( .A(n7905), .B(n7909), .ZN(n9700) );
  INV_X1 U9514 ( .A(n7906), .ZN(n7912) );
  INV_X1 U9515 ( .A(n8003), .ZN(n7907) );
  AOI211_X1 U9516 ( .C1(n7909), .C2(n7908), .A(n9846), .B(n7907), .ZN(n7911)
         );
  AOI22_X1 U9517 ( .A1(n9435), .A2(n9333), .B1(n9331), .B2(n9244), .ZN(n9190)
         );
  INV_X1 U9518 ( .A(n9190), .ZN(n7910) );
  AOI211_X1 U9519 ( .C1(n9700), .C2(n7912), .A(n7911), .B(n7910), .ZN(n9704)
         );
  NOR2_X1 U9520 ( .A1(n9831), .A2(n7913), .ZN(n9813) );
  AOI211_X1 U9521 ( .C1(n9702), .C2(n7914), .A(n9616), .B(n8009), .ZN(n9701)
         );
  NAND2_X1 U9522 ( .A1(n9701), .A2(n9828), .ZN(n7916) );
  AOI22_X1 U9523 ( .A1(n9620), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9194), .B2(
        n9830), .ZN(n7915) );
  OAI211_X1 U9524 ( .C1(n9191), .C2(n9834), .A(n7916), .B(n7915), .ZN(n7917)
         );
  AOI21_X1 U9525 ( .B1(n9700), .B2(n9813), .A(n7917), .ZN(n7918) );
  OAI21_X1 U9526 ( .B1(n9704), .B2(n9620), .A(n7918), .ZN(P1_U3279) );
  INV_X1 U9527 ( .A(n7919), .ZN(n7921) );
  NOR3_X1 U9528 ( .A1(n7922), .A2(n7921), .A3(n7920), .ZN(n7925) );
  INV_X1 U9529 ( .A(n7923), .ZN(n7924) );
  OAI21_X1 U9530 ( .B1(n7925), .B2(n7924), .A(n9307), .ZN(n7931) );
  NOR2_X1 U9531 ( .A1(n9311), .A2(n7926), .ZN(n7927) );
  AOI211_X1 U9532 ( .C1(n9313), .C2(n7929), .A(n7928), .B(n7927), .ZN(n7930)
         );
  OAI211_X1 U9533 ( .C1(n6542), .C2(n9317), .A(n7931), .B(n7930), .ZN(P1_U3224) );
  NOR2_X1 U9534 ( .A1(n7946), .A2(n7932), .ZN(n7934) );
  AOI22_X1 U9535 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8053), .B1(n8050), .B2(
        n7947), .ZN(n7935) );
  AOI21_X1 U9536 ( .B1(n7936), .B2(n7935), .A(n8049), .ZN(n7959) );
  AOI22_X1 U9537 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8050), .B1(n8053), .B2(
        n7948), .ZN(n7942) );
  NAND2_X1 U9538 ( .A1(n7938), .A2(n7937), .ZN(n7940) );
  OAI21_X1 U9539 ( .B1(n7942), .B2(n7941), .A(n8052), .ZN(n7957) );
  INV_X1 U9540 ( .A(n7943), .ZN(n7945) );
  AOI21_X1 U9541 ( .B1(n7946), .B2(n7945), .A(n7944), .ZN(n8057) );
  MUX2_X1 U9542 ( .A(n7948), .B(n7947), .S(n8811), .Z(n7949) );
  NOR2_X1 U9543 ( .A1(n7949), .A2(n8053), .ZN(n8055) );
  NAND2_X1 U9544 ( .A1(n7949), .A2(n8053), .ZN(n8056) );
  INV_X1 U9545 ( .A(n8056), .ZN(n7950) );
  NOR2_X1 U9546 ( .A1(n8055), .A2(n7950), .ZN(n7952) );
  NAND2_X1 U9547 ( .A1(n8057), .A2(n7952), .ZN(n7951) );
  OAI211_X1 U9548 ( .C1(n8057), .C2(n7952), .A(n9892), .B(n7951), .ZN(n7955)
         );
  NOR2_X1 U9549 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7953), .ZN(n8043) );
  AOI21_X1 U9550 ( .B1(n9898), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8043), .ZN(
        n7954) );
  OAI211_X1 U9551 ( .C1(n8840), .C2(n8050), .A(n7955), .B(n7954), .ZN(n7956)
         );
  AOI21_X1 U9552 ( .B1(n7957), .B2(n9904), .A(n7956), .ZN(n7958) );
  OAI21_X1 U9553 ( .B1(n7959), .B2(n9908), .A(n7958), .ZN(P2_U3194) );
  INV_X1 U9554 ( .A(n9980), .ZN(n7973) );
  XNOR2_X1 U9555 ( .A(n7963), .B(n7064), .ZN(n7964) );
  INV_X1 U9556 ( .A(n7964), .ZN(n8037) );
  OAI211_X1 U9557 ( .C1(n7965), .C2(n8037), .A(n8714), .B(n8040), .ZN(n7972)
         );
  INV_X1 U9558 ( .A(n7966), .ZN(n7970) );
  AOI21_X1 U9559 ( .B1(n8729), .B2(n8750), .A(n7967), .ZN(n7968) );
  OAI21_X1 U9560 ( .B1(n8035), .B2(n8731), .A(n7968), .ZN(n7969) );
  AOI21_X1 U9561 ( .B1(n7970), .B2(n8734), .A(n7969), .ZN(n7971) );
  OAI211_X1 U9562 ( .C1(n7973), .C2(n8738), .A(n7972), .B(n7971), .ZN(P2_U3176) );
  INV_X1 U9563 ( .A(n7974), .ZN(n8017) );
  AOI22_X1 U9564 ( .A1(n8464), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n9786), .ZN(n7975) );
  OAI21_X1 U9565 ( .B1(n8017), .B2(n9792), .A(n7975), .ZN(P1_U3333) );
  XNOR2_X1 U9566 ( .A(n7976), .B(n7981), .ZN(n9983) );
  NAND2_X1 U9567 ( .A1(n7978), .A2(n7977), .ZN(n7980) );
  AND2_X1 U9568 ( .A1(n7980), .A2(n7979), .ZN(n7982) );
  XNOR2_X1 U9569 ( .A(n7982), .B(n7981), .ZN(n7983) );
  OAI222_X1 U9570 ( .A1(n9012), .A2(n8532), .B1(n9010), .B2(n8038), .C1(n7983), 
        .C2(n9007), .ZN(n9984) );
  NAND2_X1 U9571 ( .A1(n9984), .A2(n9047), .ZN(n7986) );
  OAI22_X1 U9572 ( .A1(n9047), .A2(n7948), .B1(n8045), .B2(n9030), .ZN(n7984)
         );
  AOI21_X1 U9573 ( .B1(n9986), .B2(n4315), .A(n7984), .ZN(n7985) );
  OAI211_X1 U9574 ( .C1(n9055), .C2(n9983), .A(n7986), .B(n7985), .ZN(P2_U3221) );
  INV_X1 U9575 ( .A(n7997), .ZN(n8071) );
  NOR2_X1 U9576 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9189), .ZN(n7993) );
  NAND2_X1 U9577 ( .A1(n7997), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8067) );
  OR2_X1 U9578 ( .A1(n7997), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U9579 ( .A1(n8067), .A2(n7988), .ZN(n7990) );
  INV_X1 U9580 ( .A(n8068), .ZN(n7989) );
  AOI211_X1 U9581 ( .C1(n7991), .C2(n7990), .A(n7989), .B(n9387), .ZN(n7992)
         );
  AOI211_X1 U9582 ( .C1(n9804), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7993), .B(
        n7992), .ZN(n8000) );
  INV_X1 U9583 ( .A(n7994), .ZN(n7995) );
  AOI21_X1 U9584 ( .B1(n7996), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7995), .ZN(
        n8073) );
  XNOR2_X1 U9585 ( .A(n7997), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n8074) );
  XOR2_X1 U9586 ( .A(n8073), .B(n8074), .Z(n7998) );
  NAND2_X1 U9587 ( .A1(n9399), .A2(n7998), .ZN(n7999) );
  OAI211_X1 U9588 ( .C1(n9403), .C2(n8071), .A(n8000), .B(n7999), .ZN(P1_U3257) );
  XNOR2_X1 U9589 ( .A(n8001), .B(n8002), .ZN(n8025) );
  AOI22_X1 U9590 ( .A1(n8012), .A2(n9640), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9874), .ZN(n8011) );
  NAND2_X1 U9591 ( .A1(n8003), .A2(n8252), .ZN(n8004) );
  XNOR2_X1 U9592 ( .A(n8004), .B(n8345), .ZN(n8008) );
  OR2_X1 U9593 ( .A1(n9242), .A2(n9409), .ZN(n8006) );
  NAND2_X1 U9594 ( .A1(n9332), .A2(n9435), .ZN(n8005) );
  AND2_X1 U9595 ( .A1(n8006), .A2(n8005), .ZN(n9310) );
  INV_X1 U9596 ( .A(n9310), .ZN(n8007) );
  AOI21_X1 U9597 ( .B1(n8008), .B2(n9609), .A(n8007), .ZN(n8033) );
  OAI211_X1 U9598 ( .C1(n9318), .C2(n8009), .A(n9584), .B(n8168), .ZN(n8027)
         );
  NAND2_X1 U9599 ( .A1(n8033), .A2(n8027), .ZN(n8013) );
  NAND2_X1 U9600 ( .A1(n8013), .A2(n9876), .ZN(n8010) );
  OAI211_X1 U9601 ( .C1(n8025), .C2(n9687), .A(n8011), .B(n8010), .ZN(P1_U3537) );
  AOI22_X1 U9602 ( .A1(n8012), .A2(n9721), .B1(P1_REG0_REG_15__SCAN_IN), .B2(
        n9867), .ZN(n8015) );
  NAND2_X1 U9603 ( .A1(n8013), .A2(n9869), .ZN(n8014) );
  OAI211_X1 U9604 ( .C1(n8025), .C2(n9761), .A(n8015), .B(n8014), .ZN(P1_U3498) );
  OAI222_X1 U9605 ( .A1(n8590), .A2(n8018), .B1(n8587), .B2(n8017), .C1(
        P2_U3151), .C2(n8016), .ZN(P2_U3273) );
  INV_X1 U9606 ( .A(n5886), .ZN(n8020) );
  NAND2_X1 U9607 ( .A1(n9790), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8019) );
  OAI211_X1 U9608 ( .C1(n8020), .C2(n9792), .A(n8467), .B(n8019), .ZN(P1_U3332) );
  NAND2_X1 U9609 ( .A1(n5886), .A2(n8021), .ZN(n8023) );
  OAI211_X1 U9610 ( .C1(n8024), .C2(n8590), .A(n8023), .B(n8022), .ZN(P2_U3272) );
  INV_X1 U9611 ( .A(n8025), .ZN(n8026) );
  NAND2_X1 U9612 ( .A1(n8026), .A2(n9838), .ZN(n8032) );
  INV_X1 U9613 ( .A(n8027), .ZN(n8030) );
  AOI22_X1 U9614 ( .A1(n9620), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9314), .B2(
        n9830), .ZN(n8028) );
  OAI21_X1 U9615 ( .B1(n9318), .B2(n9834), .A(n8028), .ZN(n8029) );
  AOI21_X1 U9616 ( .B1(n8030), .B2(n9828), .A(n8029), .ZN(n8031) );
  OAI211_X1 U9617 ( .C1(n9831), .C2(n8033), .A(n8032), .B(n8031), .ZN(P1_U3278) );
  XNOR2_X1 U9618 ( .A(n9986), .B(n8564), .ZN(n8036) );
  INV_X1 U9619 ( .A(n8036), .ZN(n8034) );
  NAND2_X1 U9620 ( .A1(n8034), .A2(n8748), .ZN(n8085) );
  NAND2_X1 U9621 ( .A1(n8036), .A2(n8035), .ZN(n8083) );
  NAND2_X1 U9622 ( .A1(n8085), .A2(n8083), .ZN(n8041) );
  XOR2_X1 U9623 ( .A(n8041), .B(n8084), .Z(n8048) );
  NOR2_X1 U9624 ( .A1(n8731), .A2(n8532), .ZN(n8042) );
  AOI211_X1 U9625 ( .C1(n8729), .C2(n8749), .A(n8043), .B(n8042), .ZN(n8044)
         );
  OAI21_X1 U9626 ( .B1(n8045), .B2(n8664), .A(n8044), .ZN(n8046) );
  AOI21_X1 U9627 ( .B1(n9986), .B2(n8657), .A(n8046), .ZN(n8047) );
  OAI21_X1 U9628 ( .B1(n8048), .B2(n8724), .A(n8047), .ZN(P2_U3164) );
  AOI21_X1 U9629 ( .B1(n8107), .B2(n8051), .A(n8125), .ZN(n8066) );
  OAI21_X1 U9630 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8054), .A(n8120), .ZN(
        n8064) );
  MUX2_X1 U9631 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8811), .Z(n8130) );
  XNOR2_X1 U9632 ( .A(n8130), .B(n8124), .ZN(n8059) );
  AOI21_X1 U9633 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8058) );
  NAND2_X1 U9634 ( .A1(n8058), .A2(n8059), .ZN(n8131) );
  OAI21_X1 U9635 ( .B1(n8059), .B2(n8058), .A(n8131), .ZN(n8060) );
  AND2_X1 U9636 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8089) );
  AOI21_X1 U9637 ( .B1(n8060), .B2(n9892), .A(n8089), .ZN(n8062) );
  NAND2_X1 U9638 ( .A1(n9898), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8061) );
  OAI211_X1 U9639 ( .C1(n8840), .C2(n8129), .A(n8062), .B(n8061), .ZN(n8063)
         );
  AOI21_X1 U9640 ( .B1(n8064), .B2(n9904), .A(n8063), .ZN(n8065) );
  OAI21_X1 U9641 ( .B1(n8066), .B2(n9908), .A(n8065), .ZN(P2_U3195) );
  INV_X1 U9642 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8070) );
  INV_X1 U9643 ( .A(n8481), .ZN(n8468) );
  XNOR2_X1 U9644 ( .A(n8469), .B(n8468), .ZN(n8069) );
  NOR2_X1 U9645 ( .A1(n8070), .A2(n8069), .ZN(n8470) );
  AOI211_X1 U9646 ( .C1(n8070), .C2(n8069), .A(n8470), .B(n9387), .ZN(n8080)
         );
  INV_X1 U9647 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8072) );
  OAI22_X1 U9648 ( .A1(n8074), .A2(n8073), .B1(n8072), .B2(n8071), .ZN(n8480)
         );
  XNOR2_X1 U9649 ( .A(n8480), .B(n8468), .ZN(n8075) );
  NAND2_X1 U9650 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n8075), .ZN(n8482) );
  OAI211_X1 U9651 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n8075), .A(n9399), .B(
        n8482), .ZN(n8078) );
  NOR2_X1 U9652 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9309), .ZN(n8076) );
  AOI21_X1 U9653 ( .B1(n9804), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n8076), .ZN(
        n8077) );
  OAI211_X1 U9654 ( .C1(n9403), .C2(n8468), .A(n8078), .B(n8077), .ZN(n8079)
         );
  OR2_X1 U9655 ( .A1(n8080), .A2(n8079), .ZN(P1_U3258) );
  INV_X1 U9656 ( .A(n8081), .ZN(n8096) );
  AOI22_X1 U9657 ( .A1(n5700), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n9786), .ZN(n8082) );
  OAI21_X1 U9658 ( .B1(n8096), .B2(n9792), .A(n8082), .ZN(P1_U3331) );
  NAND2_X1 U9659 ( .A1(n8084), .A2(n8083), .ZN(n8086) );
  NAND2_X1 U9660 ( .A1(n8086), .A2(n8085), .ZN(n8536) );
  XNOR2_X1 U9661 ( .A(n8111), .B(n8564), .ZN(n8533) );
  XNOR2_X1 U9662 ( .A(n8533), .B(n8747), .ZN(n8087) );
  XNOR2_X1 U9663 ( .A(n8536), .B(n8087), .ZN(n8093) );
  NOR2_X1 U9664 ( .A1(n8731), .A2(n8539), .ZN(n8088) );
  AOI211_X1 U9665 ( .C1(n8729), .C2(n8748), .A(n8089), .B(n8088), .ZN(n8090)
         );
  OAI21_X1 U9666 ( .B1(n8112), .B2(n8664), .A(n8090), .ZN(n8091) );
  AOI21_X1 U9667 ( .B1(n8111), .B2(n8657), .A(n8091), .ZN(n8092) );
  OAI21_X1 U9668 ( .B1(n8093), .B2(n8724), .A(n8092), .ZN(P2_U3174) );
  OAI222_X1 U9669 ( .A1(n8587), .A2(n8096), .B1(P2_U3151), .B2(n8095), .C1(
        n8094), .C2(n8590), .ZN(P2_U3271) );
  XNOR2_X1 U9670 ( .A(n8097), .B(n8101), .ZN(n8118) );
  INV_X1 U9671 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8104) );
  AND2_X1 U9672 ( .A1(n8748), .A2(n9041), .ZN(n8103) );
  INV_X1 U9673 ( .A(n8098), .ZN(n8099) );
  AOI211_X1 U9674 ( .C1(n8101), .C2(n8100), .A(n9007), .B(n8099), .ZN(n8102)
         );
  AOI211_X1 U9675 ( .C1(n9043), .C2(n8746), .A(n8103), .B(n8102), .ZN(n8110)
         );
  MUX2_X1 U9676 ( .A(n8104), .B(n8110), .S(n9988), .Z(n8106) );
  NAND2_X1 U9677 ( .A1(n8111), .A2(n6505), .ZN(n8105) );
  OAI211_X1 U9678 ( .C1(n8118), .C2(n9171), .A(n8106), .B(n8105), .ZN(P2_U3429) );
  MUX2_X1 U9679 ( .A(n8107), .B(n8110), .S(n10005), .Z(n8109) );
  NAND2_X1 U9680 ( .A1(n8111), .A2(n9105), .ZN(n8108) );
  OAI211_X1 U9681 ( .C1(n8118), .C2(n9108), .A(n8109), .B(n8108), .ZN(P2_U3472) );
  INV_X1 U9682 ( .A(n8110), .ZN(n8115) );
  INV_X1 U9683 ( .A(n8111), .ZN(n8113) );
  OAI22_X1 U9684 ( .A1(n8113), .A2(n8937), .B1(n8112), .B2(n9030), .ZN(n8114)
         );
  OAI21_X1 U9685 ( .B1(n8115), .B2(n8114), .A(n9047), .ZN(n8117) );
  NAND2_X1 U9686 ( .A1(n9037), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8116) );
  OAI211_X1 U9687 ( .C1(n8118), .C2(n9055), .A(n8117), .B(n8116), .ZN(P2_U3220) );
  NAND2_X1 U9688 ( .A1(n8129), .A2(n8119), .ZN(n8121) );
  NAND2_X1 U9689 ( .A1(n8139), .A2(n5932), .ZN(n8762) );
  OAI21_X1 U9690 ( .B1(n8139), .B2(n5932), .A(n8762), .ZN(n8122) );
  XNOR2_X1 U9691 ( .A(n8761), .B(n8122), .ZN(n8142) );
  NOR2_X1 U9692 ( .A1(n8124), .A2(n8123), .ZN(n8126) );
  XNOR2_X1 U9693 ( .A(n8139), .B(n8156), .ZN(n8127) );
  AOI21_X1 U9694 ( .B1(n4400), .B2(n8127), .A(n8766), .ZN(n8128) );
  OR2_X1 U9695 ( .A1(n8128), .A2(n9908), .ZN(n8141) );
  MUX2_X1 U9696 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8811), .Z(n8770) );
  XNOR2_X1 U9697 ( .A(n8139), .B(n8770), .ZN(n8134) );
  OR2_X1 U9698 ( .A1(n8130), .A2(n8129), .ZN(n8132) );
  NAND2_X1 U9699 ( .A1(n8132), .A2(n8131), .ZN(n8133) );
  NAND2_X1 U9700 ( .A1(n8134), .A2(n8133), .ZN(n8771) );
  OAI21_X1 U9701 ( .B1(n8134), .B2(n8133), .A(n8771), .ZN(n8135) );
  NAND2_X1 U9702 ( .A1(n8135), .A2(n9892), .ZN(n8136) );
  NAND2_X1 U9703 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8605) );
  OAI211_X1 U9704 ( .C1(n9896), .C2(n8137), .A(n8136), .B(n8605), .ZN(n8138)
         );
  AOI21_X1 U9705 ( .B1(n9902), .B2(n8139), .A(n8138), .ZN(n8140) );
  OAI211_X1 U9706 ( .C1(n8142), .C2(n8877), .A(n8141), .B(n8140), .ZN(P2_U3196) );
  XOR2_X1 U9707 ( .A(n8143), .B(n8147), .Z(n8144) );
  AOI222_X1 U9708 ( .A1(n9046), .A2(n8144), .B1(n9042), .B2(n9043), .C1(n8747), 
        .C2(n9041), .ZN(n8155) );
  INV_X1 U9709 ( .A(n8155), .ZN(n8146) );
  OAI22_X1 U9710 ( .A1(n8612), .A2(n8937), .B1(n8607), .B2(n9030), .ZN(n8145)
         );
  OAI21_X1 U9711 ( .B1(n8146), .B2(n8145), .A(n9047), .ZN(n8150) );
  XNOR2_X1 U9712 ( .A(n8148), .B(n8147), .ZN(n8158) );
  AOI22_X1 U9713 ( .A1(n8158), .A2(n9035), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9037), .ZN(n8149) );
  NAND2_X1 U9714 ( .A1(n8150), .A2(n8149), .ZN(P2_U3219) );
  INV_X1 U9715 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8151) );
  MUX2_X1 U9716 ( .A(n8151), .B(n8155), .S(n9988), .Z(n8154) );
  INV_X1 U9717 ( .A(n9171), .ZN(n8152) );
  AOI22_X1 U9718 ( .A1(n8158), .A2(n8152), .B1(n6505), .B2(n8537), .ZN(n8153)
         );
  NAND2_X1 U9719 ( .A1(n8154), .A2(n8153), .ZN(P2_U3432) );
  MUX2_X1 U9720 ( .A(n8156), .B(n8155), .S(n10005), .Z(n8160) );
  INV_X1 U9721 ( .A(n9108), .ZN(n8157) );
  AOI22_X1 U9722 ( .A1(n8158), .A2(n8157), .B1(n9105), .B2(n8537), .ZN(n8159)
         );
  NAND2_X1 U9723 ( .A1(n8160), .A2(n8159), .ZN(P2_U3473) );
  XNOR2_X1 U9724 ( .A(n8161), .B(n8344), .ZN(n9696) );
  INV_X1 U9725 ( .A(n9696), .ZN(n8173) );
  XNOR2_X1 U9726 ( .A(n8162), .B(n8344), .ZN(n8163) );
  NAND2_X1 U9727 ( .A1(n8163), .A2(n9609), .ZN(n8166) );
  OAI22_X1 U9728 ( .A1(n9282), .A2(n9409), .B1(n8164), .B2(n9281), .ZN(n9235)
         );
  INV_X1 U9729 ( .A(n9235), .ZN(n8165) );
  NAND2_X1 U9730 ( .A1(n8166), .A2(n8165), .ZN(n9694) );
  INV_X1 U9731 ( .A(n9617), .ZN(n8167) );
  AOI211_X1 U9732 ( .C1(n6548), .C2(n8168), .A(n9616), .B(n8167), .ZN(n9695)
         );
  NAND2_X1 U9733 ( .A1(n9695), .A2(n9828), .ZN(n8170) );
  AOI22_X1 U9734 ( .A1(n9620), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9232), .B2(
        n9830), .ZN(n8169) );
  OAI211_X1 U9735 ( .C1(n9774), .C2(n9834), .A(n8170), .B(n8169), .ZN(n8171)
         );
  AOI21_X1 U9736 ( .B1(n9624), .B2(n9694), .A(n8171), .ZN(n8172) );
  OAI21_X1 U9737 ( .B1(n8173), .B2(n9626), .A(n8172), .ZN(P1_U3277) );
  INV_X1 U9738 ( .A(n8174), .ZN(n8179) );
  AOI22_X1 U9739 ( .A1(n8175), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9786), .ZN(n8176) );
  OAI21_X1 U9740 ( .B1(n8179), .B2(n9792), .A(n8176), .ZN(P1_U3330) );
  OAI222_X1 U9741 ( .A1(n8587), .A2(n8179), .B1(P2_U3151), .B2(n8178), .C1(
        n8177), .C2(n8590), .ZN(P2_U3270) );
  XNOR2_X1 U9742 ( .A(n8181), .B(n8180), .ZN(n8195) );
  INV_X1 U9743 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8185) );
  XNOR2_X1 U9744 ( .A(n8182), .B(n8183), .ZN(n8184) );
  AOI222_X1 U9745 ( .A1(n9046), .A2(n8184), .B1(n9023), .B2(n9043), .C1(n8746), 
        .C2(n9041), .ZN(n8190) );
  MUX2_X1 U9746 ( .A(n8185), .B(n8190), .S(n9988), .Z(n8187) );
  NAND2_X1 U9747 ( .A1(n8542), .A2(n6505), .ZN(n8186) );
  OAI211_X1 U9748 ( .C1(n8195), .C2(n9171), .A(n8187), .B(n8186), .ZN(P2_U3435) );
  MUX2_X1 U9749 ( .A(n8767), .B(n8190), .S(n10005), .Z(n8189) );
  NAND2_X1 U9750 ( .A1(n8542), .A2(n9105), .ZN(n8188) );
  OAI211_X1 U9751 ( .C1(n9108), .C2(n8195), .A(n8189), .B(n8188), .ZN(P2_U3474) );
  MUX2_X1 U9752 ( .A(n8191), .B(n8190), .S(n9047), .Z(n8194) );
  INV_X1 U9753 ( .A(n8192), .ZN(n8735) );
  AOI22_X1 U9754 ( .A1(n8542), .A2(n4315), .B1(n9051), .B2(n8735), .ZN(n8193)
         );
  OAI211_X1 U9755 ( .C1(n8195), .C2(n9055), .A(n8194), .B(n8193), .ZN(P2_U3218) );
  INV_X1 U9756 ( .A(n8196), .ZN(n8199) );
  AOI22_X1 U9757 ( .A1(n8197), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9786), .ZN(n8198) );
  OAI21_X1 U9758 ( .B1(n8199), .B2(n9792), .A(n8198), .ZN(P1_U3329) );
  OAI222_X1 U9759 ( .A1(n8590), .A2(n8201), .B1(P2_U3151), .B2(n8200), .C1(
        n8587), .C2(n8199), .ZN(P2_U3269) );
  INV_X1 U9760 ( .A(n8202), .ZN(n8499) );
  AOI22_X1 U9761 ( .A1(n8203), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n9786), .ZN(n8204) );
  OAI21_X1 U9762 ( .B1(n8499), .B2(n9792), .A(n8204), .ZN(P1_U3328) );
  INV_X1 U9763 ( .A(n8205), .ZN(n8586) );
  AOI22_X1 U9764 ( .A1(n8206), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9786), .ZN(n8207) );
  OAI21_X1 U9765 ( .B1(n8586), .B2(n9792), .A(n8207), .ZN(P1_U3327) );
  NAND2_X1 U9766 ( .A1(n8436), .A2(n8360), .ZN(n8208) );
  NAND2_X1 U9767 ( .A1(n8283), .A2(n8273), .ZN(n8363) );
  MUX2_X1 U9768 ( .A(n8208), .B(n8363), .S(n8458), .Z(n8285) );
  NAND2_X1 U9769 ( .A1(n8267), .A2(n8209), .ZN(n8426) );
  NAND2_X1 U9770 ( .A1(n8247), .A2(n8210), .ZN(n8239) );
  OR2_X1 U9771 ( .A1(n8239), .A2(n8211), .ZN(n8416) );
  INV_X1 U9772 ( .A(n8416), .ZN(n8242) );
  OAI21_X1 U9773 ( .B1(n8213), .B2(n8212), .A(n8332), .ZN(n8214) );
  NAND2_X1 U9774 ( .A1(n8214), .A2(n8223), .ZN(n8226) );
  NAND2_X1 U9775 ( .A1(n8215), .A2(n8404), .ZN(n8217) );
  NAND3_X1 U9776 ( .A1(n8217), .A2(n8216), .A3(n8332), .ZN(n8219) );
  NAND2_X1 U9777 ( .A1(n8219), .A2(n8218), .ZN(n8224) );
  NAND2_X1 U9778 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  AOI21_X1 U9779 ( .B1(n8224), .B2(n8223), .A(n8222), .ZN(n8225) );
  MUX2_X1 U9780 ( .A(n8226), .B(n8225), .S(n8458), .Z(n8230) );
  NAND2_X1 U9781 ( .A1(n8227), .A2(n8333), .ZN(n8228) );
  INV_X1 U9782 ( .A(n8458), .ZN(n8319) );
  NAND2_X1 U9783 ( .A1(n8228), .A2(n8319), .ZN(n8229) );
  NAND2_X1 U9784 ( .A1(n8230), .A2(n8229), .ZN(n8234) );
  MUX2_X1 U9785 ( .A(n8232), .B(n8231), .S(n8319), .Z(n8233) );
  NAND2_X1 U9786 ( .A1(n8234), .A2(n8233), .ZN(n8245) );
  NAND2_X1 U9787 ( .A1(n8245), .A2(n8235), .ZN(n8241) );
  AND2_X1 U9788 ( .A1(n8237), .A2(n8236), .ZN(n8238) );
  OR2_X1 U9789 ( .A1(n8239), .A2(n8238), .ZN(n8240) );
  NAND2_X1 U9790 ( .A1(n8240), .A2(n8249), .ZN(n8413) );
  AOI21_X1 U9791 ( .B1(n8242), .B2(n8241), .A(n8413), .ZN(n8250) );
  NAND2_X1 U9792 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  NAND2_X1 U9793 ( .A1(n8258), .A2(n8414), .ZN(n8255) );
  AND2_X1 U9794 ( .A1(n8252), .A2(n8251), .ZN(n8419) );
  NAND2_X1 U9795 ( .A1(n9702), .A2(n8253), .ZN(n8259) );
  INV_X1 U9796 ( .A(n8259), .ZN(n8254) );
  AOI21_X1 U9797 ( .B1(n8255), .B2(n8419), .A(n8254), .ZN(n8256) );
  NOR2_X1 U9798 ( .A1(n8426), .A2(n8256), .ZN(n8264) );
  AND2_X1 U9799 ( .A1(n8265), .A2(n8259), .ZN(n8397) );
  NAND3_X1 U9800 ( .A1(n8260), .A2(n8397), .A3(n8424), .ZN(n8261) );
  NAND3_X1 U9801 ( .A1(n8262), .A2(n8267), .A3(n8261), .ZN(n8263) );
  INV_X1 U9802 ( .A(n8265), .ZN(n8266) );
  NAND2_X1 U9803 ( .A1(n8267), .A2(n8266), .ZN(n8268) );
  NAND2_X1 U9804 ( .A1(n8268), .A2(n8424), .ZN(n8269) );
  AND2_X1 U9805 ( .A1(n8277), .A2(n8271), .ZN(n8427) );
  AND2_X1 U9806 ( .A1(n8281), .A2(n8276), .ZN(n8431) );
  NAND2_X1 U9807 ( .A1(n8272), .A2(n8431), .ZN(n8274) );
  AND2_X1 U9808 ( .A1(n8276), .A2(n8275), .ZN(n8430) );
  NAND2_X1 U9809 ( .A1(n8432), .A2(n8277), .ZN(n8278) );
  AOI21_X1 U9810 ( .B1(n8360), .B2(n8281), .A(n8319), .ZN(n8282) );
  MUX2_X1 U9811 ( .A(n8436), .B(n8283), .S(n8319), .Z(n8284) );
  OR2_X1 U9812 ( .A1(n9540), .A2(n9212), .ZN(n8286) );
  NAND2_X1 U9813 ( .A1(n8292), .A2(n8286), .ZN(n8355) );
  NAND2_X1 U9814 ( .A1(n8355), .A2(n8458), .ZN(n8287) );
  NAND2_X1 U9815 ( .A1(n8288), .A2(n9505), .ZN(n8291) );
  NAND2_X1 U9816 ( .A1(n9505), .A2(n8289), .ZN(n8364) );
  NAND2_X1 U9817 ( .A1(n8364), .A2(n8319), .ZN(n8290) );
  OR2_X1 U9818 ( .A1(n8292), .A2(n8458), .ZN(n8293) );
  MUX2_X1 U9819 ( .A(n8366), .B(n9479), .S(n8458), .Z(n8294) );
  NAND2_X1 U9820 ( .A1(n8375), .A2(n8370), .ZN(n8299) );
  AOI21_X1 U9821 ( .B1(n8295), .B2(n8359), .A(n8299), .ZN(n8296) );
  NAND2_X1 U9822 ( .A1(n9429), .A2(n8373), .ZN(n8439) );
  NOR2_X1 U9823 ( .A1(n8296), .A2(n8439), .ZN(n8297) );
  NAND2_X1 U9824 ( .A1(n9431), .A2(n8303), .ZN(n8379) );
  NAND2_X1 U9825 ( .A1(n8298), .A2(n8359), .ZN(n8302) );
  INV_X1 U9826 ( .A(n8299), .ZN(n8301) );
  INV_X1 U9827 ( .A(n8373), .ZN(n8300) );
  AOI21_X1 U9828 ( .B1(n8302), .B2(n8301), .A(n8300), .ZN(n8305) );
  INV_X1 U9829 ( .A(n8303), .ZN(n8304) );
  OAI211_X1 U9830 ( .C1(n8305), .C2(n8304), .A(n8353), .B(n9429), .ZN(n8306)
         );
  NAND2_X1 U9831 ( .A1(n9182), .A2(n8313), .ZN(n8308) );
  NAND2_X1 U9832 ( .A1(n4326), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U9833 ( .A1(n8308), .A2(n8307), .ZN(n9404) );
  NAND2_X1 U9834 ( .A1(n9404), .A2(n8309), .ZN(n8384) );
  NAND2_X1 U9835 ( .A1(n8354), .A2(n8384), .ZN(n9432) );
  NAND2_X1 U9836 ( .A1(n8588), .A2(n8313), .ZN(n8312) );
  NAND2_X1 U9837 ( .A1(n4326), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U9838 ( .A1(n9175), .A2(n8313), .ZN(n8315) );
  NAND2_X1 U9839 ( .A1(n4326), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8314) );
  INV_X1 U9840 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U9841 ( .A1(n4323), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U9842 ( .A1(n4324), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8316) );
  OAI211_X1 U9843 ( .C1(n8318), .C2(n9712), .A(n8317), .B(n8316), .ZN(n9433)
         );
  OAI211_X1 U9844 ( .C1(n9414), .C2(n8319), .A(n8320), .B(n9433), .ZN(n8322)
         );
  AOI22_X1 U9845 ( .A1(n9414), .A2(n8319), .B1(n9410), .B2(n9433), .ZN(n8321)
         );
  AND2_X1 U9846 ( .A1(n8320), .A2(n8382), .ZN(n8388) );
  OR2_X1 U9847 ( .A1(n5462), .A2(n5719), .ZN(n8324) );
  INV_X1 U9848 ( .A(n9433), .ZN(n8351) );
  NOR2_X1 U9849 ( .A1(n9414), .A2(n8351), .ZN(n8386) );
  NOR2_X1 U9850 ( .A1(n8388), .A2(n8386), .ZN(n8445) );
  INV_X1 U9851 ( .A(n9528), .ZN(n9532) );
  INV_X1 U9852 ( .A(n9612), .ZN(n8346) );
  NAND3_X1 U9853 ( .A1(n9844), .A2(n8398), .A3(n8325), .ZN(n8329) );
  NAND2_X1 U9854 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  NOR4_X1 U9855 ( .A1(n8331), .A2(n8330), .A3(n8329), .A4(n8328), .ZN(n8334)
         );
  NAND4_X1 U9856 ( .A1(n8335), .A2(n8334), .A3(n8333), .A4(n8332), .ZN(n8336)
         );
  NOR4_X1 U9857 ( .A1(n8338), .A2(n8337), .A3(n8408), .A4(n8336), .ZN(n8340)
         );
  NAND4_X1 U9858 ( .A1(n8342), .A2(n8341), .A3(n8340), .A4(n8339), .ZN(n8343)
         );
  NOR4_X1 U9859 ( .A1(n8346), .A2(n8345), .A3(n8344), .A4(n8343), .ZN(n8347)
         );
  NAND4_X1 U9860 ( .A1(n9568), .A2(n9594), .A3(n9579), .A4(n8347), .ZN(n8348)
         );
  NOR4_X1 U9861 ( .A1(n9520), .A2(n9532), .A3(n9545), .A4(n8348), .ZN(n8349)
         );
  NAND4_X1 U9862 ( .A1(n9470), .A2(n9484), .A3(n9504), .A4(n8349), .ZN(n8350)
         );
  NOR4_X1 U9863 ( .A1(n9432), .A2(n9428), .A3(n9451), .A4(n8350), .ZN(n8352)
         );
  NAND2_X1 U9864 ( .A1(n9414), .A2(n8351), .ZN(n8385) );
  NAND4_X1 U9865 ( .A1(n8445), .A2(n8352), .A3(n8448), .A4(n8385), .ZN(n8393)
         );
  AND2_X1 U9866 ( .A1(n8354), .A2(n8353), .ZN(n8440) );
  INV_X1 U9867 ( .A(n9429), .ZN(n8381) );
  NAND2_X1 U9868 ( .A1(n8355), .A2(n9505), .ZN(n8356) );
  NAND2_X1 U9869 ( .A1(n8356), .A2(n9479), .ZN(n8357) );
  NAND2_X1 U9870 ( .A1(n8357), .A2(n8366), .ZN(n8358) );
  NAND2_X1 U9871 ( .A1(n8359), .A2(n8358), .ZN(n8372) );
  INV_X1 U9872 ( .A(n8360), .ZN(n8361) );
  NOR2_X1 U9873 ( .A1(n8372), .A2(n8361), .ZN(n8396) );
  NAND4_X1 U9874 ( .A1(n8396), .A2(n8373), .A3(n8436), .A4(n8362), .ZN(n8380)
         );
  INV_X1 U9875 ( .A(n8436), .ZN(n8368) );
  INV_X1 U9876 ( .A(n8363), .ZN(n8367) );
  INV_X1 U9877 ( .A(n8364), .ZN(n8365) );
  OAI211_X1 U9878 ( .C1(n8368), .C2(n8367), .A(n8366), .B(n8365), .ZN(n8369)
         );
  INV_X1 U9879 ( .A(n8369), .ZN(n8371) );
  OAI21_X1 U9880 ( .B1(n8372), .B2(n8371), .A(n8370), .ZN(n8374) );
  NAND2_X1 U9881 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  NAND2_X1 U9882 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  AND2_X1 U9883 ( .A1(n8377), .A2(n9429), .ZN(n8378) );
  NOR2_X1 U9884 ( .A1(n8379), .A2(n8378), .ZN(n8443) );
  OAI21_X1 U9885 ( .B1(n8381), .B2(n8380), .A(n8443), .ZN(n8383) );
  AOI22_X1 U9886 ( .A1(n8440), .A2(n8383), .B1(n8382), .B2(n9414), .ZN(n8387)
         );
  AND2_X1 U9887 ( .A1(n8385), .A2(n8384), .ZN(n8444) );
  AOI22_X1 U9888 ( .A1(n8387), .A2(n8444), .B1(n8386), .B2(n9410), .ZN(n8390)
         );
  INV_X1 U9889 ( .A(n8448), .ZN(n8456) );
  INV_X1 U9890 ( .A(n8388), .ZN(n8457) );
  OAI211_X1 U9891 ( .C1(n8390), .C2(n8456), .A(n8389), .B(n8457), .ZN(n8391)
         );
  AOI21_X1 U9892 ( .B1(n8393), .B2(n8391), .A(n8455), .ZN(n8392) );
  NOR2_X1 U9893 ( .A1(n5462), .A2(n8395), .ZN(n8452) );
  INV_X1 U9894 ( .A(n8396), .ZN(n8438) );
  INV_X1 U9895 ( .A(n8397), .ZN(n8423) );
  AOI21_X1 U9896 ( .B1(n6526), .B2(n6525), .A(n8398), .ZN(n8402) );
  AND4_X1 U9897 ( .A1(n8402), .A2(n8401), .A3(n8400), .A4(n8399), .ZN(n8405)
         );
  NAND3_X1 U9898 ( .A1(n8405), .A2(n8404), .A3(n8403), .ZN(n8406) );
  NAND2_X1 U9899 ( .A1(n8407), .A2(n8406), .ZN(n8412) );
  INV_X1 U9900 ( .A(n8408), .ZN(n8411) );
  INV_X1 U9901 ( .A(n8409), .ZN(n8410) );
  AOI21_X1 U9902 ( .B1(n8412), .B2(n8411), .A(n8410), .ZN(n8417) );
  INV_X1 U9903 ( .A(n8413), .ZN(n8415) );
  OAI211_X1 U9904 ( .C1(n8417), .C2(n8416), .A(n8415), .B(n8414), .ZN(n8418)
         );
  INV_X1 U9905 ( .A(n8418), .ZN(n8421) );
  INV_X1 U9906 ( .A(n8419), .ZN(n8420) );
  NOR2_X1 U9907 ( .A1(n8421), .A2(n8420), .ZN(n8422) );
  NOR2_X1 U9908 ( .A1(n8423), .A2(n8422), .ZN(n8425) );
  OAI21_X1 U9909 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8429) );
  INV_X1 U9910 ( .A(n8427), .ZN(n8428) );
  AOI21_X1 U9911 ( .B1(n8430), .B2(n8429), .A(n8428), .ZN(n8434) );
  INV_X1 U9912 ( .A(n8431), .ZN(n8433) );
  OAI21_X1 U9913 ( .B1(n8434), .B2(n8433), .A(n8432), .ZN(n8435) );
  NAND2_X1 U9914 ( .A1(n8436), .A2(n8435), .ZN(n8437) );
  OR3_X1 U9915 ( .A1(n8439), .A2(n8438), .A3(n8437), .ZN(n8442) );
  INV_X1 U9916 ( .A(n8440), .ZN(n8441) );
  AOI21_X1 U9917 ( .B1(n8443), .B2(n8442), .A(n8441), .ZN(n8447) );
  INV_X1 U9918 ( .A(n8444), .ZN(n8446) );
  OAI21_X1 U9919 ( .B1(n8447), .B2(n8446), .A(n8445), .ZN(n8449) );
  NAND2_X1 U9920 ( .A1(n8449), .A2(n8448), .ZN(n8450) );
  MUX2_X1 U9921 ( .A(n8452), .B(n8451), .S(n8450), .Z(n8453) );
  INV_X1 U9922 ( .A(n8453), .ZN(n8460) );
  NOR3_X1 U9923 ( .A1(n8463), .A2(n8462), .A3(n8461), .ZN(n8466) );
  OAI21_X1 U9924 ( .B1(n8467), .B2(n8464), .A(P1_B_REG_SCAN_IN), .ZN(n8465) );
  NOR2_X1 U9925 ( .A1(n8469), .A2(n8468), .ZN(n8471) );
  NAND2_X1 U9926 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9366), .ZN(n8472) );
  OAI21_X1 U9927 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9366), .A(n8472), .ZN(
        n9360) );
  INV_X1 U9928 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8473) );
  XNOR2_X1 U9929 ( .A(n9375), .B(n8473), .ZN(n9374) );
  OR2_X1 U9930 ( .A1(n9375), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U9931 ( .A1(n8475), .A2(n8474), .ZN(n9390) );
  INV_X1 U9932 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9603) );
  OR2_X1 U9933 ( .A1(n9386), .A2(n9603), .ZN(n8477) );
  NAND2_X1 U9934 ( .A1(n9386), .A2(n9603), .ZN(n8476) );
  AND2_X1 U9935 ( .A1(n8477), .A2(n8476), .ZN(n9389) );
  NOR2_X1 U9936 ( .A1(n9390), .A2(n9389), .ZN(n9388) );
  AND2_X1 U9937 ( .A1(n9386), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8478) );
  INV_X1 U9938 ( .A(n8491), .ZN(n8488) );
  XNOR2_X1 U9939 ( .A(n9386), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9394) );
  INV_X1 U9940 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9691) );
  XNOR2_X1 U9941 ( .A(n9375), .B(n9691), .ZN(n9381) );
  INV_X1 U9942 ( .A(n9366), .ZN(n8484) );
  XNOR2_X1 U9943 ( .A(n9366), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U9944 ( .A1(n8481), .A2(n8480), .ZN(n8483) );
  NAND2_X1 U9945 ( .A1(n8483), .A2(n8482), .ZN(n9364) );
  NOR2_X1 U9946 ( .A1(n9363), .A2(n9364), .ZN(n9362) );
  AOI21_X1 U9947 ( .B1(n9697), .B2(n8484), .A(n9362), .ZN(n8485) );
  INV_X1 U9948 ( .A(n8485), .ZN(n9380) );
  NOR2_X1 U9949 ( .A1(n9375), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9395) );
  NOR3_X1 U9950 ( .A1(n9394), .A2(n9396), .A3(n9395), .ZN(n9393) );
  AOI21_X1 U9951 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9386), .A(n9393), .ZN(
        n8486) );
  XNOR2_X1 U9952 ( .A(n8486), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8489) );
  OAI21_X1 U9953 ( .B1(n8489), .B2(n9370), .A(n9403), .ZN(n8487) );
  AOI21_X1 U9954 ( .B1(n8488), .B2(n8490), .A(n8487), .ZN(n8493) );
  AOI22_X1 U9955 ( .A1(n8491), .A2(n8490), .B1(n9399), .B2(n8489), .ZN(n8492)
         );
  MUX2_X1 U9956 ( .A(n8493), .B(n8492), .S(n5462), .Z(n8495) );
  NAND2_X1 U9957 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n8494) );
  OAI211_X1 U9958 ( .C1(n8497), .C2(n8496), .A(n8495), .B(n8494), .ZN(P1_U3262) );
  OAI222_X1 U9959 ( .A1(n8587), .A2(n8499), .B1(n8811), .B2(P2_U3151), .C1(
        n8498), .C2(n8590), .ZN(P2_U3268) );
  OAI22_X1 U9960 ( .A1(n8501), .A2(n9601), .B1(n8500), .B2(n9624), .ZN(n8504)
         );
  NOR2_X1 U9961 ( .A1(n8502), .A2(n9586), .ZN(n8503) );
  AOI211_X1 U9962 ( .C1(n9590), .C2(n6560), .A(n8504), .B(n8503), .ZN(n8507)
         );
  OR2_X1 U9963 ( .A1(n8505), .A2(n9620), .ZN(n8506) );
  OAI211_X1 U9964 ( .C1(n8508), .C2(n9626), .A(n8507), .B(n8506), .ZN(P1_U3265) );
  NAND2_X1 U9965 ( .A1(n8510), .A2(n8509), .ZN(n9056) );
  NOR2_X1 U9966 ( .A1(n9056), .A2(n9990), .ZN(n9110) );
  AOI21_X1 U9967 ( .B1(n9990), .B2(P2_REG0_REG_30__SCAN_IN), .A(n9110), .ZN(
        n8511) );
  OAI21_X1 U9968 ( .B1(n6380), .B2(n9163), .A(n8511), .ZN(P2_U3457) );
  NAND2_X1 U9969 ( .A1(n8512), .A2(n9051), .ZN(n8526) );
  AOI21_X1 U9970 ( .B1(n8526), .B2(n9056), .A(n9037), .ZN(n8881) );
  AOI21_X1 U9971 ( .B1(n9037), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8881), .ZN(
        n8513) );
  OAI21_X1 U9972 ( .B1(n6380), .B2(n9028), .A(n8513), .ZN(P2_U3203) );
  INV_X1 U9973 ( .A(n8515), .ZN(n8516) );
  NOR2_X1 U9974 ( .A1(n8517), .A2(n8516), .ZN(n8518) );
  XNOR2_X1 U9975 ( .A(n8514), .B(n8518), .ZN(n8524) );
  INV_X1 U9976 ( .A(n8519), .ZN(n9581) );
  OAI22_X1 U9977 ( .A1(n9211), .A2(n9409), .B1(n8520), .B2(n9281), .ZN(n9576)
         );
  AOI22_X1 U9978 ( .A1(n9576), .A2(n9301), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n8521) );
  OAI21_X1 U9979 ( .B1(n9581), .B2(n9299), .A(n8521), .ZN(n8522) );
  AOI21_X1 U9980 ( .B1(n9589), .B2(n9286), .A(n8522), .ZN(n8523) );
  OAI21_X1 U9981 ( .B1(n8524), .B2(n9288), .A(n8523), .ZN(P1_U3219) );
  NAND2_X1 U9982 ( .A1(n8525), .A2(n9047), .ZN(n8530) );
  OAI21_X1 U9983 ( .B1(n9047), .B2(n8527), .A(n8526), .ZN(n8528) );
  AOI21_X1 U9984 ( .B1(n5845), .B2(n4315), .A(n8528), .ZN(n8529) );
  OAI211_X1 U9985 ( .C1(n6476), .C2(n8531), .A(n8530), .B(n8529), .ZN(P2_U3204) );
  NAND2_X1 U9986 ( .A1(n8533), .A2(n8532), .ZN(n8535) );
  INV_X1 U9987 ( .A(n8533), .ZN(n8534) );
  AOI21_X2 U9988 ( .B1(n8536), .B2(n8535), .A(n4905), .ZN(n8602) );
  XNOR2_X1 U9989 ( .A(n8537), .B(n7064), .ZN(n8538) );
  XNOR2_X1 U9990 ( .A(n8538), .B(n8539), .ZN(n8603) );
  NAND2_X1 U9991 ( .A1(n8602), .A2(n8603), .ZN(n8601) );
  INV_X1 U9992 ( .A(n8538), .ZN(n8540) );
  NAND2_X1 U9993 ( .A1(n8540), .A2(n8539), .ZN(n8541) );
  NAND2_X1 U9994 ( .A1(n8601), .A2(n8541), .ZN(n8726) );
  XNOR2_X1 U9995 ( .A(n8542), .B(n7064), .ZN(n8544) );
  XNOR2_X1 U9996 ( .A(n8544), .B(n9042), .ZN(n8725) );
  INV_X1 U9997 ( .A(n8725), .ZN(n8543) );
  NAND2_X1 U9998 ( .A1(n8544), .A2(n9042), .ZN(n8545) );
  XNOR2_X1 U9999 ( .A(n9168), .B(n7064), .ZN(n8546) );
  XNOR2_X1 U10000 ( .A(n8546), .B(n8732), .ZN(n8652) );
  XNOR2_X1 U10001 ( .A(n9100), .B(n7064), .ZN(n8547) );
  NOR2_X1 U10002 ( .A1(n8547), .A2(n9044), .ZN(n8702) );
  AOI21_X1 U10003 ( .B1(n9044), .B2(n8547), .A(n8702), .ZN(n8661) );
  NAND2_X1 U10004 ( .A1(n8662), .A2(n8661), .ZN(n8660) );
  INV_X1 U10005 ( .A(n8702), .ZN(n8548) );
  NAND2_X1 U10006 ( .A1(n8660), .A2(n8548), .ZN(n8549) );
  XNOR2_X1 U10007 ( .A(n8700), .B(n7064), .ZN(n8550) );
  XNOR2_X1 U10008 ( .A(n8550), .B(n8997), .ZN(n8701) );
  INV_X1 U10009 ( .A(n8550), .ZN(n8551) );
  NAND2_X1 U10010 ( .A1(n8551), .A2(n8997), .ZN(n8552) );
  XNOR2_X1 U10011 ( .A(n9156), .B(n7064), .ZN(n8554) );
  XNOR2_X1 U10012 ( .A(n8554), .B(n8745), .ZN(n8622) );
  XNOR2_X1 U10013 ( .A(n9089), .B(n8564), .ZN(n8553) );
  NAND2_X1 U10014 ( .A1(n8553), .A2(n8998), .ZN(n8632) );
  OAI21_X1 U10015 ( .B1(n8553), .B2(n8998), .A(n8632), .ZN(n8681) );
  AND2_X1 U10016 ( .A1(n8554), .A2(n8745), .ZN(n8680) );
  NOR2_X1 U10017 ( .A1(n8681), .A2(n8680), .ZN(n8555) );
  NAND2_X1 U10018 ( .A1(n8624), .A2(n8555), .ZN(n8631) );
  NAND2_X1 U10019 ( .A1(n8631), .A2(n8632), .ZN(n8556) );
  XNOR2_X1 U10020 ( .A(n9085), .B(n7064), .ZN(n8557) );
  XNOR2_X1 U10021 ( .A(n8557), .B(n8985), .ZN(n8633) );
  NAND2_X1 U10022 ( .A1(n8556), .A2(n8633), .ZN(n8635) );
  INV_X1 U10023 ( .A(n8557), .ZN(n8558) );
  NAND2_X1 U10024 ( .A1(n8558), .A2(n8985), .ZN(n8559) );
  XNOR2_X1 U10025 ( .A(n6457), .B(n7064), .ZN(n8561) );
  XNOR2_X1 U10026 ( .A(n8561), .B(n8742), .ZN(n8692) );
  INV_X1 U10027 ( .A(n8692), .ZN(n8560) );
  NAND2_X1 U10028 ( .A1(n8561), .A2(n8742), .ZN(n8562) );
  XNOR2_X1 U10029 ( .A(n8950), .B(n8564), .ZN(n8614) );
  NAND2_X1 U10030 ( .A1(n8614), .A2(n8958), .ZN(n8563) );
  NAND2_X1 U10031 ( .A1(n8613), .A2(n8563), .ZN(n8568) );
  INV_X1 U10032 ( .A(n8614), .ZN(n8566) );
  XNOR2_X1 U10033 ( .A(n9133), .B(n8564), .ZN(n8565) );
  NAND2_X1 U10034 ( .A1(n8565), .A2(n8946), .ZN(n8644) );
  OAI21_X1 U10035 ( .B1(n8565), .B2(n8946), .A(n8644), .ZN(n8669) );
  AOI21_X1 U10036 ( .B1(n8935), .B2(n8566), .A(n8669), .ZN(n8567) );
  XNOR2_X1 U10037 ( .A(n9127), .B(n7064), .ZN(n8569) );
  XNOR2_X1 U10038 ( .A(n8569), .B(n8717), .ZN(n8645) );
  INV_X1 U10039 ( .A(n8569), .ZN(n8570) );
  NAND2_X1 U10040 ( .A1(n8570), .A2(n8717), .ZN(n8571) );
  XNOR2_X1 U10041 ( .A(n9122), .B(n7064), .ZN(n8572) );
  NAND2_X1 U10042 ( .A1(n8712), .A2(n8713), .ZN(n8711) );
  INV_X1 U10043 ( .A(n8572), .ZN(n8573) );
  NAND2_X1 U10044 ( .A1(n8574), .A2(n8573), .ZN(n8575) );
  NAND2_X1 U10045 ( .A1(n8711), .A2(n8575), .ZN(n8592) );
  XNOR2_X1 U10046 ( .A(n9116), .B(n7064), .ZN(n8576) );
  XNOR2_X1 U10047 ( .A(n8576), .B(n8914), .ZN(n8591) );
  NAND2_X1 U10048 ( .A1(n8593), .A2(n8577), .ZN(n8579) );
  XNOR2_X1 U10049 ( .A(n8895), .B(n7064), .ZN(n8578) );
  XNOR2_X1 U10050 ( .A(n8579), .B(n8578), .ZN(n8584) );
  AOI22_X1 U10051 ( .A1(n8889), .A2(n8734), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8581) );
  NAND2_X1 U10052 ( .A1(n8914), .A2(n8729), .ZN(n8580) );
  OAI211_X1 U10053 ( .C1(n8741), .C2(n8731), .A(n8581), .B(n8580), .ZN(n8582)
         );
  AOI21_X1 U10054 ( .B1(n9062), .B2(n8657), .A(n8582), .ZN(n8583) );
  OAI21_X1 U10055 ( .B1(n8584), .B2(n8724), .A(n8583), .ZN(P2_U3160) );
  OAI222_X1 U10056 ( .A1(n8587), .A2(n8586), .B1(n6403), .B2(P2_U3151), .C1(
        n8585), .C2(n8590), .ZN(P2_U3267) );
  INV_X1 U10057 ( .A(n8588), .ZN(n9789) );
  OAI222_X1 U10058 ( .A1(n8590), .A2(n10044), .B1(n8587), .B2(n9789), .C1(
        P2_U3151), .C2(n8589), .ZN(P2_U3265) );
  INV_X1 U10059 ( .A(n9116), .ZN(n8600) );
  AOI21_X1 U10060 ( .B1(n8592), .B2(n8591), .A(n8724), .ZN(n8594) );
  NAND2_X1 U10061 ( .A1(n8594), .A2(n8593), .ZN(n8599) );
  AOI22_X1 U10062 ( .A1(n8908), .A2(n8734), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8595) );
  OAI21_X1 U10063 ( .B1(n8596), .B2(n8731), .A(n8595), .ZN(n8597) );
  AOI21_X1 U10064 ( .B1(n8729), .B2(n8924), .A(n8597), .ZN(n8598) );
  OAI211_X1 U10065 ( .C1(n8600), .C2(n8738), .A(n8599), .B(n8598), .ZN(
        P2_U3154) );
  OAI21_X1 U10066 ( .B1(n8603), .B2(n8602), .A(n8601), .ZN(n8604) );
  NAND2_X1 U10067 ( .A1(n8604), .A2(n8714), .ZN(n8611) );
  OAI21_X1 U10068 ( .B1(n8731), .B2(n8606), .A(n8605), .ZN(n8609) );
  NOR2_X1 U10069 ( .A1(n8664), .A2(n8607), .ZN(n8608) );
  AOI211_X1 U10070 ( .C1(n8729), .C2(n8747), .A(n8609), .B(n8608), .ZN(n8610)
         );
  OAI211_X1 U10071 ( .C1(n8612), .C2(n8738), .A(n8611), .B(n8610), .ZN(
        P2_U3155) );
  INV_X1 U10072 ( .A(n8613), .ZN(n8615) );
  NAND2_X1 U10073 ( .A1(n8615), .A2(n8614), .ZN(n8670) );
  OAI21_X1 U10074 ( .B1(n8615), .B2(n8614), .A(n8670), .ZN(n8616) );
  NOR2_X1 U10075 ( .A1(n8616), .A2(n8935), .ZN(n8673) );
  AOI21_X1 U10076 ( .B1(n8935), .B2(n8616), .A(n8673), .ZN(n8621) );
  AOI22_X1 U10077 ( .A1(n8923), .A2(n8686), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8618) );
  NAND2_X1 U10078 ( .A1(n8734), .A2(n8949), .ZN(n8617) );
  OAI211_X1 U10079 ( .C1(n8968), .C2(n8716), .A(n8618), .B(n8617), .ZN(n8619)
         );
  AOI21_X1 U10080 ( .B1(n8950), .B2(n8657), .A(n8619), .ZN(n8620) );
  OAI21_X1 U10081 ( .B1(n8621), .B2(n8724), .A(n8620), .ZN(P2_U3156) );
  INV_X1 U10082 ( .A(n9156), .ZN(n8630) );
  AOI21_X1 U10083 ( .B1(n8623), .B2(n8622), .A(n8724), .ZN(n8625) );
  NAND2_X1 U10084 ( .A1(n8625), .A2(n8624), .ZN(n8629) );
  NAND2_X1 U10085 ( .A1(n8729), .A2(n9024), .ZN(n8626) );
  NAND2_X1 U10086 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8870) );
  OAI211_X1 U10087 ( .C1(n8998), .C2(n8731), .A(n8626), .B(n8870), .ZN(n8627)
         );
  AOI21_X1 U10088 ( .B1(n9003), .B2(n8734), .A(n8627), .ZN(n8628) );
  OAI211_X1 U10089 ( .C1(n8630), .C2(n8738), .A(n8629), .B(n8628), .ZN(
        P2_U3159) );
  INV_X1 U10090 ( .A(n9085), .ZN(n8642) );
  INV_X1 U10091 ( .A(n8631), .ZN(n8685) );
  INV_X1 U10092 ( .A(n8632), .ZN(n8634) );
  NOR3_X1 U10093 ( .A1(n8685), .A2(n8634), .A3(n8633), .ZN(n8637) );
  INV_X1 U10094 ( .A(n8635), .ZN(n8636) );
  OAI21_X1 U10095 ( .B1(n8637), .B2(n8636), .A(n8714), .ZN(n8641) );
  AOI22_X1 U10096 ( .A1(n8742), .A2(n8686), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8638) );
  OAI21_X1 U10097 ( .B1(n8998), .B2(n8716), .A(n8638), .ZN(n8639) );
  AOI21_X1 U10098 ( .B1(n8973), .B2(n8734), .A(n8639), .ZN(n8640) );
  OAI211_X1 U10099 ( .C1(n8642), .C2(n8738), .A(n8641), .B(n8640), .ZN(
        P2_U3163) );
  INV_X1 U10100 ( .A(n9127), .ZN(n8926) );
  INV_X1 U10101 ( .A(n8643), .ZN(n8674) );
  NOR3_X1 U10102 ( .A1(n8674), .A2(n4663), .A3(n8645), .ZN(n8646) );
  OAI21_X1 U10103 ( .B1(n8646), .B2(n4348), .A(n8714), .ZN(n8651) );
  INV_X1 U10104 ( .A(n8928), .ZN(n8648) );
  AOI22_X1 U10105 ( .A1(n8923), .A2(n8729), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8647) );
  OAI21_X1 U10106 ( .B1(n8648), .B2(n8664), .A(n8647), .ZN(n8649) );
  AOI21_X1 U10107 ( .B1(n8686), .B2(n8924), .A(n8649), .ZN(n8650) );
  OAI211_X1 U10108 ( .C1(n8926), .C2(n8738), .A(n8651), .B(n8650), .ZN(
        P2_U3165) );
  XNOR2_X1 U10109 ( .A(n8653), .B(n8652), .ZN(n8659) );
  NAND2_X1 U10110 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8795) );
  OAI21_X1 U10111 ( .B1(n8731), .B2(n9009), .A(n8795), .ZN(n8654) );
  AOI21_X1 U10112 ( .B1(n8729), .B2(n9042), .A(n8654), .ZN(n8655) );
  OAI21_X1 U10113 ( .B1(n9049), .B2(n8664), .A(n8655), .ZN(n8656) );
  AOI21_X1 U10114 ( .B1(n9168), .B2(n8657), .A(n8656), .ZN(n8658) );
  OAI21_X1 U10115 ( .B1(n8659), .B2(n8724), .A(n8658), .ZN(P2_U3166) );
  INV_X1 U10116 ( .A(n9100), .ZN(n9029) );
  OAI21_X1 U10117 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8663) );
  NAND2_X1 U10118 ( .A1(n8663), .A2(n8714), .ZN(n8668) );
  NAND2_X1 U10119 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8823) );
  OAI21_X1 U10120 ( .B1(n8731), .B2(n8997), .A(n8823), .ZN(n8666) );
  NOR2_X1 U10121 ( .A1(n8664), .A2(n9031), .ZN(n8665) );
  AOI211_X1 U10122 ( .C1(n8729), .C2(n9023), .A(n8666), .B(n8665), .ZN(n8667)
         );
  OAI211_X1 U10123 ( .C1(n9029), .C2(n8738), .A(n8668), .B(n8667), .ZN(
        P2_U3168) );
  INV_X1 U10124 ( .A(n9133), .ZN(n8938) );
  INV_X1 U10125 ( .A(n8669), .ZN(n8672) );
  INV_X1 U10126 ( .A(n8670), .ZN(n8671) );
  NOR3_X1 U10127 ( .A1(n8673), .A2(n8672), .A3(n8671), .ZN(n8675) );
  OAI21_X1 U10128 ( .B1(n8675), .B2(n8674), .A(n8714), .ZN(n8679) );
  AOI22_X1 U10129 ( .A1(n8934), .A2(n8686), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8676) );
  OAI21_X1 U10130 ( .B1(n8958), .B2(n8716), .A(n8676), .ZN(n8677) );
  AOI21_X1 U10131 ( .B1(n8940), .B2(n8734), .A(n8677), .ZN(n8678) );
  OAI211_X1 U10132 ( .C1(n8938), .C2(n8738), .A(n8679), .B(n8678), .ZN(
        P2_U3169) );
  INV_X1 U10133 ( .A(n9089), .ZN(n8691) );
  INV_X1 U10134 ( .A(n8680), .ZN(n8683) );
  INV_X1 U10135 ( .A(n8681), .ZN(n8682) );
  AOI21_X1 U10136 ( .B1(n8624), .B2(n8683), .A(n8682), .ZN(n8684) );
  OAI21_X1 U10137 ( .B1(n8685), .B2(n8684), .A(n8714), .ZN(n8690) );
  AOI22_X1 U10138 ( .A1(n8686), .A2(n8743), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8687) );
  OAI21_X1 U10139 ( .B1(n9011), .B2(n8716), .A(n8687), .ZN(n8688) );
  AOI21_X1 U10140 ( .B1(n8986), .B2(n8734), .A(n8688), .ZN(n8689) );
  OAI211_X1 U10141 ( .C1(n8691), .C2(n8738), .A(n8690), .B(n8689), .ZN(
        P2_U3173) );
  AOI21_X1 U10142 ( .B1(n8693), .B2(n8692), .A(n8724), .ZN(n8695) );
  NAND2_X1 U10143 ( .A1(n8695), .A2(n8694), .ZN(n8699) );
  AOI22_X1 U10144 ( .A1(n8729), .A2(n8743), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8696) );
  OAI21_X1 U10145 ( .B1(n8958), .B2(n8731), .A(n8696), .ZN(n8697) );
  AOI21_X1 U10146 ( .B1(n8961), .B2(n8734), .A(n8697), .ZN(n8698) );
  OAI211_X1 U10147 ( .C1(n9145), .C2(n8738), .A(n8699), .B(n8698), .ZN(
        P2_U3175) );
  INV_X1 U10148 ( .A(n8660), .ZN(n8703) );
  NOR3_X1 U10149 ( .A1(n8703), .A2(n8702), .A3(n8701), .ZN(n8706) );
  INV_X1 U10150 ( .A(n8704), .ZN(n8705) );
  OAI21_X1 U10151 ( .B1(n8706), .B2(n8705), .A(n8714), .ZN(n8710) );
  NAND2_X1 U10152 ( .A1(n8729), .A2(n9044), .ZN(n8707) );
  NAND2_X1 U10153 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8843) );
  OAI211_X1 U10154 ( .C1(n9011), .C2(n8731), .A(n8707), .B(n8843), .ZN(n8708)
         );
  AOI21_X1 U10155 ( .B1(n9017), .B2(n8734), .A(n8708), .ZN(n8709) );
  OAI211_X1 U10156 ( .C1(n9164), .C2(n8738), .A(n8710), .B(n8709), .ZN(
        P2_U3178) );
  INV_X1 U10157 ( .A(n9122), .ZN(n8723) );
  OAI21_X1 U10158 ( .B1(n8713), .B2(n8712), .A(n8711), .ZN(n8715) );
  NAND2_X1 U10159 ( .A1(n8715), .A2(n8714), .ZN(n8722) );
  OAI22_X1 U10160 ( .A1(n8717), .A2(n8716), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10160), .ZN(n8720) );
  NOR2_X1 U10161 ( .A1(n8718), .A2(n8731), .ZN(n8719) );
  AOI211_X1 U10162 ( .C1(n8917), .C2(n8734), .A(n8720), .B(n8719), .ZN(n8721)
         );
  OAI211_X1 U10163 ( .C1(n8723), .C2(n8738), .A(n8722), .B(n8721), .ZN(
        P2_U3180) );
  AOI21_X1 U10164 ( .B1(n8726), .B2(n8725), .A(n8724), .ZN(n8728) );
  NAND2_X1 U10165 ( .A1(n8728), .A2(n8727), .ZN(n8737) );
  NAND2_X1 U10166 ( .A1(n8729), .A2(n8746), .ZN(n8730) );
  NAND2_X1 U10167 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8764) );
  OAI211_X1 U10168 ( .C1(n8732), .C2(n8731), .A(n8730), .B(n8764), .ZN(n8733)
         );
  AOI21_X1 U10169 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8736) );
  OAI211_X1 U10170 ( .C1(n8739), .C2(n8738), .A(n8737), .B(n8736), .ZN(
        P2_U3181) );
  MUX2_X1 U10171 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8740), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10172 ( .A(n8741), .ZN(n8884) );
  MUX2_X1 U10173 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8884), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10174 ( .A(n8904), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8841), .Z(
        P2_U3519) );
  MUX2_X1 U10175 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8914), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10176 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8924), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10177 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8934), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10178 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8923), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10179 ( .A(n8935), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8841), .Z(
        P2_U3514) );
  MUX2_X1 U10180 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8742), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10181 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8743), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10182 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8744), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10183 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8745), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10184 ( .A(n9024), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8841), .Z(
        P2_U3509) );
  MUX2_X1 U10185 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9044), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10186 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9023), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10187 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9042), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10188 ( .A(n8746), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8841), .Z(
        P2_U3505) );
  MUX2_X1 U10189 ( .A(n8747), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8841), .Z(
        P2_U3504) );
  MUX2_X1 U10190 ( .A(n8748), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8841), .Z(
        P2_U3503) );
  MUX2_X1 U10191 ( .A(n8749), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8841), .Z(
        P2_U3502) );
  MUX2_X1 U10192 ( .A(n8750), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8841), .Z(
        P2_U3501) );
  MUX2_X1 U10193 ( .A(n8751), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8841), .Z(
        P2_U3500) );
  MUX2_X1 U10194 ( .A(n8752), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8841), .Z(
        P2_U3499) );
  MUX2_X1 U10195 ( .A(n8753), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8841), .Z(
        P2_U3498) );
  MUX2_X1 U10196 ( .A(n8754), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8841), .Z(
        P2_U3497) );
  MUX2_X1 U10197 ( .A(n8755), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8841), .Z(
        P2_U3496) );
  MUX2_X1 U10198 ( .A(n8756), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8841), .Z(
        P2_U3495) );
  MUX2_X1 U10199 ( .A(n8757), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8841), .Z(
        P2_U3494) );
  MUX2_X1 U10200 ( .A(n8758), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8841), .Z(
        P2_U3493) );
  MUX2_X1 U10201 ( .A(n8759), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8841), .Z(
        P2_U3492) );
  MUX2_X1 U10202 ( .A(n8760), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8841), .Z(
        P2_U3491) );
  NOR2_X1 U10203 ( .A1(n8191), .A2(n8763), .ZN(n8799) );
  AOI21_X1 U10204 ( .B1(n8191), .B2(n8763), .A(n8799), .ZN(n8781) );
  OAI21_X1 U10205 ( .B1(n9896), .B2(n8765), .A(n8764), .ZN(n8779) );
  XNOR2_X1 U10206 ( .A(n8798), .B(n8782), .ZN(n8768) );
  NOR2_X1 U10207 ( .A1(n8767), .A2(n8768), .ZN(n8783) );
  AOI21_X1 U10208 ( .B1(n8768), .B2(n8767), .A(n8783), .ZN(n8777) );
  MUX2_X1 U10209 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8811), .Z(n8788) );
  XNOR2_X1 U10210 ( .A(n8798), .B(n8788), .ZN(n8774) );
  OR2_X1 U10211 ( .A1(n8770), .A2(n8769), .ZN(n8772) );
  NAND2_X1 U10212 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  NAND2_X1 U10213 ( .A1(n8774), .A2(n8773), .ZN(n8789) );
  OAI21_X1 U10214 ( .B1(n8774), .B2(n8773), .A(n8789), .ZN(n8775) );
  NAND2_X1 U10215 ( .A1(n8775), .A2(n9892), .ZN(n8776) );
  OAI21_X1 U10216 ( .B1(n8777), .B2(n9908), .A(n8776), .ZN(n8778) );
  AOI211_X1 U10217 ( .C1(n8798), .C2(n9902), .A(n8779), .B(n8778), .ZN(n8780)
         );
  OAI21_X1 U10218 ( .B1(n8781), .B2(n8877), .A(n8780), .ZN(P2_U3197) );
  NOR2_X1 U10219 ( .A1(n8798), .A2(n8782), .ZN(n8784) );
  XNOR2_X1 U10220 ( .A(n8806), .B(n9104), .ZN(n8785) );
  NOR2_X1 U10221 ( .A1(n8786), .A2(n8785), .ZN(n8817) );
  AOI21_X1 U10222 ( .B1(n8786), .B2(n8785), .A(n8817), .ZN(n8808) );
  MUX2_X1 U10223 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8811), .Z(n8812) );
  XNOR2_X1 U10224 ( .A(n8812), .B(n8806), .ZN(n8792) );
  OR2_X1 U10225 ( .A1(n8788), .A2(n8787), .ZN(n8790) );
  NAND2_X1 U10226 ( .A1(n8790), .A2(n8789), .ZN(n8791) );
  NAND2_X1 U10227 ( .A1(n8792), .A2(n8791), .ZN(n8813) );
  OAI21_X1 U10228 ( .B1(n8792), .B2(n8791), .A(n8813), .ZN(n8793) );
  NAND2_X1 U10229 ( .A1(n8793), .A2(n9892), .ZN(n8794) );
  OAI211_X1 U10230 ( .C1(n9896), .C2(n8796), .A(n8795), .B(n8794), .ZN(n8805)
         );
  NOR2_X1 U10231 ( .A1(n8798), .A2(n8797), .ZN(n8800) );
  NOR2_X1 U10232 ( .A1(n8800), .A2(n8799), .ZN(n8802) );
  AOI22_X1 U10233 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8806), .B1(n8818), .B2(
        n9048), .ZN(n8801) );
  NOR2_X1 U10234 ( .A1(n8802), .A2(n8801), .ZN(n8809) );
  AOI21_X1 U10235 ( .B1(n8802), .B2(n8801), .A(n8809), .ZN(n8803) );
  NOR2_X1 U10236 ( .A1(n8803), .A2(n8877), .ZN(n8804) );
  AOI211_X1 U10237 ( .C1(n9902), .C2(n8806), .A(n8805), .B(n8804), .ZN(n8807)
         );
  OAI21_X1 U10238 ( .B1(n8808), .B2(n9908), .A(n8807), .ZN(P2_U3198) );
  AOI21_X1 U10239 ( .B1(n9032), .B2(n8810), .A(n8847), .ZN(n8829) );
  MUX2_X1 U10240 ( .A(n9032), .B(n8819), .S(n8811), .Z(n8836) );
  XOR2_X1 U10241 ( .A(n8846), .B(n8836), .Z(n8816) );
  OR2_X1 U10242 ( .A1(n8812), .A2(n8818), .ZN(n8814) );
  NAND2_X1 U10243 ( .A1(n8814), .A2(n8813), .ZN(n8815) );
  NAND2_X1 U10244 ( .A1(n8816), .A2(n8815), .ZN(n8834) );
  OAI21_X1 U10245 ( .B1(n8816), .B2(n8815), .A(n8834), .ZN(n8825) );
  NOR2_X1 U10246 ( .A1(n9896), .A2(n8826), .ZN(n8827) );
  AOI21_X1 U10247 ( .B1(n9902), .B2(n8846), .A(n8827), .ZN(n8828) );
  NOR2_X1 U10248 ( .A1(n8846), .A2(n8830), .ZN(n8832) );
  NAND2_X1 U10249 ( .A1(n8849), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8858) );
  OAI21_X1 U10250 ( .B1(n8849), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8858), .ZN(
        n8833) );
  AOI21_X1 U10251 ( .B1(n4357), .B2(n8833), .A(n8860), .ZN(n8857) );
  INV_X1 U10252 ( .A(n8834), .ZN(n8835) );
  AOI21_X1 U10253 ( .B1(n8836), .B2(n8846), .A(n8835), .ZN(n8838) );
  MUX2_X1 U10254 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8811), .Z(n8837) );
  NOR2_X1 U10255 ( .A1(n8838), .A2(n8837), .ZN(n8866) );
  INV_X1 U10256 ( .A(n8866), .ZN(n8839) );
  NAND2_X1 U10257 ( .A1(n8838), .A2(n8837), .ZN(n8864) );
  NAND2_X1 U10258 ( .A1(n8839), .A2(n8864), .ZN(n8842) );
  OAI21_X1 U10259 ( .B1(n8841), .B2(n8842), .A(n8840), .ZN(n8855) );
  INV_X1 U10260 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10011) );
  NAND3_X1 U10261 ( .A1(n8842), .A2(n9892), .A3(n8849), .ZN(n8844) );
  OAI211_X1 U10262 ( .C1(n10011), .C2(n9896), .A(n8844), .B(n8843), .ZN(n8854)
         );
  NOR2_X1 U10263 ( .A1(n8846), .A2(n8845), .ZN(n8848) );
  NAND2_X1 U10264 ( .A1(n8849), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8872) );
  OAI21_X1 U10265 ( .B1(n8849), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8872), .ZN(
        n8850) );
  NOR2_X1 U10266 ( .A1(n8851), .A2(n8850), .ZN(n8874) );
  AOI21_X1 U10267 ( .B1(n8851), .B2(n8850), .A(n8874), .ZN(n8852) );
  NOR2_X1 U10268 ( .A1(n8852), .A2(n8877), .ZN(n8853) );
  OAI21_X1 U10269 ( .B1(n8857), .B2(n9908), .A(n8856), .ZN(P2_U3200) );
  INV_X1 U10270 ( .A(n8858), .ZN(n8859) );
  NOR2_X1 U10271 ( .A1(n8860), .A2(n8859), .ZN(n8861) );
  XNOR2_X1 U10272 ( .A(n8862), .B(n9092), .ZN(n8863) );
  XNOR2_X1 U10273 ( .A(n8861), .B(n8863), .ZN(n8880) );
  MUX2_X1 U10274 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9002), .S(n8862), .Z(n8875) );
  MUX2_X1 U10275 ( .A(n8863), .B(n8875), .S(n6869), .Z(n8868) );
  OAI21_X1 U10276 ( .B1(n8866), .B2(n8865), .A(n8864), .ZN(n8867) );
  XOR2_X1 U10277 ( .A(n8868), .B(n8867), .Z(n8879) );
  NAND2_X1 U10278 ( .A1(n9902), .A2(n8869), .ZN(n8871) );
  OAI211_X1 U10279 ( .C1(n4408), .C2(n9896), .A(n8871), .B(n8870), .ZN(n8878)
         );
  INV_X1 U10280 ( .A(n8872), .ZN(n8873) );
  NOR2_X1 U10281 ( .A1(n8874), .A2(n8873), .ZN(n8876) );
  AOI21_X1 U10282 ( .B1(n9037), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8881), .ZN(
        n8882) );
  OAI21_X1 U10283 ( .B1(n9112), .B2(n9028), .A(n8882), .ZN(P2_U3202) );
  XNOR2_X1 U10284 ( .A(n8883), .B(n8895), .ZN(n8888) );
  NAND2_X1 U10285 ( .A1(n8884), .A2(n9043), .ZN(n8886) );
  NAND2_X1 U10286 ( .A1(n8914), .A2(n9041), .ZN(n8885) );
  INV_X1 U10287 ( .A(n8889), .ZN(n8891) );
  OAI22_X1 U10288 ( .A1(n8891), .A2(n9030), .B1(n9047), .B2(n8890), .ZN(n8897)
         );
  INV_X1 U10289 ( .A(n8892), .ZN(n8893) );
  AOI21_X1 U10290 ( .B1(n8895), .B2(n8894), .A(n8893), .ZN(n9065) );
  NOR2_X1 U10291 ( .A1(n9065), .A2(n9055), .ZN(n8896) );
  AOI211_X1 U10292 ( .C1(n4315), .C2(n9062), .A(n8897), .B(n8896), .ZN(n8898)
         );
  OAI21_X1 U10293 ( .B1(n9064), .B2(n9037), .A(n8898), .ZN(P2_U3205) );
  XOR2_X1 U10294 ( .A(n8899), .B(n8900), .Z(n9119) );
  NOR2_X1 U10295 ( .A1(n8901), .A2(n8900), .ZN(n8903) );
  AOI22_X1 U10296 ( .A1(n8904), .A2(n9043), .B1(n9041), .B2(n8924), .ZN(n8905)
         );
  MUX2_X1 U10297 ( .A(n9115), .B(n8907), .S(n9037), .Z(n8910) );
  AOI22_X1 U10298 ( .A1(n9116), .A2(n4315), .B1(n9051), .B2(n8908), .ZN(n8909)
         );
  OAI211_X1 U10299 ( .C1(n9119), .C2(n9055), .A(n8910), .B(n8909), .ZN(
        P2_U3206) );
  XOR2_X1 U10300 ( .A(n8911), .B(n8912), .Z(n9125) );
  XNOR2_X1 U10301 ( .A(n8913), .B(n8912), .ZN(n8915) );
  AOI222_X1 U10302 ( .A1(n9046), .A2(n8915), .B1(n8914), .B2(n9043), .C1(n8934), .C2(n9041), .ZN(n9120) );
  MUX2_X1 U10303 ( .A(n8916), .B(n9120), .S(n9047), .Z(n8919) );
  AOI22_X1 U10304 ( .A1(n9122), .A2(n4315), .B1(n8917), .B2(n9051), .ZN(n8918)
         );
  OAI211_X1 U10305 ( .C1(n9125), .C2(n9055), .A(n8919), .B(n8918), .ZN(
        P2_U3207) );
  XNOR2_X1 U10306 ( .A(n8920), .B(n8922), .ZN(n9130) );
  XOR2_X1 U10307 ( .A(n8922), .B(n8921), .Z(n8925) );
  AOI222_X1 U10308 ( .A1(n9046), .A2(n8925), .B1(n8924), .B2(n9043), .C1(n8923), .C2(n9041), .ZN(n9126) );
  OAI21_X1 U10309 ( .B1(n8926), .B2(n8937), .A(n9126), .ZN(n8927) );
  NAND2_X1 U10310 ( .A1(n8927), .A2(n9047), .ZN(n8930) );
  AOI22_X1 U10311 ( .A1(n8928), .A2(n9051), .B1(n9037), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8929) );
  OAI211_X1 U10312 ( .C1(n9130), .C2(n9055), .A(n8930), .B(n8929), .ZN(
        P2_U3208) );
  XOR2_X1 U10313 ( .A(n8932), .B(n8931), .Z(n9136) );
  XNOR2_X1 U10314 ( .A(n8933), .B(n8932), .ZN(n8936) );
  AOI222_X1 U10315 ( .A1(n9046), .A2(n8936), .B1(n8935), .B2(n9041), .C1(n8934), .C2(n9043), .ZN(n9131) );
  OAI21_X1 U10316 ( .B1(n8938), .B2(n8937), .A(n9131), .ZN(n8939) );
  NAND2_X1 U10317 ( .A1(n8939), .A2(n9047), .ZN(n8942) );
  AOI22_X1 U10318 ( .A1(n8940), .A2(n9051), .B1(n9037), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8941) );
  OAI211_X1 U10319 ( .C1(n9136), .C2(n9055), .A(n8942), .B(n8941), .ZN(
        P2_U3209) );
  XNOR2_X1 U10320 ( .A(n8943), .B(n4914), .ZN(n9139) );
  XNOR2_X1 U10321 ( .A(n8944), .B(n4914), .ZN(n8945) );
  OAI222_X1 U10322 ( .A1(n9012), .A2(n8946), .B1(n9010), .B2(n8968), .C1(n9007), .C2(n8945), .ZN(n9137) );
  INV_X1 U10323 ( .A(n9137), .ZN(n8947) );
  MUX2_X1 U10324 ( .A(n8948), .B(n8947), .S(n9047), .Z(n8952) );
  AOI22_X1 U10325 ( .A1(n8950), .A2(n4315), .B1(n9051), .B2(n8949), .ZN(n8951)
         );
  OAI211_X1 U10326 ( .C1(n9139), .C2(n9055), .A(n8952), .B(n8951), .ZN(
        P2_U3210) );
  NAND2_X1 U10327 ( .A1(n8966), .A2(n8971), .ZN(n8954) );
  NAND2_X1 U10328 ( .A1(n8954), .A2(n8953), .ZN(n8956) );
  XNOR2_X1 U10329 ( .A(n8956), .B(n8955), .ZN(n8957) );
  OAI222_X1 U10330 ( .A1(n9012), .A2(n8958), .B1(n9010), .B2(n8985), .C1(n9007), .C2(n8957), .ZN(n9080) );
  INV_X1 U10331 ( .A(n9080), .ZN(n8965) );
  XNOR2_X1 U10332 ( .A(n8960), .B(n8959), .ZN(n9081) );
  AOI22_X1 U10333 ( .A1(n9037), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8961), .B2(
        n9051), .ZN(n8962) );
  OAI21_X1 U10334 ( .B1(n9145), .B2(n9028), .A(n8962), .ZN(n8963) );
  AOI21_X1 U10335 ( .B1(n9081), .B2(n9035), .A(n8963), .ZN(n8964) );
  OAI21_X1 U10336 ( .B1(n8965), .B2(n9037), .A(n8964), .ZN(P2_U3211) );
  XOR2_X1 U10337 ( .A(n8966), .B(n8971), .Z(n8967) );
  OAI222_X1 U10338 ( .A1(n9012), .A2(n8968), .B1(n9010), .B2(n8998), .C1(n9007), .C2(n8967), .ZN(n9084) );
  NAND2_X1 U10339 ( .A1(n8970), .A2(n8969), .ZN(n8972) );
  XNOR2_X1 U10340 ( .A(n8972), .B(n8971), .ZN(n9149) );
  AOI22_X1 U10341 ( .A1(n9037), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9051), .B2(
        n8973), .ZN(n8975) );
  NAND2_X1 U10342 ( .A1(n9085), .A2(n4315), .ZN(n8974) );
  OAI211_X1 U10343 ( .C1(n9149), .C2(n9055), .A(n8975), .B(n8974), .ZN(n8976)
         );
  AOI21_X1 U10344 ( .B1(n9084), .B2(n9047), .A(n8976), .ZN(n8977) );
  INV_X1 U10345 ( .A(n8977), .ZN(P2_U3212) );
  XNOR2_X1 U10346 ( .A(n8979), .B(n8978), .ZN(n9153) );
  INV_X1 U10347 ( .A(n8980), .ZN(n8981) );
  AOI21_X1 U10348 ( .B1(n8983), .B2(n8982), .A(n8981), .ZN(n8984) );
  OAI222_X1 U10349 ( .A1(n9012), .A2(n8985), .B1(n9010), .B2(n9011), .C1(n9007), .C2(n8984), .ZN(n9088) );
  NAND2_X1 U10350 ( .A1(n9088), .A2(n9047), .ZN(n8991) );
  INV_X1 U10351 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8988) );
  INV_X1 U10352 ( .A(n8986), .ZN(n8987) );
  OAI22_X1 U10353 ( .A1(n9047), .A2(n8988), .B1(n8987), .B2(n9030), .ZN(n8989)
         );
  AOI21_X1 U10354 ( .B1(n9089), .B2(n4315), .A(n8989), .ZN(n8990) );
  OAI211_X1 U10355 ( .C1(n9153), .C2(n9055), .A(n8991), .B(n8990), .ZN(
        P2_U3213) );
  XOR2_X1 U10356 ( .A(n8992), .B(n8995), .Z(n9159) );
  NAND2_X1 U10357 ( .A1(n8994), .A2(n8993), .ZN(n8996) );
  AOI21_X1 U10358 ( .B1(n8996), .B2(n8995), .A(n9007), .ZN(n9001) );
  OAI22_X1 U10359 ( .A1(n8998), .A2(n9012), .B1(n8997), .B2(n9010), .ZN(n8999)
         );
  AOI21_X1 U10360 ( .B1(n9001), .B2(n9000), .A(n8999), .ZN(n9155) );
  MUX2_X1 U10361 ( .A(n9155), .B(n9002), .S(n9037), .Z(n9005) );
  AOI22_X1 U10362 ( .A1(n9156), .A2(n4315), .B1(n9051), .B2(n9003), .ZN(n9004)
         );
  OAI211_X1 U10363 ( .C1(n9159), .C2(n9055), .A(n9005), .B(n9004), .ZN(
        P2_U3214) );
  XNOR2_X1 U10364 ( .A(n9006), .B(n9016), .ZN(n9008) );
  OAI222_X1 U10365 ( .A1(n9012), .A2(n9011), .B1(n9010), .B2(n9009), .C1(n9008), .C2(n9007), .ZN(n9095) );
  INV_X1 U10366 ( .A(n9095), .ZN(n9021) );
  INV_X1 U10367 ( .A(n9014), .ZN(n9015) );
  AOI21_X1 U10368 ( .B1(n9013), .B2(n9016), .A(n9015), .ZN(n9096) );
  AOI22_X1 U10369 ( .A1(n9037), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9051), .B2(
        n9017), .ZN(n9018) );
  OAI21_X1 U10370 ( .B1(n9164), .B2(n9028), .A(n9018), .ZN(n9019) );
  AOI21_X1 U10371 ( .B1(n9096), .B2(n9035), .A(n9019), .ZN(n9020) );
  OAI21_X1 U10372 ( .B1(n9021), .B2(n9037), .A(n9020), .ZN(P2_U3215) );
  XNOR2_X1 U10373 ( .A(n9022), .B(n9027), .ZN(n9025) );
  AOI222_X1 U10374 ( .A1(n9046), .A2(n9025), .B1(n9024), .B2(n9043), .C1(n9023), .C2(n9041), .ZN(n9103) );
  XNOR2_X1 U10375 ( .A(n9026), .B(n9027), .ZN(n9101) );
  NOR2_X1 U10376 ( .A1(n9029), .A2(n9028), .ZN(n9034) );
  OAI22_X1 U10377 ( .A1(n9047), .A2(n9032), .B1(n9031), .B2(n9030), .ZN(n9033)
         );
  AOI211_X1 U10378 ( .C1(n9101), .C2(n9035), .A(n9034), .B(n9033), .ZN(n9036)
         );
  OAI21_X1 U10379 ( .B1(n9103), .B2(n9037), .A(n9036), .ZN(P2_U3216) );
  XOR2_X1 U10380 ( .A(n9038), .B(n9040), .Z(n9172) );
  XOR2_X1 U10381 ( .A(n9039), .B(n9040), .Z(n9045) );
  AOI222_X1 U10382 ( .A1(n9046), .A2(n9045), .B1(n9044), .B2(n9043), .C1(n9042), .C2(n9041), .ZN(n9166) );
  MUX2_X1 U10383 ( .A(n9048), .B(n9166), .S(n9047), .Z(n9054) );
  INV_X1 U10384 ( .A(n9049), .ZN(n9050) );
  AOI22_X1 U10385 ( .A1(n9168), .A2(n4315), .B1(n9051), .B2(n9050), .ZN(n9053)
         );
  OAI211_X1 U10386 ( .C1(n9172), .C2(n9055), .A(n9054), .B(n9053), .ZN(
        P2_U3217) );
  NOR2_X1 U10387 ( .A1(n9056), .A2(n10003), .ZN(n9058) );
  AOI21_X1 U10388 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10003), .A(n9058), .ZN(
        n9057) );
  OAI21_X1 U10389 ( .B1(n9112), .B2(n9099), .A(n9057), .ZN(P2_U3490) );
  INV_X1 U10390 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U10391 ( .A1(n5843), .A2(n9105), .ZN(n9060) );
  INV_X1 U10392 ( .A(n9058), .ZN(n9059) );
  OAI211_X1 U10393 ( .C1(n10005), .C2(n9061), .A(n9060), .B(n9059), .ZN(
        P2_U3489) );
  NAND2_X1 U10394 ( .A1(n9062), .A2(n9987), .ZN(n9063) );
  OAI211_X1 U10395 ( .C1(n9982), .C2(n9065), .A(n9064), .B(n9063), .ZN(n9113)
         );
  MUX2_X1 U10396 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9113), .S(n10005), .Z(
        P2_U3487) );
  INV_X1 U10397 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9066) );
  MUX2_X1 U10398 ( .A(n9115), .B(n9066), .S(n10003), .Z(n9068) );
  NAND2_X1 U10399 ( .A1(n9116), .A2(n9105), .ZN(n9067) );
  OAI211_X1 U10400 ( .C1(n9119), .C2(n9108), .A(n9068), .B(n9067), .ZN(
        P2_U3486) );
  INV_X1 U10401 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9069) );
  MUX2_X1 U10402 ( .A(n9069), .B(n9120), .S(n10005), .Z(n9071) );
  NAND2_X1 U10403 ( .A1(n9122), .A2(n9105), .ZN(n9070) );
  OAI211_X1 U10404 ( .C1(n9125), .C2(n9108), .A(n9071), .B(n9070), .ZN(
        P2_U3485) );
  INV_X1 U10405 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9072) );
  MUX2_X1 U10406 ( .A(n9072), .B(n9126), .S(n10005), .Z(n9074) );
  NAND2_X1 U10407 ( .A1(n9127), .A2(n9105), .ZN(n9073) );
  OAI211_X1 U10408 ( .C1(n9108), .C2(n9130), .A(n9074), .B(n9073), .ZN(
        P2_U3484) );
  INV_X1 U10409 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9075) );
  MUX2_X1 U10410 ( .A(n9075), .B(n9131), .S(n10005), .Z(n9077) );
  NAND2_X1 U10411 ( .A1(n9133), .A2(n9105), .ZN(n9076) );
  OAI211_X1 U10412 ( .C1(n9108), .C2(n9136), .A(n9077), .B(n9076), .ZN(
        P2_U3483) );
  MUX2_X1 U10413 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9137), .S(n10005), .Z(
        n9079) );
  OAI22_X1 U10414 ( .A1(n9139), .A2(n9108), .B1(n9138), .B2(n9099), .ZN(n9078)
         );
  OR2_X1 U10415 ( .A1(n9079), .A2(n9078), .ZN(P2_U3482) );
  INV_X1 U10416 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9082) );
  AOI21_X1 U10417 ( .B1(n9949), .B2(n9081), .A(n9080), .ZN(n9142) );
  MUX2_X1 U10418 ( .A(n9082), .B(n9142), .S(n10005), .Z(n9083) );
  OAI21_X1 U10419 ( .B1(n9145), .B2(n9099), .A(n9083), .ZN(P2_U3481) );
  INV_X1 U10420 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9086) );
  AOI21_X1 U10421 ( .B1(n9987), .B2(n9085), .A(n9084), .ZN(n9146) );
  MUX2_X1 U10422 ( .A(n9086), .B(n9146), .S(n10005), .Z(n9087) );
  OAI21_X1 U10423 ( .B1(n9108), .B2(n9149), .A(n9087), .ZN(P2_U3480) );
  INV_X1 U10424 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9090) );
  AOI21_X1 U10425 ( .B1(n9987), .B2(n9089), .A(n9088), .ZN(n9150) );
  MUX2_X1 U10426 ( .A(n9090), .B(n9150), .S(n10005), .Z(n9091) );
  OAI21_X1 U10427 ( .B1(n9108), .B2(n9153), .A(n9091), .ZN(P2_U3479) );
  MUX2_X1 U10428 ( .A(n9155), .B(n9092), .S(n10003), .Z(n9094) );
  NAND2_X1 U10429 ( .A1(n9156), .A2(n9105), .ZN(n9093) );
  OAI211_X1 U10430 ( .C1(n9159), .C2(n9108), .A(n9094), .B(n9093), .ZN(
        P2_U3478) );
  AOI21_X1 U10431 ( .B1(n9096), .B2(n9949), .A(n9095), .ZN(n9160) );
  MUX2_X1 U10432 ( .A(n9097), .B(n9160), .S(n10005), .Z(n9098) );
  OAI21_X1 U10433 ( .B1(n9164), .B2(n9099), .A(n9098), .ZN(P2_U3477) );
  AOI22_X1 U10434 ( .A1(n9101), .A2(n9949), .B1(n9987), .B2(n9100), .ZN(n9102)
         );
  NAND2_X1 U10435 ( .A1(n9103), .A2(n9102), .ZN(n9165) );
  MUX2_X1 U10436 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9165), .S(n10005), .Z(
        P2_U3476) );
  MUX2_X1 U10437 ( .A(n9104), .B(n9166), .S(n10005), .Z(n9107) );
  NAND2_X1 U10438 ( .A1(n9168), .A2(n9105), .ZN(n9106) );
  OAI211_X1 U10439 ( .C1(n9172), .C2(n9108), .A(n9107), .B(n9106), .ZN(
        P2_U3475) );
  MUX2_X1 U10440 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9109), .S(n10005), .Z(
        P2_U3459) );
  AOI21_X1 U10441 ( .B1(n9990), .B2(P2_REG0_REG_31__SCAN_IN), .A(n9110), .ZN(
        n9111) );
  OAI21_X1 U10442 ( .B1(n9112), .B2(n9163), .A(n9111), .ZN(P2_U3458) );
  MUX2_X1 U10443 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9113), .S(n9988), .Z(
        P2_U3455) );
  INV_X1 U10444 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9114) );
  MUX2_X1 U10445 ( .A(n9115), .B(n9114), .S(n9990), .Z(n9118) );
  NAND2_X1 U10446 ( .A1(n9116), .A2(n6505), .ZN(n9117) );
  OAI211_X1 U10447 ( .C1(n9119), .C2(n9171), .A(n9118), .B(n9117), .ZN(
        P2_U3454) );
  INV_X1 U10448 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9121) );
  MUX2_X1 U10449 ( .A(n9121), .B(n9120), .S(n9988), .Z(n9124) );
  NAND2_X1 U10450 ( .A1(n9122), .A2(n6505), .ZN(n9123) );
  OAI211_X1 U10451 ( .C1(n9125), .C2(n9171), .A(n9124), .B(n9123), .ZN(
        P2_U3453) );
  MUX2_X1 U10452 ( .A(n10187), .B(n9126), .S(n9988), .Z(n9129) );
  NAND2_X1 U10453 ( .A1(n9127), .A2(n6505), .ZN(n9128) );
  OAI211_X1 U10454 ( .C1(n9130), .C2(n9171), .A(n9129), .B(n9128), .ZN(
        P2_U3452) );
  INV_X1 U10455 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9132) );
  MUX2_X1 U10456 ( .A(n9132), .B(n9131), .S(n9988), .Z(n9135) );
  NAND2_X1 U10457 ( .A1(n9133), .A2(n6505), .ZN(n9134) );
  OAI211_X1 U10458 ( .C1(n9136), .C2(n9171), .A(n9135), .B(n9134), .ZN(
        P2_U3451) );
  MUX2_X1 U10459 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9137), .S(n9988), .Z(n9141) );
  OAI22_X1 U10460 ( .A1(n9139), .A2(n9171), .B1(n9138), .B2(n9163), .ZN(n9140)
         );
  OR2_X1 U10461 ( .A1(n9141), .A2(n9140), .ZN(P2_U3450) );
  INV_X1 U10462 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9143) );
  MUX2_X1 U10463 ( .A(n9143), .B(n9142), .S(n9988), .Z(n9144) );
  OAI21_X1 U10464 ( .B1(n9145), .B2(n9163), .A(n9144), .ZN(P2_U3449) );
  INV_X1 U10465 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9147) );
  MUX2_X1 U10466 ( .A(n9147), .B(n9146), .S(n9988), .Z(n9148) );
  OAI21_X1 U10467 ( .B1(n9149), .B2(n9171), .A(n9148), .ZN(P2_U3448) );
  INV_X1 U10468 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9151) );
  MUX2_X1 U10469 ( .A(n9151), .B(n9150), .S(n9988), .Z(n9152) );
  OAI21_X1 U10470 ( .B1(n9153), .B2(n9171), .A(n9152), .ZN(P2_U3447) );
  INV_X1 U10471 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9154) );
  MUX2_X1 U10472 ( .A(n9155), .B(n9154), .S(n9990), .Z(n9158) );
  NAND2_X1 U10473 ( .A1(n9156), .A2(n6505), .ZN(n9157) );
  OAI211_X1 U10474 ( .C1(n9159), .C2(n9171), .A(n9158), .B(n9157), .ZN(
        P2_U3446) );
  MUX2_X1 U10475 ( .A(n9161), .B(n9160), .S(n9988), .Z(n9162) );
  OAI21_X1 U10476 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(P2_U3444) );
  MUX2_X1 U10477 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9165), .S(n9988), .Z(
        P2_U3441) );
  INV_X1 U10478 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9167) );
  MUX2_X1 U10479 ( .A(n9167), .B(n9166), .S(n9988), .Z(n9170) );
  NAND2_X1 U10480 ( .A1(n9168), .A2(n6505), .ZN(n9169) );
  OAI211_X1 U10481 ( .C1(n9172), .C2(n9171), .A(n9170), .B(n9169), .ZN(
        P2_U3438) );
  MUX2_X1 U10482 ( .A(n9174), .B(P2_D_REG_1__SCAN_IN), .S(n9173), .Z(P2_U3377)
         );
  INV_X1 U10483 ( .A(n9175), .ZN(n9785) );
  NOR4_X1 U10484 ( .A1(n9176), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9177), .ZN(n9179) );
  AOI21_X1 U10485 ( .B1(n9180), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9179), .ZN(
        n9181) );
  OAI21_X1 U10486 ( .B1(n9785), .B2(n8587), .A(n9181), .ZN(P2_U3264) );
  INV_X1 U10487 ( .A(n9182), .ZN(n9793) );
  OAI222_X1 U10488 ( .A1(n8587), .A2(n9793), .B1(n9184), .B2(P2_U3151), .C1(
        n9183), .C2(n8590), .ZN(P2_U3266) );
  NAND2_X1 U10489 ( .A1(n4397), .A2(n9186), .ZN(n9188) );
  XNOR2_X1 U10490 ( .A(n9188), .B(n9187), .ZN(n9196) );
  OAI22_X1 U10491 ( .A1(n9311), .A2(n9190), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9189), .ZN(n9193) );
  NOR2_X1 U10492 ( .A1(n9191), .A2(n9317), .ZN(n9192) );
  AOI211_X1 U10493 ( .C1(n9313), .C2(n9194), .A(n9193), .B(n9192), .ZN(n9195)
         );
  OAI21_X1 U10494 ( .B1(n9196), .B2(n9288), .A(n9195), .ZN(P1_U3215) );
  INV_X1 U10495 ( .A(n9198), .ZN(n9200) );
  NOR3_X1 U10496 ( .A1(n4910), .A2(n9200), .A3(n9199), .ZN(n9201) );
  OAI21_X1 U10497 ( .B1(n9201), .B2(n5575), .A(n9307), .ZN(n9207) );
  OR2_X1 U10498 ( .A1(n9221), .A2(n9409), .ZN(n9203) );
  NAND2_X1 U10499 ( .A1(n9324), .A2(n9435), .ZN(n9202) );
  NAND2_X1 U10500 ( .A1(n9203), .A2(n9202), .ZN(n9522) );
  OAI22_X1 U10501 ( .A1(n9524), .A2(n9299), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9204), .ZN(n9205) );
  AOI21_X1 U10502 ( .B1(n9522), .B2(n9301), .A(n9205), .ZN(n9206) );
  OAI211_X1 U10503 ( .C1(n9518), .C2(n9317), .A(n9207), .B(n9206), .ZN(
        P1_U3216) );
  OAI21_X1 U10504 ( .B1(n9210), .B2(n9209), .A(n9208), .ZN(n9216) );
  OAI22_X1 U10505 ( .A1(n9212), .A2(n9409), .B1(n9211), .B2(n9281), .ZN(n9549)
         );
  AOI22_X1 U10506 ( .A1(n9549), .A2(n9301), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9214) );
  NAND2_X1 U10507 ( .A1(n9313), .A2(n9553), .ZN(n9213) );
  OAI211_X1 U10508 ( .C1(n9745), .C2(n9317), .A(n9214), .B(n9213), .ZN(n9215)
         );
  AOI21_X1 U10509 ( .B1(n9216), .B2(n9307), .A(n9215), .ZN(n9217) );
  INV_X1 U10510 ( .A(n9217), .ZN(P1_U3223) );
  OAI21_X1 U10511 ( .B1(n9219), .B2(n9218), .A(n9291), .ZN(n9220) );
  NAND2_X1 U10512 ( .A1(n9220), .A2(n9307), .ZN(n9227) );
  OAI22_X1 U10513 ( .A1(n9222), .A2(n9409), .B1(n9221), .B2(n9281), .ZN(n9482)
         );
  INV_X1 U10514 ( .A(n9223), .ZN(n9488) );
  OAI22_X1 U10515 ( .A1(n9488), .A2(n9299), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9224), .ZN(n9225) );
  AOI21_X1 U10516 ( .B1(n9482), .B2(n9301), .A(n9225), .ZN(n9226) );
  OAI211_X1 U10517 ( .C1(n9731), .C2(n9317), .A(n9227), .B(n9226), .ZN(
        P1_U3225) );
  OAI21_X1 U10518 ( .B1(n9230), .B2(n9229), .A(n9228), .ZN(n9231) );
  NAND2_X1 U10519 ( .A1(n9231), .A2(n9307), .ZN(n9237) );
  AND2_X1 U10520 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9365) );
  INV_X1 U10521 ( .A(n9232), .ZN(n9233) );
  NOR2_X1 U10522 ( .A1(n9299), .A2(n9233), .ZN(n9234) );
  AOI211_X1 U10523 ( .C1(n9301), .C2(n9235), .A(n9365), .B(n9234), .ZN(n9236)
         );
  OAI211_X1 U10524 ( .C1(n9774), .C2(n9317), .A(n9237), .B(n9236), .ZN(
        P1_U3226) );
  OAI21_X1 U10525 ( .B1(n9240), .B2(n9239), .A(n9238), .ZN(n9241) );
  NAND2_X1 U10526 ( .A1(n9241), .A2(n9307), .ZN(n9247) );
  NOR2_X1 U10527 ( .A1(n9242), .A2(n9281), .ZN(n9243) );
  AOI21_X1 U10528 ( .B1(n9329), .B2(n9244), .A(n9243), .ZN(n9613) );
  NAND2_X1 U10529 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9376) );
  OAI21_X1 U10530 ( .B1(n9311), .B2(n9613), .A(n9376), .ZN(n9245) );
  AOI21_X1 U10531 ( .B1(n9619), .B2(n9313), .A(n9245), .ZN(n9246) );
  OAI211_X1 U10532 ( .C1(n9769), .C2(n9317), .A(n9247), .B(n9246), .ZN(
        P1_U3228) );
  NOR3_X1 U10533 ( .A1(n5575), .A2(n4597), .A3(n9249), .ZN(n9253) );
  BUF_X1 U10534 ( .A(n9250), .Z(n9251) );
  INV_X1 U10535 ( .A(n9251), .ZN(n9252) );
  OAI21_X1 U10536 ( .B1(n9253), .B2(n9252), .A(n9307), .ZN(n9259) );
  OAI22_X1 U10537 ( .A1(n9254), .A2(n9409), .B1(n9270), .B2(n9281), .ZN(n9507)
         );
  INV_X1 U10538 ( .A(n9255), .ZN(n9501) );
  OAI22_X1 U10539 ( .A1(n9501), .A2(n9299), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9256), .ZN(n9257) );
  AOI21_X1 U10540 ( .B1(n9507), .B2(n9301), .A(n9257), .ZN(n9258) );
  OAI211_X1 U10541 ( .C1(n9499), .C2(n9317), .A(n9259), .B(n9258), .ZN(
        P1_U3229) );
  OAI21_X1 U10542 ( .B1(n9262), .B2(n9261), .A(n9260), .ZN(n9266) );
  NOR2_X1 U10543 ( .A1(n9563), .A2(n9317), .ZN(n9265) );
  OAI22_X1 U10544 ( .A1(n9269), .A2(n9409), .B1(n9283), .B2(n9281), .ZN(n9570)
         );
  AOI22_X1 U10545 ( .A1(n9570), .A2(n9301), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9263) );
  OAI21_X1 U10546 ( .B1(n9564), .B2(n9299), .A(n9263), .ZN(n9264) );
  AOI211_X1 U10547 ( .C1(n9266), .C2(n9307), .A(n9265), .B(n9264), .ZN(n9267)
         );
  INV_X1 U10548 ( .A(n9267), .ZN(P1_U3233) );
  AOI21_X1 U10549 ( .B1(n9268), .B2(n9197), .A(n4910), .ZN(n9275) );
  OAI22_X1 U10550 ( .A1(n9270), .A2(n9409), .B1(n9269), .B2(n9281), .ZN(n9530)
         );
  OAI22_X1 U10551 ( .A1(n9538), .A2(n9299), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9271), .ZN(n9273) );
  NOR2_X1 U10552 ( .A1(n6597), .A2(n9317), .ZN(n9272) );
  AOI211_X1 U10553 ( .C1(n9301), .C2(n9530), .A(n9273), .B(n9272), .ZN(n9274)
         );
  OAI21_X1 U10554 ( .B1(n9275), .B2(n9288), .A(n9274), .ZN(P1_U3235) );
  INV_X1 U10555 ( .A(n9276), .ZN(n9278) );
  NAND2_X1 U10556 ( .A1(n9278), .A2(n9277), .ZN(n9279) );
  XNOR2_X1 U10557 ( .A(n9280), .B(n9279), .ZN(n9289) );
  OAI22_X1 U10558 ( .A1(n9283), .A2(n9409), .B1(n9282), .B2(n9281), .ZN(n9595)
         );
  AOI22_X1 U10559 ( .A1(n9595), .A2(n9301), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9284) );
  OAI21_X1 U10560 ( .B1(n9602), .B2(n9299), .A(n9284), .ZN(n9285) );
  AOI21_X1 U10561 ( .B1(n9684), .B2(n9286), .A(n9285), .ZN(n9287) );
  OAI21_X1 U10562 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(P1_U3238) );
  AND2_X1 U10563 ( .A1(n9291), .A2(n9290), .ZN(n9294) );
  OAI211_X1 U10564 ( .C1(n9294), .C2(n9293), .A(n9307), .B(n9292), .ZN(n9303)
         );
  OR2_X1 U10565 ( .A1(n9295), .A2(n9409), .ZN(n9297) );
  NAND2_X1 U10566 ( .A1(n9321), .A2(n9435), .ZN(n9296) );
  NAND2_X1 U10567 ( .A1(n9297), .A2(n9296), .ZN(n9474) );
  OAI22_X1 U10568 ( .A1(n9466), .A2(n9299), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9298), .ZN(n9300) );
  AOI21_X1 U10569 ( .B1(n9474), .B2(n9301), .A(n9300), .ZN(n9302) );
  OAI21_X1 U10570 ( .B1(n9306), .B2(n9305), .A(n9304), .ZN(n9308) );
  NAND2_X1 U10571 ( .A1(n9308), .A2(n9307), .ZN(n9316) );
  OAI22_X1 U10572 ( .A1(n9311), .A2(n9310), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9309), .ZN(n9312) );
  AOI21_X1 U10573 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9315) );
  OAI211_X1 U10574 ( .C1(n9318), .C2(n9317), .A(n9316), .B(n9315), .ZN(
        P1_U3241) );
  MUX2_X1 U10575 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9433), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10576 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9319), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10577 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n6558), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10578 ( .A(n9320), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9326), .Z(
        P1_U3580) );
  MUX2_X1 U10579 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9321), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10580 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9322), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10581 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9323), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10582 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9324), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10583 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9325), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10584 ( .A(n9327), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9326), .Z(
        P1_U3574) );
  MUX2_X1 U10585 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9328), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10586 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9329), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10587 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9330), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10588 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9331), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10589 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9332), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10590 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9333), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10591 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9334), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10592 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9335), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10593 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9336), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10594 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9337), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10595 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9338), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10596 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9339), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10597 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9340), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10598 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9341), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10599 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9342), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10600 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9343), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10601 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9344), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10602 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6524), .S(P1_U3973), .Z(
        P1_U3554) );
  AOI211_X1 U10603 ( .C1(n9347), .C2(n9346), .A(n9345), .B(n9387), .ZN(n9353)
         );
  INV_X1 U10604 ( .A(n9348), .ZN(n9349) );
  AOI211_X1 U10605 ( .C1(n9351), .C2(n9350), .A(n9349), .B(n9370), .ZN(n9352)
         );
  NOR2_X1 U10606 ( .A1(n9353), .A2(n9352), .ZN(n9358) );
  AOI22_X1 U10607 ( .A1(n9804), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9357) );
  NAND2_X1 U10608 ( .A1(n9367), .A2(n9354), .ZN(n9355) );
  NAND4_X1 U10609 ( .A1(n9358), .A2(n9357), .A3(n9356), .A4(n9355), .ZN(
        P1_U3245) );
  AOI211_X1 U10610 ( .C1(n9361), .C2(n9360), .A(n9359), .B(n9387), .ZN(n9373)
         );
  AOI21_X1 U10611 ( .B1(n9364), .B2(n9363), .A(n9362), .ZN(n9371) );
  AOI21_X1 U10612 ( .B1(n9804), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9365), .ZN(
        n9369) );
  NAND2_X1 U10613 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  OAI211_X1 U10614 ( .C1(n9371), .C2(n9370), .A(n9369), .B(n9368), .ZN(n9372)
         );
  OR2_X1 U10615 ( .A1(n9373), .A2(n9372), .ZN(P1_U3259) );
  XOR2_X1 U10616 ( .A(n9374), .B(n4343), .Z(n9385) );
  INV_X1 U10617 ( .A(n9375), .ZN(n9378) );
  NAND2_X1 U10618 ( .A1(n9804), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9377) );
  OAI211_X1 U10619 ( .C1(n9403), .C2(n9378), .A(n9377), .B(n9376), .ZN(n9379)
         );
  INV_X1 U10620 ( .A(n9379), .ZN(n9384) );
  NOR2_X1 U10621 ( .A1(n9381), .A2(n9380), .ZN(n9382) );
  OAI21_X1 U10622 ( .B1(n9396), .B2(n9382), .A(n9399), .ZN(n9383) );
  OAI211_X1 U10623 ( .C1(n9385), .C2(n9387), .A(n9384), .B(n9383), .ZN(
        P1_U3260) );
  INV_X1 U10624 ( .A(n9386), .ZN(n9402) );
  AND2_X1 U10625 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9392) );
  AOI211_X1 U10626 ( .C1(n9390), .C2(n9389), .A(n9388), .B(n9387), .ZN(n9391)
         );
  AOI211_X1 U10627 ( .C1(n9804), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9392), .B(
        n9391), .ZN(n9401) );
  INV_X1 U10628 ( .A(n9393), .ZN(n9398) );
  OAI21_X1 U10629 ( .B1(n9396), .B2(n9395), .A(n9394), .ZN(n9397) );
  NAND3_X1 U10630 ( .A1(n9399), .A2(n9398), .A3(n9397), .ZN(n9400) );
  OAI211_X1 U10631 ( .C1(n9403), .C2(n9402), .A(n9401), .B(n9400), .ZN(
        P1_U3261) );
  NOR2_X1 U10632 ( .A1(n9414), .A2(n9439), .ZN(n9405) );
  XOR2_X1 U10633 ( .A(n8320), .B(n9405), .Z(n9406) );
  NOR2_X1 U10634 ( .A1(n9406), .A2(n9616), .ZN(n9628) );
  NAND2_X1 U10635 ( .A1(n9628), .A2(n9828), .ZN(n9413) );
  NOR2_X1 U10636 ( .A1(n9796), .A2(n9407), .ZN(n9408) );
  NOR2_X1 U10637 ( .A1(n9409), .A2(n9408), .ZN(n9434) );
  INV_X1 U10638 ( .A(n9631), .ZN(n9411) );
  NOR2_X1 U10639 ( .A1(n9831), .A2(n9411), .ZN(n9417) );
  AOI21_X1 U10640 ( .B1(n9831), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9417), .ZN(
        n9412) );
  OAI211_X1 U10641 ( .C1(n9710), .C2(n9834), .A(n9413), .B(n9412), .ZN(
        P1_U3263) );
  XNOR2_X1 U10642 ( .A(n9414), .B(n9439), .ZN(n9415) );
  NAND2_X1 U10643 ( .A1(n9632), .A2(n9828), .ZN(n9419) );
  AND2_X1 U10644 ( .A1(n9620), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9416) );
  NOR2_X1 U10645 ( .A1(n9417), .A2(n9416), .ZN(n9418) );
  OAI211_X1 U10646 ( .C1(n9714), .C2(n9834), .A(n9419), .B(n9418), .ZN(
        P1_U3264) );
  NAND2_X1 U10647 ( .A1(n6559), .A2(n9420), .ZN(n9422) );
  NOR2_X1 U10648 ( .A1(n6559), .A2(n9420), .ZN(n9421) );
  AOI21_X1 U10649 ( .B1(n9423), .B2(n9422), .A(n9421), .ZN(n9424) );
  XNOR2_X1 U10650 ( .A(n9432), .B(n9424), .ZN(n9715) );
  NAND2_X1 U10651 ( .A1(n9715), .A2(n9838), .ZN(n9444) );
  OAI22_X1 U10652 ( .A1(n9426), .A2(n9601), .B1(n9425), .B2(n9624), .ZN(n9427)
         );
  AOI21_X1 U10653 ( .B1(n9404), .B2(n9590), .A(n9427), .ZN(n9443) );
  INV_X1 U10654 ( .A(n9428), .ZN(n9430) );
  AOI22_X1 U10655 ( .A1(n6558), .A2(n9435), .B1(n9434), .B2(n9433), .ZN(n9436)
         );
  NAND2_X1 U10656 ( .A1(n9636), .A2(n9624), .ZN(n9442) );
  AOI21_X1 U10657 ( .B1(n9404), .B2(n9438), .A(n9616), .ZN(n9440) );
  NAND2_X1 U10658 ( .A1(n9635), .A2(n9828), .ZN(n9441) );
  NAND4_X1 U10659 ( .A1(n9444), .A2(n9443), .A3(n9442), .A4(n9441), .ZN(
        P1_U3356) );
  XNOR2_X1 U10660 ( .A(n9445), .B(n9451), .ZN(n9722) );
  INV_X1 U10661 ( .A(n9722), .ZN(n9460) );
  AOI211_X1 U10662 ( .C1(n9720), .C2(n9463), .A(n9616), .B(n4340), .ZN(n9642)
         );
  NOR2_X1 U10663 ( .A1(n9446), .A2(n9834), .ZN(n9450) );
  OAI22_X1 U10664 ( .A1(n9448), .A2(n9601), .B1(n9447), .B2(n9624), .ZN(n9449)
         );
  AOI211_X1 U10665 ( .C1(n9642), .C2(n9828), .A(n9450), .B(n9449), .ZN(n9459)
         );
  OAI21_X1 U10666 ( .B1(n9471), .B2(n9452), .A(n9451), .ZN(n9453) );
  NAND3_X1 U10667 ( .A1(n9454), .A2(n9453), .A3(n9609), .ZN(n9457) );
  INV_X1 U10668 ( .A(n9455), .ZN(n9456) );
  NAND2_X1 U10669 ( .A1(n9457), .A2(n9456), .ZN(n9641) );
  NAND2_X1 U10670 ( .A1(n9641), .A2(n9624), .ZN(n9458) );
  OAI211_X1 U10671 ( .C1(n9460), .C2(n9626), .A(n9459), .B(n9458), .ZN(
        P1_U3266) );
  XOR2_X1 U10672 ( .A(n9470), .B(n9461), .Z(n9730) );
  INV_X1 U10673 ( .A(n9462), .ZN(n9490) );
  INV_X1 U10674 ( .A(n9463), .ZN(n9464) );
  AOI211_X1 U10675 ( .C1(n9648), .C2(n9490), .A(n9616), .B(n9464), .ZN(n9647)
         );
  NOR2_X1 U10676 ( .A1(n6598), .A2(n9834), .ZN(n9468) );
  OAI22_X1 U10677 ( .A1(n9466), .A2(n9601), .B1(n9465), .B2(n9624), .ZN(n9467)
         );
  AOI211_X1 U10678 ( .C1(n9647), .C2(n9828), .A(n9468), .B(n9467), .ZN(n9478)
         );
  INV_X1 U10679 ( .A(n9469), .ZN(n9473) );
  INV_X1 U10680 ( .A(n9470), .ZN(n9472) );
  AOI21_X1 U10681 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(n9476) );
  INV_X1 U10682 ( .A(n9474), .ZN(n9475) );
  OAI21_X1 U10683 ( .B1(n9476), .B2(n9846), .A(n9475), .ZN(n9646) );
  NAND2_X1 U10684 ( .A1(n9646), .A2(n9624), .ZN(n9477) );
  OAI211_X1 U10685 ( .C1(n9730), .C2(n9626), .A(n9478), .B(n9477), .ZN(
        P1_U3267) );
  INV_X1 U10686 ( .A(n9484), .ZN(n9481) );
  NAND2_X1 U10687 ( .A1(n9506), .A2(n9479), .ZN(n9480) );
  XNOR2_X1 U10688 ( .A(n9481), .B(n9480), .ZN(n9483) );
  AOI21_X1 U10689 ( .B1(n9483), .B2(n9609), .A(n9482), .ZN(n9652) );
  XNOR2_X1 U10690 ( .A(n9485), .B(n9484), .ZN(n9732) );
  INV_X1 U10691 ( .A(n9732), .ZN(n9486) );
  NAND2_X1 U10692 ( .A1(n9486), .A2(n9838), .ZN(n9495) );
  OAI22_X1 U10693 ( .A1(n9488), .A2(n9601), .B1(n9487), .B2(n9624), .ZN(n9492)
         );
  INV_X1 U10694 ( .A(n9489), .ZN(n9497) );
  OAI211_X1 U10695 ( .C1(n9497), .C2(n9731), .A(n9584), .B(n9490), .ZN(n9651)
         );
  NOR2_X1 U10696 ( .A1(n9651), .A2(n9586), .ZN(n9491) );
  AOI211_X1 U10697 ( .C1(n9590), .C2(n9493), .A(n9492), .B(n9491), .ZN(n9494)
         );
  OAI211_X1 U10698 ( .C1(n9831), .C2(n9652), .A(n9495), .B(n9494), .ZN(
        P1_U3268) );
  XOR2_X1 U10699 ( .A(n9496), .B(n9504), .Z(n9739) );
  INV_X1 U10700 ( .A(n9516), .ZN(n9498) );
  AOI211_X1 U10701 ( .C1(n6564), .C2(n9498), .A(n9616), .B(n9497), .ZN(n9655)
         );
  NOR2_X1 U10702 ( .A1(n9499), .A2(n9834), .ZN(n9503) );
  OAI22_X1 U10703 ( .A1(n9501), .A2(n9601), .B1(n9500), .B2(n9624), .ZN(n9502)
         );
  AOI211_X1 U10704 ( .C1(n9655), .C2(n9828), .A(n9503), .B(n9502), .ZN(n9512)
         );
  AOI21_X1 U10705 ( .B1(n9505), .B2(n9521), .A(n9504), .ZN(n9510) );
  NAND2_X1 U10706 ( .A1(n9506), .A2(n9609), .ZN(n9509) );
  INV_X1 U10707 ( .A(n9507), .ZN(n9508) );
  OAI21_X1 U10708 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9656) );
  NAND2_X1 U10709 ( .A1(n9656), .A2(n9624), .ZN(n9511) );
  OAI211_X1 U10710 ( .C1(n9739), .C2(n9626), .A(n9512), .B(n9511), .ZN(
        P1_U3269) );
  XOR2_X1 U10711 ( .A(n9513), .B(n9520), .Z(n9662) );
  NAND2_X1 U10712 ( .A1(n6589), .A2(n9535), .ZN(n9514) );
  NAND2_X1 U10713 ( .A1(n9514), .A2(n9584), .ZN(n9515) );
  NOR2_X1 U10714 ( .A1(n9516), .A2(n9515), .ZN(n9659) );
  OAI22_X1 U10715 ( .A1(n9518), .A2(n9834), .B1(n9517), .B2(n9624), .ZN(n9519)
         );
  AOI21_X1 U10716 ( .B1(n9659), .B2(n9828), .A(n9519), .ZN(n9527) );
  OAI21_X1 U10717 ( .B1(n4354), .B2(n4639), .A(n9521), .ZN(n9523) );
  AOI21_X1 U10718 ( .B1(n9523), .B2(n9609), .A(n9522), .ZN(n9661) );
  OAI21_X1 U10719 ( .B1(n9524), .B2(n9601), .A(n9661), .ZN(n9525) );
  NAND2_X1 U10720 ( .A1(n9525), .A2(n9624), .ZN(n9526) );
  OAI211_X1 U10721 ( .C1(n9662), .C2(n9626), .A(n9527), .B(n9526), .ZN(
        P1_U3270) );
  XNOR2_X1 U10722 ( .A(n9529), .B(n9528), .ZN(n9531) );
  AOI21_X1 U10723 ( .B1(n9531), .B2(n9609), .A(n9530), .ZN(n9664) );
  XNOR2_X1 U10724 ( .A(n9533), .B(n9532), .ZN(n9743) );
  INV_X1 U10725 ( .A(n9534), .ZN(n9552) );
  AOI21_X1 U10726 ( .B1(n9540), .B2(n9552), .A(n9616), .ZN(n9536) );
  NAND2_X1 U10727 ( .A1(n9536), .A2(n9535), .ZN(n9663) );
  OAI22_X1 U10728 ( .A1(n9538), .A2(n9601), .B1(n9537), .B2(n9624), .ZN(n9539)
         );
  AOI21_X1 U10729 ( .B1(n9540), .B2(n9590), .A(n9539), .ZN(n9541) );
  OAI21_X1 U10730 ( .B1(n9663), .B2(n9586), .A(n9541), .ZN(n9542) );
  AOI21_X1 U10731 ( .B1(n9743), .B2(n9838), .A(n9542), .ZN(n9543) );
  OAI21_X1 U10732 ( .B1(n9831), .B2(n9664), .A(n9543), .ZN(P1_U3271) );
  XNOR2_X1 U10733 ( .A(n9544), .B(n9545), .ZN(n9746) );
  NAND2_X1 U10734 ( .A1(n9546), .A2(n9545), .ZN(n9547) );
  NAND2_X1 U10735 ( .A1(n9548), .A2(n9547), .ZN(n9550) );
  AOI21_X1 U10736 ( .B1(n9550), .B2(n9609), .A(n9549), .ZN(n9668) );
  INV_X1 U10737 ( .A(n9668), .ZN(n9558) );
  INV_X1 U10738 ( .A(n9551), .ZN(n9562) );
  OAI211_X1 U10739 ( .C1(n9745), .C2(n9562), .A(n9584), .B(n9552), .ZN(n9667)
         );
  AOI22_X1 U10740 ( .A1(n9553), .A2(n9830), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9831), .ZN(n9556) );
  NAND2_X1 U10741 ( .A1(n9554), .A2(n9590), .ZN(n9555) );
  OAI211_X1 U10742 ( .C1(n9667), .C2(n9586), .A(n9556), .B(n9555), .ZN(n9557)
         );
  AOI21_X1 U10743 ( .B1(n9558), .B2(n9624), .A(n9557), .ZN(n9559) );
  OAI21_X1 U10744 ( .B1(n9746), .B2(n9626), .A(n9559), .ZN(P1_U3272) );
  XNOR2_X1 U10745 ( .A(n9560), .B(n9568), .ZN(n9753) );
  INV_X1 U10746 ( .A(n9561), .ZN(n9585) );
  AOI211_X1 U10747 ( .C1(n9673), .C2(n9585), .A(n9616), .B(n9562), .ZN(n9671)
         );
  NOR2_X1 U10748 ( .A1(n9563), .A2(n9834), .ZN(n9567) );
  OAI22_X1 U10749 ( .A1(n9624), .A2(n9565), .B1(n9564), .B2(n9601), .ZN(n9566)
         );
  AOI211_X1 U10750 ( .C1(n9671), .C2(n9828), .A(n9567), .B(n9566), .ZN(n9574)
         );
  XNOR2_X1 U10751 ( .A(n9569), .B(n9568), .ZN(n9572) );
  INV_X1 U10752 ( .A(n9570), .ZN(n9571) );
  OAI21_X1 U10753 ( .B1(n9572), .B2(n9846), .A(n9571), .ZN(n9672) );
  NAND2_X1 U10754 ( .A1(n9672), .A2(n9624), .ZN(n9573) );
  OAI211_X1 U10755 ( .C1(n9753), .C2(n9626), .A(n9574), .B(n9573), .ZN(
        P1_U3273) );
  XNOR2_X1 U10756 ( .A(n9575), .B(n9579), .ZN(n9577) );
  AOI21_X1 U10757 ( .B1(n9577), .B2(n9609), .A(n9576), .ZN(n9677) );
  XNOR2_X1 U10758 ( .A(n9578), .B(n9579), .ZN(n9755) );
  INV_X1 U10759 ( .A(n9755), .ZN(n9580) );
  NAND2_X1 U10760 ( .A1(n9580), .A2(n9838), .ZN(n9592) );
  OAI22_X1 U10761 ( .A1(n9624), .A2(n9582), .B1(n9581), .B2(n9601), .ZN(n9588)
         );
  INV_X1 U10762 ( .A(n9583), .ZN(n9600) );
  OAI211_X1 U10763 ( .C1(n9754), .C2(n9600), .A(n9585), .B(n9584), .ZN(n9676)
         );
  NOR2_X1 U10764 ( .A1(n9676), .A2(n9586), .ZN(n9587) );
  AOI211_X1 U10765 ( .C1(n9590), .C2(n9589), .A(n9588), .B(n9587), .ZN(n9591)
         );
  OAI211_X1 U10766 ( .C1(n9831), .C2(n9677), .A(n9592), .B(n9591), .ZN(
        P1_U3274) );
  OAI21_X1 U10767 ( .B1(n4393), .B2(n9594), .A(n9593), .ZN(n9596) );
  AOI21_X1 U10768 ( .B1(n9596), .B2(n9609), .A(n9595), .ZN(n9681) );
  XNOR2_X1 U10769 ( .A(n9598), .B(n9597), .ZN(n9680) );
  NAND2_X1 U10770 ( .A1(n9680), .A2(n9838), .ZN(n9607) );
  AOI211_X1 U10771 ( .C1(n9684), .C2(n9615), .A(n9616), .B(n9600), .ZN(n9683)
         );
  NOR2_X1 U10772 ( .A1(n6596), .A2(n9834), .ZN(n9605) );
  OAI22_X1 U10773 ( .A1(n9624), .A2(n9603), .B1(n9602), .B2(n9601), .ZN(n9604)
         );
  AOI211_X1 U10774 ( .C1(n9683), .C2(n9828), .A(n9605), .B(n9604), .ZN(n9606)
         );
  OAI211_X1 U10775 ( .C1(n9831), .C2(n9681), .A(n9607), .B(n9606), .ZN(
        P1_U3275) );
  XNOR2_X1 U10776 ( .A(n9608), .B(n9612), .ZN(n9764) );
  INV_X1 U10777 ( .A(n9764), .ZN(n9627) );
  OAI211_X1 U10778 ( .C1(n9612), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9614)
         );
  NAND2_X1 U10779 ( .A1(n9614), .A2(n9613), .ZN(n9689) );
  AOI211_X1 U10780 ( .C1(n9618), .C2(n9617), .A(n9616), .B(n9599), .ZN(n9690)
         );
  NAND2_X1 U10781 ( .A1(n9690), .A2(n9828), .ZN(n9622) );
  AOI22_X1 U10782 ( .A1(n9620), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9619), .B2(
        n9830), .ZN(n9621) );
  OAI211_X1 U10783 ( .C1(n9769), .C2(n9834), .A(n9622), .B(n9621), .ZN(n9623)
         );
  AOI21_X1 U10784 ( .B1(n9624), .B2(n9689), .A(n9623), .ZN(n9625) );
  OAI21_X1 U10785 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(P1_U3276) );
  INV_X1 U10786 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9629) );
  NOR2_X1 U10787 ( .A1(n9628), .A2(n9631), .ZN(n9707) );
  MUX2_X1 U10788 ( .A(n9629), .B(n9707), .S(n9876), .Z(n9630) );
  OAI21_X1 U10789 ( .B1(n9710), .B2(n9699), .A(n9630), .ZN(P1_U3553) );
  INV_X1 U10790 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9633) );
  NOR2_X1 U10791 ( .A1(n9632), .A2(n9631), .ZN(n9711) );
  MUX2_X1 U10792 ( .A(n9633), .B(n9711), .S(n9876), .Z(n9634) );
  OAI21_X1 U10793 ( .B1(n9714), .B2(n9699), .A(n9634), .ZN(P1_U3552) );
  AOI22_X1 U10794 ( .A1(n9715), .A2(n9688), .B1(n9640), .B2(n9404), .ZN(n9639)
         );
  INV_X1 U10795 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9637) );
  NOR2_X1 U10796 ( .A1(n9636), .A2(n9635), .ZN(n9716) );
  NAND2_X1 U10797 ( .A1(n9639), .A2(n9638), .ZN(P1_U3551) );
  AOI22_X1 U10798 ( .A1(n9722), .A2(n9688), .B1(n9640), .B2(n9720), .ZN(n9645)
         );
  INV_X1 U10799 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9643) );
  NOR2_X1 U10800 ( .A1(n9642), .A2(n9641), .ZN(n9723) );
  MUX2_X1 U10801 ( .A(n9643), .B(n9723), .S(n9876), .Z(n9644) );
  NAND2_X1 U10802 ( .A1(n9645), .A2(n9644), .ZN(P1_U3549) );
  INV_X1 U10803 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9649) );
  AOI211_X1 U10804 ( .C1(n9860), .C2(n9648), .A(n9647), .B(n9646), .ZN(n9727)
         );
  MUX2_X1 U10805 ( .A(n9649), .B(n9727), .S(n9876), .Z(n9650) );
  OAI21_X1 U10806 ( .B1(n9730), .B2(n9687), .A(n9650), .ZN(P1_U3548) );
  OAI22_X1 U10807 ( .A1(n9732), .A2(n9687), .B1(n9731), .B2(n9699), .ZN(n9654)
         );
  NAND2_X1 U10808 ( .A1(n9652), .A2(n9651), .ZN(n9733) );
  MUX2_X1 U10809 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9733), .S(n9876), .Z(n9653) );
  OR2_X1 U10810 ( .A1(n9654), .A2(n9653), .ZN(P1_U3547) );
  INV_X1 U10811 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9657) );
  AOI211_X1 U10812 ( .C1(n9860), .C2(n6564), .A(n9656), .B(n9655), .ZN(n9736)
         );
  MUX2_X1 U10813 ( .A(n9657), .B(n9736), .S(n9876), .Z(n9658) );
  OAI21_X1 U10814 ( .B1(n9739), .B2(n9687), .A(n9658), .ZN(P1_U3546) );
  AOI21_X1 U10815 ( .B1(n9860), .B2(n6589), .A(n9659), .ZN(n9660) );
  OAI211_X1 U10816 ( .C1(n9662), .C2(n9845), .A(n9661), .B(n9660), .ZN(n9740)
         );
  MUX2_X1 U10817 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9740), .S(n9876), .Z(
        P1_U3545) );
  OAI211_X1 U10818 ( .C1(n6597), .C2(n9853), .A(n9664), .B(n9663), .ZN(n9741)
         );
  MUX2_X1 U10819 ( .A(n9741), .B(P1_REG1_REG_22__SCAN_IN), .S(n9874), .Z(n9665) );
  AOI21_X1 U10820 ( .B1(n9743), .B2(n9688), .A(n9665), .ZN(n9666) );
  INV_X1 U10821 ( .A(n9666), .ZN(P1_U3544) );
  OAI22_X1 U10822 ( .A1(n9746), .A2(n9687), .B1(n9745), .B2(n9699), .ZN(n9670)
         );
  NAND2_X1 U10823 ( .A1(n9668), .A2(n9667), .ZN(n9747) );
  MUX2_X1 U10824 ( .A(n9747), .B(P1_REG1_REG_21__SCAN_IN), .S(n9874), .Z(n9669) );
  OR2_X1 U10825 ( .A1(n9670), .A2(n9669), .ZN(P1_U3543) );
  INV_X1 U10826 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9674) );
  AOI211_X1 U10827 ( .C1(n9860), .C2(n9673), .A(n9672), .B(n9671), .ZN(n9750)
         );
  MUX2_X1 U10828 ( .A(n9674), .B(n9750), .S(n9876), .Z(n9675) );
  OAI21_X1 U10829 ( .B1(n9753), .B2(n9687), .A(n9675), .ZN(P1_U3542) );
  OAI22_X1 U10830 ( .A1(n9755), .A2(n9687), .B1(n9754), .B2(n9699), .ZN(n9679)
         );
  NAND2_X1 U10831 ( .A1(n9677), .A2(n9676), .ZN(n9756) );
  MUX2_X1 U10832 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9756), .S(n9876), .Z(n9678) );
  OR2_X1 U10833 ( .A1(n9679), .A2(n9678), .ZN(P1_U3541) );
  INV_X1 U10834 ( .A(n9680), .ZN(n9762) );
  INV_X1 U10835 ( .A(n9681), .ZN(n9682) );
  AOI211_X1 U10836 ( .C1(n9860), .C2(n9684), .A(n9683), .B(n9682), .ZN(n9759)
         );
  MUX2_X1 U10837 ( .A(n9685), .B(n9759), .S(n9876), .Z(n9686) );
  OAI21_X1 U10838 ( .B1(n9762), .B2(n9687), .A(n9686), .ZN(P1_U3540) );
  NAND2_X1 U10839 ( .A1(n9764), .A2(n9688), .ZN(n9693) );
  NOR2_X1 U10840 ( .A1(n9690), .A2(n9689), .ZN(n9765) );
  MUX2_X1 U10841 ( .A(n9691), .B(n9765), .S(n9876), .Z(n9692) );
  OAI211_X1 U10842 ( .C1(n9769), .C2(n9699), .A(n9693), .B(n9692), .ZN(
        P1_U3539) );
  AOI211_X1 U10843 ( .C1(n9696), .C2(n9858), .A(n9695), .B(n9694), .ZN(n9770)
         );
  MUX2_X1 U10844 ( .A(n9697), .B(n9770), .S(n9876), .Z(n9698) );
  OAI21_X1 U10845 ( .B1(n9774), .B2(n9699), .A(n9698), .ZN(P1_U3538) );
  INV_X1 U10846 ( .A(n9700), .ZN(n9705) );
  AOI21_X1 U10847 ( .B1(n9860), .B2(n9702), .A(n9701), .ZN(n9703) );
  OAI211_X1 U10848 ( .C1(n9706), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9775)
         );
  MUX2_X1 U10849 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9775), .S(n9876), .Z(
        P1_U3536) );
  INV_X1 U10850 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9708) );
  MUX2_X1 U10851 ( .A(n9708), .B(n9707), .S(n9869), .Z(n9709) );
  OAI21_X1 U10852 ( .B1(n9710), .B2(n9773), .A(n9709), .ZN(P1_U3521) );
  MUX2_X1 U10853 ( .A(n9712), .B(n9711), .S(n9869), .Z(n9713) );
  OAI21_X1 U10854 ( .B1(n9714), .B2(n9773), .A(n9713), .ZN(P1_U3520) );
  AOI22_X1 U10855 ( .A1(n9715), .A2(n9763), .B1(n9721), .B2(n9404), .ZN(n9719)
         );
  INV_X1 U10856 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U10857 ( .A1(n9719), .A2(n9718), .ZN(P1_U3519) );
  AOI22_X1 U10858 ( .A1(n9722), .A2(n9763), .B1(n9721), .B2(n9720), .ZN(n9726)
         );
  INV_X1 U10859 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9724) );
  MUX2_X1 U10860 ( .A(n9724), .B(n9723), .S(n9869), .Z(n9725) );
  NAND2_X1 U10861 ( .A1(n9726), .A2(n9725), .ZN(P1_U3517) );
  INV_X1 U10862 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9728) );
  MUX2_X1 U10863 ( .A(n9728), .B(n9727), .S(n9869), .Z(n9729) );
  OAI21_X1 U10864 ( .B1(n9730), .B2(n9761), .A(n9729), .ZN(P1_U3516) );
  OAI22_X1 U10865 ( .A1(n9732), .A2(n9761), .B1(n9731), .B2(n9773), .ZN(n9735)
         );
  MUX2_X1 U10866 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9733), .S(n9869), .Z(n9734) );
  OR2_X1 U10867 ( .A1(n9735), .A2(n9734), .ZN(P1_U3515) );
  INV_X1 U10868 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9737) );
  MUX2_X1 U10869 ( .A(n9737), .B(n9736), .S(n9869), .Z(n9738) );
  OAI21_X1 U10870 ( .B1(n9739), .B2(n9761), .A(n9738), .ZN(P1_U3514) );
  MUX2_X1 U10871 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9740), .S(n9869), .Z(
        P1_U3513) );
  MUX2_X1 U10872 ( .A(n9741), .B(P1_REG0_REG_22__SCAN_IN), .S(n9867), .Z(n9742) );
  AOI21_X1 U10873 ( .B1(n9743), .B2(n9763), .A(n9742), .ZN(n9744) );
  INV_X1 U10874 ( .A(n9744), .ZN(P1_U3512) );
  OAI22_X1 U10875 ( .A1(n9746), .A2(n9761), .B1(n9745), .B2(n9773), .ZN(n9749)
         );
  MUX2_X1 U10876 ( .A(n9747), .B(P1_REG0_REG_21__SCAN_IN), .S(n9867), .Z(n9748) );
  OR2_X1 U10877 ( .A1(n9749), .A2(n9748), .ZN(P1_U3511) );
  INV_X1 U10878 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9751) );
  MUX2_X1 U10879 ( .A(n9751), .B(n9750), .S(n9869), .Z(n9752) );
  OAI21_X1 U10880 ( .B1(n9753), .B2(n9761), .A(n9752), .ZN(P1_U3510) );
  OAI22_X1 U10881 ( .A1(n9755), .A2(n9761), .B1(n9754), .B2(n9773), .ZN(n9758)
         );
  MUX2_X1 U10882 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9756), .S(n9869), .Z(n9757) );
  OR2_X1 U10883 ( .A1(n9758), .A2(n9757), .ZN(P1_U3509) );
  MUX2_X1 U10884 ( .A(n10202), .B(n9759), .S(n9869), .Z(n9760) );
  OAI21_X1 U10885 ( .B1(n9762), .B2(n9761), .A(n9760), .ZN(P1_U3507) );
  NAND2_X1 U10886 ( .A1(n9764), .A2(n9763), .ZN(n9768) );
  INV_X1 U10887 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9766) );
  MUX2_X1 U10888 ( .A(n9766), .B(n9765), .S(n9869), .Z(n9767) );
  OAI211_X1 U10889 ( .C1(n9769), .C2(n9773), .A(n9768), .B(n9767), .ZN(
        P1_U3504) );
  MUX2_X1 U10890 ( .A(n9771), .B(n9770), .S(n9869), .Z(n9772) );
  OAI21_X1 U10891 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(P1_U3501) );
  MUX2_X1 U10892 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9775), .S(n9869), .Z(
        P1_U3495) );
  MUX2_X1 U10893 ( .A(P1_D_REG_1__SCAN_IN), .B(n9778), .S(n9841), .Z(P1_U3440)
         );
  MUX2_X1 U10894 ( .A(P1_D_REG_0__SCAN_IN), .B(n9779), .S(n9841), .Z(P1_U3439)
         );
  NAND3_X1 U10895 ( .A1(n9781), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9782) );
  NOR4_X1 U10896 ( .A1(n9780), .A2(P1_IR_REG_30__SCAN_IN), .A3(
        P1_IR_REG_28__SCAN_IN), .A4(n9782), .ZN(n9783) );
  AOI21_X1 U10897 ( .B1(n9790), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9783), .ZN(
        n9784) );
  OAI21_X1 U10898 ( .B1(n9785), .B2(n9792), .A(n9784), .ZN(P1_U3324) );
  AOI22_X1 U10899 ( .A1(n9787), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9786), .ZN(n9788) );
  OAI21_X1 U10900 ( .B1(n9789), .B2(n9792), .A(n9788), .ZN(P1_U3325) );
  AOI22_X1 U10901 ( .A1(n5034), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9790), .ZN(n9791) );
  OAI21_X1 U10902 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(P1_U3326) );
  INV_X1 U10903 ( .A(n9794), .ZN(n9795) );
  MUX2_X1 U10904 ( .A(n9795), .B(n9798), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U10905 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10906 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10907 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9870) );
  AND2_X1 U10908 ( .A1(n9796), .A2(n9870), .ZN(n9800) );
  NOR2_X1 U10909 ( .A1(n9797), .A2(n9800), .ZN(n9799) );
  MUX2_X1 U10910 ( .A(n9800), .B(n9799), .S(n9798), .Z(n9803) );
  INV_X1 U10911 ( .A(n9801), .ZN(n9802) );
  OR2_X1 U10912 ( .A1(n9803), .A2(n9802), .ZN(n9806) );
  AOI22_X1 U10913 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9804), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9805) );
  OAI21_X1 U10914 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(P1_U3243) );
  AOI22_X1 U10915 ( .A1(n9831), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n9808), .B2(
        n9830), .ZN(n9809) );
  OAI21_X1 U10916 ( .B1(n9834), .B2(n9810), .A(n9809), .ZN(n9811) );
  INV_X1 U10917 ( .A(n9811), .ZN(n9816) );
  AOI22_X1 U10918 ( .A1(n9814), .A2(n9813), .B1(n9828), .B2(n9812), .ZN(n9815)
         );
  OAI211_X1 U10919 ( .C1(n9620), .C2(n9817), .A(n9816), .B(n9815), .ZN(
        P1_U3286) );
  INV_X1 U10920 ( .A(n9818), .ZN(n9823) );
  NAND2_X1 U10921 ( .A1(n9819), .A2(n9828), .ZN(n9822) );
  AOI22_X1 U10922 ( .A1(n9831), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9820), .B2(
        n9830), .ZN(n9821) );
  OAI211_X1 U10923 ( .C1(n9823), .C2(n9834), .A(n9822), .B(n9821), .ZN(n9824)
         );
  AOI21_X1 U10924 ( .B1(n9825), .B2(n9838), .A(n9824), .ZN(n9826) );
  OAI21_X1 U10925 ( .B1(n9620), .B2(n9827), .A(n9826), .ZN(P1_U3287) );
  NAND2_X1 U10926 ( .A1(n9829), .A2(n9828), .ZN(n9833) );
  AOI22_X1 U10927 ( .A1(n9831), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9830), .ZN(n9832) );
  OAI211_X1 U10928 ( .C1(n9835), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9836)
         );
  AOI21_X1 U10929 ( .B1(n9838), .B2(n9837), .A(n9836), .ZN(n9839) );
  OAI21_X1 U10930 ( .B1(n9620), .B2(n9840), .A(n9839), .ZN(P1_U3291) );
  AND2_X1 U10931 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9842), .ZN(P1_U3294) );
  INV_X1 U10932 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10169) );
  NOR2_X1 U10933 ( .A1(n9841), .A2(n10169), .ZN(P1_U3295) );
  AND2_X1 U10934 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9842), .ZN(P1_U3296) );
  AND2_X1 U10935 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9842), .ZN(P1_U3297) );
  AND2_X1 U10936 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9842), .ZN(P1_U3298) );
  AND2_X1 U10937 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9842), .ZN(P1_U3299) );
  AND2_X1 U10938 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9842), .ZN(P1_U3300) );
  AND2_X1 U10939 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9842), .ZN(P1_U3301) );
  AND2_X1 U10940 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9842), .ZN(P1_U3302) );
  AND2_X1 U10941 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9842), .ZN(P1_U3303) );
  AND2_X1 U10942 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9842), .ZN(P1_U3304) );
  AND2_X1 U10943 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9842), .ZN(P1_U3305) );
  AND2_X1 U10944 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9842), .ZN(P1_U3306) );
  INV_X1 U10945 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10183) );
  NOR2_X1 U10946 ( .A1(n9841), .A2(n10183), .ZN(P1_U3307) );
  INV_X1 U10947 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U10948 ( .A1(n9841), .A2(n10031), .ZN(P1_U3308) );
  INV_X1 U10949 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10182) );
  NOR2_X1 U10950 ( .A1(n9841), .A2(n10182), .ZN(P1_U3309) );
  AND2_X1 U10951 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9842), .ZN(P1_U3310) );
  AND2_X1 U10952 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9842), .ZN(P1_U3311) );
  AND2_X1 U10953 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9842), .ZN(P1_U3312) );
  AND2_X1 U10954 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9842), .ZN(P1_U3313) );
  AND2_X1 U10955 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9842), .ZN(P1_U3314) );
  AND2_X1 U10956 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9842), .ZN(P1_U3315) );
  AND2_X1 U10957 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9842), .ZN(P1_U3316) );
  AND2_X1 U10958 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9842), .ZN(P1_U3317) );
  AND2_X1 U10959 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9842), .ZN(P1_U3318) );
  AND2_X1 U10960 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9842), .ZN(P1_U3319) );
  AND2_X1 U10961 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9842), .ZN(P1_U3320) );
  AND2_X1 U10962 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9842), .ZN(P1_U3321) );
  AND2_X1 U10963 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9842), .ZN(P1_U3322) );
  AND2_X1 U10964 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9842), .ZN(P1_U3323) );
  INV_X1 U10965 ( .A(n9843), .ZN(n9848) );
  AOI21_X1 U10966 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9847) );
  AOI211_X1 U10967 ( .C1(n9850), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9871)
         );
  INV_X1 U10968 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10969 ( .A1(n9869), .A2(n9871), .B1(n9851), .B2(n9867), .ZN(
        P1_U3453) );
  OAI21_X1 U10970 ( .B1(n6525), .B2(n9853), .A(n9852), .ZN(n9855) );
  AOI211_X1 U10971 ( .C1(n9858), .C2(n9856), .A(n9855), .B(n9854), .ZN(n9873)
         );
  INV_X1 U10972 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U10973 ( .A1(n9869), .A2(n9873), .B1(n9857), .B2(n9867), .ZN(
        P1_U3456) );
  NAND2_X1 U10974 ( .A1(n9859), .A2(n9858), .ZN(n9866) );
  NAND2_X1 U10975 ( .A1(n9861), .A2(n9860), .ZN(n9862) );
  AND2_X1 U10976 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  INV_X1 U10977 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U10978 ( .A1(n9869), .A2(n9875), .B1(n9868), .B2(n9867), .ZN(
        P1_U3477) );
  AOI22_X1 U10979 ( .A1(n9876), .A2(n9871), .B1(n9870), .B2(n9874), .ZN(
        P1_U3522) );
  AOI22_X1 U10980 ( .A1(n9876), .A2(n9873), .B1(n9872), .B2(n9874), .ZN(
        P1_U3523) );
  AOI22_X1 U10981 ( .A1(n9876), .A2(n9875), .B1(n6915), .B2(n9874), .ZN(
        P1_U3530) );
  INV_X1 U10982 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U10983 ( .A1(n9878), .A2(n9877), .ZN(n9879) );
  NAND2_X1 U10984 ( .A1(n9880), .A2(n9879), .ZN(n9881) );
  NAND2_X1 U10985 ( .A1(n9904), .A2(n9881), .ZN(n9887) );
  NAND2_X1 U10986 ( .A1(n9882), .A2(n5959), .ZN(n9883) );
  NAND2_X1 U10987 ( .A1(n9884), .A2(n9883), .ZN(n9885) );
  NAND2_X1 U10988 ( .A1(n8821), .A2(n9885), .ZN(n9886) );
  OAI211_X1 U10989 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9888), .A(n9887), .B(
        n9886), .ZN(n9889) );
  AOI21_X1 U10990 ( .B1(n6897), .B2(n9902), .A(n9889), .ZN(n9895) );
  XOR2_X1 U10991 ( .A(n9891), .B(n9890), .Z(n9893) );
  NAND2_X1 U10992 ( .A1(n9893), .A2(n9892), .ZN(n9894) );
  OAI211_X1 U10993 ( .C1(n10200), .C2(n9896), .A(n9895), .B(n9894), .ZN(
        P2_U3183) );
  AOI21_X1 U10994 ( .B1(n9898), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9897), .ZN(
        n9918) );
  OAI21_X1 U10995 ( .B1(n9901), .B2(n9900), .A(n9899), .ZN(n9905) );
  AOI22_X1 U10996 ( .A1(n9905), .A2(n9904), .B1(n9903), .B2(n9902), .ZN(n9917)
         );
  AOI21_X1 U10997 ( .B1(n9907), .B2(n9906), .A(n4403), .ZN(n9909) );
  OR2_X1 U10998 ( .A1(n9909), .A2(n9908), .ZN(n9916) );
  AOI21_X1 U10999 ( .B1(n9912), .B2(n9911), .A(n9910), .ZN(n9914) );
  OR2_X1 U11000 ( .A1(n9914), .A2(n9913), .ZN(n9915) );
  NAND4_X1 U11001 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(
        P2_U3190) );
  INV_X1 U11002 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9924) );
  INV_X1 U11003 ( .A(n9919), .ZN(n9923) );
  OAI22_X1 U11004 ( .A1(n9921), .A2(n9982), .B1(n9920), .B2(n9955), .ZN(n9922)
         );
  NOR2_X1 U11005 ( .A1(n9923), .A2(n9922), .ZN(n9991) );
  AOI22_X1 U11006 ( .A1(n9990), .A2(n9924), .B1(n9991), .B2(n9988), .ZN(
        P2_U3393) );
  INV_X1 U11007 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9932) );
  INV_X1 U11008 ( .A(n9925), .ZN(n9929) );
  OAI22_X1 U11009 ( .A1(n9927), .A2(n9971), .B1(n9926), .B2(n9955), .ZN(n9928)
         );
  AOI211_X1 U11010 ( .C1(n9931), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9992)
         );
  AOI22_X1 U11011 ( .A1(n9990), .A2(n9932), .B1(n9992), .B2(n9988), .ZN(
        P2_U3396) );
  INV_X1 U11012 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9937) );
  OAI21_X1 U11013 ( .B1(n9934), .B2(n9955), .A(n9933), .ZN(n9935) );
  AOI21_X1 U11014 ( .B1(n9936), .B2(n9949), .A(n9935), .ZN(n9993) );
  AOI22_X1 U11015 ( .A1(n9990), .A2(n9937), .B1(n9993), .B2(n9988), .ZN(
        P2_U3399) );
  INV_X1 U11016 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9943) );
  INV_X1 U11017 ( .A(n9938), .ZN(n9942) );
  OAI21_X1 U11018 ( .B1(n9940), .B2(n9955), .A(n9939), .ZN(n9941) );
  AOI21_X1 U11019 ( .B1(n9942), .B2(n9949), .A(n9941), .ZN(n9994) );
  AOI22_X1 U11020 ( .A1(n9990), .A2(n9943), .B1(n9994), .B2(n9988), .ZN(
        P2_U3402) );
  INV_X1 U11021 ( .A(n9944), .ZN(n9948) );
  OAI21_X1 U11022 ( .B1(n9946), .B2(n9955), .A(n9945), .ZN(n9947) );
  AOI21_X1 U11023 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9995) );
  AOI22_X1 U11024 ( .A1(n9990), .A2(n6030), .B1(n9995), .B2(n9988), .ZN(
        P2_U3405) );
  INV_X1 U11025 ( .A(n9950), .ZN(n9954) );
  OAI22_X1 U11026 ( .A1(n9952), .A2(n9982), .B1(n9951), .B2(n9955), .ZN(n9953)
         );
  NOR2_X1 U11027 ( .A1(n9954), .A2(n9953), .ZN(n9996) );
  AOI22_X1 U11028 ( .A1(n9990), .A2(n5948), .B1(n9996), .B2(n9988), .ZN(
        P2_U3408) );
  OAI22_X1 U11029 ( .A1(n9957), .A2(n9971), .B1(n9956), .B2(n9955), .ZN(n9958)
         );
  NOR2_X1 U11030 ( .A1(n9959), .A2(n9958), .ZN(n9998) );
  AOI22_X1 U11031 ( .A1(n9990), .A2(n6069), .B1(n9998), .B2(n9988), .ZN(
        P2_U3411) );
  INV_X1 U11032 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9965) );
  NOR2_X1 U11033 ( .A1(n9960), .A2(n9982), .ZN(n9963) );
  INV_X1 U11034 ( .A(n9961), .ZN(n9962) );
  AOI211_X1 U11035 ( .C1(n9987), .C2(n9964), .A(n9963), .B(n9962), .ZN(n9999)
         );
  AOI22_X1 U11036 ( .A1(n9990), .A2(n9965), .B1(n9999), .B2(n9988), .ZN(
        P2_U3414) );
  INV_X1 U11037 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9970) );
  NOR2_X1 U11038 ( .A1(n9966), .A2(n9971), .ZN(n9968) );
  AOI211_X1 U11039 ( .C1(n9987), .C2(n9969), .A(n9968), .B(n9967), .ZN(n10000)
         );
  AOI22_X1 U11040 ( .A1(n9990), .A2(n9970), .B1(n10000), .B2(n9988), .ZN(
        P2_U3417) );
  INV_X1 U11041 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9976) );
  NOR2_X1 U11042 ( .A1(n9972), .A2(n9971), .ZN(n9974) );
  AOI211_X1 U11043 ( .C1(n9987), .C2(n9975), .A(n9974), .B(n9973), .ZN(n10001)
         );
  AOI22_X1 U11044 ( .A1(n9990), .A2(n9976), .B1(n10001), .B2(n9988), .ZN(
        P2_U3420) );
  INV_X1 U11045 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U11046 ( .A1(n9977), .A2(n9982), .ZN(n9979) );
  AOI211_X1 U11047 ( .C1(n9987), .C2(n9980), .A(n9979), .B(n9978), .ZN(n10002)
         );
  AOI22_X1 U11048 ( .A1(n9990), .A2(n9981), .B1(n10002), .B2(n9988), .ZN(
        P2_U3423) );
  INV_X1 U11049 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9989) );
  NOR2_X1 U11050 ( .A1(n9983), .A2(n9982), .ZN(n9985) );
  AOI211_X1 U11051 ( .C1(n9987), .C2(n9986), .A(n9985), .B(n9984), .ZN(n10004)
         );
  AOI22_X1 U11052 ( .A1(n9990), .A2(n9989), .B1(n10004), .B2(n9988), .ZN(
        P2_U3426) );
  AOI22_X1 U11053 ( .A1(n10005), .A2(n9991), .B1(n5959), .B2(n10003), .ZN(
        P2_U3460) );
  AOI22_X1 U11054 ( .A1(n10005), .A2(n9992), .B1(n5981), .B2(n10003), .ZN(
        P2_U3461) );
  AOI22_X1 U11055 ( .A1(n10005), .A2(n9993), .B1(n5995), .B2(n10003), .ZN(
        P2_U3462) );
  AOI22_X1 U11056 ( .A1(n10005), .A2(n9994), .B1(n6013), .B2(n10003), .ZN(
        P2_U3463) );
  AOI22_X1 U11057 ( .A1(n10005), .A2(n9995), .B1(n6026), .B2(n10003), .ZN(
        P2_U3464) );
  AOI22_X1 U11058 ( .A1(n10005), .A2(n9996), .B1(n7162), .B2(n10003), .ZN(
        P2_U3465) );
  AOI22_X1 U11059 ( .A1(n10005), .A2(n9998), .B1(n9997), .B2(n10003), .ZN(
        P2_U3466) );
  AOI22_X1 U11060 ( .A1(n10005), .A2(n9999), .B1(n7594), .B2(n10003), .ZN(
        P2_U3467) );
  AOI22_X1 U11061 ( .A1(n10005), .A2(n10000), .B1(n7601), .B2(n10003), .ZN(
        P2_U3468) );
  AOI22_X1 U11062 ( .A1(n10005), .A2(n10001), .B1(n7729), .B2(n10003), .ZN(
        P2_U3469) );
  AOI22_X1 U11063 ( .A1(n10005), .A2(n10002), .B1(n6102), .B2(n10003), .ZN(
        P2_U3470) );
  AOI22_X1 U11064 ( .A1(n10005), .A2(n10004), .B1(n7947), .B2(n10003), .ZN(
        P2_U3471) );
  NOR2_X1 U11065 ( .A1(n10007), .A2(n10006), .ZN(n10008) );
  XNOR2_X1 U11066 ( .A(n10008), .B(n10200), .ZN(ADD_1068_U5) );
  XOR2_X1 U11067 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11068 ( .A1(n10010), .A2(n10009), .ZN(n10012) );
  XNOR2_X1 U11069 ( .A(n10012), .B(n10011), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11070 ( .A(n10014), .B(n10013), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11071 ( .A(n10016), .B(n10015), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11072 ( .A(n10018), .B(n10017), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11073 ( .A(n10020), .B(n10019), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11074 ( .A(n10022), .B(n10021), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11075 ( .A(n10024), .B(n10023), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11076 ( .A(n10026), .B(n10025), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11077 ( .A(n10028), .B(n10027), .ZN(ADD_1068_U63) );
  NAND2_X1 U11078 ( .A1(n10029), .A2(P2_D_REG_9__SCAN_IN), .ZN(n10219) );
  INV_X1 U11079 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10032) );
  AOI22_X1 U11080 ( .A1(n10032), .A2(keyinput93), .B1(keyinput89), .B2(n10031), 
        .ZN(n10030) );
  OAI221_X1 U11081 ( .B1(n10032), .B2(keyinput93), .C1(n10031), .C2(keyinput89), .A(n10030), .ZN(n10042) );
  INV_X1 U11082 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10034) );
  AOI22_X1 U11083 ( .A1(n10034), .A2(keyinput98), .B1(keyinput67), .B2(n10171), 
        .ZN(n10033) );
  OAI221_X1 U11084 ( .B1(n10034), .B2(keyinput98), .C1(n10171), .C2(keyinput67), .A(n10033), .ZN(n10041) );
  AOI22_X1 U11085 ( .A1(n6276), .A2(keyinput76), .B1(n10158), .B2(keyinput118), 
        .ZN(n10035) );
  OAI221_X1 U11086 ( .B1(n6276), .B2(keyinput76), .C1(n10158), .C2(keyinput118), .A(n10035), .ZN(n10040) );
  AOI22_X1 U11087 ( .A1(n10038), .A2(keyinput121), .B1(n10037), .B2(
        keyinput127), .ZN(n10036) );
  OAI221_X1 U11088 ( .B1(n10038), .B2(keyinput121), .C1(n10037), .C2(
        keyinput127), .A(n10036), .ZN(n10039) );
  NOR4_X1 U11089 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n10079) );
  AOI22_X1 U11090 ( .A1(n6013), .A2(keyinput78), .B1(keyinput117), .B2(n10044), 
        .ZN(n10043) );
  OAI221_X1 U11091 ( .B1(n6013), .B2(keyinput78), .C1(n10044), .C2(keyinput117), .A(n10043), .ZN(n10055) );
  INV_X1 U11092 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11093 ( .A1(n10047), .A2(keyinput90), .B1(keyinput74), .B2(n10046), 
        .ZN(n10045) );
  OAI221_X1 U11094 ( .B1(n10047), .B2(keyinput90), .C1(n10046), .C2(keyinput74), .A(n10045), .ZN(n10054) );
  INV_X1 U11095 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n10199) );
  INV_X1 U11096 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10049) );
  AOI22_X1 U11097 ( .A1(n10199), .A2(keyinput86), .B1(n10049), .B2(keyinput111), .ZN(n10048) );
  OAI221_X1 U11098 ( .B1(n10199), .B2(keyinput86), .C1(n10049), .C2(
        keyinput111), .A(n10048), .ZN(n10053) );
  XNOR2_X1 U11099 ( .A(P1_REG0_REG_15__SCAN_IN), .B(keyinput105), .ZN(n10051)
         );
  XNOR2_X1 U11100 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput72), .ZN(n10050) );
  NAND2_X1 U11101 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  NOR4_X1 U11102 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        n10078) );
  AOI22_X1 U11103 ( .A1(n10057), .A2(keyinput77), .B1(n10161), .B2(keyinput73), 
        .ZN(n10056) );
  OAI221_X1 U11104 ( .B1(n10057), .B2(keyinput77), .C1(n10161), .C2(keyinput73), .A(n10056), .ZN(n10064) );
  AOI22_X1 U11105 ( .A1(n10169), .A2(keyinput95), .B1(n10188), .B2(keyinput87), 
        .ZN(n10058) );
  OAI221_X1 U11106 ( .B1(n10169), .B2(keyinput95), .C1(n10188), .C2(keyinput87), .A(n10058), .ZN(n10063) );
  INV_X1 U11107 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U11108 ( .A1(n9603), .A2(keyinput81), .B1(keyinput123), .B2(n10203), 
        .ZN(n10059) );
  OAI221_X1 U11109 ( .B1(n9603), .B2(keyinput81), .C1(n10203), .C2(keyinput123), .A(n10059), .ZN(n10062) );
  AOI22_X1 U11110 ( .A1(n4938), .A2(keyinput113), .B1(keyinput88), .B2(n5018), 
        .ZN(n10060) );
  OAI221_X1 U11111 ( .B1(n4938), .B2(keyinput113), .C1(n5018), .C2(keyinput88), 
        .A(n10060), .ZN(n10061) );
  NOR4_X1 U11112 ( .A1(n10064), .A2(n10063), .A3(n10062), .A4(n10061), .ZN(
        n10077) );
  AOI22_X1 U11113 ( .A1(n8907), .A2(keyinput97), .B1(keyinput99), .B2(n10183), 
        .ZN(n10065) );
  OAI221_X1 U11114 ( .B1(n8907), .B2(keyinput97), .C1(n10183), .C2(keyinput99), 
        .A(n10065), .ZN(n10075) );
  INV_X1 U11115 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11116 ( .A1(n7240), .A2(keyinput103), .B1(n10155), .B2(keyinput68), 
        .ZN(n10066) );
  OAI221_X1 U11117 ( .B1(n7240), .B2(keyinput103), .C1(n10155), .C2(keyinput68), .A(n10066), .ZN(n10074) );
  AOI22_X1 U11118 ( .A1(n10069), .A2(keyinput66), .B1(n10068), .B2(keyinput102), .ZN(n10067) );
  OAI221_X1 U11119 ( .B1(n10069), .B2(keyinput66), .C1(n10068), .C2(
        keyinput102), .A(n10067), .ZN(n10073) );
  XOR2_X1 U11120 ( .A(n9189), .B(keyinput84), .Z(n10071) );
  XNOR2_X1 U11121 ( .A(SI_3_), .B(keyinput85), .ZN(n10070) );
  NAND2_X1 U11122 ( .A1(n10071), .A2(n10070), .ZN(n10072) );
  NOR4_X1 U11123 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n10076) );
  AND4_X1 U11124 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10217) );
  OAI22_X1 U11125 ( .A1(P2_D_REG_12__SCAN_IN), .A2(keyinput94), .B1(
        P2_REG0_REG_6__SCAN_IN), .B2(keyinput107), .ZN(n10080) );
  AOI221_X1 U11126 ( .B1(P2_D_REG_12__SCAN_IN), .B2(keyinput94), .C1(
        keyinput107), .C2(P2_REG0_REG_6__SCAN_IN), .A(n10080), .ZN(n10087) );
  OAI22_X1 U11127 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(keyinput104), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(keyinput83), .ZN(n10081) );
  AOI221_X1 U11128 ( .B1(P2_IR_REG_16__SCAN_IN), .B2(keyinput104), .C1(
        keyinput83), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n10081), .ZN(n10086) );
  OAI22_X1 U11129 ( .A1(P2_D_REG_31__SCAN_IN), .A2(keyinput65), .B1(
        keyinput116), .B2(P2_ADDR_REG_14__SCAN_IN), .ZN(n10082) );
  AOI221_X1 U11130 ( .B1(P2_D_REG_31__SCAN_IN), .B2(keyinput65), .C1(
        P2_ADDR_REG_14__SCAN_IN), .C2(keyinput116), .A(n10082), .ZN(n10085) );
  OAI22_X1 U11131 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput82), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput114), .ZN(n10083) );
  AOI221_X1 U11132 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput82), .C1(
        keyinput114), .C2(P1_IR_REG_15__SCAN_IN), .A(n10083), .ZN(n10084) );
  NAND4_X1 U11133 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        n10117) );
  OAI22_X1 U11134 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(keyinput115), .B1(
        P1_REG0_REG_30__SCAN_IN), .B2(keyinput75), .ZN(n10088) );
  AOI221_X1 U11135 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(keyinput115), .C1(
        keyinput75), .C2(P1_REG0_REG_30__SCAN_IN), .A(n10088), .ZN(n10095) );
  OAI22_X1 U11136 ( .A1(P1_D_REG_16__SCAN_IN), .A2(keyinput91), .B1(
        P2_ADDR_REG_8__SCAN_IN), .B2(keyinput122), .ZN(n10089) );
  AOI221_X1 U11137 ( .B1(P1_D_REG_16__SCAN_IN), .B2(keyinput91), .C1(
        keyinput122), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10089), .ZN(n10094) );
  OAI22_X1 U11138 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(keyinput106), .B1(
        P1_REG0_REG_18__SCAN_IN), .B2(keyinput112), .ZN(n10090) );
  AOI221_X1 U11139 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(keyinput106), .C1(
        keyinput112), .C2(P1_REG0_REG_18__SCAN_IN), .A(n10090), .ZN(n10093) );
  OAI22_X1 U11140 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput100), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(keyinput119), .ZN(n10091) );
  AOI221_X1 U11141 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput100), .C1(
        keyinput119), .C2(P1_DATAO_REG_25__SCAN_IN), .A(n10091), .ZN(n10092)
         );
  NAND4_X1 U11142 ( .A1(n10095), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n10116) );
  OAI22_X1 U11143 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput96), .B1(
        keyinput80), .B2(P2_REG2_REG_15__SCAN_IN), .ZN(n10096) );
  AOI221_X1 U11144 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput96), .C1(
        P2_REG2_REG_15__SCAN_IN), .C2(keyinput80), .A(n10096), .ZN(n10105) );
  OAI22_X1 U11145 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput110), .B1(
        P1_REG2_REG_27__SCAN_IN), .B2(keyinput108), .ZN(n10097) );
  AOI221_X1 U11146 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput110), .C1(
        keyinput108), .C2(P1_REG2_REG_27__SCAN_IN), .A(n10097), .ZN(n10104) );
  INV_X1 U11147 ( .A(keyinput125), .ZN(n10098) );
  XNOR2_X1 U11148 ( .A(n10098), .B(P1_IR_REG_27__SCAN_IN), .ZN(n10102) );
  XNOR2_X1 U11149 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput124), .ZN(n10101) );
  XNOR2_X1 U11150 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput101), .ZN(n10100) );
  XNOR2_X1 U11151 ( .A(keyinput109), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n10099)
         );
  AND4_X1 U11152 ( .A1(n10102), .A2(n10101), .A3(n10100), .A4(n10099), .ZN(
        n10103) );
  NAND3_X1 U11153 ( .A1(n10105), .A2(n10104), .A3(n10103), .ZN(n10115) );
  OAI22_X1 U11154 ( .A1(SI_18_), .A2(keyinput64), .B1(keyinput71), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n10106) );
  AOI221_X1 U11155 ( .B1(SI_18_), .B2(keyinput64), .C1(P1_REG2_REG_24__SCAN_IN), .C2(keyinput71), .A(n10106), .ZN(n10113) );
  OAI22_X1 U11156 ( .A1(SI_27_), .A2(keyinput79), .B1(P2_REG0_REG_25__SCAN_IN), 
        .B2(keyinput69), .ZN(n10107) );
  AOI221_X1 U11157 ( .B1(SI_27_), .B2(keyinput79), .C1(keyinput69), .C2(
        P2_REG0_REG_25__SCAN_IN), .A(n10107), .ZN(n10112) );
  OAI22_X1 U11158 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput126), .B1(
        P2_REG0_REG_7__SCAN_IN), .B2(keyinput92), .ZN(n10108) );
  AOI221_X1 U11159 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput126), .C1(
        keyinput92), .C2(P2_REG0_REG_7__SCAN_IN), .A(n10108), .ZN(n10111) );
  OAI22_X1 U11160 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput70), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput120), .ZN(n10109) );
  AOI221_X1 U11161 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput70), .C1(
        keyinput120), .C2(P1_IR_REG_2__SCAN_IN), .A(n10109), .ZN(n10110) );
  NAND4_X1 U11162 ( .A1(n10113), .A2(n10112), .A3(n10111), .A4(n10110), .ZN(
        n10114) );
  NOR4_X1 U11163 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10216) );
  AOI22_X1 U11164 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput60), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(keyinput55), .ZN(n10118) );
  OAI221_X1 U11165 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput60), .C1(
        P1_DATAO_REG_25__SCAN_IN), .C2(keyinput55), .A(n10118), .ZN(n10125) );
  AOI22_X1 U11166 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(keyinput57), .B1(
        P1_REG2_REG_20__SCAN_IN), .B2(keyinput51), .ZN(n10119) );
  OAI221_X1 U11167 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(keyinput57), .C1(
        P1_REG2_REG_20__SCAN_IN), .C2(keyinput51), .A(n10119), .ZN(n10124) );
  AOI22_X1 U11168 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(keyinput20), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput36), .ZN(n10120) );
  OAI221_X1 U11169 ( .B1(P1_REG3_REG_14__SCAN_IN), .B2(keyinput20), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput36), .A(n10120), .ZN(n10123) );
  AOI22_X1 U11170 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(keyinput7), .B1(
        P2_REG2_REG_15__SCAN_IN), .B2(keyinput16), .ZN(n10121) );
  OAI221_X1 U11171 ( .B1(P1_REG2_REG_24__SCAN_IN), .B2(keyinput7), .C1(
        P2_REG2_REG_15__SCAN_IN), .C2(keyinput16), .A(n10121), .ZN(n10122) );
  NOR4_X1 U11172 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10153) );
  AOI22_X1 U11173 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(keyinput11), .B1(
        P1_REG1_REG_9__SCAN_IN), .B2(keyinput26), .ZN(n10126) );
  OAI221_X1 U11174 ( .B1(P1_REG0_REG_30__SCAN_IN), .B2(keyinput11), .C1(
        P1_REG1_REG_9__SCAN_IN), .C2(keyinput26), .A(n10126), .ZN(n10133) );
  AOI22_X1 U11175 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput61), .B1(
        P2_REG0_REG_7__SCAN_IN), .B2(keyinput28), .ZN(n10127) );
  OAI221_X1 U11176 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput61), .C1(
        P2_REG0_REG_7__SCAN_IN), .C2(keyinput28), .A(n10127), .ZN(n10132) );
  AOI22_X1 U11177 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput38), .B1(
        P2_IR_REG_27__SCAN_IN), .B2(keyinput29), .ZN(n10128) );
  OAI221_X1 U11178 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput38), .C1(
        P2_IR_REG_27__SCAN_IN), .C2(keyinput29), .A(n10128), .ZN(n10131) );
  AOI22_X1 U11179 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput53), .B1(
        P1_D_REG_17__SCAN_IN), .B2(keyinput25), .ZN(n10129) );
  OAI221_X1 U11180 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput53), .C1(
        P1_D_REG_17__SCAN_IN), .C2(keyinput25), .A(n10129), .ZN(n10130) );
  NOR4_X1 U11181 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10152) );
  AOI22_X1 U11182 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput24), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput32), .ZN(n10134) );
  OAI221_X1 U11183 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput24), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput32), .A(n10134), .ZN(n10141) );
  AOI22_X1 U11184 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(keyinput34), .B1(
        P2_IR_REG_28__SCAN_IN), .B2(keyinput37), .ZN(n10135) );
  OAI221_X1 U11185 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(keyinput34), .C1(
        P2_IR_REG_28__SCAN_IN), .C2(keyinput37), .A(n10135), .ZN(n10140) );
  AOI22_X1 U11186 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(keyinput10), .B1(
        P2_ADDR_REG_14__SCAN_IN), .B2(keyinput52), .ZN(n10136) );
  OAI221_X1 U11187 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(keyinput10), .C1(
        P2_ADDR_REG_14__SCAN_IN), .C2(keyinput52), .A(n10136), .ZN(n10139) );
  AOI22_X1 U11188 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(keyinput42), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(keyinput13), .ZN(n10137) );
  OAI221_X1 U11189 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(keyinput42), .C1(
        P2_REG1_REG_0__SCAN_IN), .C2(keyinput13), .A(n10137), .ZN(n10138) );
  NOR4_X1 U11190 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10151) );
  AOI22_X1 U11191 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(keyinput44), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput47), .ZN(n10142) );
  OAI221_X1 U11192 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(keyinput44), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput47), .A(n10142), .ZN(n10149) );
  AOI22_X1 U11193 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(keyinput39), .B1(
        P2_D_REG_31__SCAN_IN), .B2(keyinput1), .ZN(n10143) );
  OAI221_X1 U11194 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(keyinput39), .C1(
        P2_D_REG_31__SCAN_IN), .C2(keyinput1), .A(n10143), .ZN(n10148) );
  AOI22_X1 U11195 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput8), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput18), .ZN(n10144) );
  OAI221_X1 U11196 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput8), .C1(
        P1_DATAO_REG_21__SCAN_IN), .C2(keyinput18), .A(n10144), .ZN(n10147) );
  AOI22_X1 U11197 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput6), .B1(
        P2_REG2_REG_27__SCAN_IN), .B2(keyinput33), .ZN(n10145) );
  OAI221_X1 U11198 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput6), .C1(
        P2_REG2_REG_27__SCAN_IN), .C2(keyinput33), .A(n10145), .ZN(n10146) );
  NOR4_X1 U11199 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10150) );
  NAND4_X1 U11200 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10215) );
  AOI22_X1 U11201 ( .A1(n10155), .A2(keyinput4), .B1(keyinput17), .B2(n9603), 
        .ZN(n10154) );
  OAI221_X1 U11202 ( .B1(n10155), .B2(keyinput4), .C1(n9603), .C2(keyinput17), 
        .A(n10154), .ZN(n10167) );
  AOI22_X1 U11203 ( .A1(n10158), .A2(keyinput54), .B1(keyinput30), .B2(n10157), 
        .ZN(n10156) );
  OAI221_X1 U11204 ( .B1(n10158), .B2(keyinput54), .C1(n10157), .C2(keyinput30), .A(n10156), .ZN(n10166) );
  AOI22_X1 U11205 ( .A1(n10161), .A2(keyinput9), .B1(keyinput46), .B2(n10160), 
        .ZN(n10159) );
  OAI221_X1 U11206 ( .B1(n10161), .B2(keyinput9), .C1(n10160), .C2(keyinput46), 
        .A(n10159), .ZN(n10165) );
  XNOR2_X1 U11207 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput40), .ZN(n10163) );
  XNOR2_X1 U11208 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(keyinput63), .ZN(n10162)
         );
  NAND2_X1 U11209 ( .A1(n10163), .A2(n10162), .ZN(n10164) );
  NOR4_X1 U11210 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10213) );
  AOI22_X1 U11211 ( .A1(n6276), .A2(keyinput12), .B1(n10169), .B2(keyinput31), 
        .ZN(n10168) );
  OAI221_X1 U11212 ( .B1(n6276), .B2(keyinput12), .C1(n10169), .C2(keyinput31), 
        .A(n10168), .ZN(n10180) );
  AOI22_X1 U11213 ( .A1(n10171), .A2(keyinput3), .B1(n6013), .B2(keyinput14), 
        .ZN(n10170) );
  OAI221_X1 U11214 ( .B1(n10171), .B2(keyinput3), .C1(n6013), .C2(keyinput14), 
        .A(n10170), .ZN(n10179) );
  AOI22_X1 U11215 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput2), .B1(
        P1_REG0_REG_15__SCAN_IN), .B2(keyinput41), .ZN(n10172) );
  OAI221_X1 U11216 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput2), .C1(
        P1_REG0_REG_15__SCAN_IN), .C2(keyinput41), .A(n10172), .ZN(n10177) );
  XNOR2_X1 U11217 ( .A(n10173), .B(keyinput62), .ZN(n10176) );
  INV_X1 U11218 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10174) );
  XNOR2_X1 U11219 ( .A(n10174), .B(keyinput58), .ZN(n10175) );
  OR3_X1 U11220 ( .A1(n10177), .A2(n10176), .A3(n10175), .ZN(n10178) );
  NOR3_X1 U11221 ( .A1(n10180), .A2(n10179), .A3(n10178), .ZN(n10212) );
  AOI22_X1 U11222 ( .A1(n10183), .A2(keyinput35), .B1(keyinput27), .B2(n10182), 
        .ZN(n10181) );
  OAI221_X1 U11223 ( .B1(n10183), .B2(keyinput35), .C1(n10182), .C2(keyinput27), .A(n10181), .ZN(n10194) );
  AOI22_X1 U11224 ( .A1(n10185), .A2(keyinput15), .B1(keyinput56), .B2(n4614), 
        .ZN(n10184) );
  OAI221_X1 U11225 ( .B1(n10185), .B2(keyinput15), .C1(n4614), .C2(keyinput56), 
        .A(n10184), .ZN(n10193) );
  AOI22_X1 U11226 ( .A1(n10188), .A2(keyinput23), .B1(keyinput5), .B2(n10187), 
        .ZN(n10186) );
  OAI221_X1 U11227 ( .B1(n10188), .B2(keyinput23), .C1(n10187), .C2(keyinput5), 
        .A(n10186), .ZN(n10192) );
  XNOR2_X1 U11228 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput49), .ZN(n10190)
         );
  XNOR2_X1 U11229 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput50), .ZN(n10189) );
  NAND2_X1 U11230 ( .A1(n10190), .A2(n10189), .ZN(n10191) );
  NOR4_X1 U11231 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n10211) );
  AOI22_X1 U11232 ( .A1(n10197), .A2(keyinput0), .B1(n10196), .B2(keyinput45), 
        .ZN(n10195) );
  OAI221_X1 U11233 ( .B1(n10197), .B2(keyinput0), .C1(n10196), .C2(keyinput45), 
        .A(n10195), .ZN(n10209) );
  AOI22_X1 U11234 ( .A1(n10200), .A2(keyinput19), .B1(n10199), .B2(keyinput22), 
        .ZN(n10198) );
  OAI221_X1 U11235 ( .B1(n10200), .B2(keyinput19), .C1(n10199), .C2(keyinput22), .A(n10198), .ZN(n10208) );
  AOI22_X1 U11236 ( .A1(n10203), .A2(keyinput59), .B1(n10202), .B2(keyinput48), 
        .ZN(n10201) );
  OAI221_X1 U11237 ( .B1(n10203), .B2(keyinput59), .C1(n10202), .C2(keyinput48), .A(n10201), .ZN(n10207) );
  XOR2_X1 U11238 ( .A(n5948), .B(keyinput43), .Z(n10205) );
  XNOR2_X1 U11239 ( .A(SI_3_), .B(keyinput21), .ZN(n10204) );
  NAND2_X1 U11240 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  NOR4_X1 U11241 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10210) );
  NAND4_X1 U11242 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        n10214) );
  AOI211_X1 U11243 ( .C1(n10217), .C2(n10216), .A(n10215), .B(n10214), .ZN(
        n10218) );
  XNOR2_X1 U11244 ( .A(n10219), .B(n10218), .ZN(P2_U3256) );
  XNOR2_X1 U11245 ( .A(n10221), .B(n10220), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11246 ( .A(n10223), .B(n10222), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11247 ( .A(n10225), .B(n10224), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11248 ( .A(n10227), .B(n10226), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11249 ( .A(n10229), .B(n10228), .ZN(ADD_1068_U48) );
  XOR2_X1 U11250 ( .A(n10231), .B(n10230), .Z(ADD_1068_U54) );
  XOR2_X1 U11251 ( .A(n10233), .B(n10232), .Z(ADD_1068_U53) );
  XNOR2_X1 U11252 ( .A(n10235), .B(n10234), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4841 ( .A(n5145), .Z(n5657) );
  OAI21_X1 U4873 ( .B1(n7135), .B2(n7240), .A(n7134), .ZN(n7154) );
  NOR2_X2 U4888 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5987) );
  CLKBUF_X1 U4904 ( .A(n5982), .Z(n6185) );
  XNOR2_X1 U5097 ( .A(n5001), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5700) );
endmodule

