

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778;

  INV_X4 U2246 ( .A(n2886), .ZN(n2861) );
  INV_X2 U2247 ( .A(n2875), .ZN(n2839) );
  NAND2_X1 U2248 ( .A1(n2409), .A2(n2408), .ZN(n4366) );
  XNOR2_X1 U2249 ( .A(n2376), .B(n2375), .ZN(n2408) );
  CLKBUF_X2 U2250 ( .A(n2570), .Z(n2802) );
  BUF_X1 U2252 ( .A(n2512), .Z(n2570) );
  AND2_X2 U2253 ( .A1(n2402), .A2(n2421), .ZN(n2858) );
  INV_X1 U2254 ( .A(n2839), .ZN(n2837) );
  NOR2_X1 U2255 ( .A1(n3002), .A2(n2026), .ZN(n2284) );
  OAI21_X1 U2256 ( .B1(n2269), .B2(n3756), .A(n2095), .ZN(n4008) );
  NOR2_X2 U2257 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2437)
         );
  INV_X1 U2258 ( .A(n3299), .ZN(n2966) );
  NAND2_X1 U2259 ( .A1(n3190), .A2(n3191), .ZN(n3189) );
  CLKBUF_X2 U2260 ( .A(n2510), .Z(n3750) );
  INV_X1 U2261 ( .A(n2451), .ZN(n2467) );
  AND2_X1 U2262 ( .A1(n2175), .A2(n2071), .ZN(n2500) );
  AND2_X1 U2263 ( .A1(n2878), .A2(n2867), .ZN(n4038) );
  NOR2_X2 U2264 ( .A1(n2353), .A2(n3531), .ZN(n4312) );
  NAND2_X1 U2265 ( .A1(n2405), .A2(IR_REG_31__SCAN_IN), .ZN(n2406) );
  AOI211_X1 U2266 ( .C1(n4349), .C2(n4255), .A(n4041), .B(n4040), .ZN(n4042)
         );
  XNOR2_X1 U2267 ( .A(n2406), .B(IR_REG_22__SCAN_IN), .ZN(n4487) );
  AND4_X1 U2268 ( .A1(n2720), .A2(n2359), .A3(n2358), .A4(n2357), .ZN(n2004)
         );
  INV_X2 U2269 ( .A(n2958), .ZN(n2955) );
  NOR2_X2 U2270 ( .A1(n3341), .A2(n3492), .ZN(n3360) );
  NAND2_X2 U2271 ( .A1(n2092), .A2(n2091), .ZN(n2090) );
  OAI22_X2 U2272 ( .A1(n4145), .A2(n2996), .B1(n2995), .B2(n4160), .ZN(n4130)
         );
  XNOR2_X2 U2273 ( .A(n3324), .B(n3236), .ZN(n3235) );
  NAND2_X2 U2274 ( .A1(n3233), .A2(n2346), .ZN(n3324) );
  NAND4_X2 U2275 ( .A1(n2435), .A2(n2432), .A3(n2431), .A4(n2433), .ZN(n2958)
         );
  OAI21_X1 U2276 ( .B1(n4008), .B2(n4007), .A(n4006), .ZN(n4009) );
  AND2_X1 U2277 ( .A1(n2858), .A2(n4366), .ZN(n2005) );
  AOI21_X2 U2278 ( .B1(n4094), .B2(n3001), .A(n2347), .ZN(n4078) );
  NAND2_X2 U2279 ( .A1(n4113), .A2(n3000), .ZN(n4094) );
  XNOR2_X2 U2280 ( .A(n3084), .B(n2479), .ZN(n3922) );
  NAND2_X1 U2281 ( .A1(n2408), .A2(n4488), .ZN(n2402) );
  NAND2_X1 U2282 ( .A1(n3662), .A2(n2814), .ZN(n3517) );
  OR2_X1 U2283 ( .A1(n3183), .A2(n3184), .ZN(n3185) );
  NAND2_X1 U2284 ( .A1(n3819), .A2(n3822), .ZN(n3777) );
  NAND2_X1 U2285 ( .A1(n3007), .A2(n3166), .ZN(n3165) );
  BUF_X2 U2286 ( .A(n3749), .Z(n3754) );
  NAND2_X1 U2287 ( .A1(n2944), .A2(n3807), .ZN(n3149) );
  INV_X1 U2288 ( .A(n2457), .ZN(n2636) );
  NAND2_X1 U2289 ( .A1(n2175), .A2(n2345), .ZN(n2498) );
  NOR2_X1 U2290 ( .A1(n4342), .A2(n4341), .ZN(n4347) );
  AND2_X1 U2291 ( .A1(n4350), .A2(n2070), .ZN(n2069) );
  AND2_X1 U2292 ( .A1(n2105), .A2(n2104), .ZN(n4350) );
  NAND2_X1 U2293 ( .A1(n4061), .A2(n2267), .ZN(n2095) );
  AOI21_X1 U2294 ( .B1(n3517), .B2(n3461), .A(n3460), .ZN(n3615) );
  NAND2_X1 U2295 ( .A1(n4531), .A2(n3947), .ZN(n3948) );
  NAND2_X1 U2296 ( .A1(n3026), .A2(n3852), .ZN(n4206) );
  OR2_X1 U2297 ( .A1(n4352), .A2(n4366), .ZN(n2070) );
  NAND2_X1 U2298 ( .A1(n4533), .A2(n4532), .ZN(n4531) );
  OAI21_X1 U2299 ( .B1(n2008), .B2(n2276), .A(n2030), .ZN(n2275) );
  OAI21_X1 U2300 ( .B1(n4071), .B2(n4070), .A(n4069), .ZN(n4437) );
  NAND2_X1 U2301 ( .A1(n4124), .A2(n2318), .ZN(n4086) );
  XNOR2_X1 U2302 ( .A(n2080), .B(n4492), .ZN(n3939) );
  NAND2_X1 U2303 ( .A1(n2941), .A2(n2940), .ZN(n4774) );
  OR2_X1 U2304 ( .A1(n4504), .A2(n2052), .ZN(n2080) );
  AND2_X1 U2305 ( .A1(n2836), .A2(n2835), .ZN(n4048) );
  NAND2_X1 U2306 ( .A1(n2857), .A2(n2856), .ZN(n4065) );
  NAND2_X1 U2307 ( .A1(n2824), .A2(n2823), .ZN(n4102) );
  INV_X1 U2308 ( .A(n4201), .ZN(n2993) );
  NAND2_X1 U2309 ( .A1(n2798), .A2(REG3_REG_23__SCAN_IN), .ZN(n2818) );
  AND2_X1 U2310 ( .A1(n2750), .A2(n2749), .ZN(n4190) );
  AND2_X1 U2311 ( .A1(n2963), .A2(n2962), .ZN(n3443) );
  NAND2_X1 U2312 ( .A1(n3159), .A2(n3158), .ZN(n3161) );
  CLKBUF_X1 U2313 ( .A(n3010), .Z(n3813) );
  BUF_X1 U2314 ( .A(n3007), .Z(n3778) );
  NAND2_X1 U2315 ( .A1(n3145), .A2(REG1_REG_8__SCAN_IN), .ZN(n3159) );
  AND2_X1 U2316 ( .A1(n3818), .A2(n3815), .ZN(n3782) );
  XNOR2_X1 U2317 ( .A(n3155), .B(n4497), .ZN(n3145) );
  CLKBUF_X1 U2318 ( .A(n3901), .Z(n2064) );
  AND2_X1 U2319 ( .A1(n3224), .A2(n3169), .ZN(n3211) );
  INV_X1 U2320 ( .A(n3452), .ZN(n2317) );
  NAND2_X1 U2321 ( .A1(n2087), .A2(n2093), .ZN(n3155) );
  OR2_X2 U2322 ( .A1(n3204), .A2(n3169), .ZN(n3009) );
  NAND4_X2 U2323 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(n3896)
         );
  CLKBUF_X1 U2324 ( .A(n3204), .Z(n2058) );
  NAND4_X1 U2325 ( .A1(n2471), .A2(n2469), .A3(n2470), .A4(n2468), .ZN(n3899)
         );
  NAND2_X1 U2326 ( .A1(n2221), .A2(n2399), .ZN(n3204) );
  NAND4_X2 U2327 ( .A1(n2455), .A2(n2454), .A3(n2453), .A4(n2452), .ZN(n3900)
         );
  INV_X1 U2328 ( .A(n2954), .ZN(n3203) );
  INV_X1 U2329 ( .A(n2510), .ZN(n2805) );
  AND2_X2 U2330 ( .A1(n2397), .A2(n4483), .ZN(n2510) );
  NAND2_X1 U2331 ( .A1(n2388), .A2(IR_REG_31__SCAN_IN), .ZN(n2389) );
  AND2_X1 U2332 ( .A1(n2379), .A2(n2405), .ZN(n4488) );
  OR2_X1 U2333 ( .A1(n2931), .A2(n2167), .ZN(n2396) );
  AOI21_X1 U2334 ( .B1(n2170), .B2(n2172), .A(n2167), .ZN(n2166) );
  NOR2_X2 U2335 ( .A1(n2908), .A2(n2340), .ZN(n2931) );
  XNOR2_X1 U2336 ( .A(n2521), .B(IR_REG_6__SCAN_IN), .ZN(n4498) );
  NOR2_X1 U2337 ( .A1(n2498), .A2(n2305), .ZN(n2304) );
  AND2_X1 U2338 ( .A1(n2374), .A2(n2174), .ZN(n2173) );
  CLKBUF_X1 U2339 ( .A(n3912), .Z(n2103) );
  AND3_X1 U2340 ( .A1(n2004), .A2(n2372), .A3(n2365), .ZN(n2307) );
  AND2_X1 U2341 ( .A1(n2364), .A2(n2363), .ZN(n2365) );
  AND4_X1 U2342 ( .A1(n2360), .A2(n2362), .A3(n2361), .A4(n4635), .ZN(n2372)
         );
  OR2_X1 U2343 ( .A1(n2437), .A2(n2167), .ZN(n2439) );
  NAND2_X1 U2344 ( .A1(n2306), .A2(n2910), .ZN(n2305) );
  NOR2_X1 U2345 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2357)
         );
  INV_X1 U2346 ( .A(IR_REG_23__SCAN_IN), .ZN(n2910) );
  NOR2_X1 U2347 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2359)
         );
  NOR2_X1 U2348 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2358)
         );
  NOR2_X1 U2349 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2361)
         );
  NOR2_X1 U2350 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2362)
         );
  NOR2_X1 U2351 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2360)
         );
  CLKBUF_X1 U2352 ( .A(IR_REG_7__SCAN_IN), .Z(n4669) );
  NOR2_X1 U2353 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2345)
         );
  INV_X1 U2354 ( .A(IR_REG_6__SCAN_IN), .ZN(n4635) );
  NOR2_X2 U2355 ( .A1(n2488), .A2(n4634), .ZN(n2513) );
  NOR2_X4 U2356 ( .A1(n3210), .A2(n3288), .ZN(n3453) );
  OR2_X2 U2357 ( .A1(n3374), .A2(n3632), .ZN(n2353) );
  AOI21_X1 U2358 ( .B1(n2294), .B2(n2293), .A(n2034), .ZN(n2292) );
  INV_X1 U2359 ( .A(n2297), .ZN(n2293) );
  INV_X1 U2360 ( .A(IR_REG_19__SCAN_IN), .ZN(n2403) );
  AOI21_X1 U2361 ( .B1(n3851), .B2(n2266), .A(n2987), .ZN(n2265) );
  NOR2_X1 U2362 ( .A1(n2980), .A2(n2256), .ZN(n2255) );
  INV_X1 U2363 ( .A(n2149), .ZN(n2148) );
  AND2_X1 U2364 ( .A1(n2421), .A2(n4488), .ZN(n2176) );
  NAND2_X1 U2365 ( .A1(n4050), .A2(n4037), .ZN(n3870) );
  AND2_X1 U2366 ( .A1(n3955), .A2(REG1_REG_15__SCAN_IN), .ZN(n2101) );
  AND2_X1 U2367 ( .A1(n2959), .A2(n3279), .ZN(n2961) );
  NOR2_X1 U2368 ( .A1(n3900), .A2(n3288), .ZN(n2960) );
  AND2_X1 U2369 ( .A1(n2231), .A2(n3779), .ZN(n2230) );
  INV_X1 U2370 ( .A(n2171), .ZN(n2170) );
  OAI21_X1 U2371 ( .B1(n2173), .B2(n2172), .A(n2403), .ZN(n2171) );
  AND4_X1 U2372 ( .A1(n2373), .A2(n2701), .A3(n4694), .A4(n4753), .ZN(n2374)
         );
  AND2_X1 U2373 ( .A1(n3652), .A2(n2343), .ZN(n2342) );
  INV_X1 U2374 ( .A(n3651), .ZN(n2343) );
  AND2_X1 U2375 ( .A1(n3754), .A2(DATAI_21_), .ZN(n3569) );
  NAND2_X1 U2376 ( .A1(n3215), .A2(n3214), .ZN(n2322) );
  INV_X1 U2377 ( .A(n2943), .ZN(n2928) );
  INV_X1 U2378 ( .A(n2802), .ZN(n2868) );
  INV_X1 U2379 ( .A(n2490), .ZN(n2529) );
  INV_X2 U2380 ( .A(n2529), .ZN(n3751) );
  NAND2_X1 U2381 ( .A1(n2398), .A2(n2397), .ZN(n2490) );
  NAND2_X1 U2382 ( .A1(n3917), .A2(n3093), .ZN(n3094) );
  XNOR2_X1 U2383 ( .A(n3097), .B(n3096), .ZN(n3928) );
  NAND2_X1 U2384 ( .A1(n3967), .A2(n2197), .ZN(n4545) );
  OR2_X1 U2385 ( .A1(n4491), .A2(REG1_REG_17__SCAN_IN), .ZN(n2197) );
  AOI21_X1 U2386 ( .B1(n2194), .B2(n2193), .A(n2196), .ZN(n2192) );
  INV_X1 U2387 ( .A(n3960), .ZN(n2193) );
  NAND2_X1 U2388 ( .A1(n2282), .A2(n3005), .ZN(n2277) );
  INV_X1 U2389 ( .A(n2275), .ZN(n2274) );
  NAND2_X1 U2390 ( .A1(n3754), .A2(DATAI_25_), .ZN(n4070) );
  OR2_X1 U2391 ( .A1(n2408), .A2(n3149), .ZN(n4289) );
  NOR2_X2 U2392 ( .A1(n4086), .A2(n3469), .ZN(n4068) );
  INV_X1 U2393 ( .A(n3713), .ZN(n4055) );
  MUX2_X1 U2394 ( .A(n3979), .B(n2751), .S(n3754), .Z(n4181) );
  AND2_X1 U2395 ( .A1(n2345), .A2(n2306), .ZN(n2071) );
  INV_X1 U2396 ( .A(n2588), .ZN(n2151) );
  INV_X1 U2397 ( .A(n2016), .ZN(n2266) );
  NAND2_X1 U2398 ( .A1(n3204), .A2(n3169), .ZN(n3810) );
  INV_X1 U2399 ( .A(IR_REG_17__SCAN_IN), .ZN(n4694) );
  INV_X1 U2400 ( .A(n2461), .ZN(n2888) );
  OAI21_X1 U2401 ( .B1(n2332), .B2(n2330), .A(n3672), .ZN(n2329) );
  INV_X1 U2402 ( .A(n2612), .ZN(n2327) );
  NAND2_X1 U2403 ( .A1(n2612), .A2(n2331), .ZN(n2330) );
  INV_X1 U2404 ( .A(n3671), .ZN(n2331) );
  INV_X1 U2405 ( .A(n2326), .ZN(n2325) );
  OAI21_X1 U2406 ( .B1(n2332), .B2(n2327), .A(n3671), .ZN(n2326) );
  OAI22_X1 U2407 ( .A1(n2715), .A2(n2164), .B1(n2714), .B2(n3589), .ZN(n2163)
         );
  INV_X1 U2408 ( .A(n3508), .ZN(n2164) );
  OR2_X1 U2409 ( .A1(n3642), .A2(n2046), .ZN(n2336) );
  INV_X1 U2410 ( .A(n3526), .ZN(n2332) );
  AOI21_X1 U2411 ( .B1(n2161), .B2(n2715), .A(n2158), .ZN(n2157) );
  INV_X1 U2412 ( .A(n3605), .ZN(n2158) );
  INV_X1 U2413 ( .A(n4483), .ZN(n2398) );
  OR2_X1 U2414 ( .A1(n2490), .A2(n2412), .ZN(n2416) );
  INV_X1 U2415 ( .A(n3984), .ZN(n4022) );
  INV_X1 U2416 ( .A(n3003), .ZN(n2279) );
  NAND2_X1 U2417 ( .A1(n2352), .A2(n2351), .ZN(n2296) );
  AND2_X1 U2418 ( .A1(n2042), .A2(n2984), .ZN(n2219) );
  AND2_X1 U2419 ( .A1(n2254), .A2(n2257), .ZN(n2253) );
  OR2_X1 U2420 ( .A1(n3897), .A2(n3702), .ZN(n2969) );
  NAND2_X1 U2421 ( .A1(n2085), .A2(n2084), .ZN(n3825) );
  INV_X1 U2422 ( .A(n2970), .ZN(n2084) );
  INV_X1 U2423 ( .A(n3896), .ZN(n2085) );
  NAND2_X1 U2424 ( .A1(n3896), .A2(n2970), .ZN(n3828) );
  NAND2_X1 U2425 ( .A1(n2964), .A2(n2317), .ZN(n3819) );
  AND2_X1 U2426 ( .A1(n4487), .A2(n4488), .ZN(n3070) );
  INV_X1 U2427 ( .A(n4487), .ZN(n2944) );
  INV_X1 U2428 ( .A(IR_REG_28__SCAN_IN), .ZN(n2394) );
  INV_X1 U2429 ( .A(IR_REG_21__SCAN_IN), .ZN(n2364) );
  INV_X1 U2430 ( .A(IR_REG_25__SCAN_IN), .ZN(n2381) );
  CLKBUF_X1 U2431 ( .A(n2908), .Z(n2909) );
  OR2_X1 U2432 ( .A1(n2851), .A2(n2850), .ZN(n2866) );
  NAND2_X1 U2433 ( .A1(n2098), .A2(REG3_REG_13__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U2434 ( .A1(n2146), .A2(n2147), .ZN(n3527) );
  OR2_X1 U2435 ( .A1(n2149), .A2(n2036), .ZN(n2147) );
  INV_X1 U2436 ( .A(n3901), .ZN(n3181) );
  INV_X1 U2437 ( .A(n4070), .ZN(n3469) );
  NAND2_X1 U2438 ( .A1(n3509), .A2(n2165), .ZN(n2162) );
  INV_X1 U2439 ( .A(n2163), .ZN(n2160) );
  INV_X1 U2440 ( .A(n2800), .ZN(n2798) );
  NAND2_X1 U2441 ( .A1(n3489), .A2(n3488), .ZN(n2334) );
  INV_X1 U2442 ( .A(n2152), .ZN(n3639) );
  OAI21_X1 U2443 ( .B1(n3509), .B2(n2156), .A(n2153), .ZN(n2152) );
  NAND2_X1 U2444 ( .A1(n2757), .A2(n2161), .ZN(n2156) );
  NOR2_X1 U2445 ( .A1(n2756), .A2(n2154), .ZN(n2153) );
  AND2_X1 U2446 ( .A1(n2770), .A2(n2769), .ZN(n3642) );
  NAND2_X1 U2447 ( .A1(n3663), .A2(n3664), .ZN(n3662) );
  NAND2_X1 U2448 ( .A1(n2333), .A2(n2332), .ZN(n3528) );
  INV_X1 U2449 ( .A(n3527), .ZN(n2333) );
  OR2_X1 U2450 ( .A1(n2570), .A2(n3493), .ZN(n2536) );
  OR2_X1 U2451 ( .A1(n2570), .A2(n3323), .ZN(n2492) );
  NAND2_X1 U2452 ( .A1(n4483), .A2(n4482), .ZN(n2512) );
  NAND2_X1 U2453 ( .A1(n2467), .A2(REG2_REG_3__SCAN_IN), .ZN(n2453) );
  XNOR2_X1 U2454 ( .A(n4503), .B(n2199), .ZN(n3434) );
  INV_X1 U2455 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2199) );
  OAI211_X1 U2456 ( .C1(n2198), .C2(REG2_REG_1__SCAN_IN), .A(n3436), .B(n2183), 
        .ZN(n3914) );
  NAND2_X1 U2457 ( .A1(n2198), .A2(REG2_REG_1__SCAN_IN), .ZN(n2183) );
  NAND2_X1 U2458 ( .A1(n2198), .A2(REG2_REG_1__SCAN_IN), .ZN(n3913) );
  NAND2_X1 U2459 ( .A1(n2106), .A2(n3095), .ZN(n3097) );
  NAND2_X1 U2460 ( .A1(n3105), .A2(REG2_REG_3__SCAN_IN), .ZN(n2106) );
  NAND2_X1 U2461 ( .A1(n2124), .A2(n2123), .ZN(n2122) );
  AND2_X1 U2462 ( .A1(n2123), .A2(n4498), .ZN(n2121) );
  NAND2_X1 U2463 ( .A1(n3142), .A2(n3141), .ZN(n3152) );
  NAND2_X1 U2464 ( .A1(n2208), .A2(REG2_REG_7__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U2465 ( .A1(n3144), .A2(n2530), .ZN(n2093) );
  AND2_X1 U2466 ( .A1(n2206), .A2(n2006), .ZN(n2088) );
  INV_X1 U2467 ( .A(n2132), .ZN(n2131) );
  OAI22_X1 U2468 ( .A1(n2140), .A2(n2133), .B1(n4495), .B2(n2044), .ZN(n2132)
         );
  NAND2_X1 U2469 ( .A1(n3236), .A2(n2134), .ZN(n2133) );
  INV_X1 U2470 ( .A(n3229), .ZN(n2134) );
  AOI21_X1 U2471 ( .B1(n3329), .B2(n2012), .A(n2128), .ZN(n2181) );
  AOI21_X1 U2472 ( .B1(n2138), .B2(n2137), .A(n2136), .ZN(n2128) );
  NAND2_X1 U2473 ( .A1(n2178), .A2(n4495), .ZN(n2136) );
  INV_X1 U2474 ( .A(n2130), .ZN(n2138) );
  OAI21_X1 U2475 ( .B1(n2140), .B2(n3229), .A(n2044), .ZN(n2130) );
  NAND2_X1 U2476 ( .A1(n3153), .A2(n2045), .ZN(n2137) );
  INV_X1 U2477 ( .A(n3327), .ZN(n2215) );
  NAND2_X1 U2478 ( .A1(n4494), .A2(REG1_REG_11__SCAN_IN), .ZN(n2091) );
  NAND2_X1 U2479 ( .A1(n2080), .A2(n2212), .ZN(n2211) );
  NAND2_X1 U2480 ( .A1(n4528), .A2(n3958), .ZN(n3959) );
  INV_X1 U2481 ( .A(n4543), .ZN(n2195) );
  NOR2_X1 U2482 ( .A1(n3756), .A2(n3872), .ZN(n2267) );
  INV_X1 U2483 ( .A(n2284), .ZN(n2283) );
  NAND2_X1 U2484 ( .A1(n2270), .A2(n2268), .ZN(n4032) );
  INV_X1 U2485 ( .A(n2271), .ZN(n2268) );
  NAND2_X1 U2486 ( .A1(n2097), .A2(REG3_REG_25__SCAN_IN), .ZN(n2851) );
  NAND2_X1 U2487 ( .A1(n2100), .A2(n2054), .ZN(n2789) );
  AND2_X1 U2488 ( .A1(n4153), .A2(n4138), .ZN(n2997) );
  AND2_X1 U2489 ( .A1(n4118), .A2(n3569), .ZN(n2083) );
  NOR2_X1 U2490 ( .A1(n2993), .A2(n2298), .ZN(n2297) );
  INV_X1 U2491 ( .A(n2351), .ZN(n2298) );
  NAND2_X1 U2492 ( .A1(n2300), .A2(n2302), .ZN(n2299) );
  OR2_X1 U2493 ( .A1(n4182), .A2(n2802), .ZN(n2750) );
  INV_X1 U2494 ( .A(n2014), .ZN(n2300) );
  INV_X1 U2495 ( .A(n2099), .ZN(n2693) );
  NAND2_X1 U2496 ( .A1(n2260), .A2(n2258), .ZN(n4222) );
  AOI21_X1 U2497 ( .B1(n2262), .B2(n2264), .A(n2259), .ZN(n2258) );
  INV_X1 U2498 ( .A(n3739), .ZN(n2259) );
  NAND2_X1 U2499 ( .A1(n2217), .A2(n3839), .ZN(n4317) );
  AND2_X1 U2500 ( .A1(n3420), .A2(n3843), .ZN(n4316) );
  CLKBUF_X1 U2501 ( .A(n3372), .Z(n3373) );
  NAND2_X1 U2502 ( .A1(n2244), .A2(n2245), .ZN(n3263) );
  AOI21_X1 U2503 ( .B1(n2248), .B2(n2251), .A(n2246), .ZN(n2245) );
  INV_X1 U2504 ( .A(n3821), .ZN(n2246) );
  NOR2_X1 U2505 ( .A1(n2961), .A2(n2960), .ZN(n2962) );
  AND2_X1 U2506 ( .A1(n2959), .A2(n3197), .ZN(n2957) );
  NAND2_X1 U2507 ( .A1(n3778), .A2(n2028), .ZN(n2227) );
  AND2_X1 U2508 ( .A1(n3881), .A2(n3037), .ZN(n4330) );
  AND2_X1 U2509 ( .A1(n3070), .A2(n3904), .ZN(n4293) );
  OR2_X1 U2510 ( .A1(n3039), .A2(n3904), .ZN(n4320) );
  INV_X1 U2511 ( .A(n3900), .ZN(n3446) );
  NAND2_X1 U2512 ( .A1(n4017), .A2(n4016), .ZN(n4342) );
  INV_X1 U2513 ( .A(n4015), .ZN(n4016) );
  NAND2_X1 U2514 ( .A1(n4010), .A2(n4268), .ZN(n4017) );
  OAI21_X1 U2515 ( .B1(n4014), .B2(n4320), .A(n4013), .ZN(n4015) );
  NOR2_X1 U2516 ( .A1(n3621), .A2(n2320), .ZN(n2318) );
  NAND2_X1 U2517 ( .A1(n2895), .A2(n2894), .ZN(n3064) );
  NAND2_X1 U2518 ( .A1(n2341), .A2(n2394), .ZN(n2340) );
  INV_X1 U2519 ( .A(n2393), .ZN(n2341) );
  NAND2_X1 U2520 ( .A1(n3475), .A2(IR_REG_31__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U2521 ( .A1(n2382), .A2(n2381), .ZN(n2388) );
  INV_X1 U2522 ( .A(n2384), .ZN(n2382) );
  OR2_X1 U2523 ( .A1(n2378), .A2(IR_REG_21__SCAN_IN), .ZN(n2405) );
  INV_X1 U2524 ( .A(IR_REG_20__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U2525 ( .A1(n2168), .A2(n2166), .ZN(n2376) );
  NAND2_X1 U2526 ( .A1(n2668), .A2(n2374), .ZN(n2740) );
  INV_X1 U2527 ( .A(IR_REG_16__SCAN_IN), .ZN(n4753) );
  INV_X1 U2528 ( .A(IR_REG_4__SCAN_IN), .ZN(n2475) );
  OAI21_X1 U2529 ( .B1(n3712), .B2(n3710), .A(n3708), .ZN(n3500) );
  NAND2_X1 U2530 ( .A1(n3749), .A2(DATAI_23_), .ZN(n4105) );
  NAND2_X1 U2531 ( .A1(n3189), .A2(n2449), .ZN(n3215) );
  NOR2_X1 U2532 ( .A1(n3500), .A2(n3499), .ZN(n2953) );
  INV_X1 U2533 ( .A(n4118), .ZN(n4153) );
  OR2_X1 U2534 ( .A1(n2928), .A2(n2913), .ZN(n3719) );
  INV_X1 U2535 ( .A(n3689), .ZN(n3731) );
  INV_X1 U2536 ( .A(n3716), .ZN(n3728) );
  INV_X1 U2537 ( .A(n4014), .ZN(n4035) );
  NAND2_X1 U2538 ( .A1(n2796), .A2(n2795), .ZN(n3891) );
  NAND4_X1 U2539 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n3894)
         );
  NOR2_X1 U2540 ( .A1(n3134), .A2(n3133), .ZN(n3132) );
  XNOR2_X1 U2541 ( .A(n3152), .B(n3156), .ZN(n3153) );
  NAND2_X1 U2542 ( .A1(n4547), .A2(n4535), .ZN(n4551) );
  XNOR2_X1 U2543 ( .A(n2404), .B(n2403), .ZN(n3979) );
  NAND2_X1 U2544 ( .A1(n2169), .A2(IR_REG_31__SCAN_IN), .ZN(n2404) );
  AND2_X1 U2545 ( .A1(n4576), .A2(REG1_REG_18__SCAN_IN), .ZN(n2102) );
  XNOR2_X1 U2546 ( .A(n2086), .B(n2018), .ZN(n4354) );
  NAND2_X1 U2547 ( .A1(n4435), .A2(n4416), .ZN(n2062) );
  NAND2_X1 U2548 ( .A1(n4416), .A2(n4602), .ZN(n4419) );
  OR2_X1 U2549 ( .A1(n4437), .A2(n4480), .ZN(n2082) );
  NOR2_X1 U2550 ( .A1(n2242), .A2(n3016), .ZN(n2241) );
  INV_X1 U2551 ( .A(n3824), .ZN(n2242) );
  NOR2_X1 U2552 ( .A1(n2626), .A2(n2625), .ZN(n2098) );
  NAND2_X1 U2553 ( .A1(n2150), .A2(n2025), .ZN(n2149) );
  OR2_X1 U2554 ( .A1(n2019), .A2(n2151), .ZN(n2150) );
  INV_X1 U2555 ( .A(IR_REG_27__SCAN_IN), .ZN(n2367) );
  AND2_X1 U2556 ( .A1(n2757), .A2(n2155), .ZN(n2154) );
  INV_X1 U2557 ( .A(n2157), .ZN(n2155) );
  NAND2_X1 U2558 ( .A1(n2356), .A2(n2755), .ZN(n2756) );
  INV_X1 U2559 ( .A(n3542), .ZN(n2755) );
  INV_X1 U2560 ( .A(n2858), .ZN(n2885) );
  NOR2_X1 U2561 ( .A1(n3509), .A2(n3508), .ZN(n3591) );
  INV_X1 U2562 ( .A(n3330), .ZN(n2178) );
  OAI21_X1 U2563 ( .B1(n2011), .B2(n2043), .A(n2143), .ZN(n2142) );
  INV_X1 U2564 ( .A(n4508), .ZN(n2143) );
  NAND3_X1 U2565 ( .A1(n2186), .A2(n2184), .A3(n2053), .ZN(n3957) );
  INV_X1 U2566 ( .A(n3005), .ZN(n2276) );
  OAI21_X1 U2567 ( .B1(n3872), .B2(n3771), .A(n3760), .ZN(n2271) );
  OR2_X1 U2568 ( .A1(n3891), .A2(n4125), .ZN(n4098) );
  AOI21_X1 U2569 ( .B1(n2292), .B2(n2295), .A(n2301), .ZN(n2290) );
  NOR2_X1 U2570 ( .A1(n2744), .A2(n2743), .ZN(n2100) );
  NOR2_X1 U2571 ( .A1(n2678), .A2(n2677), .ZN(n2099) );
  AOI21_X1 U2572 ( .B1(n2265), .B2(n2263), .A(n2032), .ZN(n2262) );
  INV_X1 U2573 ( .A(n3851), .ZN(n2263) );
  INV_X1 U2574 ( .A(n2265), .ZN(n2264) );
  OAI21_X1 U2575 ( .B1(n3421), .B2(n2266), .A(n3851), .ZN(n4266) );
  NAND2_X1 U2576 ( .A1(n2261), .A2(n2265), .ZN(n4265) );
  NAND2_X1 U2577 ( .A1(n3421), .A2(n3851), .ZN(n2261) );
  INV_X1 U2578 ( .A(n2098), .ZN(n2647) );
  OR2_X1 U2579 ( .A1(n2572), .A2(n2571), .ZN(n2591) );
  INV_X1 U2580 ( .A(n3829), .ZN(n2236) );
  INV_X1 U2581 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2552) );
  OR2_X1 U2582 ( .A1(n2553), .A2(n2552), .ZN(n2572) );
  AOI21_X1 U2583 ( .B1(n2241), .B2(n3836), .A(n2239), .ZN(n2238) );
  INV_X1 U2584 ( .A(n3828), .ZN(n2239) );
  INV_X1 U2585 ( .A(n2241), .ZN(n2240) );
  INV_X1 U2586 ( .A(n3263), .ZN(n3015) );
  NOR2_X1 U2587 ( .A1(n2250), .A2(n2249), .ZN(n2248) );
  NOR2_X1 U2588 ( .A1(n3819), .A2(n2251), .ZN(n2249) );
  INV_X1 U2589 ( .A(n3835), .ZN(n2250) );
  INV_X1 U2590 ( .A(n3822), .ZN(n2251) );
  NAND2_X1 U2591 ( .A1(n3778), .A2(n3009), .ZN(n2229) );
  NOR2_X1 U2592 ( .A1(n2311), .A2(n4022), .ZN(n2310) );
  INV_X1 U2593 ( .A(n2312), .ZN(n2311) );
  NOR2_X1 U2594 ( .A1(n4001), .A2(n3501), .ZN(n2312) );
  NOR2_X1 U2595 ( .A1(n4251), .A2(n4233), .ZN(n2315) );
  NOR2_X1 U2596 ( .A1(n3582), .A2(n4327), .ZN(n2308) );
  INV_X1 U2597 ( .A(IR_REG_26__SCAN_IN), .ZN(n2391) );
  INV_X1 U2598 ( .A(IR_REG_24__SCAN_IN), .ZN(n4693) );
  INV_X1 U2599 ( .A(IR_REG_3__SCAN_IN), .ZN(n2472) );
  OR2_X1 U2600 ( .A1(n2660), .A2(n2659), .ZN(n2678) );
  NOR2_X1 U2601 ( .A1(n2328), .A2(n2325), .ZN(n2324) );
  AOI22_X1 U2602 ( .A1(n2328), .A2(n2330), .B1(n2325), .B2(n2327), .ZN(n2323)
         );
  INV_X1 U2603 ( .A(n2329), .ZN(n2328) );
  AND2_X1 U2604 ( .A1(n3754), .A2(DATAI_24_), .ZN(n3621) );
  AND2_X1 U2605 ( .A1(n3517), .A2(n3459), .ZN(n3616) );
  OR2_X1 U2606 ( .A1(n2426), .A2(n2422), .ZN(n3221) );
  NOR2_X1 U2607 ( .A1(n3639), .A2(n3640), .ZN(n3638) );
  NAND2_X1 U2608 ( .A1(n2336), .A2(n2337), .ZN(n2335) );
  XNOR2_X1 U2609 ( .A(n2407), .B(n2886), .ZN(n2429) );
  OAI21_X1 U2610 ( .B1(n3509), .B2(n2159), .A(n2157), .ZN(n3686) );
  AND2_X1 U2611 ( .A1(n3058), .A2(n3253), .ZN(n2943) );
  OR2_X1 U2612 ( .A1(n2512), .A2(n3196), .ZN(n2432) );
  AND3_X1 U2613 ( .A1(n2223), .A2(n2225), .A3(n2222), .ZN(n2221) );
  NAND2_X1 U2614 ( .A1(n2398), .A2(n2224), .ZN(n2223) );
  NAND2_X1 U2615 ( .A1(n2418), .A2(n2417), .ZN(n3901) );
  OR2_X1 U2616 ( .A1(n2570), .A2(n3123), .ZN(n2417) );
  AND3_X1 U2617 ( .A1(n2416), .A2(n2414), .A3(n2415), .ZN(n2418) );
  NAND2_X1 U2618 ( .A1(n2127), .A2(n4498), .ZN(n2124) );
  NAND2_X1 U2619 ( .A1(n2007), .A2(n2355), .ZN(n2206) );
  AND2_X1 U2620 ( .A1(n3235), .A2(REG1_REG_10__SCAN_IN), .ZN(n3326) );
  AND2_X1 U2621 ( .A1(n2181), .A2(n2180), .ZN(n3934) );
  NAND2_X1 U2622 ( .A1(n4494), .A2(REG2_REG_11__SCAN_IN), .ZN(n2180) );
  NAND2_X1 U2623 ( .A1(n2090), .A2(n4493), .ZN(n2065) );
  NAND2_X1 U2624 ( .A1(n2145), .A2(n2144), .ZN(n3952) );
  NAND2_X1 U2625 ( .A1(n4514), .A2(n4301), .ZN(n2144) );
  OAI21_X1 U2626 ( .B1(n3934), .B2(n2011), .A(n2141), .ZN(n2145) );
  INV_X1 U2627 ( .A(n2142), .ZN(n2141) );
  NAND2_X1 U2628 ( .A1(n3953), .A2(n2185), .ZN(n2184) );
  INV_X1 U2629 ( .A(n4516), .ZN(n2185) );
  OR2_X1 U2630 ( .A1(n3937), .A2(n2187), .ZN(n2186) );
  OR2_X1 U2631 ( .A1(n4516), .A2(n2662), .ZN(n2187) );
  INV_X1 U2632 ( .A(n4521), .ZN(n2078) );
  XNOR2_X1 U2633 ( .A(n3957), .B(n4579), .ZN(n4530) );
  NAND2_X1 U2634 ( .A1(n4530), .A2(n4529), .ZN(n4528) );
  INV_X1 U2635 ( .A(IR_REG_18__SCAN_IN), .ZN(n2174) );
  OR2_X1 U2636 ( .A1(n2020), .A2(n2286), .ZN(n2281) );
  NAND2_X1 U2637 ( .A1(n2282), .A2(n2279), .ZN(n2278) );
  AND2_X1 U2638 ( .A1(n3004), .A2(n2023), .ZN(n2286) );
  AND2_X1 U2639 ( .A1(n2866), .A2(n2852), .ZN(n4056) );
  NOR2_X1 U2640 ( .A1(n4061), .A2(n3748), .ZN(n4045) );
  INV_X1 U2641 ( .A(n2097), .ZN(n2830) );
  NAND2_X1 U2642 ( .A1(n2234), .A2(n3789), .ZN(n4080) );
  AND2_X1 U2643 ( .A1(n4097), .A2(n4096), .ZN(n4116) );
  AND2_X1 U2644 ( .A1(n2808), .A2(n2807), .ZN(n4120) );
  OR2_X1 U2645 ( .A1(n4107), .A2(n2802), .ZN(n2808) );
  NAND2_X1 U2646 ( .A1(n2788), .A2(REG3_REG_22__SCAN_IN), .ZN(n2800) );
  INV_X1 U2647 ( .A(n2789), .ZN(n2788) );
  INV_X1 U2648 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2743) );
  INV_X1 U2649 ( .A(n2100), .ZN(n2772) );
  AND2_X1 U2650 ( .A1(n2739), .A2(n2738), .ZN(n4175) );
  OR2_X1 U2651 ( .A1(n4197), .A2(n2802), .ZN(n2739) );
  OR2_X1 U2652 ( .A1(n2716), .A2(n4719), .ZN(n2733) );
  NAND2_X1 U2653 ( .A1(n2731), .A2(REG3_REG_18__SCAN_IN), .ZN(n2744) );
  INV_X1 U2654 ( .A(n2733), .ZN(n2731) );
  AND3_X1 U2655 ( .A1(n2700), .A2(n2699), .A3(n2698), .ZN(n4208) );
  NAND2_X1 U2656 ( .A1(n2099), .A2(REG3_REG_16__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U2657 ( .A1(n2590), .A2(REG3_REG_10__SCAN_IN), .ZN(n2626) );
  INV_X1 U2658 ( .A(n2591), .ZN(n2590) );
  NAND2_X1 U2659 ( .A1(n2252), .A2(n2253), .ZN(n4309) );
  NAND2_X1 U2660 ( .A1(n2218), .A2(n3830), .ZN(n3405) );
  INV_X1 U2661 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2531) );
  OR2_X1 U2662 ( .A1(n2532), .A2(n2531), .ZN(n2553) );
  NAND2_X1 U2663 ( .A1(n2243), .A2(n3824), .ZN(n3336) );
  NAND2_X1 U2664 ( .A1(n3015), .A2(n3014), .ZN(n2243) );
  CLKBUF_X1 U2665 ( .A(n3267), .Z(n3293) );
  NAND2_X1 U2666 ( .A1(n2247), .A2(n3822), .ZN(n3294) );
  NAND2_X1 U2667 ( .A1(n3013), .A2(n3819), .ZN(n2247) );
  NAND2_X1 U2668 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2488) );
  NAND2_X1 U2669 ( .A1(n3453), .A2(n3452), .ZN(n3451) );
  NOR2_X1 U2670 ( .A1(n2958), .A2(n3203), .ZN(n3279) );
  INV_X1 U2671 ( .A(n4320), .ZN(n4223) );
  NAND2_X1 U2672 ( .A1(n2200), .A2(n2107), .ZN(n3169) );
  NAND2_X1 U2673 ( .A1(n2636), .A2(n2201), .ZN(n2107) );
  AND2_X1 U2674 ( .A1(n3901), .A2(n3008), .ZN(n3166) );
  AND2_X1 U2675 ( .A1(n3177), .A2(n3047), .ZN(n3252) );
  NAND2_X1 U2676 ( .A1(n3181), .A2(n3008), .ZN(n3809) );
  INV_X1 U2677 ( .A(n4289), .ZN(n4326) );
  AND2_X1 U2678 ( .A1(n3754), .A2(DATAI_28_), .ZN(n4001) );
  NAND2_X1 U2679 ( .A1(n4053), .A2(n2312), .ZN(n4021) );
  NAND2_X1 U2680 ( .A1(n4053), .A2(n4037), .ZN(n4036) );
  NAND2_X1 U2681 ( .A1(n4124), .A2(n2319), .ZN(n4085) );
  AND2_X1 U2682 ( .A1(n4124), .A2(n4125), .ZN(n4368) );
  NOR2_X2 U2683 ( .A1(n4159), .A2(n3569), .ZN(n4124) );
  NOR2_X1 U2684 ( .A1(n4216), .A2(n4193), .ZN(n4196) );
  NAND2_X1 U2685 ( .A1(n2315), .A2(n4207), .ZN(n4216) );
  INV_X1 U2686 ( .A(n2315), .ZN(n4393) );
  NAND2_X1 U2687 ( .A1(n4312), .A2(n2308), .ZN(n4296) );
  NAND2_X1 U2688 ( .A1(n4312), .A2(n4311), .ZN(n4310) );
  NAND3_X1 U2689 ( .A1(n3453), .A2(n2966), .A3(n2316), .ZN(n3341) );
  NOR2_X1 U2690 ( .A1(n2317), .A2(n3702), .ZN(n2316) );
  AND2_X1 U2691 ( .A1(n4562), .A2(n2944), .ZN(n4595) );
  NAND2_X1 U2692 ( .A1(n2384), .A2(n2387), .ZN(n2892) );
  XNOR2_X1 U2693 ( .A(n2911), .B(n2910), .ZN(n3069) );
  OR2_X1 U2694 ( .A1(n2722), .A2(IR_REG_14__SCAN_IN), .ZN(n2686) );
  INV_X1 U2695 ( .A(IR_REG_15__SCAN_IN), .ZN(n2701) );
  INV_X1 U2696 ( .A(IR_REG_11__SCAN_IN), .ZN(n2632) );
  OR3_X1 U2697 ( .A1(n2578), .A2(IR_REG_8__SCAN_IN), .A3(n4669), .ZN(n2597) );
  INV_X1 U2698 ( .A(n2970), .ZN(n3492) );
  AND2_X1 U2699 ( .A1(n2916), .A2(n3726), .ZN(n2917) );
  NAND2_X1 U2700 ( .A1(n2334), .A2(n2551), .ZN(n3554) );
  INV_X1 U2701 ( .A(n3169), .ZN(n2956) );
  NOR2_X1 U2702 ( .A1(n3638), .A2(n3642), .ZN(n3568) );
  NAND2_X1 U2703 ( .A1(n2162), .A2(n2160), .ZN(n3608) );
  INV_X1 U2704 ( .A(n3243), .ZN(n2321) );
  NAND2_X1 U2705 ( .A1(n2334), .A2(n2019), .ZN(n3627) );
  INV_X1 U2706 ( .A(DATAI_0_), .ZN(n2303) );
  AND2_X1 U2707 ( .A1(n3754), .A2(DATAI_20_), .ZN(n4150) );
  NAND2_X1 U2708 ( .A1(n3749), .A2(DATAI_22_), .ZN(n4125) );
  NAND2_X1 U2709 ( .A1(n3528), .A2(n2612), .ZN(n3674) );
  INV_X1 U2710 ( .A(n3719), .ZN(n3726) );
  OR2_X1 U2711 ( .A1(n4073), .A2(n2802), .ZN(n2836) );
  NAND2_X1 U2712 ( .A1(n2943), .A2(n3885), .ZN(n3716) );
  OR2_X1 U2713 ( .A1(n2847), .A2(n2846), .ZN(n2848) );
  NAND2_X1 U2714 ( .A1(n2873), .A2(n2872), .ZN(n4050) );
  INV_X1 U2715 ( .A(n4048), .ZN(n4082) );
  INV_X1 U2716 ( .A(n4120), .ZN(n3890) );
  NAND2_X1 U2717 ( .A1(n2778), .A2(n2777), .ZN(n4118) );
  INV_X1 U2718 ( .A(n4190), .ZN(n4151) );
  INV_X1 U2719 ( .A(n4175), .ZN(n4210) );
  INV_X1 U2720 ( .A(n4208), .ZN(n4243) );
  OR2_X1 U2721 ( .A1(n2685), .A2(n2684), .ZN(n4264) );
  NAND4_X1 U2722 ( .A1(n2652), .A2(n2651), .A3(n2650), .A4(n2649), .ZN(n4261)
         );
  OR2_X1 U2723 ( .A1(n2451), .A2(n2534), .ZN(n2535) );
  AND3_X1 U2724 ( .A1(n2519), .A2(n2518), .A3(n2041), .ZN(n2063) );
  OR2_X1 U2725 ( .A1(n3751), .A2(n2511), .ZN(n2520) );
  OR2_X1 U2726 ( .A1(n2451), .A2(n3298), .ZN(n2496) );
  NOR2_X1 U2727 ( .A1(n2805), .A2(n2493), .ZN(n2494) );
  OR2_X1 U2728 ( .A1(n2490), .A2(n2450), .ZN(n2454) );
  CLKBUF_X1 U2729 ( .A(n2958), .Z(n2436) );
  INV_X1 U2730 ( .A(n2198), .ZN(n2201) );
  NAND2_X1 U2731 ( .A1(n3092), .A2(n2182), .ZN(n3917) );
  NAND2_X1 U2732 ( .A1(n3913), .A2(n3914), .ZN(n2182) );
  XNOR2_X1 U2733 ( .A(n3094), .B(n3107), .ZN(n3105) );
  AOI21_X1 U2734 ( .B1(n3928), .B2(REG2_REG_4__SCAN_IN), .A(n3098), .ZN(n3134)
         );
  NAND2_X1 U2735 ( .A1(n2205), .A2(n2204), .ZN(n2210) );
  INV_X1 U2736 ( .A(n2355), .ZN(n2204) );
  NAND2_X1 U2737 ( .A1(n2116), .A2(n2114), .ZN(n3142) );
  NAND2_X1 U2738 ( .A1(n2117), .A2(n2120), .ZN(n2113) );
  AOI21_X1 U2739 ( .B1(n3153), .B2(REG2_REG_8__SCAN_IN), .A(n2139), .ZN(n3230)
         );
  INV_X1 U2740 ( .A(n2140), .ZN(n2139) );
  NAND2_X1 U2741 ( .A1(n3157), .A2(n4497), .ZN(n3158) );
  NAND2_X1 U2742 ( .A1(n2035), .A2(n2129), .ZN(n3329) );
  NAND2_X1 U2743 ( .A1(n3153), .A2(n2047), .ZN(n2135) );
  AOI21_X1 U2744 ( .B1(n3329), .B2(REG2_REG_10__SCAN_IN), .A(n2179), .ZN(n3331) );
  AOI21_X1 U2745 ( .B1(n2138), .B2(n2137), .A(n3236), .ZN(n2179) );
  NAND2_X1 U2746 ( .A1(n3325), .A2(n2215), .ZN(n2213) );
  NOR2_X1 U2747 ( .A1(n3326), .A2(n3325), .ZN(n3328) );
  XNOR2_X1 U2748 ( .A(n2633), .B(n2632), .ZN(n3395) );
  XNOR2_X1 U2749 ( .A(n3934), .B(n2089), .ZN(n3936) );
  XNOR2_X1 U2750 ( .A(n2090), .B(n2089), .ZN(n3399) );
  NAND2_X1 U2751 ( .A1(n3399), .A2(REG1_REG_12__SCAN_IN), .ZN(n3938) );
  AOI21_X1 U2752 ( .B1(n3934), .B2(n2043), .A(n2011), .ZN(n4510) );
  OR2_X1 U2753 ( .A1(n3937), .A2(n2662), .ZN(n2189) );
  XNOR2_X1 U2754 ( .A(n3952), .B(n4492), .ZN(n3937) );
  NAND2_X1 U2755 ( .A1(n2186), .A2(n2184), .ZN(n4515) );
  NAND2_X1 U2756 ( .A1(n4542), .A2(n4543), .ZN(n2111) );
  NAND2_X1 U2757 ( .A1(n3974), .A2(n3973), .ZN(n4542) );
  AOI21_X1 U2758 ( .B1(n3974), .B2(n2194), .A(n4541), .ZN(n2110) );
  INV_X1 U2759 ( .A(n4548), .ZN(n4540) );
  AOI21_X1 U2760 ( .B1(n2191), .B2(n2194), .A(n2190), .ZN(n3976) );
  INV_X1 U2761 ( .A(n2192), .ZN(n2190) );
  NOR2_X1 U2762 ( .A1(n3125), .A2(n3099), .ZN(n4537) );
  INV_X1 U2763 ( .A(n2096), .ZN(n3487) );
  OAI21_X1 U2764 ( .B1(n3038), .B2(n4330), .A(n3043), .ZN(n2096) );
  AOI21_X1 U2765 ( .B1(n4035), .B2(n4293), .A(n4034), .ZN(n2104) );
  OR2_X1 U2766 ( .A1(n4033), .A2(n4330), .ZN(n2105) );
  NAND2_X1 U2767 ( .A1(n2014), .A2(n2297), .ZN(n2291) );
  AND2_X1 U2768 ( .A1(n2299), .A2(n2297), .ZN(n4203) );
  CLKBUF_X1 U2769 ( .A(n3425), .Z(n3426) );
  OAI21_X1 U2770 ( .B1(n3373), .B2(n2021), .A(n2979), .ZN(n3403) );
  CLKBUF_X1 U2771 ( .A(n3354), .Z(n3355) );
  OR2_X1 U2772 ( .A1(n3340), .A2(n4366), .ZN(n4315) );
  AND2_X1 U2773 ( .A1(n4570), .A2(n3273), .ZN(n4255) );
  INV_X1 U2774 ( .A(n4255), .ZN(n4143) );
  INV_X1 U2775 ( .A(n4566), .ZN(n4313) );
  AND2_X1 U2776 ( .A1(n2408), .A2(n4490), .ZN(n4562) );
  AND2_X1 U2777 ( .A1(n4570), .A2(n3255), .ZN(n4568) );
  XOR2_X1 U2778 ( .A(n3987), .B(n3990), .Z(n4424) );
  NAND2_X1 U2779 ( .A1(n3064), .A2(n3177), .ZN(n4573) );
  NOR2_X1 U2780 ( .A1(n2340), .A2(IR_REG_29__SCAN_IN), .ZN(n2338) );
  INV_X1 U2781 ( .A(IR_REG_30__SCAN_IN), .ZN(n3476) );
  INV_X1 U2782 ( .A(n2397), .ZN(n4482) );
  INV_X1 U2783 ( .A(n3904), .ZN(n4484) );
  MUX2_X1 U2784 ( .A(IR_REG_31__SCAN_IN), .B(n2380), .S(IR_REG_25__SCAN_IN), 
        .Z(n2383) );
  INV_X1 U2785 ( .A(n2892), .ZN(n4486) );
  NAND2_X1 U2786 ( .A1(n3069), .A2(STATE_REG_SCAN_IN), .ZN(n4574) );
  INV_X1 U2787 ( .A(n3979), .ZN(n4490) );
  XNOR2_X1 U2788 ( .A(n2741), .B(IR_REG_18__SCAN_IN), .ZN(n4576) );
  AND2_X1 U2789 ( .A1(n2724), .A2(n2740), .ZN(n4491) );
  INV_X1 U2790 ( .A(n3096), .ZN(n2479) );
  XNOR2_X1 U2791 ( .A(n2473), .B(IR_REG_3__SCAN_IN), .ZN(n4500) );
  NAND2_X1 U2792 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2177)
         );
  OR3_X1 U2793 ( .A1(n3521), .A2(n3520), .A3(n3719), .ZN(n3525) );
  NAND2_X1 U2794 ( .A1(n2112), .A2(n2108), .ZN(U3258) );
  AOI21_X1 U2795 ( .B1(n2111), .B2(n2110), .A(n2109), .ZN(n2108) );
  INV_X1 U2796 ( .A(n4552), .ZN(n2112) );
  OAI21_X1 U2797 ( .B1(n4554), .B2(n4743), .A(n4553), .ZN(n2109) );
  NAND2_X1 U2798 ( .A1(n2068), .A2(n2067), .ZN(U3545) );
  NAND2_X1 U2799 ( .A1(n4334), .A2(REG1_REG_27__SCAN_IN), .ZN(n2067) );
  AND2_X1 U2800 ( .A1(n2074), .A2(n2073), .ZN(n2072) );
  NAND2_X1 U2801 ( .A1(n4334), .A2(REG1_REG_26__SCAN_IN), .ZN(n2073) );
  OR2_X1 U2802 ( .A1(n4434), .A2(n4419), .ZN(n2074) );
  OR2_X1 U2803 ( .A1(n4437), .A2(n4419), .ZN(n2081) );
  NAND2_X1 U2804 ( .A1(n2062), .A2(n2061), .ZN(n4358) );
  NAND2_X1 U2805 ( .A1(n4334), .A2(n4357), .ZN(n2061) );
  MUX2_X1 U2806 ( .A(n4361), .B(n4438), .S(n4416), .Z(n4362) );
  OAI21_X1 U2807 ( .B1(n4433), .B2(n4610), .A(n2066), .ZN(U3512) );
  AND2_X1 U2808 ( .A1(n2094), .A2(n2050), .ZN(n2066) );
  OR2_X1 U2809 ( .A1(n4434), .A2(n4480), .ZN(n2094) );
  AND2_X1 U2810 ( .A1(n2082), .A2(n2051), .ZN(n2075) );
  NAND2_X1 U2811 ( .A1(n2060), .A2(n4425), .ZN(n2059) );
  INV_X1 U2812 ( .A(n4440), .ZN(n2060) );
  NAND2_X1 U2813 ( .A1(n2208), .A2(REG1_REG_7__SCAN_IN), .ZN(n2006) );
  OR2_X1 U2814 ( .A1(n2031), .A2(n4498), .ZN(n2007) );
  AND2_X1 U2815 ( .A1(n2278), .A2(n2281), .ZN(n2008) );
  OR2_X1 U2816 ( .A1(n3640), .A2(n3564), .ZN(n2009) );
  INV_X1 U2817 ( .A(n2295), .ZN(n2294) );
  OAI21_X1 U2818 ( .B1(n2993), .B2(n2296), .A(n2033), .ZN(n2295) );
  INV_X1 U2819 ( .A(n3789), .ZN(n2233) );
  AND2_X1 U2820 ( .A1(n2308), .A2(n4298), .ZN(n2010) );
  AND2_X1 U2821 ( .A1(n2089), .A2(n3935), .ZN(n2011) );
  INV_X1 U2822 ( .A(n3144), .ZN(n2208) );
  AND2_X1 U2823 ( .A1(n2178), .A2(REG2_REG_10__SCAN_IN), .ZN(n2012) );
  INV_X1 U2824 ( .A(n4492), .ZN(n2212) );
  NAND2_X1 U2825 ( .A1(n2566), .A2(n2567), .ZN(n2013) );
  AND2_X1 U2826 ( .A1(n4229), .A2(n2992), .ZN(n2014) );
  NAND2_X1 U2827 ( .A1(n4196), .A2(n4181), .ZN(n4158) );
  AND2_X1 U2828 ( .A1(n3938), .A2(n2065), .ZN(n2015) );
  AND2_X1 U2829 ( .A1(n4284), .A2(n3022), .ZN(n2016) );
  OR2_X1 U2830 ( .A1(n2209), .A2(n2207), .ZN(n2017) );
  XOR2_X1 U2831 ( .A(n4065), .B(n4055), .Z(n2018) );
  AND2_X1 U2832 ( .A1(n2013), .A2(n2551), .ZN(n2019) );
  NOR2_X1 U2833 ( .A1(n4065), .A2(n3713), .ZN(n2020) );
  NAND2_X1 U2834 ( .A1(n2220), .A2(n2984), .ZN(n4282) );
  AND2_X1 U2835 ( .A1(n3894), .A2(n3632), .ZN(n2021) );
  AND2_X1 U2836 ( .A1(n2291), .A2(n2294), .ZN(n2022) );
  XNOR2_X1 U2837 ( .A(n2560), .B(IR_REG_8__SCAN_IN), .ZN(n4497) );
  INV_X1 U2838 ( .A(n3872), .ZN(n2272) );
  INV_X1 U2839 ( .A(n2715), .ZN(n2165) );
  OR2_X1 U2840 ( .A1(n4048), .A2(n4070), .ZN(n2023) );
  NOR2_X1 U2841 ( .A1(n3801), .A2(n2233), .ZN(n2232) );
  AND2_X1 U2842 ( .A1(n2299), .A2(n2351), .ZN(n2024) );
  OR2_X1 U2843 ( .A1(n2587), .A2(n3628), .ZN(n2025) );
  AND2_X1 U2844 ( .A1(n4048), .A2(n4070), .ZN(n2026) );
  INV_X1 U2845 ( .A(n2161), .ZN(n2159) );
  NOR2_X1 U2846 ( .A1(n2163), .A2(n3604), .ZN(n2161) );
  AND2_X1 U2847 ( .A1(n2269), .A2(n2270), .ZN(n2027) );
  AND2_X1 U2848 ( .A1(n3009), .A2(n3813), .ZN(n2028) );
  NAND2_X1 U2849 ( .A1(n2314), .A2(n2313), .ZN(n2029) );
  OR2_X1 U2850 ( .A1(n3041), .A2(n4037), .ZN(n2030) );
  AND2_X1 U2851 ( .A1(n2209), .A2(REG1_REG_6__SCAN_IN), .ZN(n2031) );
  AND2_X1 U2852 ( .A1(n4082), .A2(n4070), .ZN(n3748) );
  OR2_X1 U2853 ( .A1(n2385), .A2(IR_REG_24__SCAN_IN), .ZN(n2384) );
  OR2_X1 U2854 ( .A1(n4246), .A2(n3025), .ZN(n2032) );
  INV_X1 U2855 ( .A(n3564), .ZN(n2337) );
  AND2_X1 U2856 ( .A1(n2787), .A2(n2786), .ZN(n3564) );
  NAND2_X1 U2857 ( .A1(n2559), .A2(n2541), .ZN(n3144) );
  NOR2_X1 U2858 ( .A1(n4031), .A2(n2271), .ZN(n2269) );
  NAND2_X1 U2859 ( .A1(n4175), .A2(n2994), .ZN(n2033) );
  NOR2_X1 U2860 ( .A1(n4190), .A2(n4181), .ZN(n2034) );
  INV_X1 U2861 ( .A(n2282), .ZN(n2280) );
  NOR2_X1 U2862 ( .A1(n2020), .A2(n2283), .ZN(n2282) );
  NOR2_X1 U2863 ( .A1(n4151), .A2(n3547), .ZN(n2301) );
  AND2_X1 U2864 ( .A1(n2135), .A2(n2131), .ZN(n2035) );
  INV_X1 U2865 ( .A(n2127), .ZN(n2125) );
  NAND2_X1 U2866 ( .A1(n4499), .A2(REG2_REG_5__SCAN_IN), .ZN(n2127) );
  AND2_X1 U2867 ( .A1(n2588), .A2(n3488), .ZN(n2036) );
  OR2_X1 U2868 ( .A1(n2017), .A2(n2355), .ZN(n2037) );
  INV_X1 U2869 ( .A(n2987), .ZN(n4267) );
  AND2_X1 U2870 ( .A1(n2010), .A2(n4273), .ZN(n2038) );
  AND2_X1 U2871 ( .A1(n2189), .A2(n2188), .ZN(n2039) );
  AND2_X1 U2872 ( .A1(n2215), .A2(REG1_REG_10__SCAN_IN), .ZN(n2040) );
  NAND2_X1 U2873 ( .A1(n2510), .A2(REG1_REG_6__SCAN_IN), .ZN(n2041) );
  INV_X1 U2874 ( .A(IR_REG_5__SCAN_IN), .ZN(n2306) );
  OR2_X1 U2875 ( .A1(n4261), .A2(n3656), .ZN(n2042) );
  INV_X1 U2876 ( .A(n3002), .ZN(n2288) );
  INV_X1 U2877 ( .A(IR_REG_31__SCAN_IN), .ZN(n2167) );
  INV_X1 U2878 ( .A(IR_REG_31__SCAN_IN), .ZN(n2172) );
  NAND2_X2 U2879 ( .A1(n4313), .A2(n3254), .ZN(n4570) );
  INV_X1 U2880 ( .A(n4498), .ZN(n2209) );
  OR2_X1 U2881 ( .A1(n2089), .A2(n3935), .ZN(n2043) );
  OR2_X1 U2882 ( .A1(n3232), .A2(n3228), .ZN(n2044) );
  NOR2_X1 U2883 ( .A1(n3229), .A2(n3363), .ZN(n2045) );
  AND2_X1 U2884 ( .A1(n4312), .A2(n2038), .ZN(n4248) );
  XNOR2_X1 U2885 ( .A(n2635), .B(IR_REG_12__SCAN_IN), .ZN(n4493) );
  INV_X1 U2886 ( .A(n4493), .ZN(n2089) );
  NAND2_X1 U2887 ( .A1(n2383), .A2(n2388), .ZN(n2891) );
  NAND2_X1 U2888 ( .A1(n2322), .A2(n2465), .ZN(n3242) );
  AND2_X1 U2889 ( .A1(n2785), .A2(n2784), .ZN(n2046) );
  NOR2_X1 U2890 ( .A1(n4158), .A2(n4150), .ZN(n3055) );
  NAND2_X1 U2891 ( .A1(n4312), .A2(n2010), .ZN(n2309) );
  AND2_X1 U2892 ( .A1(n2045), .A2(n3236), .ZN(n2047) );
  INV_X1 U2893 ( .A(n2352), .ZN(n2302) );
  XNOR2_X1 U2894 ( .A(n2704), .B(n4753), .ZN(n4579) );
  NAND2_X1 U2895 ( .A1(n2954), .A2(n3211), .ZN(n3210) );
  AND3_X1 U2896 ( .A1(n3453), .A2(n2966), .A3(n3452), .ZN(n2048) );
  NAND2_X1 U2897 ( .A1(n4322), .A2(n4586), .ZN(n4411) );
  NAND2_X1 U2898 ( .A1(n3749), .A2(DATAI_27_), .ZN(n4037) );
  AND3_X1 U2899 ( .A1(n2203), .A2(n2206), .A3(n2202), .ZN(n2049) );
  OR2_X1 U2900 ( .A1(n4612), .A2(n4645), .ZN(n2050) );
  OR2_X1 U2901 ( .A1(n4612), .A2(n4436), .ZN(n2051) );
  OAI21_X1 U2902 ( .B1(n3132), .B2(n2125), .A(n4498), .ZN(n2126) );
  AND2_X1 U2903 ( .A1(n4582), .A2(REG1_REG_13__SCAN_IN), .ZN(n2052) );
  NAND2_X1 U2904 ( .A1(n3955), .A2(REG2_REG_15__SCAN_IN), .ZN(n2053) );
  AND2_X1 U2905 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2054) );
  OR2_X1 U2906 ( .A1(n2909), .A2(n2393), .ZN(n2055) );
  INV_X1 U2907 ( .A(n2320), .ZN(n2319) );
  NAND2_X1 U2908 ( .A1(n4105), .A2(n4125), .ZN(n2320) );
  OR2_X1 U2909 ( .A1(n4540), .A2(n2201), .ZN(n2056) );
  AND2_X1 U2910 ( .A1(n2113), .A2(n2126), .ZN(n2057) );
  INV_X1 U2911 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4634) );
  INV_X1 U2912 ( .A(n3236), .ZN(n4495) );
  AND2_X1 U2913 ( .A1(n2195), .A2(n3973), .ZN(n2194) );
  INV_X1 U2914 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2207) );
  INV_X1 U2915 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2226) );
  NAND2_X1 U2916 ( .A1(n2988), .A2(n2987), .ZN(n4258) );
  NOR2_X1 U2917 ( .A1(n2998), .A2(n2997), .ZN(n4114) );
  NOR2_X1 U2918 ( .A1(n2495), .A2(n2494), .ZN(n2497) );
  AOI21_X1 U2919 ( .B1(n4247), .B2(n2991), .A(n2990), .ZN(n4232) );
  NAND2_X2 U2920 ( .A1(n3825), .A2(n3828), .ZN(n3790) );
  NAND2_X1 U2921 ( .A1(n2955), .A2(n3203), .ZN(n3010) );
  NAND2_X1 U2922 ( .A1(n2307), .A2(n2500), .ZN(n2908) );
  NAND2_X2 U2923 ( .A1(n2063), .A2(n2520), .ZN(n3897) );
  NAND2_X1 U2924 ( .A1(n3372), .A2(n2255), .ZN(n2252) );
  NAND2_X1 U2925 ( .A1(n3443), .A2(n3777), .ZN(n3444) );
  XNOR2_X2 U2926 ( .A(n2395), .B(n3476), .ZN(n2397) );
  NAND2_X1 U2927 ( .A1(n4439), .A2(n2059), .ZN(U3510) );
  INV_X1 U2928 ( .A(n2979), .ZN(n2256) );
  NAND2_X1 U2929 ( .A1(n2255), .A2(n2021), .ZN(n2254) );
  OR2_X2 U2930 ( .A1(n4483), .A2(n2397), .ZN(n2451) );
  OR3_X1 U2931 ( .A1(n4345), .A2(n4344), .A3(n4604), .ZN(n4348) );
  NAND2_X1 U2932 ( .A1(n3425), .A2(n2983), .ZN(n2220) );
  NAND2_X1 U2933 ( .A1(n3444), .A2(n2965), .ZN(n3267) );
  NAND2_X1 U2934 ( .A1(n2220), .A2(n2219), .ZN(n2986) );
  NOR2_X1 U2935 ( .A1(n2397), .A2(n3091), .ZN(n2224) );
  NOR2_X2 U2936 ( .A1(n4519), .A2(n2101), .ZN(n3946) );
  AND2_X2 U2937 ( .A1(n2079), .A2(n2078), .ZN(n4519) );
  NAND3_X1 U2938 ( .A1(n3165), .A2(n3198), .A3(n2957), .ZN(n2963) );
  INV_X1 U2939 ( .A(n2273), .ZN(n3999) );
  OAI21_X1 U2940 ( .B1(n3267), .B2(n3269), .A(n2972), .ZN(n2975) );
  INV_X1 U2941 ( .A(IR_REG_2__SCAN_IN), .ZN(n2438) );
  NAND3_X1 U2942 ( .A1(n2252), .A2(n2253), .A3(n2981), .ZN(n4307) );
  NAND2_X1 U2943 ( .A1(n2287), .A2(n2023), .ZN(n2086) );
  NAND2_X1 U2944 ( .A1(n4114), .A2(n4115), .ZN(n4113) );
  NAND2_X1 U2945 ( .A1(n4432), .A2(n4416), .ZN(n2068) );
  NAND2_X1 U2946 ( .A1(n4351), .A2(n2069), .ZN(n4432) );
  OAI21_X1 U2947 ( .B1(n4078), .B2(n2280), .A(n2008), .ZN(n4029) );
  INV_X1 U2948 ( .A(n3445), .ZN(n3013) );
  NAND2_X1 U2949 ( .A1(n4147), .A2(n3743), .ZN(n2216) );
  NAND2_X2 U2950 ( .A1(n3036), .A2(n3800), .ZN(n4061) );
  NAND2_X2 U2951 ( .A1(n4317), .A2(n3843), .ZN(n3421) );
  NAND2_X1 U2952 ( .A1(n2986), .A2(n2985), .ZN(n4260) );
  OAI21_X1 U2953 ( .B1(n4433), .B2(n4334), .A(n2072), .ZN(U3544) );
  NAND2_X1 U2954 ( .A1(n2285), .A2(n2284), .ZN(n2287) );
  NAND2_X1 U2955 ( .A1(n2076), .A2(n2075), .ZN(U3511) );
  OR2_X1 U2956 ( .A1(n4435), .A2(n4610), .ZN(n2076) );
  XNOR2_X1 U2957 ( .A(n2077), .B(n4062), .ZN(n4356) );
  NAND2_X1 U2958 ( .A1(n2285), .A2(n2288), .ZN(n2077) );
  INV_X1 U2959 ( .A(n2079), .ZN(n4520) );
  NAND2_X1 U2960 ( .A1(n3945), .A2(n2211), .ZN(n2079) );
  NAND2_X1 U2961 ( .A1(n4358), .A2(n2081), .ZN(U3543) );
  AOI22_X2 U2962 ( .A1(n3104), .A2(REG1_REG_3__SCAN_IN), .B1(n3083), .B2(n4500), .ZN(n3084) );
  NAND2_X1 U2963 ( .A1(n3939), .A2(REG1_REG_14__SCAN_IN), .ZN(n3945) );
  NOR2_X1 U2964 ( .A1(n2015), .A2(n4505), .ZN(n4504) );
  NAND2_X1 U2965 ( .A1(n3948), .A2(n3949), .ZN(n3967) );
  AOI22_X2 U2966 ( .A1(n3922), .A2(REG1_REG_4__SCAN_IN), .B1(n2479), .B2(n3085), .ZN(n3131) );
  INV_X1 U2967 ( .A(n3398), .ZN(n2092) );
  XNOR2_X1 U2968 ( .A(n3946), .B(n2705), .ZN(n4533) );
  NOR2_X1 U2969 ( .A1(n4130), .A2(n2083), .ZN(n2998) );
  NAND2_X1 U2970 ( .A1(n4258), .A2(n2989), .ZN(n4247) );
  NAND3_X1 U2971 ( .A1(n2203), .A2(n2202), .A3(n2088), .ZN(n2087) );
  NOR2_X1 U2972 ( .A1(n4550), .A2(n2102), .ZN(n3969) );
  XNOR2_X1 U2973 ( .A(n3082), .B(n4500), .ZN(n3104) );
  NOR2_X1 U2974 ( .A1(n4545), .A2(n4544), .ZN(n4550) );
  NOR2_X2 U2975 ( .A1(n3131), .A2(n3130), .ZN(n3129) );
  OR2_X2 U2976 ( .A1(n3129), .A2(n2037), .ZN(n2203) );
  NAND2_X1 U2977 ( .A1(n3010), .A2(n3816), .ZN(n3198) );
  NAND2_X1 U2978 ( .A1(n2307), .A2(n2304), .ZN(n2385) );
  NAND2_X1 U2979 ( .A1(n2513), .A2(REG3_REG_6__SCAN_IN), .ZN(n2532) );
  INV_X2 U2980 ( .A(n4050), .ZN(n3041) );
  NOR2_X2 U2981 ( .A1(n2818), .A2(n3619), .ZN(n2097) );
  NAND2_X1 U2982 ( .A1(n3129), .A2(n2007), .ZN(n2202) );
  MUX2_X1 U2983 ( .A(n3091), .B(REG2_REG_1__SCAN_IN), .S(n4503), .Z(n3438) );
  AOI21_X1 U2984 ( .B1(n2115), .B2(n2126), .A(n3115), .ZN(n2114) );
  INV_X1 U2985 ( .A(n2120), .ZN(n2115) );
  NAND2_X1 U2986 ( .A1(n2126), .A2(n2118), .ZN(n2116) );
  INV_X1 U2987 ( .A(n2118), .ZN(n2117) );
  OAI21_X1 U2988 ( .B1(n2122), .B2(n3132), .A(REG2_REG_6__SCAN_IN), .ZN(n2118)
         );
  OAI211_X1 U2989 ( .C1(n3132), .C2(n2124), .A(n2123), .B(n2119), .ZN(n3114)
         );
  NAND2_X1 U2990 ( .A1(n3132), .A2(n2209), .ZN(n2119) );
  NAND2_X1 U2991 ( .A1(n3132), .A2(n2121), .ZN(n2120) );
  NAND2_X1 U2992 ( .A1(n2125), .A2(n2209), .ZN(n2123) );
  NAND3_X1 U2993 ( .A1(n2137), .A2(n2138), .A3(n4495), .ZN(n2129) );
  NAND2_X1 U2994 ( .A1(n3152), .A2(n4497), .ZN(n2140) );
  NAND3_X1 U2995 ( .A1(n2528), .A2(n2527), .A3(n2148), .ZN(n2146) );
  NAND2_X1 U2996 ( .A1(n2528), .A2(n2527), .ZN(n3489) );
  NAND2_X1 U2997 ( .A1(n2668), .A2(n2170), .ZN(n2168) );
  NAND2_X1 U2998 ( .A1(n2668), .A2(n2173), .ZN(n2169) );
  INV_X1 U2999 ( .A(n2456), .ZN(n2175) );
  NAND2_X2 U3000 ( .A1(n2408), .A2(n2176), .ZN(n2875) );
  INV_X2 U3001 ( .A(n2875), .ZN(n2767) );
  XNOR2_X2 U3002 ( .A(IR_REG_1__SCAN_IN), .B(n2177), .ZN(n4503) );
  INV_X1 U3003 ( .A(n2181), .ZN(n3396) );
  INV_X1 U3004 ( .A(n2189), .ZN(n3954) );
  INV_X1 U3005 ( .A(n3953), .ZN(n2188) );
  INV_X1 U3006 ( .A(n3959), .ZN(n2191) );
  NAND2_X1 U3007 ( .A1(n3959), .A2(n3960), .ZN(n3974) );
  AND2_X1 U3008 ( .A1(n4576), .A2(REG2_REG_18__SCAN_IN), .ZN(n2196) );
  BUF_X1 U3009 ( .A(n4503), .Z(n2198) );
  NAND2_X1 U3010 ( .A1(n2457), .A2(n2371), .ZN(n2200) );
  NAND3_X1 U3011 ( .A1(n3442), .A2(n3441), .A3(n2056), .ZN(U3241) );
  INV_X1 U3012 ( .A(n3129), .ZN(n2205) );
  XNOR2_X1 U3013 ( .A(n2210), .B(n2209), .ZN(n3112) );
  NAND2_X1 U3014 ( .A1(n3235), .A2(n2040), .ZN(n2214) );
  NAND2_X1 U3015 ( .A1(n2214), .A2(n2213), .ZN(n3398) );
  NAND2_X2 U3016 ( .A1(n2216), .A2(n3859), .ZN(n4131) );
  OR2_X2 U3017 ( .A1(n4206), .A2(n3855), .ZN(n4147) );
  NAND2_X1 U3018 ( .A1(n3405), .A2(n3842), .ZN(n2217) );
  NAND2_X1 U3019 ( .A1(n3019), .A2(n3018), .ZN(n2218) );
  XNOR2_X2 U3020 ( .A(n2396), .B(IR_REG_29__SCAN_IN), .ZN(n4483) );
  NAND3_X1 U3021 ( .A1(n2398), .A2(n2397), .A3(REG0_REG_1__SCAN_IN), .ZN(n2222) );
  NAND3_X1 U3022 ( .A1(n4482), .A2(n4483), .A3(REG3_REG_1__SCAN_IN), .ZN(n2225) );
  OAI211_X1 U3023 ( .C1(n2230), .C2(n2228), .A(n3782), .B(n2227), .ZN(n3012)
         );
  INV_X1 U3024 ( .A(n3813), .ZN(n2228) );
  NAND2_X1 U3025 ( .A1(n3200), .A2(n3813), .ZN(n3283) );
  NAND2_X1 U3026 ( .A1(n2230), .A2(n2229), .ZN(n3200) );
  OAI21_X1 U3027 ( .B1(n3778), .B2(n3809), .A(n3009), .ZN(n3201) );
  NAND2_X1 U3028 ( .A1(n3009), .A2(n3809), .ZN(n2231) );
  NAND2_X1 U3029 ( .A1(n2234), .A2(n2232), .ZN(n3036) );
  NAND2_X1 U3030 ( .A1(n3034), .A2(n3746), .ZN(n2234) );
  OAI21_X1 U3031 ( .B1(n3015), .B2(n2240), .A(n2238), .ZN(n3356) );
  NAND2_X1 U3032 ( .A1(n2237), .A2(n2235), .ZN(n3017) );
  AOI21_X1 U3033 ( .B1(n2238), .B2(n2240), .A(n2236), .ZN(n2235) );
  NAND2_X1 U3034 ( .A1(n3015), .A2(n2238), .ZN(n2237) );
  NAND2_X1 U3035 ( .A1(n3013), .A2(n2248), .ZN(n2244) );
  OR2_X1 U3036 ( .A1(n4321), .A2(n3021), .ZN(n2257) );
  NAND2_X1 U3037 ( .A1(n3421), .A2(n2262), .ZN(n2260) );
  NAND2_X1 U3038 ( .A1(n4061), .A2(n2272), .ZN(n2270) );
  NAND2_X1 U3039 ( .A1(n4078), .A2(n3003), .ZN(n2285) );
  OAI21_X2 U3040 ( .B1(n4078), .B2(n2277), .A(n2274), .ZN(n2273) );
  NAND2_X1 U3041 ( .A1(n2014), .A2(n2292), .ZN(n2289) );
  NAND2_X1 U3042 ( .A1(n2289), .A2(n2290), .ZN(n4145) );
  MUX2_X1 U3043 ( .A(n4627), .B(n2303), .S(n2457), .Z(n3224) );
  INV_X1 U3044 ( .A(n2309), .ZN(n4297) );
  NAND2_X1 U3045 ( .A1(n4053), .A2(n2310), .ZN(n2314) );
  INV_X1 U3046 ( .A(n2314), .ZN(n4020) );
  NAND2_X1 U3047 ( .A1(n4021), .A2(n4022), .ZN(n2313) );
  NAND2_X1 U3048 ( .A1(n2956), .A2(n3204), .ZN(n3197) );
  NAND3_X1 U3049 ( .A1(n2322), .A2(n2465), .A3(n2321), .ZN(n3244) );
  OAI21_X2 U3050 ( .B1(n3527), .B2(n2324), .A(n2323), .ZN(n3579) );
  OAI21_X2 U3051 ( .B1(n3639), .B2(n2009), .A(n2335), .ZN(n3663) );
  NAND2_X1 U3052 ( .A1(n2339), .A2(n2338), .ZN(n3475) );
  INV_X1 U3053 ( .A(n2908), .ZN(n2339) );
  OAI22_X2 U3054 ( .A1(n3654), .A2(n2342), .B1(n3652), .B2(n2343), .ZN(n3509)
         );
  OAI21_X1 U3055 ( .B1(n4551), .B2(n4550), .A(n4549), .ZN(n4552) );
  CLKBUF_X1 U3056 ( .A(n4229), .Z(n4230) );
  NAND2_X1 U3057 ( .A1(n2369), .A2(n2368), .ZN(n2370) );
  OR2_X1 U3058 ( .A1(n3088), .A2(n2367), .ZN(n2368) );
  INV_X1 U3059 ( .A(n3155), .ZN(n3157) );
  NAND2_X1 U3060 ( .A1(n4248), .A2(n4249), .ZN(n4251) );
  NAND2_X1 U3061 ( .A1(n4545), .A2(n4544), .ZN(n4547) );
  INV_X1 U3062 ( .A(n3224), .ZN(n3008) );
  NAND2_X1 U3063 ( .A1(n4020), .A2(n3991), .ZN(n3990) );
  OAI21_X1 U3064 ( .B1(n2029), .B2(n4366), .A(n2348), .ZN(n4341) );
  MUX2_X1 U3065 ( .A(n4500), .B(DATAI_3_), .S(n2457), .Z(n3288) );
  INV_X2 U3066 ( .A(n4610), .ZN(n4612) );
  INV_X1 U3067 ( .A(n4619), .ZN(n4334) );
  OR2_X1 U3068 ( .A1(n4612), .A2(REG0_REG_28__SCAN_IN), .ZN(n2344) );
  OR2_X1 U3069 ( .A1(n3232), .A2(n3231), .ZN(n2346) );
  AND2_X1 U3070 ( .A1(n3890), .A2(n3035), .ZN(n2347) );
  OR3_X1 U3071 ( .A1(n4343), .A2(n4344), .A3(n4604), .ZN(n2348) );
  OR2_X1 U3072 ( .A1(n3480), .A2(n4480), .ZN(n2349) );
  OR2_X1 U3073 ( .A1(n3480), .A2(n4419), .ZN(n2350) );
  NAND2_X1 U3074 ( .A1(n4224), .A2(n4214), .ZN(n2351) );
  NOR2_X1 U3075 ( .A1(n4224), .A2(n4214), .ZN(n2352) );
  INV_X1 U3076 ( .A(n3891), .ZN(n4133) );
  NAND2_X1 U3077 ( .A1(n2394), .A2(IR_REG_27__SCAN_IN), .ZN(n2354) );
  INV_X1 U3078 ( .A(n3898), .ZN(n2967) );
  AND2_X1 U3079 ( .A1(n4499), .A2(REG1_REG_5__SCAN_IN), .ZN(n2355) );
  OR3_X1 U3080 ( .A1(n3541), .A2(n3539), .A3(n3684), .ZN(n2356) );
  INV_X1 U3081 ( .A(IR_REG_22__SCAN_IN), .ZN(n2363) );
  AND2_X1 U3082 ( .A1(n4098), .A2(n4096), .ZN(n3863) );
  AND2_X1 U3083 ( .A1(n3268), .A2(n2969), .ZN(n2971) );
  INV_X1 U3084 ( .A(n4316), .ZN(n2981) );
  AND2_X1 U3085 ( .A1(n2971), .A2(n3790), .ZN(n2972) );
  OR2_X1 U3086 ( .A1(n2713), .A2(n2712), .ZN(n2711) );
  INV_X1 U3087 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U3088 ( .A1(n2510), .A2(REG1_REG_0__SCAN_IN), .ZN(n2414) );
  INV_X1 U3089 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3971) );
  INV_X1 U3090 ( .A(n3557), .ZN(n3054) );
  INV_X1 U3091 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2659) );
  AND2_X1 U3092 ( .A1(n2707), .A2(n2708), .ZN(n3508) );
  AND2_X1 U3093 ( .A1(n2754), .A2(n2753), .ZN(n3541) );
  INV_X1 U3094 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2677) );
  AND2_X1 U3095 ( .A1(n3518), .A2(n3519), .ZN(n2814) );
  OR2_X1 U3096 ( .A1(n2837), .A2(n2926), .ZN(n2934) );
  OR2_X1 U3097 ( .A1(n3482), .A2(n2802), .ZN(n2884) );
  INV_X1 U3098 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4719) );
  OR2_X1 U3099 ( .A1(n4019), .A2(n2802), .ZN(n2941) );
  NAND2_X1 U3100 ( .A1(n3891), .A2(n2999), .ZN(n3000) );
  AND2_X1 U3101 ( .A1(n3071), .A2(n3754), .ZN(n3086) );
  NAND2_X1 U3102 ( .A1(n2943), .A2(n2935), .ZN(n3689) );
  CLKBUF_X2 U3103 ( .A(n2451), .Z(n2680) );
  AND2_X1 U3104 ( .A1(n3097), .A2(n2479), .ZN(n3098) );
  AND2_X1 U3105 ( .A1(n3324), .A2(n4495), .ZN(n3325) );
  NAND2_X1 U3106 ( .A1(n3087), .A2(n3086), .ZN(n3125) );
  INV_X1 U3107 ( .A(n4488), .ZN(n3807) );
  AND2_X1 U3108 ( .A1(n3754), .A2(DATAI_26_), .ZN(n3713) );
  INV_X1 U3109 ( .A(n3729), .ZN(n4249) );
  INV_X1 U3110 ( .A(n4595), .ZN(n4586) );
  OR2_X1 U3111 ( .A1(n3177), .A2(n3884), .ZN(n3087) );
  AND2_X1 U3112 ( .A1(n2830), .A2(n2819), .ZN(n4089) );
  NAND2_X1 U3113 ( .A1(n2929), .A2(n3176), .ZN(n3733) );
  NOR2_X1 U3114 ( .A1(n3125), .A2(n4484), .ZN(n4548) );
  AOI21_X1 U3115 ( .B1(n4774), .B2(n4293), .A(n3042), .ZN(n3043) );
  INV_X1 U3116 ( .A(n4330), .ZN(n4268) );
  INV_X1 U3117 ( .A(n4315), .ZN(n4557) );
  NAND2_X1 U3118 ( .A1(n4334), .A2(n3051), .ZN(n3052) );
  OAI22_X1 U3119 ( .A1(n3064), .A2(D_REG_0__SCAN_IN), .B1(n4486), .B2(n2894), 
        .ZN(n3251) );
  INV_X1 U3120 ( .A(n3621), .ZN(n4087) );
  INV_X1 U3121 ( .A(n4366), .ZN(n4602) );
  AND2_X1 U3122 ( .A1(n2421), .A2(n3067), .ZN(n3177) );
  AND2_X1 U3123 ( .A1(n3087), .A2(n3072), .ZN(n4527) );
  INV_X1 U3124 ( .A(n3733), .ZN(n3695) );
  NAND2_X1 U3125 ( .A1(n2763), .A2(n2762), .ZN(n4177) );
  INV_X1 U3126 ( .A(n4537), .ZN(n4541) );
  INV_X1 U3127 ( .A(n4535), .ZN(n4546) );
  INV_X1 U3128 ( .A(n4570), .ZN(n4280) );
  INV_X1 U3129 ( .A(n4570), .ZN(n4276) );
  INV_X1 U3130 ( .A(n4568), .ZN(n4306) );
  INV_X2 U3131 ( .A(n4334), .ZN(n4416) );
  NOR2_X1 U3132 ( .A1(n3059), .A2(n3251), .ZN(n4619) );
  NAND2_X1 U3133 ( .A1(n4612), .A2(n4602), .ZN(n4480) );
  OR2_X1 U3134 ( .A1(n3059), .A2(n3058), .ZN(n4610) );
  INV_X1 U3135 ( .A(n4574), .ZN(n3067) );
  INV_X1 U3136 ( .A(n3907), .ZN(U4043) );
  INV_X2 U3137 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3138 ( .A(DATAI_1_), .ZN(n2371) );
  NOR2_X2 U3139 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2720)
         );
  NAND2_X1 U3140 ( .A1(n2437), .A2(n2438), .ZN(n2456) );
  NAND3_X1 U3141 ( .A1(n2381), .A2(n4693), .A3(n2391), .ZN(n2366) );
  OAI21_X2 U3142 ( .B1(n2385), .B2(n2366), .A(IR_REG_31__SCAN_IN), .ZN(n3088)
         );
  NAND2_X1 U3143 ( .A1(n3088), .A2(n2394), .ZN(n2369) );
  NAND2_X2 U3144 ( .A1(n2370), .A2(n2354), .ZN(n2457) );
  NOR2_X1 U3146 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2373)
         );
  NAND2_X1 U3147 ( .A1(n2668), .A2(n2004), .ZN(n2378) );
  NAND2_X1 U31480 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2377) );
  MUX2_X1 U31490 ( .A(IR_REG_31__SCAN_IN), .B(n2377), .S(IR_REG_21__SCAN_IN), 
        .Z(n2379) );
  NAND2_X1 U3150 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3151 ( .A1(n2385), .A2(IR_REG_31__SCAN_IN), .ZN(n2386) );
  MUX2_X1 U3152 ( .A(IR_REG_31__SCAN_IN), .B(n2386), .S(IR_REG_24__SCAN_IN), 
        .Z(n2387) );
  NOR2_X1 U3153 ( .A1(n2891), .A2(n2892), .ZN(n2390) );
  XNOR2_X2 U3154 ( .A(n2389), .B(IR_REG_26__SCAN_IN), .ZN(n2894) );
  NAND2_X2 U3155 ( .A1(n2390), .A2(n2894), .ZN(n2421) );
  NAND2_X1 U3156 ( .A1(n2956), .A2(n2858), .ZN(n2401) );
  NOR2_X1 U3157 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2392)
         );
  NAND4_X1 U3158 ( .A1(n2392), .A2(n4693), .A3(n2910), .A4(n2391), .ZN(n2393)
         );
  NAND2_X1 U3159 ( .A1(n2510), .A2(REG1_REG_1__SCAN_IN), .ZN(n2399) );
  INV_X1 U3160 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3091) );
  INV_X1 U3161 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3256) );
  NAND2_X1 U3162 ( .A1(n2058), .A2(n2767), .ZN(n2400) );
  NAND2_X1 U3163 ( .A1(n2401), .A2(n2400), .ZN(n2407) );
  NAND2_X1 U3164 ( .A1(n3979), .A2(n4487), .ZN(n2925) );
  NAND2_X4 U3165 ( .A1(n2402), .A2(n2925), .ZN(n2886) );
  INV_X1 U3166 ( .A(n3149), .ZN(n2409) );
  AND2_X2 U3167 ( .A1(n2858), .A2(n4366), .ZN(n2461) );
  NAND2_X1 U3168 ( .A1(n2005), .A2(n2058), .ZN(n2411) );
  NAND2_X1 U3169 ( .A1(n2956), .A2(n2767), .ZN(n2410) );
  NAND2_X1 U3170 ( .A1(n2411), .A2(n2410), .ZN(n2428) );
  XNOR2_X1 U3171 ( .A(n2429), .B(n2428), .ZN(n3183) );
  INV_X1 U3172 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2412) );
  INV_X1 U3173 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2413) );
  OR2_X1 U3174 ( .A1(n2451), .A2(n2413), .ZN(n2415) );
  INV_X1 U3175 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U3176 ( .A1(n2064), .A2(n2767), .ZN(n2420) );
  NAND2_X1 U3177 ( .A1(n3008), .A2(n2858), .ZN(n2419) );
  NAND2_X1 U3178 ( .A1(n2420), .A2(n2419), .ZN(n2426) );
  INV_X1 U3179 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U3180 ( .A1(n2421), .A2(n4638), .ZN(n2422) );
  NAND2_X1 U3181 ( .A1(n2005), .A2(n2064), .ZN(n2425) );
  INV_X1 U3182 ( .A(IR_REG_0__SCAN_IN), .ZN(n4627) );
  NOR2_X1 U3183 ( .A1(n2421), .A2(n4627), .ZN(n2423) );
  AOI21_X1 U3184 ( .B1(n2839), .B2(n3008), .A(n2423), .ZN(n2424) );
  NAND2_X1 U3185 ( .A1(n2425), .A2(n2424), .ZN(n3220) );
  INV_X1 U3186 ( .A(n2426), .ZN(n2427) );
  AOI22_X1 U3187 ( .A1(n3221), .A2(n3220), .B1(n2427), .B2(n2861), .ZN(n3184)
         );
  NAND2_X1 U3188 ( .A1(n2429), .A2(n2428), .ZN(n2430) );
  AND2_X2 U3189 ( .A1(n3185), .A2(n2430), .ZN(n3190) );
  NAND2_X1 U3190 ( .A1(n2510), .A2(REG1_REG_2__SCAN_IN), .ZN(n2433) );
  INV_X1 U3191 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3196) );
  INV_X1 U3192 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3090) );
  OR2_X1 U3193 ( .A1(n2451), .A2(n3090), .ZN(n2431) );
  INV_X1 U3194 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2434) );
  OR2_X1 U3195 ( .A1(n2490), .A2(n2434), .ZN(n2435) );
  NAND2_X1 U3196 ( .A1(n2436), .A2(n2767), .ZN(n2442) );
  XNOR2_X2 U3197 ( .A(n2439), .B(n2438), .ZN(n3912) );
  INV_X1 U3198 ( .A(DATAI_2_), .ZN(n2440) );
  MUX2_X1 U3199 ( .A(n2103), .B(n2440), .S(n2457), .Z(n2954) );
  NAND2_X1 U3200 ( .A1(n3203), .A2(n2858), .ZN(n2441) );
  NAND2_X1 U3201 ( .A1(n2442), .A2(n2441), .ZN(n2443) );
  XNOR2_X1 U3202 ( .A(n2443), .B(n2861), .ZN(n2448) );
  NAND2_X1 U3203 ( .A1(n2461), .A2(n2436), .ZN(n2445) );
  NAND2_X1 U3204 ( .A1(n3203), .A2(n2839), .ZN(n2444) );
  NAND2_X1 U3205 ( .A1(n2445), .A2(n2444), .ZN(n2446) );
  XNOR2_X1 U3206 ( .A(n2448), .B(n2446), .ZN(n3191) );
  INV_X1 U3207 ( .A(n2446), .ZN(n2447) );
  NAND2_X1 U3208 ( .A1(n2448), .A2(n2447), .ZN(n2449) );
  NAND2_X1 U3209 ( .A1(n2510), .A2(REG1_REG_3__SCAN_IN), .ZN(n2455) );
  INV_X1 U32100 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2450) );
  OR2_X1 U32110 ( .A1(n2512), .A2(REG3_REG_3__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U32120 ( .A1(n3900), .A2(n2839), .ZN(n2459) );
  NAND2_X1 U32130 ( .A1(n2456), .A2(IR_REG_31__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U32140 ( .A1(n3288), .A2(n2858), .ZN(n2458) );
  NAND2_X1 U32150 ( .A1(n2459), .A2(n2458), .ZN(n2460) );
  XNOR2_X1 U32160 ( .A(n2460), .B(n2886), .ZN(n2462) );
  AOI22_X1 U32170 ( .A1(n2461), .A2(n3900), .B1(n2839), .B2(n3288), .ZN(n2463)
         );
  XNOR2_X1 U32180 ( .A(n2462), .B(n2463), .ZN(n3214) );
  INV_X1 U32190 ( .A(n2462), .ZN(n2464) );
  NAND2_X1 U32200 ( .A1(n2464), .A2(n2463), .ZN(n2465) );
  NAND2_X1 U32210 ( .A1(n2510), .A2(REG1_REG_4__SCAN_IN), .ZN(n2471) );
  INV_X1 U32220 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2466) );
  OR2_X1 U32230 ( .A1(n2490), .A2(n2466), .ZN(n2470) );
  OAI21_X1 U32240 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2488), .ZN(n3454) );
  OR2_X1 U32250 ( .A1(n2512), .A2(n3454), .ZN(n2469) );
  INV_X1 U32260 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3927) );
  OR2_X1 U32270 ( .A1(n2451), .A2(n3927), .ZN(n2468) );
  NAND2_X1 U32280 ( .A1(n3899), .A2(n2839), .ZN(n2481) );
  INV_X4 U32290 ( .A(n2636), .ZN(n3749) );
  NAND2_X1 U32300 ( .A1(n2473), .A2(n2472), .ZN(n2474) );
  NAND2_X1 U32310 ( .A1(n2474), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  XNOR2_X1 U32320 ( .A(n2476), .B(n2475), .ZN(n3096) );
  INV_X1 U32330 ( .A(DATAI_4_), .ZN(n2477) );
  NAND2_X1 U32340 ( .A1(n2457), .A2(n2477), .ZN(n2478) );
  OAI21_X2 U32350 ( .B1(n3749), .B2(n2479), .A(n2478), .ZN(n3452) );
  NAND2_X1 U32360 ( .A1(n2317), .A2(n2858), .ZN(n2480) );
  NAND2_X1 U32370 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  XNOR2_X1 U32380 ( .A(n2482), .B(n2886), .ZN(n2486) );
  NAND2_X1 U32390 ( .A1(n2461), .A2(n3899), .ZN(n2484) );
  NAND2_X1 U32400 ( .A1(n2317), .A2(n2839), .ZN(n2483) );
  NAND2_X1 U32410 ( .A1(n2484), .A2(n2483), .ZN(n2485) );
  XNOR2_X1 U32420 ( .A(n2486), .B(n2485), .ZN(n3243) );
  NAND2_X1 U32430 ( .A1(n2486), .A2(n2485), .ZN(n2487) );
  NAND2_X1 U32440 ( .A1(n3244), .A2(n2487), .ZN(n3317) );
  INV_X1 U32450 ( .A(n2513), .ZN(n2515) );
  NAND2_X1 U32460 ( .A1(n2488), .A2(n4634), .ZN(n2489) );
  NAND2_X1 U32470 ( .A1(n2515), .A2(n2489), .ZN(n3323) );
  NAND2_X1 U32480 ( .A1(n2529), .A2(REG0_REG_5__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U32490 ( .A1(n2492), .A2(n2491), .ZN(n2495) );
  INV_X1 U32500 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2493) );
  INV_X1 U32510 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3298) );
  NAND2_X2 U32520 ( .A1(n2497), .A2(n2496), .ZN(n3898) );
  NAND2_X1 U32530 ( .A1(n3898), .A2(n2839), .ZN(n2504) );
  NAND2_X1 U32540 ( .A1(n2498), .A2(IR_REG_31__SCAN_IN), .ZN(n2499) );
  MUX2_X1 U32550 ( .A(IR_REG_31__SCAN_IN), .B(n2499), .S(IR_REG_5__SCAN_IN), 
        .Z(n2502) );
  INV_X1 U32560 ( .A(n2500), .ZN(n2501) );
  AND2_X1 U32570 ( .A1(n2502), .A2(n2501), .ZN(n4499) );
  MUX2_X1 U32580 ( .A(n4499), .B(DATAI_5_), .S(n3749), .Z(n3299) );
  NAND2_X1 U32590 ( .A1(n3299), .A2(n2858), .ZN(n2503) );
  NAND2_X1 U32600 ( .A1(n2504), .A2(n2503), .ZN(n2505) );
  XNOR2_X1 U32610 ( .A(n2505), .B(n2886), .ZN(n2506) );
  AOI22_X1 U32620 ( .A1(n2461), .A2(n3898), .B1(n2767), .B2(n3299), .ZN(n2507)
         );
  XNOR2_X1 U32630 ( .A(n2506), .B(n2507), .ZN(n3316) );
  NAND2_X1 U32640 ( .A1(n3317), .A2(n3316), .ZN(n3315) );
  INV_X1 U32650 ( .A(n2506), .ZN(n2508) );
  OR2_X1 U32660 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  NAND2_X1 U32670 ( .A1(n3315), .A2(n2509), .ZN(n3699) );
  INV_X1 U32680 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2511) );
  INV_X1 U32690 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U32700 ( .A1(n2515), .A2(n2514), .ZN(n2516) );
  NAND2_X1 U32710 ( .A1(n2532), .A2(n2516), .ZN(n3274) );
  OR2_X1 U32720 ( .A1(n2570), .A2(n3274), .ZN(n2519) );
  INV_X1 U32730 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2517) );
  OR2_X1 U32740 ( .A1(n2451), .A2(n2517), .ZN(n2518) );
  NAND2_X1 U32750 ( .A1(n2461), .A2(n3897), .ZN(n2523) );
  OR2_X1 U32760 ( .A1(n2500), .A2(n2167), .ZN(n2521) );
  MUX2_X1 U32770 ( .A(n4498), .B(DATAI_6_), .S(n3749), .Z(n3702) );
  NAND2_X1 U32780 ( .A1(n2839), .A2(n3702), .ZN(n2522) );
  NAND2_X1 U32790 ( .A1(n2523), .A2(n2522), .ZN(n3696) );
  NAND2_X1 U32800 ( .A1(n3897), .A2(n2839), .ZN(n2525) );
  NAND2_X1 U32810 ( .A1(n3702), .A2(n2858), .ZN(n2524) );
  NAND2_X1 U32820 ( .A1(n2525), .A2(n2524), .ZN(n2526) );
  XNOR2_X1 U32830 ( .A(n2526), .B(n2886), .ZN(n3697) );
  OAI21_X1 U32840 ( .B1(n3699), .B2(n3696), .A(n3697), .ZN(n2528) );
  NAND2_X1 U32850 ( .A1(n3699), .A2(n3696), .ZN(n2527) );
  NAND2_X1 U32860 ( .A1(n2529), .A2(REG0_REG_7__SCAN_IN), .ZN(n2538) );
  INV_X1 U32870 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2530) );
  OR2_X1 U32880 ( .A1(n2805), .A2(n2530), .ZN(n2537) );
  NAND2_X1 U32890 ( .A1(n2532), .A2(n2531), .ZN(n2533) );
  NAND2_X1 U32900 ( .A1(n2553), .A2(n2533), .ZN(n3493) );
  INV_X1 U32910 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U32920 ( .A1(n3896), .A2(n2839), .ZN(n2544) );
  NAND2_X1 U32930 ( .A1(n2500), .A2(n4635), .ZN(n2578) );
  NAND2_X1 U32940 ( .A1(n2578), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  INV_X1 U32950 ( .A(n4669), .ZN(n2539) );
  NAND2_X1 U32960 ( .A1(n2540), .A2(n2539), .ZN(n2559) );
  OR2_X1 U32970 ( .A1(n2540), .A2(n2539), .ZN(n2541) );
  INV_X1 U32980 ( .A(DATAI_7_), .ZN(n2542) );
  MUX2_X1 U32990 ( .A(n3144), .B(n2542), .S(n3749), .Z(n2970) );
  NAND2_X1 U33000 ( .A1(n3492), .A2(n2858), .ZN(n2543) );
  NAND2_X1 U33010 ( .A1(n2544), .A2(n2543), .ZN(n2545) );
  XNOR2_X1 U33020 ( .A(n2545), .B(n2861), .ZN(n2548) );
  NAND2_X1 U33030 ( .A1(n2461), .A2(n3896), .ZN(n2547) );
  NAND2_X1 U33040 ( .A1(n3492), .A2(n2839), .ZN(n2546) );
  NAND2_X1 U33050 ( .A1(n2547), .A2(n2546), .ZN(n2549) );
  XNOR2_X1 U33060 ( .A(n2548), .B(n2549), .ZN(n3488) );
  INV_X1 U33070 ( .A(n2548), .ZN(n2550) );
  NAND2_X1 U33080 ( .A1(n2550), .A2(n2549), .ZN(n2551) );
  NAND2_X1 U33090 ( .A1(n2936), .A2(REG0_REG_8__SCAN_IN), .ZN(n2558) );
  INV_X1 U33100 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4716) );
  OR2_X1 U33110 ( .A1(n2805), .A2(n4716), .ZN(n2557) );
  NAND2_X1 U33120 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  NAND2_X1 U33130 ( .A1(n2572), .A2(n2554), .ZN(n3558) );
  OR2_X1 U33140 ( .A1(n2802), .A2(n3558), .ZN(n2556) );
  INV_X1 U33150 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3363) );
  OR2_X1 U33160 ( .A1(n2680), .A2(n3363), .ZN(n2555) );
  NAND4_X1 U33170 ( .A1(n2558), .A2(n2557), .A3(n2556), .A4(n2555), .ZN(n3895)
         );
  NAND2_X1 U33180 ( .A1(n3895), .A2(n2839), .ZN(n2562) );
  NAND2_X1 U33190 ( .A1(n2559), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  MUX2_X1 U33200 ( .A(n4497), .B(DATAI_8_), .S(n3749), .Z(n3557) );
  NAND2_X1 U33210 ( .A1(n3557), .A2(n2858), .ZN(n2561) );
  NAND2_X1 U33220 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  XNOR2_X1 U33230 ( .A(n2563), .B(n2886), .ZN(n2566) );
  NAND2_X1 U33240 ( .A1(n2461), .A2(n3895), .ZN(n2565) );
  NAND2_X1 U33250 ( .A1(n2767), .A2(n3557), .ZN(n2564) );
  NAND2_X1 U33260 ( .A1(n2565), .A2(n2564), .ZN(n2567) );
  INV_X1 U33270 ( .A(n2566), .ZN(n2569) );
  INV_X1 U33280 ( .A(n2567), .ZN(n2568) );
  NAND2_X1 U33290 ( .A1(n2569), .A2(n2568), .ZN(n3626) );
  NAND2_X1 U33300 ( .A1(n3750), .A2(REG1_REG_9__SCAN_IN), .ZN(n2577) );
  INV_X1 U33310 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4668) );
  OR2_X1 U33320 ( .A1(n3751), .A2(n4668), .ZN(n2576) );
  NAND2_X1 U33330 ( .A1(n2572), .A2(n2571), .ZN(n2573) );
  NAND2_X1 U33340 ( .A1(n2591), .A2(n2573), .ZN(n3376) );
  OR2_X1 U33350 ( .A1(n2802), .A2(n3376), .ZN(n2575) );
  INV_X1 U33360 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3228) );
  OR2_X1 U33370 ( .A1(n2680), .A2(n3228), .ZN(n2574) );
  NAND2_X1 U33380 ( .A1(n3894), .A2(n2839), .ZN(n2581) );
  NAND2_X1 U33390 ( .A1(n2597), .A2(IR_REG_31__SCAN_IN), .ZN(n2579) );
  XNOR2_X1 U33400 ( .A(n2579), .B(IR_REG_9__SCAN_IN), .ZN(n4496) );
  MUX2_X1 U33410 ( .A(n4496), .B(DATAI_9_), .S(n3749), .Z(n3632) );
  NAND2_X1 U33420 ( .A1(n3632), .A2(n2858), .ZN(n2580) );
  NAND2_X1 U33430 ( .A1(n2581), .A2(n2580), .ZN(n2582) );
  XNOR2_X1 U33440 ( .A(n2582), .B(n2886), .ZN(n2586) );
  INV_X1 U33450 ( .A(n2586), .ZN(n2583) );
  AOI22_X1 U33460 ( .A1(n2461), .A2(n3894), .B1(n2839), .B2(n3632), .ZN(n2585)
         );
  NAND2_X1 U33470 ( .A1(n2583), .A2(n2585), .ZN(n2584) );
  AND2_X1 U33480 ( .A1(n3626), .A2(n2584), .ZN(n2588) );
  INV_X1 U33490 ( .A(n2584), .ZN(n2587) );
  XNOR2_X1 U33500 ( .A(n2586), .B(n2585), .ZN(n3628) );
  NAND2_X1 U33510 ( .A1(n3750), .A2(REG1_REG_10__SCAN_IN), .ZN(n2596) );
  INV_X1 U33520 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2589) );
  OR2_X1 U3353 ( .A1(n3751), .A2(n2589), .ZN(n2595) );
  INV_X1 U33540 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4678) );
  NAND2_X1 U3355 ( .A1(n2591), .A2(n4678), .ZN(n2592) );
  NAND2_X1 U3356 ( .A1(n2626), .A2(n2592), .ZN(n3532) );
  OR2_X1 U3357 ( .A1(n2802), .A2(n3532), .ZN(n2594) );
  INV_X1 U3358 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3409) );
  OR2_X1 U3359 ( .A1(n2680), .A2(n3409), .ZN(n2593) );
  NAND4_X1 U3360 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n3677)
         );
  NAND2_X1 U3361 ( .A1(n3677), .A2(n2839), .ZN(n2606) );
  INV_X1 U3362 ( .A(n2597), .ZN(n2599) );
  INV_X1 U3363 ( .A(IR_REG_9__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U3364 ( .A1(n2599), .A2(n2598), .ZN(n2601) );
  NAND2_X1 U3365 ( .A1(n2601), .A2(IR_REG_31__SCAN_IN), .ZN(n2600) );
  MUX2_X1 U3366 ( .A(IR_REG_31__SCAN_IN), .B(n2600), .S(IR_REG_10__SCAN_IN), 
        .Z(n2604) );
  INV_X1 U3367 ( .A(n2601), .ZN(n2603) );
  INV_X1 U3368 ( .A(IR_REG_10__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U3369 ( .A1(n2603), .A2(n2602), .ZN(n2618) );
  NAND2_X1 U3370 ( .A1(n2604), .A2(n2618), .ZN(n3236) );
  MUX2_X1 U3371 ( .A(n4495), .B(DATAI_10_), .S(n3754), .Z(n3531) );
  NAND2_X1 U3372 ( .A1(n3531), .A2(n2858), .ZN(n2605) );
  NAND2_X1 U3373 ( .A1(n2606), .A2(n2605), .ZN(n2607) );
  XNOR2_X1 U3374 ( .A(n2607), .B(n2861), .ZN(n2608) );
  AOI22_X1 U3375 ( .A1(n2461), .A2(n3677), .B1(n2839), .B2(n3531), .ZN(n2609)
         );
  XNOR2_X1 U3376 ( .A(n2608), .B(n2609), .ZN(n3526) );
  INV_X1 U3377 ( .A(n2608), .ZN(n2611) );
  INV_X1 U3378 ( .A(n2609), .ZN(n2610) );
  NAND2_X1 U3379 ( .A1(n2611), .A2(n2610), .ZN(n2612) );
  NAND2_X1 U3380 ( .A1(n3750), .A2(REG1_REG_11__SCAN_IN), .ZN(n2617) );
  INV_X1 U3381 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4478) );
  OR2_X1 U3382 ( .A1(n3751), .A2(n4478), .ZN(n2616) );
  INV_X1 U3383 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4730) );
  XNOR2_X1 U3384 ( .A(n2626), .B(n4730), .ZN(n4314) );
  OR2_X1 U3385 ( .A1(n2802), .A2(n4314), .ZN(n2615) );
  INV_X1 U3386 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2613) );
  OR2_X1 U3387 ( .A1(n2680), .A2(n2613), .ZN(n2614) );
  NAND4_X1 U3388 ( .A1(n2617), .A2(n2616), .A3(n2615), .A4(n2614), .ZN(n3893)
         );
  NAND2_X1 U3389 ( .A1(n2461), .A2(n3893), .ZN(n2621) );
  NAND2_X1 U3390 ( .A1(n2618), .A2(IR_REG_31__SCAN_IN), .ZN(n2633) );
  INV_X1 U3391 ( .A(DATAI_11_), .ZN(n2619) );
  MUX2_X1 U3392 ( .A(n3395), .B(n2619), .S(n3749), .Z(n4311) );
  INV_X1 U3393 ( .A(n4311), .ZN(n4327) );
  NAND2_X1 U3394 ( .A1(n4327), .A2(n2767), .ZN(n2620) );
  NAND2_X1 U3395 ( .A1(n2621), .A2(n2620), .ZN(n3671) );
  NAND2_X1 U3396 ( .A1(n3893), .A2(n2839), .ZN(n2623) );
  NAND2_X1 U3397 ( .A1(n4327), .A2(n2858), .ZN(n2622) );
  NAND2_X1 U3398 ( .A1(n2623), .A2(n2622), .ZN(n2624) );
  XNOR2_X1 U3399 ( .A(n2624), .B(n2886), .ZN(n3672) );
  NAND2_X1 U3400 ( .A1(n3750), .A2(REG1_REG_12__SCAN_IN), .ZN(n2631) );
  INV_X1 U3401 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4474) );
  OR2_X1 U3402 ( .A1(n3751), .A2(n4474), .ZN(n2630) );
  INV_X1 U3403 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4731) );
  OAI21_X1 U3404 ( .B1(n2626), .B2(n4730), .A(n4731), .ZN(n2627) );
  NAND2_X1 U3405 ( .A1(REG3_REG_11__SCAN_IN), .A2(REG3_REG_12__SCAN_IN), .ZN(
        n2625) );
  NAND2_X1 U3406 ( .A1(n2627), .A2(n2647), .ZN(n3429) );
  OR2_X1 U3407 ( .A1(n2802), .A2(n3429), .ZN(n2629) );
  INV_X1 U3408 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3935) );
  OR2_X1 U3409 ( .A1(n2680), .A2(n3935), .ZN(n2628) );
  NAND4_X1 U3410 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n3892)
         );
  NAND2_X1 U3411 ( .A1(n3892), .A2(n2767), .ZN(n2638) );
  NAND2_X1 U3412 ( .A1(n2633), .A2(n2632), .ZN(n2634) );
  NAND2_X1 U3413 ( .A1(n2634), .A2(IR_REG_31__SCAN_IN), .ZN(n2635) );
  MUX2_X1 U3414 ( .A(DATAI_12_), .B(n4493), .S(n2636), .Z(n3582) );
  NAND2_X1 U3415 ( .A1(n3582), .A2(n2858), .ZN(n2637) );
  NAND2_X1 U3416 ( .A1(n2638), .A2(n2637), .ZN(n2639) );
  XNOR2_X1 U3417 ( .A(n2639), .B(n2886), .ZN(n2642) );
  NAND2_X1 U3418 ( .A1(n2461), .A2(n3892), .ZN(n2641) );
  NAND2_X1 U3419 ( .A1(n3582), .A2(n2839), .ZN(n2640) );
  NAND2_X1 U3420 ( .A1(n2641), .A2(n2640), .ZN(n2643) );
  AND2_X1 U3421 ( .A1(n2642), .A2(n2643), .ZN(n3575) );
  INV_X1 U3422 ( .A(n2642), .ZN(n2645) );
  INV_X1 U3423 ( .A(n2643), .ZN(n2644) );
  NAND2_X1 U3424 ( .A1(n2645), .A2(n2644), .ZN(n3576) );
  OAI21_X2 U3425 ( .B1(n3579), .B2(n3575), .A(n3576), .ZN(n3654) );
  NAND2_X1 U3426 ( .A1(n2936), .A2(REG0_REG_13__SCAN_IN), .ZN(n2652) );
  INV_X1 U3427 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4620) );
  OR2_X1 U3428 ( .A1(n2805), .A2(n4620), .ZN(n2651) );
  INV_X1 U3429 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U3430 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  NAND2_X1 U3431 ( .A1(n2660), .A2(n2648), .ZN(n4300) );
  OR2_X1 U3432 ( .A1(n2802), .A2(n4300), .ZN(n2650) );
  INV_X1 U3433 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4301) );
  OR2_X1 U3434 ( .A1(n2680), .A2(n4301), .ZN(n2649) );
  NAND2_X1 U3435 ( .A1(n4261), .A2(n2839), .ZN(n2655) );
  OR2_X1 U3436 ( .A1(n2668), .A2(n2172), .ZN(n2653) );
  XNOR2_X1 U3437 ( .A(n2653), .B(IR_REG_13__SCAN_IN), .ZN(n4582) );
  MUX2_X1 U3438 ( .A(n4582), .B(DATAI_13_), .S(n3749), .Z(n3656) );
  NAND2_X1 U3439 ( .A1(n3656), .A2(n2858), .ZN(n2654) );
  NAND2_X1 U3440 ( .A1(n2655), .A2(n2654), .ZN(n2656) );
  XNOR2_X1 U3441 ( .A(n2656), .B(n2861), .ZN(n3652) );
  NAND2_X1 U3442 ( .A1(n2461), .A2(n4261), .ZN(n2658) );
  NAND2_X1 U3443 ( .A1(n2839), .A2(n3656), .ZN(n2657) );
  NAND2_X1 U3444 ( .A1(n2658), .A2(n2657), .ZN(n3651) );
  NAND2_X1 U3445 ( .A1(n2660), .A2(n2659), .ZN(n2661) );
  AND2_X1 U3446 ( .A1(n2678), .A2(n2661), .ZN(n4275) );
  NAND2_X1 U3447 ( .A1(n2868), .A2(n4275), .ZN(n2666) );
  INV_X1 U3448 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4403) );
  OR2_X1 U3449 ( .A1(n2805), .A2(n4403), .ZN(n2665) );
  INV_X1 U3450 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4640) );
  OR2_X1 U3451 ( .A1(n3751), .A2(n4640), .ZN(n2664) );
  INV_X1 U3452 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2662) );
  OR2_X1 U3453 ( .A1(n2680), .A2(n2662), .ZN(n2663) );
  NAND4_X1 U3454 ( .A1(n2666), .A2(n2665), .A3(n2664), .A4(n2663), .ZN(n4292)
         );
  NAND2_X1 U3455 ( .A1(n4292), .A2(n2839), .ZN(n2673) );
  INV_X1 U3456 ( .A(IR_REG_13__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3457 ( .A1(n2668), .A2(n2667), .ZN(n2722) );
  NAND2_X1 U34580 ( .A1(n2722), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  INV_X1 U34590 ( .A(IR_REG_14__SCAN_IN), .ZN(n2669) );
  XNOR2_X1 U3460 ( .A(n2670), .B(n2669), .ZN(n4492) );
  INV_X1 U3461 ( .A(DATAI_14_), .ZN(n2671) );
  MUX2_X1 U3462 ( .A(n4492), .B(n2671), .S(n3754), .Z(n4273) );
  INV_X1 U3463 ( .A(n4273), .ZN(n3512) );
  NAND2_X1 U3464 ( .A1(n3512), .A2(n2858), .ZN(n2672) );
  NAND2_X1 U3465 ( .A1(n2673), .A2(n2672), .ZN(n2674) );
  XNOR2_X1 U3466 ( .A(n2674), .B(n2886), .ZN(n2707) );
  NAND2_X1 U34670 ( .A1(n2461), .A2(n4292), .ZN(n2676) );
  NAND2_X1 U3468 ( .A1(n3512), .A2(n2839), .ZN(n2675) );
  NAND2_X1 U34690 ( .A1(n2676), .A2(n2675), .ZN(n2708) );
  NAND2_X1 U3470 ( .A1(n2678), .A2(n2677), .ZN(n2679) );
  NAND2_X1 U34710 ( .A1(n2693), .A2(n2679), .ZN(n3732) );
  INV_X1 U3472 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2681) );
  OR2_X1 U34730 ( .A1(n2680), .A2(n2681), .ZN(n2682) );
  OAI21_X1 U3474 ( .B1(n3732), .B2(n2802), .A(n2682), .ZN(n2685) );
  INV_X1 U34750 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4399) );
  INV_X1 U3476 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4463) );
  OR2_X1 U34770 ( .A1(n3751), .A2(n4463), .ZN(n2683) );
  OAI21_X1 U3478 ( .B1(n2805), .B2(n4399), .A(n2683), .ZN(n2684) );
  NAND2_X1 U34790 ( .A1(n2461), .A2(n4264), .ZN(n2688) );
  NAND2_X1 U3480 ( .A1(n2686), .A2(IR_REG_31__SCAN_IN), .ZN(n2702) );
  XNOR2_X1 U34810 ( .A(n2702), .B(IR_REG_15__SCAN_IN), .ZN(n3955) );
  MUX2_X1 U3482 ( .A(n3955), .B(DATAI_15_), .S(n3754), .Z(n3729) );
  NAND2_X1 U34830 ( .A1(n2767), .A2(n3729), .ZN(n2687) );
  NAND2_X1 U3484 ( .A1(n2688), .A2(n2687), .ZN(n3724) );
  NAND2_X1 U34850 ( .A1(n4264), .A2(n2767), .ZN(n2690) );
  NAND2_X1 U3486 ( .A1(n3729), .A2(n2858), .ZN(n2689) );
  NAND2_X1 U34870 ( .A1(n2690), .A2(n2689), .ZN(n2691) );
  XNOR2_X1 U3488 ( .A(n2691), .B(n2886), .ZN(n3592) );
  INV_X1 U34890 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2692) );
  NAND2_X1 U3490 ( .A1(n2693), .A2(n2692), .ZN(n2694) );
  NAND2_X1 U34910 ( .A1(n2716), .A2(n2694), .ZN(n4234) );
  OR2_X1 U3492 ( .A1(n4234), .A2(n2802), .ZN(n2700) );
  INV_X1 U34930 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4532) );
  OR2_X1 U3494 ( .A1(n2805), .A2(n4532), .ZN(n2697) );
  INV_X1 U34950 ( .A(REG0_REG_16__SCAN_IN), .ZN(n2695) );
  OR2_X1 U3496 ( .A1(n3751), .A2(n2695), .ZN(n2696) );
  AND2_X1 U34970 ( .A1(n2697), .A2(n2696), .ZN(n2699) );
  NAND2_X1 U3498 ( .A1(n2467), .A2(REG2_REG_16__SCAN_IN), .ZN(n2698) );
  NAND2_X1 U34990 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  NAND2_X1 U3500 ( .A1(n2703), .A2(IR_REG_31__SCAN_IN), .ZN(n2704) );
  INV_X1 U35010 ( .A(n4579), .ZN(n2705) );
  MUX2_X1 U3502 ( .A(n2705), .B(DATAI_16_), .S(n3749), .Z(n4233) );
  INV_X1 U35030 ( .A(n4233), .ZN(n4226) );
  OAI22_X1 U3504 ( .A1(n4208), .A2(n2837), .B1(n2885), .B2(n4226), .ZN(n2706)
         );
  XNOR2_X1 U35050 ( .A(n2706), .B(n2886), .ZN(n2713) );
  OAI22_X1 U35060 ( .A1(n4208), .A2(n2888), .B1(n2837), .B2(n4226), .ZN(n2712)
         );
  INV_X1 U35070 ( .A(n2707), .ZN(n2710) );
  INV_X1 U35080 ( .A(n2708), .ZN(n2709) );
  NAND2_X1 U35090 ( .A1(n2710), .A2(n2709), .ZN(n3507) );
  OAI211_X1 U35100 ( .C1(n3724), .C2(n3592), .A(n2711), .B(n3507), .ZN(n2715)
         );
  INV_X1 U35110 ( .A(n2711), .ZN(n3589) );
  AND2_X1 U35120 ( .A1(n2713), .A2(n2712), .ZN(n3588) );
  AOI21_X1 U35130 ( .B1(n3724), .B2(n3592), .A(n3588), .ZN(n2714) );
  NAND2_X1 U35140 ( .A1(n2716), .A2(n4719), .ZN(n2717) );
  NAND2_X1 U35150 ( .A1(n2733), .A2(n2717), .ZN(n3610) );
  AOI22_X1 U35160 ( .A1(n3750), .A2(REG1_REG_17__SCAN_IN), .B1(n2936), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2719) );
  OR2_X1 U35170 ( .A1(n2680), .A2(n3971), .ZN(n2718) );
  OAI211_X1 U35180 ( .C1(n3610), .C2(n2802), .A(n2719), .B(n2718), .ZN(n4224)
         );
  NAND2_X1 U35190 ( .A1(n4224), .A2(n2839), .ZN(n2726) );
  NAND2_X1 U35200 ( .A1(n2720), .A2(n4753), .ZN(n2721) );
  OAI21_X1 U35210 ( .B1(n2722), .B2(n2721), .A(IR_REG_31__SCAN_IN), .ZN(n2723)
         );
  MUX2_X1 U35220 ( .A(IR_REG_31__SCAN_IN), .B(n2723), .S(IR_REG_17__SCAN_IN), 
        .Z(n2724) );
  MUX2_X1 U35230 ( .A(n4491), .B(DATAI_17_), .S(n3754), .Z(n4214) );
  NAND2_X1 U35240 ( .A1(n4214), .A2(n2858), .ZN(n2725) );
  NAND2_X1 U35250 ( .A1(n2726), .A2(n2725), .ZN(n2727) );
  XNOR2_X1 U35260 ( .A(n2727), .B(n2861), .ZN(n2730) );
  AND2_X1 U35270 ( .A1(n2767), .A2(n4214), .ZN(n2728) );
  AOI21_X1 U35280 ( .B1(n4224), .B2(n2461), .A(n2728), .ZN(n2729) );
  NOR2_X1 U35290 ( .A1(n2730), .A2(n2729), .ZN(n3604) );
  NAND2_X1 U35300 ( .A1(n2730), .A2(n2729), .ZN(n3605) );
  INV_X1 U35310 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U35320 ( .A1(n2733), .A2(n2732), .ZN(n2734) );
  NAND2_X1 U35330 ( .A1(n2744), .A2(n2734), .ZN(n4197) );
  INV_X1 U35340 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3965) );
  NAND2_X1 U35350 ( .A1(n2467), .A2(REG2_REG_18__SCAN_IN), .ZN(n2736) );
  NAND2_X1 U35360 ( .A1(n2936), .A2(REG0_REG_18__SCAN_IN), .ZN(n2735) );
  OAI211_X1 U35370 ( .C1(n2805), .C2(n3965), .A(n2736), .B(n2735), .ZN(n2737)
         );
  INV_X1 U35380 ( .A(n2737), .ZN(n2738) );
  NAND2_X1 U35390 ( .A1(n2740), .A2(IR_REG_31__SCAN_IN), .ZN(n2741) );
  MUX2_X1 U35400 ( .A(n4576), .B(DATAI_18_), .S(n3754), .Z(n4193) );
  INV_X1 U35410 ( .A(n4193), .ZN(n2994) );
  OAI22_X1 U35420 ( .A1(n4175), .A2(n2888), .B1(n2837), .B2(n2994), .ZN(n3539)
         );
  OAI22_X1 U35430 ( .A1(n4175), .A2(n2837), .B1(n2885), .B2(n2994), .ZN(n2742)
         );
  XNOR2_X1 U35440 ( .A(n2742), .B(n2886), .ZN(n3684) );
  NAND2_X1 U35450 ( .A1(n2744), .A2(n2743), .ZN(n2745) );
  NAND2_X1 U35460 ( .A1(n2772), .A2(n2745), .ZN(n4182) );
  INV_X1 U35470 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4183) );
  NAND2_X1 U35480 ( .A1(n3750), .A2(REG1_REG_19__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U35490 ( .A1(n2936), .A2(REG0_REG_19__SCAN_IN), .ZN(n2746) );
  OAI211_X1 U35500 ( .C1(n4183), .C2(n2680), .A(n2747), .B(n2746), .ZN(n2748)
         );
  INV_X1 U35510 ( .A(n2748), .ZN(n2749) );
  INV_X1 U35520 ( .A(DATAI_19_), .ZN(n2751) );
  OAI22_X1 U35530 ( .A1(n4190), .A2(n2837), .B1(n2885), .B2(n4181), .ZN(n2752)
         );
  XNOR2_X1 U35540 ( .A(n2752), .B(n2886), .ZN(n2754) );
  OAI22_X1 U35550 ( .A1(n4190), .A2(n2888), .B1(n2837), .B2(n4181), .ZN(n2753)
         );
  AOI21_X1 U35560 ( .B1(n3539), .B2(n3684), .A(n3541), .ZN(n2757) );
  NOR2_X1 U35570 ( .A1(n2754), .A2(n2753), .ZN(n3542) );
  XNOR2_X1 U35580 ( .A(n2772), .B(REG3_REG_20__SCAN_IN), .ZN(n4162) );
  NAND2_X1 U35590 ( .A1(n4162), .A2(n2868), .ZN(n2763) );
  INV_X1 U35600 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2760) );
  NAND2_X1 U35610 ( .A1(n3750), .A2(REG1_REG_20__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U35620 ( .A1(n2936), .A2(REG0_REG_20__SCAN_IN), .ZN(n2758) );
  OAI211_X1 U35630 ( .C1(n2760), .C2(n2680), .A(n2759), .B(n2758), .ZN(n2761)
         );
  INV_X1 U35640 ( .A(n2761), .ZN(n2762) );
  NAND2_X1 U35650 ( .A1(n4177), .A2(n2839), .ZN(n2765) );
  NAND2_X1 U35660 ( .A1(n2858), .A2(n4150), .ZN(n2764) );
  NAND2_X1 U35670 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  XNOR2_X1 U35680 ( .A(n2766), .B(n2861), .ZN(n2770) );
  INV_X1 U35690 ( .A(n4150), .ZN(n4160) );
  NOR2_X1 U35700 ( .A1(n2875), .A2(n4160), .ZN(n2768) );
  AOI21_X1 U35710 ( .B1(n4177), .B2(n2461), .A(n2768), .ZN(n2769) );
  NOR2_X1 U35720 ( .A1(n2770), .A2(n2769), .ZN(n3640) );
  INV_X1 U35730 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3645) );
  INV_X1 U35740 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2771) );
  OAI21_X1 U35750 ( .B1(n2772), .B2(n3645), .A(n2771), .ZN(n2773) );
  AND2_X1 U35760 ( .A1(n2789), .A2(n2773), .ZN(n4139) );
  NAND2_X1 U35770 ( .A1(n4139), .A2(n2868), .ZN(n2778) );
  INV_X1 U35780 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U35790 ( .A1(n3750), .A2(REG1_REG_21__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U35800 ( .A1(n2467), .A2(REG2_REG_21__SCAN_IN), .ZN(n2774) );
  OAI211_X1 U35810 ( .C1(n3751), .C2(n4718), .A(n2775), .B(n2774), .ZN(n2776)
         );
  INV_X1 U3582 ( .A(n2776), .ZN(n2777) );
  NAND2_X1 U3583 ( .A1(n4118), .A2(n2839), .ZN(n2780) );
  NAND2_X1 U3584 ( .A1(n2858), .A2(n3569), .ZN(n2779) );
  NAND2_X1 U3585 ( .A1(n2780), .A2(n2779), .ZN(n2781) );
  XNOR2_X1 U3586 ( .A(n2781), .B(n2886), .ZN(n2787) );
  INV_X1 U3587 ( .A(n2787), .ZN(n2785) );
  NAND2_X1 U3588 ( .A1(n4118), .A2(n2461), .ZN(n2783) );
  INV_X1 U3589 ( .A(n3569), .ZN(n4138) );
  OR2_X1 U3590 ( .A1(n2837), .A2(n4138), .ZN(n2782) );
  NAND2_X1 U3591 ( .A1(n2783), .A2(n2782), .ZN(n2786) );
  INV_X1 U3592 ( .A(n2786), .ZN(n2784) );
  INV_X1 U3593 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U3594 ( .A1(n2789), .A2(n4654), .ZN(n2790) );
  AND2_X1 U3595 ( .A1(n2800), .A2(n2790), .ZN(n4123) );
  NAND2_X1 U3596 ( .A1(n4123), .A2(n2868), .ZN(n2796) );
  INV_X1 U3597 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U3598 ( .A1(n3750), .A2(REG1_REG_22__SCAN_IN), .ZN(n2792) );
  NAND2_X1 U3599 ( .A1(n2936), .A2(REG0_REG_22__SCAN_IN), .ZN(n2791) );
  OAI211_X1 U3600 ( .C1(n2793), .C2(n2680), .A(n2792), .B(n2791), .ZN(n2794)
         );
  INV_X1 U3601 ( .A(n2794), .ZN(n2795) );
  OAI22_X1 U3602 ( .A1(n4133), .A2(n2888), .B1(n2837), .B2(n4125), .ZN(n2811)
         );
  OAI22_X1 U3603 ( .A1(n4133), .A2(n2837), .B1(n2885), .B2(n4125), .ZN(n2797)
         );
  XNOR2_X1 U3604 ( .A(n2797), .B(n2886), .ZN(n2810) );
  XOR2_X1 U3605 ( .A(n2811), .B(n2810), .Z(n3664) );
  INV_X1 U3606 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2799) );
  NAND2_X1 U3607 ( .A1(n2800), .A2(n2799), .ZN(n2801) );
  NAND2_X1 U3608 ( .A1(n2818), .A2(n2801), .ZN(n4107) );
  INV_X1 U3609 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4681) );
  NAND2_X1 U3610 ( .A1(n2467), .A2(REG2_REG_23__SCAN_IN), .ZN(n2804) );
  INV_X1 U3611 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4759) );
  OR2_X1 U3612 ( .A1(n3751), .A2(n4759), .ZN(n2803) );
  OAI211_X1 U3613 ( .C1(n2805), .C2(n4681), .A(n2804), .B(n2803), .ZN(n2806)
         );
  INV_X1 U3614 ( .A(n2806), .ZN(n2807) );
  OAI22_X1 U3615 ( .A1(n4120), .A2(n2837), .B1(n2885), .B2(n4105), .ZN(n2809)
         );
  XNOR2_X1 U3616 ( .A(n2809), .B(n2861), .ZN(n2815) );
  OAI22_X1 U3617 ( .A1(n4120), .A2(n2888), .B1(n2837), .B2(n4105), .ZN(n2816)
         );
  XNOR2_X1 U3618 ( .A(n2815), .B(n2816), .ZN(n3518) );
  INV_X1 U3619 ( .A(n2810), .ZN(n2813) );
  INV_X1 U3620 ( .A(n2811), .ZN(n2812) );
  NAND2_X1 U3621 ( .A1(n2813), .A2(n2812), .ZN(n3519) );
  INV_X1 U3622 ( .A(n2815), .ZN(n2817) );
  NAND2_X1 U3623 ( .A1(n2817), .A2(n2816), .ZN(n3461) );
  INV_X1 U3624 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3619) );
  NAND2_X1 U3625 ( .A1(n2818), .A2(n3619), .ZN(n2819) );
  NAND2_X1 U3626 ( .A1(n4089), .A2(n2868), .ZN(n2824) );
  INV_X1 U3627 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U3628 ( .A1(n3750), .A2(REG1_REG_24__SCAN_IN), .ZN(n2821) );
  INV_X1 U3629 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4758) );
  OR2_X1 U3630 ( .A1(n3751), .A2(n4758), .ZN(n2820) );
  OAI211_X1 U3631 ( .C1(n4685), .C2(n2680), .A(n2821), .B(n2820), .ZN(n2822)
         );
  INV_X1 U3632 ( .A(n2822), .ZN(n2823) );
  NOR2_X1 U3633 ( .A1(n2875), .A2(n4087), .ZN(n2825) );
  AOI21_X1 U3634 ( .B1(n4102), .B2(n2461), .A(n2825), .ZN(n3460) );
  NAND2_X1 U3635 ( .A1(n3461), .A2(n3460), .ZN(n3458) );
  NAND2_X1 U3636 ( .A1(n4102), .A2(n2767), .ZN(n2827) );
  NAND2_X1 U3637 ( .A1(n2858), .A2(n3621), .ZN(n2826) );
  NAND2_X1 U3638 ( .A1(n2827), .A2(n2826), .ZN(n2828) );
  XNOR2_X1 U3639 ( .A(n2828), .B(n2861), .ZN(n3463) );
  NAND2_X1 U3640 ( .A1(n3461), .A2(n3463), .ZN(n2841) );
  INV_X1 U3641 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2829) );
  NAND2_X1 U3642 ( .A1(n2830), .A2(n2829), .ZN(n2831) );
  NAND2_X1 U3643 ( .A1(n2851), .A2(n2831), .ZN(n4073) );
  INV_X1 U3644 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4072) );
  NAND2_X1 U3645 ( .A1(n3750), .A2(REG1_REG_25__SCAN_IN), .ZN(n2833) );
  NAND2_X1 U3646 ( .A1(n2936), .A2(REG0_REG_25__SCAN_IN), .ZN(n2832) );
  OAI211_X1 U3647 ( .C1(n4072), .C2(n2680), .A(n2833), .B(n2832), .ZN(n2834)
         );
  INV_X1 U3648 ( .A(n2834), .ZN(n2835) );
  OAI22_X1 U3649 ( .A1(n4048), .A2(n2837), .B1(n2885), .B2(n4070), .ZN(n2838)
         );
  XOR2_X1 U3650 ( .A(n2886), .B(n2838), .Z(n3466) );
  NOR2_X1 U3651 ( .A1(n2837), .A2(n4070), .ZN(n2840) );
  AOI21_X1 U3652 ( .B1(n4082), .B2(n2461), .A(n2840), .ZN(n3465) );
  NOR2_X1 U3653 ( .A1(n3466), .A2(n3465), .ZN(n3464) );
  AOI21_X1 U3654 ( .B1(n3458), .B2(n2841), .A(n3464), .ZN(n2849) );
  INV_X1 U3655 ( .A(n3465), .ZN(n2845) );
  NAND2_X1 U3656 ( .A1(n3463), .A2(n3460), .ZN(n2843) );
  INV_X1 U3657 ( .A(n3466), .ZN(n2842) );
  AOI21_X1 U3658 ( .B1(n2845), .B2(n2843), .A(n2842), .ZN(n2847) );
  INV_X1 U3659 ( .A(n3463), .ZN(n3617) );
  INV_X1 U3660 ( .A(n3460), .ZN(n2844) );
  NOR3_X1 U3661 ( .A1(n2845), .A2(n3617), .A3(n2844), .ZN(n2846) );
  AOI21_X2 U3662 ( .B1(n3517), .B2(n2849), .A(n2848), .ZN(n3712) );
  INV_X1 U3663 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2850) );
  NAND2_X1 U3664 ( .A1(n2851), .A2(n2850), .ZN(n2852) );
  NAND2_X1 U3665 ( .A1(n4056), .A2(n2868), .ZN(n2857) );
  INV_X1 U3666 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4684) );
  NAND2_X1 U3667 ( .A1(n3750), .A2(REG1_REG_26__SCAN_IN), .ZN(n2854) );
  INV_X1 U3668 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4645) );
  OR2_X1 U3669 ( .A1(n3751), .A2(n4645), .ZN(n2853) );
  OAI211_X1 U3670 ( .C1(n4684), .C2(n2680), .A(n2854), .B(n2853), .ZN(n2855)
         );
  INV_X1 U3671 ( .A(n2855), .ZN(n2856) );
  NAND2_X1 U3672 ( .A1(n4065), .A2(n2839), .ZN(n2860) );
  NAND2_X1 U3673 ( .A1(n2858), .A2(n3713), .ZN(n2859) );
  NAND2_X1 U3674 ( .A1(n2860), .A2(n2859), .ZN(n2862) );
  XNOR2_X1 U3675 ( .A(n2862), .B(n2861), .ZN(n2865) );
  NOR2_X1 U3676 ( .A1(n2837), .A2(n4055), .ZN(n2863) );
  AOI21_X1 U3677 ( .B1(n4065), .B2(n2005), .A(n2863), .ZN(n2864) );
  NOR2_X1 U3678 ( .A1(n2865), .A2(n2864), .ZN(n3710) );
  NAND2_X1 U3679 ( .A1(n2865), .A2(n2864), .ZN(n3708) );
  INV_X1 U3680 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4692) );
  OR2_X2 U3681 ( .A1(n2866), .A2(n4692), .ZN(n2878) );
  NAND2_X1 U3682 ( .A1(n2866), .A2(n4692), .ZN(n2867) );
  NAND2_X1 U3683 ( .A1(n4038), .A2(n2868), .ZN(n2873) );
  INV_X1 U3684 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U3685 ( .A1(n3750), .A2(REG1_REG_27__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U3686 ( .A1(n2936), .A2(REG0_REG_27__SCAN_IN), .ZN(n2869) );
  OAI211_X1 U3687 ( .C1(n4633), .C2(n2680), .A(n2870), .B(n2869), .ZN(n2871)
         );
  INV_X1 U3688 ( .A(n2871), .ZN(n2872) );
  OAI22_X1 U3689 ( .A1(n3041), .A2(n2837), .B1(n4037), .B2(n2885), .ZN(n2874)
         );
  XNOR2_X1 U3690 ( .A(n2874), .B(n2886), .ZN(n2915) );
  OAI22_X1 U3691 ( .A1(n3041), .A2(n2888), .B1(n2875), .B2(n4037), .ZN(n2914)
         );
  XNOR2_X1 U3692 ( .A(n2915), .B(n2914), .ZN(n3499) );
  INV_X1 U3693 ( .A(n2878), .ZN(n2876) );
  NAND2_X1 U3694 ( .A1(n2876), .A2(REG3_REG_28__SCAN_IN), .ZN(n4019) );
  INV_X1 U3695 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U3696 ( .A1(n2878), .A2(n2877), .ZN(n2879) );
  NAND2_X1 U3697 ( .A1(n4019), .A2(n2879), .ZN(n3482) );
  INV_X1 U3698 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U3699 ( .A1(n3750), .A2(REG1_REG_28__SCAN_IN), .ZN(n2881) );
  NAND2_X1 U3700 ( .A1(n2936), .A2(REG0_REG_28__SCAN_IN), .ZN(n2880) );
  OAI211_X1 U3701 ( .C1(n3481), .C2(n2680), .A(n2881), .B(n2880), .ZN(n2882)
         );
  INV_X1 U3702 ( .A(n2882), .ZN(n2883) );
  AND2_X2 U3703 ( .A1(n2884), .A2(n2883), .ZN(n4014) );
  INV_X1 U3704 ( .A(n4001), .ZN(n3040) );
  OAI22_X1 U3705 ( .A1(n4014), .A2(n2837), .B1(n2885), .B2(n3040), .ZN(n2887)
         );
  XNOR2_X1 U3706 ( .A(n2887), .B(n2886), .ZN(n2890) );
  OAI22_X1 U3707 ( .A1(n4014), .A2(n2888), .B1(n2837), .B2(n3040), .ZN(n2889)
         );
  XNOR2_X1 U3708 ( .A(n2890), .B(n2889), .ZN(n2916) );
  INV_X1 U3709 ( .A(n2916), .ZN(n2919) );
  NAND2_X1 U3710 ( .A1(n2891), .A2(B_REG_SCAN_IN), .ZN(n2893) );
  MUX2_X1 U3711 ( .A(n2893), .B(B_REG_SCAN_IN), .S(n4486), .Z(n2895) );
  INV_X1 U3712 ( .A(n3251), .ZN(n3058) );
  INV_X1 U3713 ( .A(n3064), .ZN(n2907) );
  NOR4_X1 U3714 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2899) );
  NOR4_X1 U3715 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2898) );
  NOR4_X1 U3716 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2897) );
  NOR4_X1 U3717 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2896) );
  NAND4_X1 U3718 ( .A1(n2899), .A2(n2898), .A3(n2897), .A4(n2896), .ZN(n2904)
         );
  NOR2_X1 U3719 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_15__SCAN_IN), .ZN(n4649)
         );
  NOR4_X1 U3720 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2902) );
  NOR4_X1 U3721 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2901) );
  NOR4_X1 U3722 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2900) );
  NAND4_X1 U3723 ( .A1(n4649), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(n2903)
         );
  NOR2_X1 U3724 ( .A1(n2904), .A2(n2903), .ZN(n3045) );
  NAND2_X1 U3725 ( .A1(n3045), .A2(D_REG_1__SCAN_IN), .ZN(n2906) );
  INV_X1 U3726 ( .A(n2894), .ZN(n2905) );
  NAND2_X1 U3727 ( .A1(n2905), .A2(n2891), .ZN(n3046) );
  INV_X1 U3728 ( .A(n3046), .ZN(n3068) );
  AOI21_X1 U3729 ( .B1(n2907), .B2(n2906), .A(n3068), .ZN(n3253) );
  INV_X1 U3730 ( .A(n3070), .ZN(n3039) );
  OAI211_X1 U3731 ( .C1(n3149), .C2(n3979), .A(n4289), .B(n3039), .ZN(n2920)
         );
  INV_X1 U3732 ( .A(n2920), .ZN(n2912) );
  NAND2_X1 U3733 ( .A1(n2909), .A2(IR_REG_31__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U3734 ( .A1(n2912), .A2(n3177), .ZN(n2913) );
  NAND2_X1 U3735 ( .A1(n2915), .A2(n2914), .ZN(n2918) );
  NAND3_X1 U3736 ( .A1(n2919), .A2(n3726), .A3(n2918), .ZN(n2952) );
  NAND2_X1 U3737 ( .A1(n2953), .A2(n2917), .ZN(n2951) );
  NOR3_X1 U3738 ( .A1(n2919), .A2(n3719), .A3(n2918), .ZN(n2949) );
  NAND2_X1 U3739 ( .A1(n2920), .A2(n4289), .ZN(n2921) );
  NAND2_X1 U3740 ( .A1(n2928), .A2(n2921), .ZN(n2923) );
  NAND2_X1 U3741 ( .A1(n2408), .A2(n3979), .ZN(n2922) );
  NAND2_X1 U3742 ( .A1(n2922), .A2(n3070), .ZN(n3047) );
  NAND2_X1 U3743 ( .A1(n2923), .A2(n3047), .ZN(n3179) );
  NAND2_X1 U3744 ( .A1(n2421), .A2(n3069), .ZN(n2924) );
  OAI21_X1 U3745 ( .B1(n3179), .B2(n2924), .A(STATE_REG_SCAN_IN), .ZN(n2929)
         );
  OR2_X1 U3746 ( .A1(n2925), .A2(n4574), .ZN(n2926) );
  INV_X1 U3747 ( .A(n2934), .ZN(n2927) );
  NAND2_X1 U3748 ( .A1(n2928), .A2(n2927), .ZN(n3176) );
  NAND2_X1 U3749 ( .A1(n2055), .A2(IR_REG_31__SCAN_IN), .ZN(n2930) );
  MUX2_X1 U3750 ( .A(IR_REG_31__SCAN_IN), .B(n2930), .S(IR_REG_28__SCAN_IN), 
        .Z(n2933) );
  INV_X1 U3751 ( .A(n2931), .ZN(n2932) );
  NAND2_X1 U3752 ( .A1(n2933), .A2(n2932), .ZN(n3904) );
  NOR2_X1 U3753 ( .A1(n2934), .A2(n3904), .ZN(n3885) );
  NOR2_X1 U3754 ( .A1(n2934), .A2(n4484), .ZN(n2935) );
  INV_X1 U3755 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U3756 ( .A1(n3750), .A2(REG1_REG_29__SCAN_IN), .ZN(n2938) );
  NAND2_X1 U3757 ( .A1(n2936), .A2(REG0_REG_29__SCAN_IN), .ZN(n2937) );
  OAI211_X1 U3758 ( .C1(n4023), .C2(n2680), .A(n2938), .B(n2937), .ZN(n2939)
         );
  INV_X1 U3759 ( .A(n2939), .ZN(n2940) );
  AOI22_X1 U3760 ( .A1(n4050), .A2(n3728), .B1(n3731), .B2(n4774), .ZN(n2947)
         );
  AND2_X1 U3761 ( .A1(n3177), .A2(n4326), .ZN(n2942) );
  NAND2_X1 U3762 ( .A1(n2943), .A2(n2942), .ZN(n2945) );
  AND3_X1 U3763 ( .A1(n4595), .A2(n3177), .A3(n3807), .ZN(n4566) );
  NAND2_X2 U3764 ( .A1(n2945), .A2(n4313), .ZN(n3730) );
  AOI22_X1 U3765 ( .A1(n3730), .A2(n4001), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2946) );
  OAI211_X1 U3766 ( .C1(n3695), .C2(n3482), .A(n2947), .B(n2946), .ZN(n2948)
         );
  NOR2_X1 U3767 ( .A1(n2949), .A2(n2948), .ZN(n2950) );
  OAI211_X1 U3768 ( .C1(n2953), .C2(n2952), .A(n2951), .B(n2950), .ZN(U3217)
         );
  NAND2_X1 U3769 ( .A1(n3009), .A2(n3810), .ZN(n3007) );
  NAND2_X1 U3770 ( .A1(n2958), .A2(n2954), .ZN(n3816) );
  NAND2_X1 U3771 ( .A1(n3900), .A2(n3288), .ZN(n2959) );
  INV_X1 U3772 ( .A(n3899), .ZN(n2964) );
  NAND2_X1 U3773 ( .A1(n3899), .A2(n3452), .ZN(n3822) );
  NAND2_X1 U3774 ( .A1(n3899), .A2(n2317), .ZN(n2965) );
  AND2_X1 U3775 ( .A1(n3898), .A2(n3299), .ZN(n3269) );
  NAND2_X1 U3776 ( .A1(n2967), .A2(n2966), .ZN(n3268) );
  INV_X1 U3777 ( .A(n3702), .ZN(n2968) );
  AND2_X1 U3778 ( .A1(n3897), .A2(n3702), .ZN(n2973) );
  AOI22_X1 U3779 ( .A1(n3790), .A2(n2973), .B1(n3492), .B2(n3896), .ZN(n2974)
         );
  NAND2_X1 U3780 ( .A1(n2975), .A2(n2974), .ZN(n3354) );
  OR2_X1 U3781 ( .A1(n3557), .A2(n3895), .ZN(n2976) );
  NAND2_X1 U3782 ( .A1(n3354), .A2(n2976), .ZN(n2978) );
  NAND2_X1 U3783 ( .A1(n3895), .A2(n3557), .ZN(n2977) );
  NAND2_X1 U3784 ( .A1(n2978), .A2(n2977), .ZN(n3372) );
  OR2_X1 U3785 ( .A1(n3632), .A2(n3894), .ZN(n2979) );
  NOR2_X1 U3786 ( .A1(n3677), .A2(n3531), .ZN(n2980) );
  INV_X1 U3787 ( .A(n3677), .ZN(n4321) );
  INV_X1 U3788 ( .A(n3531), .ZN(n3021) );
  OR2_X1 U3789 ( .A1(n4311), .A2(n3893), .ZN(n3420) );
  NAND2_X1 U3790 ( .A1(n3893), .A2(n4311), .ZN(n3843) );
  OR2_X1 U3791 ( .A1(n4327), .A2(n3893), .ZN(n2982) );
  NAND2_X1 U3792 ( .A1(n4307), .A2(n2982), .ZN(n3425) );
  NAND2_X1 U3793 ( .A1(n3892), .A2(n3582), .ZN(n2983) );
  INV_X1 U3794 ( .A(n3892), .ZN(n4319) );
  INV_X1 U3795 ( .A(n3582), .ZN(n3427) );
  NAND2_X1 U3796 ( .A1(n4319), .A2(n3427), .ZN(n2984) );
  NAND2_X1 U3797 ( .A1(n4261), .A2(n3656), .ZN(n2985) );
  INV_X1 U3798 ( .A(n4260), .ZN(n2988) );
  OR2_X1 U3799 ( .A1(n4292), .A2(n4273), .ZN(n4239) );
  NAND2_X1 U3800 ( .A1(n4292), .A2(n4273), .ZN(n3738) );
  NAND2_X1 U3801 ( .A1(n4239), .A2(n3738), .ZN(n2987) );
  INV_X1 U3802 ( .A(n4292), .ZN(n4241) );
  NAND2_X1 U3803 ( .A1(n4241), .A2(n4273), .ZN(n2989) );
  NAND2_X1 U3804 ( .A1(n4264), .A2(n3729), .ZN(n2991) );
  NOR2_X1 U3805 ( .A1(n4264), .A2(n3729), .ZN(n2990) );
  NAND2_X1 U3806 ( .A1(n4208), .A2(n4233), .ZN(n3856) );
  NAND2_X1 U3807 ( .A1(n4243), .A2(n4226), .ZN(n3852) );
  NAND2_X1 U3808 ( .A1(n3856), .A2(n3852), .ZN(n4231) );
  NAND2_X1 U3809 ( .A1(n4232), .A2(n4231), .ZN(n4229) );
  NAND2_X1 U3810 ( .A1(n4243), .A2(n4233), .ZN(n2992) );
  NAND2_X1 U3811 ( .A1(n4175), .A2(n4193), .ZN(n4171) );
  NAND2_X1 U3812 ( .A1(n4210), .A2(n2994), .ZN(n4172) );
  NAND2_X1 U3813 ( .A1(n4171), .A2(n4172), .ZN(n4201) );
  INV_X1 U3814 ( .A(n4181), .ZN(n3547) );
  NOR2_X1 U3815 ( .A1(n4177), .A2(n4150), .ZN(n2996) );
  INV_X1 U3816 ( .A(n4177), .ZN(n2995) );
  NAND2_X1 U3817 ( .A1(n3891), .A2(n4125), .ZN(n3032) );
  NAND2_X1 U3818 ( .A1(n4098), .A2(n3032), .ZN(n4115) );
  INV_X1 U3819 ( .A(n4125), .ZN(n2999) );
  NAND2_X1 U3820 ( .A1(n4120), .A2(n4105), .ZN(n3001) );
  INV_X1 U3821 ( .A(n4105), .ZN(n3035) );
  NAND2_X1 U3822 ( .A1(n4102), .A2(n3621), .ZN(n3003) );
  NOR2_X1 U3823 ( .A1(n4102), .A2(n3621), .ZN(n3002) );
  NAND2_X1 U3824 ( .A1(n4065), .A2(n3713), .ZN(n3004) );
  NAND2_X1 U3825 ( .A1(n3041), .A2(n4037), .ZN(n3005) );
  NAND2_X1 U3826 ( .A1(n4014), .A2(n4001), .ZN(n4006) );
  NAND2_X1 U3827 ( .A1(n4035), .A2(n3040), .ZN(n4005) );
  NAND2_X1 U3828 ( .A1(n4006), .A2(n4005), .ZN(n4000) );
  XNOR2_X1 U3829 ( .A(n3999), .B(n4000), .ZN(n3479) );
  XNOR2_X1 U3830 ( .A(n2402), .B(n4487), .ZN(n3006) );
  NAND2_X1 U3831 ( .A1(n3006), .A2(n3979), .ZN(n4322) );
  NAND2_X1 U3832 ( .A1(n3479), .A2(n4411), .ZN(n3044) );
  INV_X1 U3833 ( .A(n3198), .ZN(n3779) );
  INV_X1 U3834 ( .A(n3288), .ZN(n3011) );
  OR2_X1 U3835 ( .A1(n3011), .A2(n3900), .ZN(n3818) );
  NAND2_X1 U3836 ( .A1(n3900), .A2(n3011), .ZN(n3815) );
  NAND2_X1 U3837 ( .A1(n3012), .A2(n3818), .ZN(n3445) );
  OR2_X1 U3838 ( .A1(n2966), .A2(n3898), .ZN(n3835) );
  NAND2_X1 U3839 ( .A1(n3898), .A2(n2966), .ZN(n3821) );
  AND2_X1 U3840 ( .A1(n3897), .A2(n2968), .ZN(n3836) );
  INV_X1 U3841 ( .A(n3836), .ZN(n3014) );
  OR2_X1 U3842 ( .A1(n2968), .A2(n3897), .ZN(n3824) );
  INV_X1 U3843 ( .A(n3825), .ZN(n3016) );
  OR2_X1 U3844 ( .A1(n3054), .A2(n3895), .ZN(n3829) );
  NAND2_X1 U3845 ( .A1(n3895), .A2(n3054), .ZN(n3827) );
  NAND2_X1 U3846 ( .A1(n3017), .A2(n3827), .ZN(n3368) );
  INV_X1 U3847 ( .A(n3368), .ZN(n3019) );
  INV_X1 U3848 ( .A(n3632), .ZN(n3020) );
  AND2_X1 U3849 ( .A1(n3894), .A2(n3020), .ZN(n3838) );
  INV_X1 U3850 ( .A(n3838), .ZN(n3018) );
  OR2_X1 U3851 ( .A1(n3020), .A2(n3894), .ZN(n3830) );
  NAND2_X1 U3852 ( .A1(n3677), .A2(n3021), .ZN(n3842) );
  NAND2_X1 U3853 ( .A1(n4321), .A2(n3531), .ZN(n3839) );
  NAND2_X1 U3854 ( .A1(n3892), .A2(n3427), .ZN(n4284) );
  INV_X1 U3855 ( .A(n3656), .ZN(n4298) );
  NAND2_X1 U3856 ( .A1(n4261), .A2(n4298), .ZN(n3022) );
  NAND2_X1 U3857 ( .A1(n4319), .A2(n3582), .ZN(n4283) );
  NAND2_X1 U3858 ( .A1(n4283), .A2(n3420), .ZN(n3024) );
  NOR2_X1 U3859 ( .A1(n4261), .A2(n4298), .ZN(n3023) );
  AOI21_X1 U3860 ( .B1(n3024), .B2(n2016), .A(n3023), .ZN(n3851) );
  INV_X1 U3861 ( .A(n4264), .ZN(n3599) );
  NAND2_X1 U3862 ( .A1(n3599), .A2(n3729), .ZN(n3740) );
  NAND2_X1 U3863 ( .A1(n4264), .A2(n4249), .ZN(n3739) );
  NAND2_X1 U3864 ( .A1(n3740), .A2(n3739), .ZN(n4246) );
  INV_X1 U3865 ( .A(n4239), .ZN(n3025) );
  INV_X1 U3866 ( .A(n4231), .ZN(n3776) );
  NAND2_X1 U3867 ( .A1(n4222), .A2(n3776), .ZN(n3026) );
  NAND2_X1 U3868 ( .A1(n4151), .A2(n4181), .ZN(n3027) );
  AND2_X1 U3869 ( .A1(n3027), .A2(n4172), .ZN(n3030) );
  INV_X1 U3870 ( .A(n4214), .ZN(n4207) );
  NAND2_X1 U3871 ( .A1(n4224), .A2(n4207), .ZN(n4167) );
  NAND2_X1 U3872 ( .A1(n3030), .A2(n4167), .ZN(n3855) );
  OR2_X1 U3873 ( .A1(n4224), .A2(n4207), .ZN(n4169) );
  NAND2_X1 U3874 ( .A1(n4171), .A2(n4169), .ZN(n3029) );
  NOR2_X1 U3875 ( .A1(n4151), .A2(n4181), .ZN(n3028) );
  AOI21_X1 U3876 ( .B1(n3030), .B2(n3029), .A(n3028), .ZN(n4146) );
  OR2_X1 U3877 ( .A1(n4177), .A2(n4160), .ZN(n3031) );
  AND2_X1 U3878 ( .A1(n4146), .A2(n3031), .ZN(n3743) );
  NAND2_X1 U3879 ( .A1(n4177), .A2(n4160), .ZN(n3859) );
  NAND2_X1 U3880 ( .A1(n4153), .A2(n3569), .ZN(n4096) );
  NAND2_X1 U3881 ( .A1(n4131), .A2(n3863), .ZN(n3034) );
  NAND2_X1 U3882 ( .A1(n3890), .A2(n4105), .ZN(n3788) );
  NAND2_X1 U3883 ( .A1(n3788), .A2(n3032), .ZN(n3862) );
  AND2_X1 U3884 ( .A1(n4118), .A2(n4138), .ZN(n4095) );
  AND2_X1 U3885 ( .A1(n4098), .A2(n4095), .ZN(n3033) );
  NOR2_X1 U3886 ( .A1(n3862), .A2(n3033), .ZN(n3746) );
  NAND2_X1 U3887 ( .A1(n4120), .A2(n3035), .ZN(n3789) );
  NOR2_X1 U3888 ( .A1(n4102), .A2(n4087), .ZN(n3801) );
  NAND2_X1 U3889 ( .A1(n4102), .A2(n4087), .ZN(n3800) );
  NAND2_X1 U3890 ( .A1(n4048), .A2(n3469), .ZN(n4043) );
  OAI21_X1 U3891 ( .B1(n4065), .B2(n4055), .A(n4043), .ZN(n3872) );
  NAND2_X1 U3892 ( .A1(n4065), .A2(n4055), .ZN(n3760) );
  INV_X1 U3893 ( .A(n4037), .ZN(n3501) );
  NAND2_X1 U3894 ( .A1(n3041), .A2(n3501), .ZN(n3763) );
  NAND2_X1 U3895 ( .A1(n3763), .A2(n3870), .ZN(n4031) );
  INV_X1 U3896 ( .A(n3763), .ZN(n3756) );
  XOR2_X1 U3897 ( .A(n4000), .B(n4008), .Z(n3038) );
  INV_X1 U3898 ( .A(n2408), .ZN(n4489) );
  NAND2_X1 U3899 ( .A1(n4489), .A2(n4488), .ZN(n3881) );
  NAND2_X1 U3900 ( .A1(n4490), .A2(n4487), .ZN(n3037) );
  OAI22_X1 U3901 ( .A1(n3041), .A2(n4320), .B1(n4289), .B2(n3040), .ZN(n3042)
         );
  NAND2_X1 U3902 ( .A1(n3044), .A2(n3487), .ZN(n3060) );
  OR2_X1 U3903 ( .A1(n3064), .A2(n3045), .ZN(n3050) );
  OAI21_X1 U3904 ( .B1(n3064), .B2(D_REG_1__SCAN_IN), .A(n3046), .ZN(n3049) );
  NAND2_X1 U3905 ( .A1(n4595), .A2(n3807), .ZN(n3048) );
  NAND4_X1 U3906 ( .A1(n3050), .A2(n3049), .A3(n3252), .A4(n3048), .ZN(n3059)
         );
  OR2_X1 U3907 ( .A1(n3060), .A2(n4334), .ZN(n3053) );
  INV_X1 U3908 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3909 ( .A1(n3053), .A2(n3052), .ZN(n3057) );
  NAND2_X1 U3910 ( .A1(n3360), .A2(n3054), .ZN(n3374) );
  INV_X1 U3911 ( .A(n3055), .ZN(n4159) );
  AND2_X2 U3912 ( .A1(n4068), .A2(n4055), .ZN(n4053) );
  NAND2_X1 U3913 ( .A1(n4036), .A2(n4001), .ZN(n3056) );
  NAND2_X1 U3914 ( .A1(n4021), .A2(n3056), .ZN(n3480) );
  NAND2_X1 U3915 ( .A1(n3057), .A2(n2350), .ZN(U3546) );
  OR2_X1 U3916 ( .A1(n3060), .A2(n4610), .ZN(n3061) );
  NAND2_X1 U3917 ( .A1(n3061), .A2(n2344), .ZN(n3062) );
  NAND2_X1 U3918 ( .A1(n3062), .A2(n2349), .ZN(U3514) );
  OR2_X2 U3919 ( .A1(n2421), .A2(n4574), .ZN(n3907) );
  NAND2_X1 U3920 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3063) );
  OAI21_X1 U3921 ( .B1(n2891), .B2(U3149), .A(n3063), .ZN(U3327) );
  INV_X1 U3922 ( .A(D_REG_0__SCAN_IN), .ZN(n3066) );
  NOR3_X1 U3923 ( .A1(n2894), .A2(n4486), .A3(n4574), .ZN(n3065) );
  AOI21_X1 U3924 ( .B1(n4573), .B2(n3066), .A(n3065), .ZN(U3458) );
  INV_X1 U3925 ( .A(D_REG_1__SCAN_IN), .ZN(n4755) );
  AOI22_X1 U3926 ( .A1(n4573), .A2(n4755), .B1(n3068), .B2(n3067), .ZN(U3459)
         );
  NOR2_X1 U3927 ( .A1(n3069), .A2(U3149), .ZN(n3884) );
  NAND2_X1 U3928 ( .A1(n3070), .A2(n3069), .ZN(n3071) );
  INV_X1 U3929 ( .A(n3086), .ZN(n3072) );
  NOR2_X1 U3930 ( .A1(n4527), .A2(U4043), .ZN(U3148) );
  INV_X1 U3931 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4740) );
  NAND2_X1 U3932 ( .A1(n4243), .A2(U4043), .ZN(n3073) );
  OAI21_X1 U3933 ( .B1(U4043), .B2(n4740), .A(n3073), .ZN(U3566) );
  INV_X1 U3934 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U3935 ( .A1(n3677), .A2(U4043), .ZN(n3074) );
  OAI21_X1 U3936 ( .B1(U4043), .B2(n4704), .A(n3074), .ZN(U3560) );
  INV_X1 U3937 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U3938 ( .A1(n2058), .A2(U4043), .ZN(n3075) );
  OAI21_X1 U3939 ( .B1(U4043), .B2(n4703), .A(n3075), .ZN(U3551) );
  INV_X1 U3940 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4739) );
  INV_X1 U3941 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3078) );
  NAND2_X1 U3942 ( .A1(n3750), .A2(REG1_REG_31__SCAN_IN), .ZN(n3077) );
  INV_X1 U3943 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4420) );
  OR2_X1 U3944 ( .A1(n3751), .A2(n4420), .ZN(n3076) );
  OAI211_X1 U3945 ( .C1(n2680), .C2(n3078), .A(n3077), .B(n3076), .ZN(n3986)
         );
  NAND2_X1 U3946 ( .A1(n3986), .A2(U4043), .ZN(n3079) );
  OAI21_X1 U3947 ( .B1(U4043), .B2(n4739), .A(n3079), .ZN(U3581) );
  XNOR2_X1 U3948 ( .A(n3912), .B(REG1_REG_2__SCAN_IN), .ZN(n3909) );
  AND2_X1 U3949 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3435)
         );
  NAND2_X1 U3950 ( .A1(n3434), .A2(n3435), .ZN(n3081) );
  NAND2_X1 U3951 ( .A1(n2198), .A2(REG1_REG_1__SCAN_IN), .ZN(n3080) );
  NAND2_X1 U3952 ( .A1(n3081), .A2(n3080), .ZN(n3910) );
  INV_X1 U3953 ( .A(n3912), .ZN(n4501) );
  AOI22_X1 U3954 ( .A1(n3909), .A2(n3910), .B1(n4501), .B2(REG1_REG_2__SCAN_IN), .ZN(n3082) );
  INV_X1 U3955 ( .A(n3082), .ZN(n3083) );
  INV_X1 U3956 ( .A(n3084), .ZN(n3085) );
  MUX2_X1 U3957 ( .A(n2493), .B(REG1_REG_5__SCAN_IN), .S(n4499), .Z(n3130) );
  XNOR2_X1 U3958 ( .A(n3112), .B(REG1_REG_6__SCAN_IN), .ZN(n3103) );
  XNOR2_X1 U3959 ( .A(n3088), .B(IR_REG_27__SCAN_IN), .ZN(n4485) );
  NOR2_X2 U3960 ( .A1(n3125), .A2(n4485), .ZN(n4535) );
  AND2_X1 U3961 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3701) );
  INV_X1 U3962 ( .A(n4527), .ZN(n4554) );
  INV_X1 U3963 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4679) );
  NOR2_X1 U3964 ( .A1(n4554), .A2(n4679), .ZN(n3089) );
  AOI211_X1 U3965 ( .C1(n4548), .C2(n4498), .A(n3701), .B(n3089), .ZN(n3102)
         );
  MUX2_X1 U3966 ( .A(n3090), .B(REG2_REG_2__SCAN_IN), .S(n2103), .Z(n3092) );
  AND2_X1 U3967 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3436)
         );
  NAND2_X1 U3968 ( .A1(n4501), .A2(REG2_REG_2__SCAN_IN), .ZN(n3093) );
  INV_X1 U3969 ( .A(n4500), .ZN(n3107) );
  NAND2_X1 U3970 ( .A1(n3094), .A2(n4500), .ZN(n3095) );
  MUX2_X1 U3971 ( .A(n3298), .B(REG2_REG_5__SCAN_IN), .S(n4499), .Z(n3133) );
  XOR2_X1 U3972 ( .A(REG2_REG_6__SCAN_IN), .B(n3114), .Z(n3100) );
  NAND2_X1 U3973 ( .A1(n4485), .A2(n4484), .ZN(n3099) );
  NAND2_X1 U3974 ( .A1(n3100), .A2(n4537), .ZN(n3101) );
  OAI211_X1 U3975 ( .C1(n3103), .C2(n4546), .A(n3102), .B(n3101), .ZN(U3246)
         );
  XNOR2_X1 U3976 ( .A(n3104), .B(REG1_REG_3__SCAN_IN), .ZN(n3111) );
  INV_X1 U3977 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3289) );
  XNOR2_X1 U3978 ( .A(n3105), .B(n3289), .ZN(n3109) );
  AOI22_X1 U3979 ( .A1(n4527), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3106) );
  OAI21_X1 U3980 ( .B1(n4540), .B2(n3107), .A(n3106), .ZN(n3108) );
  AOI21_X1 U3981 ( .B1(n4537), .B2(n3109), .A(n3108), .ZN(n3110) );
  OAI21_X1 U3982 ( .B1(n3111), .B2(n4546), .A(n3110), .ZN(U3243) );
  XNOR2_X1 U3983 ( .A(n3144), .B(n2530), .ZN(n3113) );
  XNOR2_X1 U3984 ( .A(n2049), .B(n3113), .ZN(n3120) );
  MUX2_X1 U3985 ( .A(REG2_REG_7__SCAN_IN), .B(n2534), .S(n3144), .Z(n3115) );
  AOI21_X1 U3986 ( .B1(n2057), .B2(n3115), .A(n4541), .ZN(n3118) );
  AND2_X1 U3987 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3491) );
  AOI21_X1 U3988 ( .B1(n4527), .B2(ADDR_REG_7__SCAN_IN), .A(n3491), .ZN(n3116)
         );
  OAI21_X1 U3989 ( .B1(n4540), .B2(n3144), .A(n3116), .ZN(n3117) );
  AOI21_X1 U3990 ( .B1(n3118), .B2(n3142), .A(n3117), .ZN(n3119) );
  OAI21_X1 U3991 ( .B1(n3120), .B2(n4546), .A(n3119), .ZN(U3247) );
  OAI21_X1 U3992 ( .B1(n4485), .B2(REG1_REG_0__SCAN_IN), .A(n4627), .ZN(n3122)
         );
  INV_X1 U3993 ( .A(n4485), .ZN(n3121) );
  OAI21_X1 U3994 ( .B1(n3121), .B2(REG2_REG_0__SCAN_IN), .A(n4484), .ZN(n3908)
         );
  MUX2_X1 U3995 ( .A(n3122), .B(n4627), .S(n3908), .Z(n3124) );
  OAI22_X1 U3996 ( .A1(n3125), .A2(n3124), .B1(STATE_REG_SCAN_IN), .B2(n3123), 
        .ZN(n3127) );
  NOR3_X1 U3997 ( .A1(n4546), .A2(REG1_REG_0__SCAN_IN), .A3(n4627), .ZN(n3126)
         );
  AOI211_X1 U3998 ( .C1(n4527), .C2(ADDR_REG_0__SCAN_IN), .A(n3127), .B(n3126), 
        .ZN(n3128) );
  INV_X1 U3999 ( .A(n3128), .ZN(U3240) );
  AOI211_X1 U4000 ( .C1(n3131), .C2(n3130), .A(n3129), .B(n4546), .ZN(n3139)
         );
  AOI211_X1 U4001 ( .C1(n3134), .C2(n3133), .A(n3132), .B(n4541), .ZN(n3138)
         );
  INV_X1 U4002 ( .A(n4499), .ZN(n3136) );
  NOR2_X1 U4003 ( .A1(STATE_REG_SCAN_IN), .A2(n4634), .ZN(n3320) );
  AOI21_X1 U4004 ( .B1(n4527), .B2(ADDR_REG_5__SCAN_IN), .A(n3320), .ZN(n3135)
         );
  OAI21_X1 U4005 ( .B1(n4540), .B2(n3136), .A(n3135), .ZN(n3137) );
  OR3_X1 U4006 ( .A1(n3139), .A2(n3138), .A3(n3137), .ZN(U3245) );
  INV_X1 U4007 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4756) );
  NAND2_X1 U4008 ( .A1(n4151), .A2(U4043), .ZN(n3140) );
  OAI21_X1 U4009 ( .B1(U4043), .B2(n4756), .A(n3140), .ZN(U3569) );
  XNOR2_X1 U4010 ( .A(n3153), .B(REG2_REG_8__SCAN_IN), .ZN(n3148) );
  AND2_X1 U4011 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n3556) );
  INV_X1 U4012 ( .A(n4497), .ZN(n3156) );
  NOR2_X1 U4013 ( .A1(n4540), .A2(n3156), .ZN(n3143) );
  AOI211_X1 U4014 ( .C1(n4527), .C2(ADDR_REG_8__SCAN_IN), .A(n3556), .B(n3143), 
        .ZN(n3147) );
  OAI211_X1 U4015 ( .C1(n3145), .C2(REG1_REG_8__SCAN_IN), .A(n3159), .B(n4535), 
        .ZN(n3146) );
  OAI211_X1 U4016 ( .C1(n3148), .C2(n4541), .A(n3147), .B(n3146), .ZN(U3248)
         );
  NAND2_X1 U4017 ( .A1(n2064), .A2(n3224), .ZN(n3811) );
  NAND2_X1 U4018 ( .A1(n3809), .A2(n3811), .ZN(n4567) );
  NOR2_X1 U4019 ( .A1(n3224), .A2(n3149), .ZN(n4565) );
  INV_X1 U4020 ( .A(n2058), .ZN(n3223) );
  INV_X1 U4021 ( .A(n4293), .ZN(n4318) );
  INV_X1 U4022 ( .A(n4322), .ZN(n3208) );
  OAI21_X1 U4023 ( .B1(n3208), .B2(n4268), .A(n4567), .ZN(n3150) );
  OAI21_X1 U4024 ( .B1(n3223), .B2(n4318), .A(n3150), .ZN(n4563) );
  AOI211_X1 U4025 ( .C1(n4595), .C2(n4567), .A(n4565), .B(n4563), .ZN(n4584)
         );
  NAND2_X1 U4026 ( .A1(n4334), .A2(REG1_REG_0__SCAN_IN), .ZN(n3151) );
  OAI21_X1 U4027 ( .B1(n4584), .B2(n4334), .A(n3151), .ZN(U3518) );
  XNOR2_X1 U4028 ( .A(n4496), .B(REG2_REG_9__SCAN_IN), .ZN(n3229) );
  XNOR2_X1 U4029 ( .A(n3230), .B(n3229), .ZN(n3164) );
  AND2_X1 U4030 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3631) );
  INV_X1 U4031 ( .A(n4496), .ZN(n3232) );
  NOR2_X1 U4032 ( .A1(n4540), .A2(n3232), .ZN(n3154) );
  AOI211_X1 U4033 ( .C1(n4527), .C2(ADDR_REG_9__SCAN_IN), .A(n3631), .B(n3154), 
        .ZN(n3163) );
  XNOR2_X1 U4034 ( .A(n3232), .B(REG1_REG_9__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U4035 ( .A1(n3161), .A2(n3160), .ZN(n3233) );
  OAI211_X1 U4036 ( .C1(n3161), .C2(n3160), .A(n3233), .B(n4535), .ZN(n3162)
         );
  OAI211_X1 U4037 ( .C1(n3164), .C2(n4541), .A(n3163), .B(n3162), .ZN(U3249)
         );
  AOI21_X1 U4038 ( .B1(n3008), .B2(n2956), .A(n3211), .ZN(n3261) );
  OAI21_X1 U4039 ( .B1(n3778), .B2(n3166), .A(n3165), .ZN(n3257) );
  NOR2_X1 U4040 ( .A1(n3257), .A2(n4586), .ZN(n3174) );
  NAND2_X1 U4041 ( .A1(n2064), .A2(n4223), .ZN(n3168) );
  NAND2_X1 U4042 ( .A1(n2436), .A2(n4293), .ZN(n3167) );
  OAI211_X1 U40430 ( .C1(n3169), .C2(n4289), .A(n3168), .B(n3167), .ZN(n3170)
         );
  INV_X1 U4044 ( .A(n3170), .ZN(n3173) );
  XNOR2_X1 U4045 ( .A(n3778), .B(n3809), .ZN(n3171) );
  NAND2_X1 U4046 ( .A1(n3171), .A2(n4268), .ZN(n3172) );
  OAI211_X1 U4047 ( .C1(n3257), .C2(n4322), .A(n3173), .B(n3172), .ZN(n3258)
         );
  AOI211_X1 U4048 ( .C1(n4602), .C2(n3261), .A(n3174), .B(n3258), .ZN(n4585)
         );
  NAND2_X1 U4049 ( .A1(n4334), .A2(REG1_REG_1__SCAN_IN), .ZN(n3175) );
  OAI21_X1 U4050 ( .B1(n4585), .B2(n4334), .A(n3175), .ZN(U3519) );
  INV_X1 U4051 ( .A(n3176), .ZN(n3180) );
  INV_X1 U4052 ( .A(n3177), .ZN(n3178) );
  NOR3_X1 U4053 ( .A1(n3180), .A2(n3179), .A3(n3178), .ZN(n3222) );
  OAI22_X1 U4054 ( .A1(n3181), .A2(n3716), .B1(n3689), .B2(n2955), .ZN(n3182)
         );
  AOI21_X1 U4055 ( .B1(n2956), .B2(n3730), .A(n3182), .ZN(n3188) );
  AOI21_X1 U4056 ( .B1(n3183), .B2(n3184), .A(n3719), .ZN(n3186) );
  NAND2_X1 U4057 ( .A1(n3186), .A2(n3185), .ZN(n3187) );
  OAI211_X1 U4058 ( .C1(n3222), .C2(n3256), .A(n3188), .B(n3187), .ZN(U3219)
         );
  OAI21_X1 U4059 ( .B1(n3191), .B2(n3190), .A(n3189), .ZN(n3192) );
  NAND2_X1 U4060 ( .A1(n3192), .A2(n3726), .ZN(n3195) );
  OAI22_X1 U4061 ( .A1(n3446), .A2(n3689), .B1(n3716), .B2(n3223), .ZN(n3193)
         );
  AOI21_X1 U4062 ( .B1(n3203), .B2(n3730), .A(n3193), .ZN(n3194) );
  OAI211_X1 U4063 ( .C1(n3222), .C2(n3196), .A(n3195), .B(n3194), .ZN(U3234)
         );
  AND2_X1 U4064 ( .A1(n3165), .A2(n3197), .ZN(n3199) );
  NAND2_X1 U4065 ( .A1(n3199), .A2(n3198), .ZN(n3281) );
  OAI21_X1 U4066 ( .B1(n3199), .B2(n3198), .A(n3281), .ZN(n4558) );
  INV_X1 U4067 ( .A(n4558), .ZN(n3209) );
  OAI21_X1 U4068 ( .B1(n3779), .B2(n3201), .A(n3200), .ZN(n3202) );
  NAND2_X1 U4069 ( .A1(n3202), .A2(n4268), .ZN(n3206) );
  AOI22_X1 U4070 ( .A1(n4223), .A2(n2058), .B1(n3203), .B2(n4326), .ZN(n3205)
         );
  OAI211_X1 U4071 ( .C1(n3446), .C2(n4318), .A(n3206), .B(n3205), .ZN(n3207)
         );
  AOI21_X1 U4072 ( .B1(n3208), .B2(n4558), .A(n3207), .ZN(n4561) );
  OAI21_X1 U4073 ( .B1(n3209), .B2(n4586), .A(n4561), .ZN(n3305) );
  OAI21_X1 U4074 ( .B1(n3211), .B2(n2954), .A(n3210), .ZN(n4555) );
  OAI22_X1 U4075 ( .A1(n4480), .A2(n4555), .B1(n4612), .B2(n2434), .ZN(n3212)
         );
  AOI21_X1 U4076 ( .B1(n3305), .B2(n4612), .A(n3212), .ZN(n3213) );
  INV_X1 U4077 ( .A(n3213), .ZN(U3471) );
  XOR2_X1 U4078 ( .A(n3215), .B(n3214), .Z(n3219) );
  INV_X1 U4079 ( .A(n3899), .ZN(n3318) );
  OAI22_X1 U4080 ( .A1(n2955), .A2(n3716), .B1(n3689), .B2(n3318), .ZN(n3217)
         );
  MUX2_X1 U4081 ( .A(n3733), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3216) );
  AOI211_X1 U4082 ( .C1(n3288), .C2(n3730), .A(n3217), .B(n3216), .ZN(n3218)
         );
  OAI21_X1 U4083 ( .B1(n3219), .B2(n3719), .A(n3218), .ZN(U3215) );
  XNOR2_X1 U4084 ( .A(n3221), .B(n3220), .ZN(n3902) );
  INV_X1 U4085 ( .A(n3222), .ZN(n3226) );
  INV_X1 U4086 ( .A(n3730), .ZN(n3666) );
  OAI22_X1 U4087 ( .A1(n3666), .A2(n3224), .B1(n3223), .B2(n3689), .ZN(n3225)
         );
  AOI21_X1 U4088 ( .B1(n3226), .B2(REG3_REG_0__SCAN_IN), .A(n3225), .ZN(n3227)
         );
  OAI21_X1 U4089 ( .B1(n3719), .B2(n3902), .A(n3227), .ZN(U3229) );
  XNOR2_X1 U4090 ( .A(n3329), .B(REG2_REG_10__SCAN_IN), .ZN(n3240) );
  INV_X1 U4091 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3231) );
  INV_X1 U4092 ( .A(n3326), .ZN(n3234) );
  OAI211_X1 U4093 ( .C1(REG1_REG_10__SCAN_IN), .C2(n3235), .A(n3234), .B(n4535), .ZN(n3239) );
  AND2_X1 U4094 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3530) );
  NOR2_X1 U4095 ( .A1(n4540), .A2(n3236), .ZN(n3237) );
  AOI211_X1 U4096 ( .C1(n4527), .C2(ADDR_REG_10__SCAN_IN), .A(n3530), .B(n3237), .ZN(n3238) );
  OAI211_X1 U4097 ( .C1(n3240), .C2(n4541), .A(n3239), .B(n3238), .ZN(U3250)
         );
  INV_X1 U4098 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U4099 ( .A1(n4102), .A2(U4043), .ZN(n3241) );
  OAI21_X1 U4100 ( .B1(U4043), .B2(n4752), .A(n3241), .ZN(U3574) );
  AOI21_X1 U4101 ( .B1(n3242), .B2(n3243), .A(n3719), .ZN(n3245) );
  NAND2_X1 U4102 ( .A1(n3245), .A2(n3244), .ZN(n3250) );
  NAND2_X1 U4103 ( .A1(n3730), .A2(n2317), .ZN(n3246) );
  OAI21_X1 U4104 ( .B1(n3446), .B2(n3716), .A(n3246), .ZN(n3248) );
  NAND2_X1 U4105 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3925) );
  OAI21_X1 U4106 ( .B1(n3689), .B2(n2967), .A(n3925), .ZN(n3247) );
  NOR2_X1 U4107 ( .A1(n3248), .A2(n3247), .ZN(n3249) );
  OAI211_X1 U4108 ( .C1(n3695), .C2(n3454), .A(n3250), .B(n3249), .ZN(U3227)
         );
  NAND3_X1 U4109 ( .A1(n3253), .A2(n3252), .A3(n3251), .ZN(n3254) );
  NAND2_X1 U4110 ( .A1(n4570), .A2(n3979), .ZN(n3340) );
  OR2_X1 U4111 ( .A1(n2402), .A2(n3979), .ZN(n3272) );
  INV_X1 U4112 ( .A(n3272), .ZN(n3255) );
  OAI22_X1 U4113 ( .A1(n4306), .A2(n3257), .B1(n3256), .B2(n4313), .ZN(n3260)
         );
  MUX2_X1 U4114 ( .A(n3258), .B(REG2_REG_1__SCAN_IN), .S(n4276), .Z(n3259) );
  AOI211_X1 U4115 ( .C1(n4557), .C2(n3261), .A(n3260), .B(n3259), .ZN(n3262)
         );
  INV_X1 U4116 ( .A(n3262), .ZN(U3289) );
  AND2_X1 U4117 ( .A1(n3014), .A2(n3824), .ZN(n3792) );
  XNOR2_X1 U4118 ( .A(n3263), .B(n3792), .ZN(n3266) );
  AOI22_X1 U4119 ( .A1(n3896), .A2(n4293), .B1(n4326), .B2(n3702), .ZN(n3265)
         );
  NAND2_X1 U4120 ( .A1(n3898), .A2(n4223), .ZN(n3264) );
  OAI211_X1 U4121 ( .C1(n3266), .C2(n4330), .A(n3265), .B(n3264), .ZN(n3307)
         );
  INV_X1 U4122 ( .A(n3307), .ZN(n3278) );
  NAND2_X1 U4123 ( .A1(n3293), .A2(n3268), .ZN(n3271) );
  INV_X1 U4124 ( .A(n3269), .ZN(n3270) );
  NAND2_X1 U4125 ( .A1(n3271), .A2(n3270), .ZN(n3344) );
  XNOR2_X1 U4126 ( .A(n3344), .B(n3792), .ZN(n3308) );
  NAND2_X1 U4127 ( .A1(n4322), .A2(n3272), .ZN(n3273) );
  OAI21_X1 U4128 ( .B1(n2048), .B2(n2968), .A(n3341), .ZN(n3311) );
  INV_X1 U4129 ( .A(n3274), .ZN(n3703) );
  AOI22_X1 U4130 ( .A1(n4276), .A2(REG2_REG_6__SCAN_IN), .B1(n3703), .B2(n4566), .ZN(n3275) );
  OAI21_X1 U4131 ( .B1(n3311), .B2(n4315), .A(n3275), .ZN(n3276) );
  AOI21_X1 U4132 ( .B1(n3308), .B2(n4255), .A(n3276), .ZN(n3277) );
  OAI21_X1 U4133 ( .B1(n3278), .B2(n4280), .A(n3277), .ZN(U3284) );
  INV_X1 U4134 ( .A(n3279), .ZN(n3280) );
  NAND2_X1 U4135 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  XNOR2_X1 U4136 ( .A(n3282), .B(n3782), .ZN(n4587) );
  XNOR2_X1 U4137 ( .A(n3283), .B(n3782), .ZN(n3286) );
  AOI22_X1 U4138 ( .A1(n3899), .A2(n4293), .B1(n4326), .B2(n3288), .ZN(n3284)
         );
  OAI21_X1 U4139 ( .B1(n2955), .B2(n4320), .A(n3284), .ZN(n3285) );
  AOI21_X1 U4140 ( .B1(n3286), .B2(n4268), .A(n3285), .ZN(n3287) );
  OAI21_X1 U4141 ( .B1(n4587), .B2(n4322), .A(n3287), .ZN(n4588) );
  NAND2_X1 U4142 ( .A1(n4588), .A2(n4570), .ZN(n3292) );
  AOI21_X1 U4143 ( .B1(n3288), .B2(n3210), .A(n3453), .ZN(n4590) );
  OAI22_X1 U4144 ( .A1(n4570), .A2(n3289), .B1(REG3_REG_3__SCAN_IN), .B2(n4313), .ZN(n3290) );
  AOI21_X1 U4145 ( .B1(n4590), .B2(n4557), .A(n3290), .ZN(n3291) );
  OAI211_X1 U4146 ( .C1(n4587), .C2(n4306), .A(n3292), .B(n3291), .ZN(U3287)
         );
  AND2_X1 U4147 ( .A1(n3835), .A2(n3821), .ZN(n3785) );
  XOR2_X1 U4148 ( .A(n3293), .B(n3785), .Z(n4597) );
  XOR2_X1 U4149 ( .A(n3294), .B(n3785), .Z(n3297) );
  AOI22_X1 U4150 ( .A1(n3897), .A2(n4293), .B1(n4326), .B2(n3299), .ZN(n3295)
         );
  OAI21_X1 U4151 ( .B1(n3318), .B2(n4320), .A(n3295), .ZN(n3296) );
  AOI21_X1 U4152 ( .B1(n3297), .B2(n4268), .A(n3296), .ZN(n4598) );
  MUX2_X1 U4153 ( .A(n4598), .B(n3298), .S(n4276), .Z(n3302) );
  AOI21_X1 U4154 ( .B1(n3299), .B2(n3451), .A(n2048), .ZN(n4601) );
  INV_X1 U4155 ( .A(n3323), .ZN(n3300) );
  AOI22_X1 U4156 ( .A1(n4601), .A2(n4557), .B1(n3300), .B2(n4566), .ZN(n3301)
         );
  OAI211_X1 U4157 ( .C1(n4143), .C2(n4597), .A(n3302), .B(n3301), .ZN(U3285)
         );
  INV_X1 U4158 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3303) );
  OAI22_X1 U4159 ( .A1(n4419), .A2(n4555), .B1(n4416), .B2(n3303), .ZN(n3304)
         );
  AOI21_X1 U4160 ( .B1(n3305), .B2(n4416), .A(n3304), .ZN(n3306) );
  INV_X1 U4161 ( .A(n3306), .ZN(U3520) );
  AOI21_X1 U4162 ( .B1(n3308), .B2(n4411), .A(n3307), .ZN(n3314) );
  OAI22_X1 U4163 ( .A1(n3311), .A2(n4419), .B1(n4416), .B2(n2207), .ZN(n3309)
         );
  INV_X1 U4164 ( .A(n3309), .ZN(n3310) );
  OAI21_X1 U4165 ( .B1(n3314), .B2(n4334), .A(n3310), .ZN(U3524) );
  OAI22_X1 U4166 ( .A1(n3311), .A2(n4480), .B1(n4612), .B2(n2511), .ZN(n3312)
         );
  INV_X1 U4167 ( .A(n3312), .ZN(n3313) );
  OAI21_X1 U4168 ( .B1(n3314), .B2(n4610), .A(n3313), .ZN(U3479) );
  OAI211_X1 U4169 ( .C1(n3317), .C2(n3316), .A(n3315), .B(n3726), .ZN(n3322)
         );
  OAI22_X1 U4170 ( .A1(n3666), .A2(n2966), .B1(n3318), .B2(n3716), .ZN(n3319)
         );
  AOI211_X1 U4171 ( .C1(n3731), .C2(n3897), .A(n3320), .B(n3319), .ZN(n3321)
         );
  OAI211_X1 U4172 ( .C1(n3695), .C2(n3323), .A(n3322), .B(n3321), .ZN(U3224)
         );
  INV_X1 U4173 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4417) );
  XNOR2_X1 U4174 ( .A(n3395), .B(n4417), .ZN(n3327) );
  AOI211_X1 U4175 ( .C1(n3328), .C2(n3327), .A(n4546), .B(n3398), .ZN(n3335)
         );
  MUX2_X1 U4176 ( .A(REG2_REG_11__SCAN_IN), .B(n2613), .S(n3395), .Z(n3330) );
  AOI211_X1 U4177 ( .C1(n3331), .C2(n3330), .A(n4541), .B(n3396), .ZN(n3334)
         );
  AND2_X1 U4178 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3676) );
  AOI21_X1 U4179 ( .B1(n4527), .B2(ADDR_REG_11__SCAN_IN), .A(n3676), .ZN(n3332) );
  OAI21_X1 U4180 ( .B1(n4540), .B2(n3395), .A(n3332), .ZN(n3333) );
  OR3_X1 U4181 ( .A1(n3335), .A2(n3334), .A3(n3333), .ZN(U3251) );
  XNOR2_X1 U4182 ( .A(n3336), .B(n3790), .ZN(n3339) );
  AOI22_X1 U4183 ( .A1(n4223), .A2(n3897), .B1(n3492), .B2(n4326), .ZN(n3338)
         );
  NAND2_X1 U4184 ( .A1(n3895), .A2(n4293), .ZN(n3337) );
  OAI211_X1 U4185 ( .C1(n3339), .C2(n4330), .A(n3338), .B(n3337), .ZN(n4606)
         );
  INV_X1 U4186 ( .A(n4606), .ZN(n3353) );
  INV_X1 U4187 ( .A(n3340), .ZN(n4200) );
  NAND2_X1 U4188 ( .A1(n3341), .A2(n3492), .ZN(n3342) );
  NAND2_X1 U4189 ( .A1(n3342), .A2(n4602), .ZN(n3343) );
  NOR2_X1 U4190 ( .A1(n3360), .A2(n3343), .ZN(n4607) );
  OAI22_X1 U4191 ( .A1(n4570), .A2(n2534), .B1(n3493), .B2(n4313), .ZN(n3351)
         );
  INV_X1 U4192 ( .A(n3344), .ZN(n3347) );
  INV_X1 U4193 ( .A(n3897), .ZN(n3346) );
  AOI21_X1 U4194 ( .B1(n3344), .B2(n3897), .A(n3702), .ZN(n3345) );
  AOI21_X1 U4195 ( .B1(n3347), .B2(n3346), .A(n3345), .ZN(n3348) );
  NOR2_X1 U4196 ( .A1(n3348), .A2(n3790), .ZN(n4605) );
  NAND2_X1 U4197 ( .A1(n3348), .A2(n3790), .ZN(n4608) );
  INV_X1 U4198 ( .A(n4608), .ZN(n3349) );
  NOR3_X1 U4199 ( .A1(n4605), .A2(n3349), .A3(n4143), .ZN(n3350) );
  AOI211_X1 U4200 ( .C1(n4200), .C2(n4607), .A(n3351), .B(n3350), .ZN(n3352)
         );
  OAI21_X1 U4201 ( .B1(n4276), .B2(n3353), .A(n3352), .ZN(U3283) );
  AND2_X1 U4202 ( .A1(n3829), .A2(n3827), .ZN(n3791) );
  XNOR2_X1 U4203 ( .A(n3355), .B(n3791), .ZN(n3383) );
  INV_X1 U4204 ( .A(n3383), .ZN(n3367) );
  XNOR2_X1 U4205 ( .A(n3356), .B(n3791), .ZN(n3359) );
  AOI22_X1 U4206 ( .A1(n3894), .A2(n4293), .B1(n4326), .B2(n3557), .ZN(n3358)
         );
  NAND2_X1 U4207 ( .A1(n3896), .A2(n4223), .ZN(n3357) );
  OAI211_X1 U4208 ( .C1(n3359), .C2(n4330), .A(n3358), .B(n3357), .ZN(n3382)
         );
  NAND2_X1 U4209 ( .A1(n3382), .A2(n4570), .ZN(n3366) );
  INV_X1 U4210 ( .A(n3360), .ZN(n3362) );
  INV_X1 U4211 ( .A(n3374), .ZN(n3361) );
  AOI21_X1 U4212 ( .B1(n3557), .B2(n3362), .A(n3361), .ZN(n3385) );
  OAI22_X1 U4213 ( .A1(n4570), .A2(n3363), .B1(n3558), .B2(n4313), .ZN(n3364)
         );
  AOI21_X1 U4214 ( .B1(n3385), .B2(n4557), .A(n3364), .ZN(n3365) );
  OAI211_X1 U4215 ( .C1(n4143), .C2(n3367), .A(n3366), .B(n3365), .ZN(U3282)
         );
  AND2_X1 U4216 ( .A1(n3018), .A2(n3830), .ZN(n3793) );
  XNOR2_X1 U4217 ( .A(n3368), .B(n3793), .ZN(n3371) );
  AOI22_X1 U4218 ( .A1(n3677), .A2(n4293), .B1(n4326), .B2(n3632), .ZN(n3370)
         );
  NAND2_X1 U4219 ( .A1(n3895), .A2(n4223), .ZN(n3369) );
  OAI211_X1 U4220 ( .C1(n3371), .C2(n4330), .A(n3370), .B(n3369), .ZN(n3388)
         );
  INV_X1 U4221 ( .A(n3388), .ZN(n3381) );
  XNOR2_X1 U4222 ( .A(n3373), .B(n3793), .ZN(n3389) );
  NAND2_X1 U4223 ( .A1(n3374), .A2(n3632), .ZN(n3375) );
  AND2_X1 U4224 ( .A1(n2353), .A2(n3375), .ZN(n3391) );
  INV_X1 U4225 ( .A(n3391), .ZN(n3378) );
  INV_X1 U4226 ( .A(n3376), .ZN(n3633) );
  AOI22_X1 U4227 ( .A1(n4276), .A2(REG2_REG_9__SCAN_IN), .B1(n3633), .B2(n4566), .ZN(n3377) );
  OAI21_X1 U4228 ( .B1(n3378), .B2(n4315), .A(n3377), .ZN(n3379) );
  AOI21_X1 U4229 ( .B1(n4255), .B2(n3389), .A(n3379), .ZN(n3380) );
  OAI21_X1 U4230 ( .B1(n3381), .B2(n4276), .A(n3380), .ZN(U3281) );
  AOI21_X1 U4231 ( .B1(n3383), .B2(n4411), .A(n3382), .ZN(n3387) );
  INV_X1 U4232 ( .A(n4419), .ZN(n4337) );
  AOI22_X1 U4233 ( .A1(n3385), .A2(n4337), .B1(REG1_REG_8__SCAN_IN), .B2(n4334), .ZN(n3384) );
  OAI21_X1 U4234 ( .B1(n3387), .B2(n4334), .A(n3384), .ZN(U3526) );
  INV_X1 U4235 ( .A(n4480), .ZN(n4425) );
  AOI22_X1 U4236 ( .A1(n3385), .A2(n4425), .B1(REG0_REG_8__SCAN_IN), .B2(n4610), .ZN(n3386) );
  OAI21_X1 U4237 ( .B1(n3387), .B2(n4610), .A(n3386), .ZN(U3483) );
  AOI21_X1 U4238 ( .B1(n3389), .B2(n4411), .A(n3388), .ZN(n3393) );
  AOI22_X1 U4239 ( .A1(n3391), .A2(n4425), .B1(REG0_REG_9__SCAN_IN), .B2(n4610), .ZN(n3390) );
  OAI21_X1 U4240 ( .B1(n3393), .B2(n4610), .A(n3390), .ZN(U3485) );
  AOI22_X1 U4241 ( .A1(n3391), .A2(n4337), .B1(REG1_REG_9__SCAN_IN), .B2(n4334), .ZN(n3392) );
  OAI21_X1 U4242 ( .B1(n3393), .B2(n4334), .A(n3392), .ZN(U3527) );
  INV_X1 U4243 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U4244 ( .A1(n4035), .A2(U4043), .ZN(n3394) );
  OAI21_X1 U4245 ( .B1(n4702), .B2(U4043), .A(n3394), .ZN(U3578) );
  INV_X1 U4246 ( .A(n3395), .ZN(n4494) );
  XOR2_X1 U4247 ( .A(REG2_REG_12__SCAN_IN), .B(n3936), .Z(n3402) );
  AND2_X1 U4248 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3581) );
  NOR2_X1 U4249 ( .A1(n4540), .A2(n2089), .ZN(n3397) );
  AOI211_X1 U4250 ( .C1(n4527), .C2(ADDR_REG_12__SCAN_IN), .A(n3581), .B(n3397), .ZN(n3401) );
  OAI211_X1 U4251 ( .C1(n3399), .C2(REG1_REG_12__SCAN_IN), .A(n3938), .B(n4535), .ZN(n3400) );
  OAI211_X1 U4252 ( .C1(n3402), .C2(n4541), .A(n3401), .B(n3400), .ZN(U3252)
         );
  AND2_X1 U4253 ( .A1(n3839), .A2(n3842), .ZN(n3784) );
  INV_X1 U4254 ( .A(n3784), .ZN(n3404) );
  XNOR2_X1 U4255 ( .A(n3403), .B(n3404), .ZN(n3415) );
  INV_X1 U4256 ( .A(n3415), .ZN(n3413) );
  XOR2_X1 U4257 ( .A(n3784), .B(n3405), .Z(n3408) );
  AOI22_X1 U4258 ( .A1(n3894), .A2(n4223), .B1(n4326), .B2(n3531), .ZN(n3407)
         );
  NAND2_X1 U4259 ( .A1(n3893), .A2(n4293), .ZN(n3406) );
  OAI211_X1 U4260 ( .C1(n3408), .C2(n4330), .A(n3407), .B(n3406), .ZN(n3414)
         );
  NAND2_X1 U4261 ( .A1(n3414), .A2(n4570), .ZN(n3412) );
  AOI21_X1 U4262 ( .B1(n3531), .B2(n2353), .A(n4312), .ZN(n3417) );
  OAI22_X1 U4263 ( .A1(n4570), .A2(n3409), .B1(n3532), .B2(n4313), .ZN(n3410)
         );
  AOI21_X1 U4264 ( .B1(n3417), .B2(n4557), .A(n3410), .ZN(n3411) );
  OAI211_X1 U4265 ( .C1(n3413), .C2(n4143), .A(n3412), .B(n3411), .ZN(U3280)
         );
  AOI21_X1 U4266 ( .B1(n4411), .B2(n3415), .A(n3414), .ZN(n3419) );
  AOI22_X1 U4267 ( .A1(n3417), .A2(n4425), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4610), .ZN(n3416) );
  OAI21_X1 U4268 ( .B1(n3419), .B2(n4610), .A(n3416), .ZN(U3487) );
  AOI22_X1 U4269 ( .A1(n3417), .A2(n4337), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4334), .ZN(n3418) );
  OAI21_X1 U4270 ( .B1(n3419), .B2(n4334), .A(n3418), .ZN(U3528) );
  NAND2_X1 U4271 ( .A1(n3421), .A2(n3420), .ZN(n4286) );
  NAND2_X1 U4272 ( .A1(n4283), .A2(n4284), .ZN(n3794) );
  XNOR2_X1 U4273 ( .A(n4286), .B(n3794), .ZN(n3424) );
  AOI22_X1 U4274 ( .A1(n4223), .A2(n3893), .B1(n4261), .B2(n4293), .ZN(n3423)
         );
  NAND2_X1 U4275 ( .A1(n3582), .A2(n4326), .ZN(n3422) );
  OAI211_X1 U4276 ( .C1(n3424), .C2(n4330), .A(n3423), .B(n3422), .ZN(n4409)
         );
  INV_X1 U4277 ( .A(n4409), .ZN(n3433) );
  XNOR2_X1 U4278 ( .A(n3426), .B(n3794), .ZN(n4410) );
  INV_X1 U4279 ( .A(n4310), .ZN(n3428) );
  OAI21_X1 U4280 ( .B1(n3428), .B2(n3427), .A(n4296), .ZN(n4476) );
  INV_X1 U4281 ( .A(n3429), .ZN(n3583) );
  AOI22_X1 U4282 ( .A1(n4276), .A2(REG2_REG_12__SCAN_IN), .B1(n3583), .B2(
        n4566), .ZN(n3430) );
  OAI21_X1 U4283 ( .B1(n4476), .B2(n4315), .A(n3430), .ZN(n3431) );
  AOI21_X1 U4284 ( .B1(n4410), .B2(n4255), .A(n3431), .ZN(n3432) );
  OAI21_X1 U4285 ( .B1(n3433), .B2(n4280), .A(n3432), .ZN(U3278) );
  XOR2_X1 U4286 ( .A(n3435), .B(n3434), .Z(n3440) );
  INV_X1 U4287 ( .A(n3436), .ZN(n3905) );
  INV_X1 U4288 ( .A(n3914), .ZN(n3437) );
  AOI211_X1 U4289 ( .C1(n3905), .C2(n3438), .A(n3437), .B(n4541), .ZN(n3439)
         );
  AOI21_X1 U4290 ( .B1(n4535), .B2(n3440), .A(n3439), .ZN(n3442) );
  AOI22_X1 U4291 ( .A1(n4527), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3441) );
  OAI21_X1 U4292 ( .B1(n3443), .B2(n3777), .A(n3444), .ZN(n4591) );
  XNOR2_X1 U4293 ( .A(n3777), .B(n3445), .ZN(n3450) );
  OAI22_X1 U4294 ( .A1(n3446), .A2(n4320), .B1(n4289), .B2(n3452), .ZN(n3448)
         );
  NOR2_X1 U4295 ( .A1(n4591), .A2(n4322), .ZN(n3447) );
  AOI211_X1 U4296 ( .C1(n4293), .C2(n3898), .A(n3448), .B(n3447), .ZN(n3449)
         );
  OAI21_X1 U4297 ( .B1(n4330), .B2(n3450), .A(n3449), .ZN(n4593) );
  OAI211_X1 U4298 ( .C1(n3453), .C2(n3452), .A(n3451), .B(n4602), .ZN(n4592)
         );
  OAI22_X1 U4299 ( .A1(n4592), .A2(n4490), .B1(n4313), .B2(n3454), .ZN(n3455)
         );
  OAI21_X1 U4300 ( .B1(n4593), .B2(n3455), .A(n4570), .ZN(n3457) );
  NAND2_X1 U4301 ( .A1(n4276), .A2(REG2_REG_4__SCAN_IN), .ZN(n3456) );
  OAI211_X1 U4302 ( .C1(n4591), .C2(n4306), .A(n3457), .B(n3456), .ZN(U3286)
         );
  INV_X1 U4303 ( .A(n3458), .ZN(n3459) );
  INV_X1 U4304 ( .A(n3615), .ZN(n3462) );
  OAI21_X1 U4305 ( .B1(n3616), .B2(n3463), .A(n3462), .ZN(n3468) );
  AOI21_X1 U4306 ( .B1(n3466), .B2(n3465), .A(n3464), .ZN(n3467) );
  XNOR2_X1 U4307 ( .A(n3468), .B(n3467), .ZN(n3474) );
  NOR2_X1 U4308 ( .A1(n4073), .A2(n3695), .ZN(n3472) );
  INV_X1 U4309 ( .A(n4102), .ZN(n4063) );
  AOI22_X1 U4310 ( .A1(n3730), .A2(n3469), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3470) );
  OAI21_X1 U4311 ( .B1(n4063), .B2(n3716), .A(n3470), .ZN(n3471) );
  AOI211_X1 U4312 ( .C1(n3731), .C2(n4065), .A(n3472), .B(n3471), .ZN(n3473)
         );
  OAI21_X1 U4313 ( .B1(n3474), .B2(n3719), .A(n3473), .ZN(U3222) );
  NAND3_X1 U4314 ( .A1(n3476), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3478) );
  INV_X1 U4315 ( .A(DATAI_31_), .ZN(n3477) );
  OAI22_X1 U4316 ( .A1(n3475), .A2(n3478), .B1(STATE_REG_SCAN_IN), .B2(n3477), 
        .ZN(U3321) );
  NAND2_X1 U4317 ( .A1(n3479), .A2(n4255), .ZN(n3486) );
  INV_X1 U4318 ( .A(n3480), .ZN(n3484) );
  OAI22_X1 U4319 ( .A1(n3482), .A2(n4313), .B1(n3481), .B2(n4570), .ZN(n3483)
         );
  AOI21_X1 U4320 ( .B1(n3484), .B2(n4557), .A(n3483), .ZN(n3485) );
  OAI211_X1 U4321 ( .C1(n3487), .C2(n4276), .A(n3486), .B(n3485), .ZN(U3262)
         );
  XOR2_X1 U4322 ( .A(n3489), .B(n3488), .Z(n3490) );
  NAND2_X1 U4323 ( .A1(n3490), .A2(n3726), .ZN(n3498) );
  AOI21_X1 U4324 ( .B1(n3731), .B2(n3895), .A(n3491), .ZN(n3497) );
  AOI22_X1 U4325 ( .A1(n3728), .A2(n3897), .B1(n3730), .B2(n3492), .ZN(n3496)
         );
  INV_X1 U4326 ( .A(n3493), .ZN(n3494) );
  NAND2_X1 U4327 ( .A1(n3733), .A2(n3494), .ZN(n3495) );
  NAND4_X1 U4328 ( .A1(n3498), .A2(n3497), .A3(n3496), .A4(n3495), .ZN(U3210)
         );
  XNOR2_X1 U4329 ( .A(n3500), .B(n3499), .ZN(n3506) );
  INV_X1 U4330 ( .A(n4065), .ZN(n4030) );
  AOI22_X1 U4331 ( .A1(n3730), .A2(n3501), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3502) );
  OAI21_X1 U4332 ( .B1(n4030), .B2(n3716), .A(n3502), .ZN(n3504) );
  NOR2_X1 U4333 ( .A1(n4014), .A2(n3689), .ZN(n3503) );
  AOI211_X1 U4334 ( .C1(n4038), .C2(n3733), .A(n3504), .B(n3503), .ZN(n3505)
         );
  OAI21_X1 U4335 ( .B1(n3506), .B2(n3719), .A(n3505), .ZN(U3211) );
  INV_X1 U4336 ( .A(n3507), .ZN(n3590) );
  NOR2_X1 U4337 ( .A1(n3590), .A2(n3508), .ZN(n3510) );
  XOR2_X1 U4338 ( .A(n3510), .B(n3509), .Z(n3511) );
  NAND2_X1 U4339 ( .A1(n3511), .A2(n3726), .ZN(n3516) );
  AND2_X1 U4340 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n3940) );
  AOI21_X1 U4341 ( .B1(n3728), .B2(n4261), .A(n3940), .ZN(n3515) );
  AOI22_X1 U4342 ( .A1(n3731), .A2(n4264), .B1(n3730), .B2(n3512), .ZN(n3514)
         );
  NAND2_X1 U4343 ( .A1(n3733), .A2(n4275), .ZN(n3513) );
  NAND4_X1 U4344 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(U3212)
         );
  INV_X1 U4345 ( .A(n3517), .ZN(n3521) );
  AOI21_X1 U4346 ( .B1(n3662), .B2(n3519), .A(n3518), .ZN(n3520) );
  AOI22_X1 U4347 ( .A1(n3891), .A2(n3728), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3522) );
  OAI21_X1 U4348 ( .B1(n3666), .B2(n4105), .A(n3522), .ZN(n3523) );
  AOI21_X1 U4349 ( .B1(n3731), .B2(n4102), .A(n3523), .ZN(n3524) );
  OAI211_X1 U4350 ( .C1(n3695), .C2(n4107), .A(n3525), .B(n3524), .ZN(U3213)
         );
  AOI21_X1 U4351 ( .B1(n3527), .B2(n3526), .A(n3719), .ZN(n3529) );
  NAND2_X1 U4352 ( .A1(n3529), .A2(n3528), .ZN(n3537) );
  AOI21_X1 U4353 ( .B1(n3728), .B2(n3894), .A(n3530), .ZN(n3536) );
  AOI22_X1 U4354 ( .A1(n3731), .A2(n3893), .B1(n3730), .B2(n3531), .ZN(n3535)
         );
  INV_X1 U4355 ( .A(n3532), .ZN(n3533) );
  NAND2_X1 U4356 ( .A1(n3733), .A2(n3533), .ZN(n3534) );
  NAND4_X1 U4357 ( .A1(n3537), .A2(n3536), .A3(n3535), .A4(n3534), .ZN(U3214)
         );
  INV_X1 U4358 ( .A(n3686), .ZN(n3540) );
  INV_X1 U4359 ( .A(n3539), .ZN(n3683) );
  NAND2_X1 U4360 ( .A1(n3686), .A2(n3683), .ZN(n3538) );
  AOI22_X1 U4361 ( .A1(n3540), .A2(n3539), .B1(n3538), .B2(n3684), .ZN(n3544)
         );
  NOR2_X1 U4362 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  XNOR2_X1 U4363 ( .A(n3544), .B(n3543), .ZN(n3545) );
  NAND2_X1 U4364 ( .A1(n3545), .A2(n3726), .ZN(n3552) );
  NAND2_X1 U4365 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3978) );
  INV_X1 U4366 ( .A(n3978), .ZN(n3546) );
  AOI21_X1 U4367 ( .B1(n4177), .B2(n3731), .A(n3546), .ZN(n3551) );
  AOI22_X1 U4368 ( .A1(n3728), .A2(n4210), .B1(n3730), .B2(n3547), .ZN(n3550)
         );
  INV_X1 U4369 ( .A(n4182), .ZN(n3548) );
  NAND2_X1 U4370 ( .A1(n3733), .A2(n3548), .ZN(n3549) );
  NAND4_X1 U4371 ( .A1(n3552), .A2(n3551), .A3(n3550), .A4(n3549), .ZN(U3216)
         );
  NAND2_X1 U4372 ( .A1(n2013), .A2(n3626), .ZN(n3553) );
  XNOR2_X1 U4373 ( .A(n3554), .B(n3553), .ZN(n3555) );
  NAND2_X1 U4374 ( .A1(n3555), .A2(n3726), .ZN(n3563) );
  AOI21_X1 U4375 ( .B1(n3728), .B2(n3896), .A(n3556), .ZN(n3562) );
  AOI22_X1 U4376 ( .A1(n3731), .A2(n3894), .B1(n3730), .B2(n3557), .ZN(n3561)
         );
  INV_X1 U4377 ( .A(n3558), .ZN(n3559) );
  NAND2_X1 U4378 ( .A1(n3733), .A2(n3559), .ZN(n3560) );
  NAND4_X1 U4379 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(U3218)
         );
  NOR2_X1 U4380 ( .A1(n2046), .A2(n3564), .ZN(n3567) );
  INV_X1 U4381 ( .A(n3642), .ZN(n3565) );
  AOI211_X1 U4382 ( .C1(n3639), .C2(n3565), .A(n3640), .B(n3567), .ZN(n3566)
         );
  AOI211_X1 U4383 ( .C1(n3568), .C2(n3567), .A(n3719), .B(n3566), .ZN(n3574)
         );
  INV_X1 U4384 ( .A(n4139), .ZN(n3572) );
  AOI22_X1 U4385 ( .A1(n3891), .A2(n3731), .B1(n3569), .B2(n3730), .ZN(n3571)
         );
  AOI22_X1 U4386 ( .A1(n4177), .A2(n3728), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3570) );
  OAI211_X1 U4387 ( .C1(n3695), .C2(n3572), .A(n3571), .B(n3570), .ZN(n3573)
         );
  OR2_X1 U4388 ( .A1(n3574), .A2(n3573), .ZN(U3220) );
  INV_X1 U4389 ( .A(n3575), .ZN(n3577) );
  NAND2_X1 U4390 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  XNOR2_X1 U4391 ( .A(n3579), .B(n3578), .ZN(n3580) );
  NAND2_X1 U4392 ( .A1(n3580), .A2(n3726), .ZN(n3587) );
  AOI21_X1 U4393 ( .B1(n3728), .B2(n3893), .A(n3581), .ZN(n3586) );
  AOI22_X1 U4394 ( .A1(n3731), .A2(n4261), .B1(n3730), .B2(n3582), .ZN(n3585)
         );
  NAND2_X1 U4395 ( .A1(n3733), .A2(n3583), .ZN(n3584) );
  NAND4_X1 U4396 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(U3221)
         );
  NOR2_X1 U4397 ( .A1(n3589), .A2(n3588), .ZN(n3596) );
  INV_X1 U4398 ( .A(n3724), .ZN(n3594) );
  NOR2_X1 U4399 ( .A1(n3591), .A2(n3590), .ZN(n3593) );
  NAND2_X1 U4400 ( .A1(n3593), .A2(n3592), .ZN(n3722) );
  NOR2_X1 U4401 ( .A1(n3593), .A2(n3592), .ZN(n3721) );
  AOI21_X1 U4402 ( .B1(n3594), .B2(n3722), .A(n3721), .ZN(n3595) );
  XOR2_X1 U4403 ( .A(n3596), .B(n3595), .Z(n3597) );
  NAND2_X1 U4404 ( .A1(n3597), .A2(n3726), .ZN(n3603) );
  INV_X1 U4405 ( .A(n4224), .ZN(n3690) );
  NAND2_X1 U4406 ( .A1(n3730), .A2(n4233), .ZN(n3598) );
  OAI21_X1 U4407 ( .B1(n3690), .B2(n3689), .A(n3598), .ZN(n3601) );
  NAND2_X1 U4408 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4525) );
  OAI21_X1 U4409 ( .B1(n3716), .B2(n3599), .A(n4525), .ZN(n3600) );
  NOR2_X1 U4410 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  OAI211_X1 U4411 ( .C1(n3695), .C2(n4234), .A(n3603), .B(n3602), .ZN(U3223)
         );
  INV_X1 U4412 ( .A(n3604), .ZN(n3606) );
  NAND2_X1 U4413 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  XNOR2_X1 U4414 ( .A(n3608), .B(n3607), .ZN(n3609) );
  NAND2_X1 U4415 ( .A1(n3609), .A2(n3726), .ZN(n3614) );
  AND2_X1 U4416 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3951) );
  AOI21_X1 U4417 ( .B1(n3728), .B2(n4243), .A(n3951), .ZN(n3613) );
  AOI22_X1 U4418 ( .A1(n3731), .A2(n4210), .B1(n3730), .B2(n4214), .ZN(n3612)
         );
  INV_X1 U4419 ( .A(n3610), .ZN(n4217) );
  NAND2_X1 U4420 ( .A1(n3733), .A2(n4217), .ZN(n3611) );
  NAND4_X1 U4421 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(U3225)
         );
  NOR2_X1 U4422 ( .A1(n3616), .A2(n3615), .ZN(n3618) );
  XNOR2_X1 U4423 ( .A(n3618), .B(n3617), .ZN(n3625) );
  OAI22_X1 U4424 ( .A1(n4120), .A2(n3716), .B1(STATE_REG_SCAN_IN), .B2(n3619), 
        .ZN(n3620) );
  AOI21_X1 U4425 ( .B1(n3621), .B2(n3730), .A(n3620), .ZN(n3622) );
  OAI21_X1 U4426 ( .B1(n4048), .B2(n3689), .A(n3622), .ZN(n3623) );
  AOI21_X1 U4427 ( .B1(n4089), .B2(n3733), .A(n3623), .ZN(n3624) );
  OAI21_X1 U4428 ( .B1(n3625), .B2(n3719), .A(n3624), .ZN(U3226) );
  NAND2_X1 U4429 ( .A1(n3627), .A2(n3626), .ZN(n3629) );
  XNOR2_X1 U4430 ( .A(n3629), .B(n3628), .ZN(n3630) );
  NAND2_X1 U4431 ( .A1(n3630), .A2(n3726), .ZN(n3637) );
  AOI21_X1 U4432 ( .B1(n3731), .B2(n3677), .A(n3631), .ZN(n3636) );
  AOI22_X1 U4433 ( .A1(n3728), .A2(n3895), .B1(n3730), .B2(n3632), .ZN(n3635)
         );
  NAND2_X1 U4434 ( .A1(n3733), .A2(n3633), .ZN(n3634) );
  NAND4_X1 U4435 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(U3228)
         );
  INV_X1 U4436 ( .A(n3638), .ZN(n3643) );
  OAI21_X1 U4437 ( .B1(n3640), .B2(n3642), .A(n3639), .ZN(n3641) );
  OAI21_X1 U4438 ( .B1(n3643), .B2(n3642), .A(n3641), .ZN(n3644) );
  NAND2_X1 U4439 ( .A1(n3644), .A2(n3726), .ZN(n3650) );
  OAI22_X1 U4440 ( .A1(n4190), .A2(n3716), .B1(STATE_REG_SCAN_IN), .B2(n3645), 
        .ZN(n3646) );
  INV_X1 U4441 ( .A(n3646), .ZN(n3649) );
  AOI22_X1 U4442 ( .A1(n4118), .A2(n3731), .B1(n4150), .B2(n3730), .ZN(n3648)
         );
  NAND2_X1 U4443 ( .A1(n3733), .A2(n4162), .ZN(n3647) );
  NAND4_X1 U4444 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(U3230)
         );
  XNOR2_X1 U4445 ( .A(n3652), .B(n3651), .ZN(n3653) );
  XNOR2_X1 U4446 ( .A(n3654), .B(n3653), .ZN(n3655) );
  NAND2_X1 U4447 ( .A1(n3655), .A2(n3726), .ZN(n3661) );
  AND2_X1 U4448 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4507) );
  AOI21_X1 U4449 ( .B1(n3728), .B2(n3892), .A(n4507), .ZN(n3660) );
  AOI22_X1 U4450 ( .A1(n3731), .A2(n4292), .B1(n3730), .B2(n3656), .ZN(n3659)
         );
  INV_X1 U4451 ( .A(n4300), .ZN(n3657) );
  NAND2_X1 U4452 ( .A1(n3733), .A2(n3657), .ZN(n3658) );
  NAND4_X1 U4453 ( .A1(n3661), .A2(n3660), .A3(n3659), .A4(n3658), .ZN(U3231)
         );
  OAI21_X1 U4454 ( .B1(n3664), .B2(n3663), .A(n3662), .ZN(n3665) );
  NAND2_X1 U4455 ( .A1(n3665), .A2(n3726), .ZN(n3670) );
  OAI22_X1 U4456 ( .A1(n4153), .A2(n3716), .B1(n3666), .B2(n4125), .ZN(n3668)
         );
  OAI22_X1 U4457 ( .A1(n4120), .A2(n3689), .B1(STATE_REG_SCAN_IN), .B2(n4654), 
        .ZN(n3667) );
  AOI211_X1 U4458 ( .C1(n4123), .C2(n3733), .A(n3668), .B(n3667), .ZN(n3669)
         );
  NAND2_X1 U4459 ( .A1(n3670), .A2(n3669), .ZN(U3232) );
  XNOR2_X1 U4460 ( .A(n3672), .B(n3671), .ZN(n3673) );
  XNOR2_X1 U4461 ( .A(n3674), .B(n3673), .ZN(n3675) );
  NAND2_X1 U4462 ( .A1(n3675), .A2(n3726), .ZN(n3682) );
  AOI21_X1 U4463 ( .B1(n3728), .B2(n3677), .A(n3676), .ZN(n3681) );
  AOI22_X1 U4464 ( .A1(n3731), .A2(n3892), .B1(n3730), .B2(n4327), .ZN(n3680)
         );
  INV_X1 U4465 ( .A(n4314), .ZN(n3678) );
  NAND2_X1 U4466 ( .A1(n3733), .A2(n3678), .ZN(n3679) );
  NAND4_X1 U4467 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(U3233)
         );
  XNOR2_X1 U4468 ( .A(n3684), .B(n3683), .ZN(n3685) );
  XNOR2_X1 U4469 ( .A(n3686), .B(n3685), .ZN(n3687) );
  NAND2_X1 U4470 ( .A1(n3687), .A2(n3726), .ZN(n3694) );
  NAND2_X1 U4471 ( .A1(n3730), .A2(n4193), .ZN(n3688) );
  OAI21_X1 U4472 ( .B1(n4190), .B2(n3689), .A(n3688), .ZN(n3692) );
  NAND2_X1 U4473 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4553) );
  OAI21_X1 U4474 ( .B1(n3716), .B2(n3690), .A(n4553), .ZN(n3691) );
  NOR2_X1 U4475 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  OAI211_X1 U4476 ( .C1(n3695), .C2(n4197), .A(n3694), .B(n3693), .ZN(U3235)
         );
  XNOR2_X1 U4477 ( .A(n3697), .B(n3696), .ZN(n3698) );
  XNOR2_X1 U4478 ( .A(n3699), .B(n3698), .ZN(n3700) );
  NAND2_X1 U4479 ( .A1(n3700), .A2(n3726), .ZN(n3707) );
  AOI21_X1 U4480 ( .B1(n3731), .B2(n3896), .A(n3701), .ZN(n3706) );
  AOI22_X1 U4481 ( .A1(n3728), .A2(n3898), .B1(n3730), .B2(n3702), .ZN(n3705)
         );
  NAND2_X1 U4482 ( .A1(n3733), .A2(n3703), .ZN(n3704) );
  NAND4_X1 U4483 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(U3236)
         );
  INV_X1 U4484 ( .A(n3708), .ZN(n3709) );
  NOR2_X1 U4485 ( .A1(n3710), .A2(n3709), .ZN(n3711) );
  XNOR2_X1 U4486 ( .A(n3712), .B(n3711), .ZN(n3720) );
  AOI22_X1 U4487 ( .A1(n3730), .A2(n3713), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3715) );
  NAND2_X1 U4488 ( .A1(n4056), .A2(n3733), .ZN(n3714) );
  OAI211_X1 U4489 ( .C1(n4048), .C2(n3716), .A(n3715), .B(n3714), .ZN(n3717)
         );
  AOI21_X1 U4490 ( .B1(n4050), .B2(n3731), .A(n3717), .ZN(n3718) );
  OAI21_X1 U4491 ( .B1(n3720), .B2(n3719), .A(n3718), .ZN(U3237) );
  INV_X1 U4492 ( .A(n3721), .ZN(n3723) );
  NAND2_X1 U4493 ( .A1(n3723), .A2(n3722), .ZN(n3725) );
  XNOR2_X1 U4494 ( .A(n3725), .B(n3724), .ZN(n3727) );
  NAND2_X1 U4495 ( .A1(n3727), .A2(n3726), .ZN(n3737) );
  AND2_X1 U4496 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4518) );
  AOI21_X1 U4497 ( .B1(n3728), .B2(n4292), .A(n4518), .ZN(n3736) );
  AOI22_X1 U4498 ( .A1(n3731), .A2(n4243), .B1(n3730), .B2(n3729), .ZN(n3735)
         );
  INV_X1 U4499 ( .A(n3732), .ZN(n4252) );
  NAND2_X1 U4500 ( .A1(n3733), .A2(n4252), .ZN(n3734) );
  NAND4_X1 U4501 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(U3238)
         );
  NAND2_X1 U4502 ( .A1(n3740), .A2(n4239), .ZN(n3847) );
  NAND2_X1 U4503 ( .A1(n3739), .A2(n3738), .ZN(n3832) );
  NAND2_X1 U4504 ( .A1(n3832), .A2(n3740), .ZN(n3848) );
  OAI21_X1 U4505 ( .B1(n4266), .B2(n3847), .A(n3848), .ZN(n3742) );
  INV_X1 U4506 ( .A(n3852), .ZN(n3741) );
  AOI211_X1 U4507 ( .C1(n3742), .C2(n3856), .A(n3741), .B(n3855), .ZN(n3744)
         );
  INV_X1 U4508 ( .A(n3743), .ZN(n3860) );
  OAI21_X1 U4509 ( .B1(n3744), .B2(n3860), .A(n3859), .ZN(n3745) );
  NAND2_X1 U4510 ( .A1(n3745), .A2(n3863), .ZN(n3747) );
  OR2_X1 U4511 ( .A1(n3801), .A2(n2233), .ZN(n3866) );
  AOI21_X1 U4512 ( .B1(n3747), .B2(n3746), .A(n3866), .ZN(n3758) );
  INV_X1 U4513 ( .A(n3748), .ZN(n3771) );
  NAND2_X1 U4514 ( .A1(n3771), .A2(n3800), .ZN(n3867) );
  NAND2_X1 U4515 ( .A1(n3754), .A2(DATAI_29_), .ZN(n3984) );
  NAND2_X1 U4516 ( .A1(n3749), .A2(DATAI_31_), .ZN(n3987) );
  NAND2_X1 U4517 ( .A1(n3986), .A2(n3987), .ZN(n3875) );
  INV_X1 U4518 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3998) );
  NAND2_X1 U4519 ( .A1(n3750), .A2(REG1_REG_30__SCAN_IN), .ZN(n3753) );
  INV_X1 U4520 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4430) );
  OR2_X1 U4521 ( .A1(n3751), .A2(n4430), .ZN(n3752) );
  OAI211_X1 U4522 ( .C1(n2680), .C2(n3998), .A(n3753), .B(n3752), .ZN(n4012)
         );
  NAND2_X1 U4523 ( .A1(n3754), .A2(DATAI_30_), .ZN(n3991) );
  OR2_X1 U4524 ( .A1(n4012), .A2(n3991), .ZN(n3755) );
  AND2_X1 U4525 ( .A1(n3875), .A2(n3755), .ZN(n3775) );
  OAI21_X1 U4526 ( .B1(n4774), .B2(n3984), .A(n3775), .ZN(n3764) );
  NOR3_X1 U4527 ( .A1(n3764), .A2(n3756), .A3(n3872), .ZN(n3757) );
  OAI211_X1 U4528 ( .C1(n3758), .C2(n3867), .A(n3757), .B(n4006), .ZN(n3768)
         );
  NAND2_X1 U4529 ( .A1(n4774), .A2(n3984), .ZN(n3759) );
  NAND2_X1 U4530 ( .A1(n4005), .A2(n3759), .ZN(n3762) );
  INV_X1 U4531 ( .A(n3760), .ZN(n3761) );
  OR2_X1 U4532 ( .A1(n3762), .A2(n3761), .ZN(n3869) );
  AOI21_X1 U4533 ( .B1(n4006), .B2(n3763), .A(n3762), .ZN(n3765) );
  NOR2_X1 U4534 ( .A1(n3765), .A2(n3764), .ZN(n3876) );
  OAI21_X1 U4535 ( .B1(n4031), .B2(n3869), .A(n3876), .ZN(n3767) );
  INV_X1 U4536 ( .A(n3986), .ZN(n3766) );
  INV_X1 U4537 ( .A(n3991), .ZN(n3993) );
  AOI22_X1 U4538 ( .A1(n3768), .A2(n3767), .B1(n3766), .B2(n3993), .ZN(n3770)
         );
  NAND2_X1 U4539 ( .A1(n4012), .A2(n3991), .ZN(n3773) );
  AOI21_X1 U4540 ( .B1(n3773), .B2(n3986), .A(n3987), .ZN(n3769) );
  NOR2_X1 U4541 ( .A1(n3770), .A2(n3769), .ZN(n3882) );
  INV_X1 U4542 ( .A(n4000), .ZN(n3806) );
  INV_X1 U4543 ( .A(n4031), .ZN(n4028) );
  NAND2_X1 U4544 ( .A1(n3771), .A2(n4043), .ZN(n4062) );
  INV_X1 U4545 ( .A(n4095), .ZN(n3858) );
  NAND2_X1 U4546 ( .A1(n3858), .A2(n4096), .ZN(n4132) );
  OR2_X1 U4547 ( .A1(n3986), .A2(n3987), .ZN(n3772) );
  NAND2_X1 U4548 ( .A1(n3773), .A2(n3772), .ZN(n3874) );
  INV_X1 U4549 ( .A(n3874), .ZN(n3774) );
  NAND4_X1 U4550 ( .A1(n3776), .A2(n4316), .A3(n3775), .A4(n3774), .ZN(n3787)
         );
  INV_X1 U4551 ( .A(n3777), .ZN(n3781) );
  INV_X1 U4552 ( .A(n3778), .ZN(n3780) );
  AND4_X1 U4553 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3783)
         );
  NAND4_X1 U4554 ( .A1(n2993), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(n3786)
         );
  NOR4_X1 U4555 ( .A1(n4115), .A2(n4132), .A3(n3787), .A4(n3786), .ZN(n3799)
         );
  NAND2_X1 U4556 ( .A1(n3789), .A2(n3788), .ZN(n4099) );
  INV_X1 U4557 ( .A(n4099), .ZN(n3798) );
  XNOR2_X1 U4558 ( .A(n4190), .B(n4181), .ZN(n4180) );
  NAND2_X1 U4559 ( .A1(n4169), .A2(n4167), .ZN(n4213) );
  OR4_X1 U4560 ( .A1(n4213), .A2(n4567), .A3(n3790), .A4(n4246), .ZN(n3796) );
  NAND4_X1 U4561 ( .A1(n3793), .A2(n3792), .A3(n4267), .A4(n3791), .ZN(n3795)
         );
  XNOR2_X1 U4562 ( .A(n4261), .B(n4298), .ZN(n4287) );
  NOR4_X1 U4563 ( .A1(n3796), .A2(n3795), .A3(n4287), .A4(n3794), .ZN(n3797)
         );
  NAND4_X1 U4564 ( .A1(n3799), .A2(n3798), .A3(n4180), .A4(n3797), .ZN(n3804)
         );
  INV_X1 U4565 ( .A(n3800), .ZN(n3802) );
  OR2_X1 U4566 ( .A1(n3802), .A2(n3801), .ZN(n4079) );
  XNOR2_X1 U4567 ( .A(n4177), .B(n4150), .ZN(n4148) );
  INV_X1 U4568 ( .A(n4148), .ZN(n3803) );
  NOR4_X1 U4569 ( .A1(n4062), .A2(n3804), .A3(n4079), .A4(n3803), .ZN(n3805)
         );
  NAND4_X1 U4570 ( .A1(n3806), .A2(n4028), .A3(n2018), .A4(n3805), .ZN(n3808)
         );
  XNOR2_X1 U4571 ( .A(n4774), .B(n3984), .ZN(n4344) );
  OAI21_X1 U4572 ( .B1(n3808), .B2(n4344), .A(n3807), .ZN(n3879) );
  INV_X1 U4573 ( .A(n3809), .ZN(n3812) );
  OAI211_X1 U4574 ( .C1(n3812), .C2(n4488), .A(n3811), .B(n3810), .ZN(n3814)
         );
  NAND3_X1 U4575 ( .A1(n3814), .A2(n3009), .A3(n3813), .ZN(n3817) );
  NAND3_X1 U4576 ( .A1(n3817), .A2(n3816), .A3(n3815), .ZN(n3820) );
  NAND3_X1 U4577 ( .A1(n3820), .A2(n3819), .A3(n3818), .ZN(n3823) );
  NAND4_X1 U4578 ( .A1(n3823), .A2(n3822), .A3(n3014), .A4(n3821), .ZN(n3826)
         );
  AND3_X1 U4579 ( .A1(n3826), .A2(n3825), .A3(n3824), .ZN(n3831) );
  NAND2_X1 U4580 ( .A1(n3828), .A2(n3827), .ZN(n3837) );
  OAI211_X1 U4581 ( .C1(n3831), .C2(n3837), .A(n3830), .B(n3829), .ZN(n3834)
         );
  INV_X1 U4582 ( .A(n3832), .ZN(n3833) );
  NAND3_X1 U4583 ( .A1(n3834), .A2(n3833), .A3(n3018), .ZN(n3846) );
  NOR4_X1 U4584 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3841)
         );
  INV_X1 U4585 ( .A(n3839), .ZN(n3840) );
  OAI21_X1 U4586 ( .B1(n3841), .B2(n3840), .A(n3848), .ZN(n3845) );
  NAND3_X1 U4587 ( .A1(n2016), .A2(n3843), .A3(n3842), .ZN(n3844) );
  AOI21_X1 U4588 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(n3854) );
  INV_X1 U4589 ( .A(n3847), .ZN(n3850) );
  INV_X1 U4590 ( .A(n3848), .ZN(n3849) );
  AOI21_X1 U4591 ( .B1(n3851), .B2(n3850), .A(n3849), .ZN(n3853) );
  OAI21_X1 U4592 ( .B1(n3854), .B2(n3853), .A(n3852), .ZN(n3857) );
  AOI21_X1 U4593 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n3861) );
  OAI211_X1 U4594 ( .C1(n3861), .C2(n3860), .A(n3859), .B(n3858), .ZN(n3864)
         );
  AOI21_X1 U4595 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3865) );
  INV_X1 U4596 ( .A(n3865), .ZN(n3868) );
  AOI21_X1 U4597 ( .B1(n3868), .B2(n2232), .A(n3867), .ZN(n3873) );
  INV_X1 U4598 ( .A(n3869), .ZN(n3871) );
  OAI211_X1 U4599 ( .C1(n3873), .C2(n3872), .A(n3871), .B(n3870), .ZN(n3877)
         );
  AOI22_X1 U4600 ( .A1(n3877), .A2(n3876), .B1(n3875), .B2(n3874), .ZN(n3878)
         );
  MUX2_X1 U4601 ( .A(n3879), .B(n3878), .S(n2408), .Z(n3880) );
  OAI21_X1 U4602 ( .B1(n3882), .B2(n3881), .A(n3880), .ZN(n3883) );
  XNOR2_X1 U4603 ( .A(n3883), .B(n3979), .ZN(n3889) );
  INV_X1 U4604 ( .A(n3884), .ZN(n3888) );
  NAND2_X1 U4605 ( .A1(n3885), .A2(n4485), .ZN(n3886) );
  OAI211_X1 U4606 ( .C1(n4487), .C2(n3888), .A(n3886), .B(B_REG_SCAN_IN), .ZN(
        n3887) );
  OAI21_X1 U4607 ( .B1(n3889), .B2(n3888), .A(n3887), .ZN(U3239) );
  MUX2_X1 U4608 ( .A(n4012), .B(DATAO_REG_30__SCAN_IN), .S(n3907), .Z(U3580)
         );
  MUX2_X1 U4609 ( .A(n4050), .B(DATAO_REG_27__SCAN_IN), .S(n3907), .Z(U3577)
         );
  MUX2_X1 U4610 ( .A(n4065), .B(DATAO_REG_26__SCAN_IN), .S(n3907), .Z(U3576)
         );
  MUX2_X1 U4611 ( .A(n4082), .B(DATAO_REG_25__SCAN_IN), .S(n3907), .Z(U3575)
         );
  MUX2_X1 U4612 ( .A(n3890), .B(DATAO_REG_23__SCAN_IN), .S(n3907), .Z(U3573)
         );
  MUX2_X1 U4613 ( .A(n3891), .B(DATAO_REG_22__SCAN_IN), .S(n3907), .Z(U3572)
         );
  MUX2_X1 U4614 ( .A(n4118), .B(DATAO_REG_21__SCAN_IN), .S(n3907), .Z(U3571)
         );
  MUX2_X1 U4615 ( .A(n4177), .B(DATAO_REG_20__SCAN_IN), .S(n3907), .Z(U3570)
         );
  MUX2_X1 U4616 ( .A(n4210), .B(DATAO_REG_18__SCAN_IN), .S(n3907), .Z(U3568)
         );
  MUX2_X1 U4617 ( .A(n4224), .B(DATAO_REG_17__SCAN_IN), .S(n3907), .Z(U3567)
         );
  MUX2_X1 U4618 ( .A(n4264), .B(DATAO_REG_15__SCAN_IN), .S(n3907), .Z(U3565)
         );
  MUX2_X1 U4619 ( .A(n4292), .B(DATAO_REG_14__SCAN_IN), .S(n3907), .Z(U3564)
         );
  MUX2_X1 U4620 ( .A(n4261), .B(DATAO_REG_13__SCAN_IN), .S(n3907), .Z(U3563)
         );
  MUX2_X1 U4621 ( .A(n3892), .B(DATAO_REG_12__SCAN_IN), .S(n3907), .Z(U3562)
         );
  MUX2_X1 U4622 ( .A(n3893), .B(DATAO_REG_11__SCAN_IN), .S(n3907), .Z(U3561)
         );
  MUX2_X1 U4623 ( .A(n3894), .B(DATAO_REG_9__SCAN_IN), .S(n3907), .Z(U3559) );
  MUX2_X1 U4624 ( .A(n3895), .B(DATAO_REG_8__SCAN_IN), .S(n3907), .Z(U3558) );
  MUX2_X1 U4625 ( .A(n3896), .B(DATAO_REG_7__SCAN_IN), .S(n3907), .Z(U3557) );
  MUX2_X1 U4626 ( .A(n3897), .B(DATAO_REG_6__SCAN_IN), .S(n3907), .Z(U3556) );
  MUX2_X1 U4627 ( .A(n3898), .B(DATAO_REG_5__SCAN_IN), .S(n3907), .Z(U3555) );
  MUX2_X1 U4628 ( .A(n3899), .B(DATAO_REG_4__SCAN_IN), .S(n3907), .Z(U3554) );
  MUX2_X1 U4629 ( .A(n3900), .B(DATAO_REG_3__SCAN_IN), .S(n3907), .Z(U3553) );
  MUX2_X1 U4630 ( .A(n2436), .B(DATAO_REG_2__SCAN_IN), .S(n3907), .Z(U3552) );
  MUX2_X1 U4631 ( .A(n2064), .B(DATAO_REG_0__SCAN_IN), .S(n3907), .Z(U3550) );
  NOR2_X1 U4632 ( .A1(n3902), .A2(n4485), .ZN(n3903) );
  AOI211_X1 U4633 ( .C1(n4485), .C2(n3905), .A(n3904), .B(n3903), .ZN(n3906)
         );
  AOI211_X1 U4634 ( .C1(n4627), .C2(n3908), .A(n3907), .B(n3906), .ZN(n3923)
         );
  INV_X1 U4635 ( .A(n3923), .ZN(n3921) );
  AOI22_X1 U4636 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4527), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3920) );
  XOR2_X1 U4637 ( .A(n3910), .B(n3909), .Z(n3911) );
  AOI22_X1 U4638 ( .A1(n4501), .A2(n4548), .B1(n4535), .B2(n3911), .ZN(n3919)
         );
  MUX2_X1 U4639 ( .A(REG2_REG_2__SCAN_IN), .B(n3090), .S(n2103), .Z(n3915) );
  NAND3_X1 U4640 ( .A1(n3915), .A2(n3914), .A3(n3913), .ZN(n3916) );
  NAND3_X1 U4641 ( .A1(n4537), .A2(n3917), .A3(n3916), .ZN(n3918) );
  NAND4_X1 U4642 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(U3242)
         );
  XOR2_X1 U4643 ( .A(n3922), .B(REG1_REG_4__SCAN_IN), .Z(n3924) );
  AOI21_X1 U4644 ( .B1(n4535), .B2(n3924), .A(n3923), .ZN(n3933) );
  NAND2_X1 U4645 ( .A1(n4527), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3932) );
  INV_X1 U4646 ( .A(n3925), .ZN(n3926) );
  AOI21_X1 U4647 ( .B1(n4548), .B2(n2479), .A(n3926), .ZN(n3931) );
  XNOR2_X1 U4648 ( .A(n3928), .B(n3927), .ZN(n3929) );
  NAND2_X1 U4649 ( .A1(n4537), .A2(n3929), .ZN(n3930) );
  NAND4_X1 U4650 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(U3244)
         );
  INV_X1 U4651 ( .A(n4582), .ZN(n4514) );
  NOR2_X1 U4652 ( .A1(n4301), .A2(n4514), .ZN(n4508) );
  AOI211_X1 U4653 ( .C1(n2662), .C2(n3937), .A(n4541), .B(n3954), .ZN(n3944)
         );
  AOI22_X1 U4654 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4514), .B1(n4582), .B2(
        n4620), .ZN(n4505) );
  OAI211_X1 U4655 ( .C1(n3939), .C2(REG1_REG_14__SCAN_IN), .A(n3945), .B(n4535), .ZN(n3942) );
  AOI21_X1 U4656 ( .B1(n4527), .B2(ADDR_REG_14__SCAN_IN), .A(n3940), .ZN(n3941) );
  OAI211_X1 U4657 ( .C1(n4540), .C2(n4492), .A(n3942), .B(n3941), .ZN(n3943)
         );
  OR2_X1 U4658 ( .A1(n3944), .A2(n3943), .ZN(U3254) );
  XOR2_X1 U4659 ( .A(REG1_REG_17__SCAN_IN), .B(n4491), .Z(n3949) );
  INV_X1 U4660 ( .A(n3955), .ZN(n4581) );
  AOI22_X1 U4661 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4581), .B1(n3955), .B2(
        n4399), .ZN(n4521) );
  NAND2_X1 U4662 ( .A1(n3946), .A2(n4579), .ZN(n3947) );
  OAI21_X1 U4663 ( .B1(n3949), .B2(n3948), .A(n3967), .ZN(n3950) );
  AOI22_X1 U4664 ( .A1(n4491), .A2(n4548), .B1(n4535), .B2(n3950), .ZN(n3964)
         );
  AOI21_X1 U4665 ( .B1(n4527), .B2(ADDR_REG_17__SCAN_IN), .A(n3951), .ZN(n3963) );
  XNOR2_X1 U4666 ( .A(n4491), .B(n3971), .ZN(n3960) );
  NOR2_X1 U4667 ( .A1(n3952), .A2(n4492), .ZN(n3953) );
  AOI22_X1 U4668 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4581), .B1(n3955), .B2(
        n2681), .ZN(n4516) );
  INV_X1 U4669 ( .A(n3957), .ZN(n3956) );
  NAND2_X1 U4670 ( .A1(n3956), .A2(n4579), .ZN(n3958) );
  INV_X1 U4671 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4529) );
  OAI21_X1 U4672 ( .B1(n3960), .B2(n3959), .A(n3974), .ZN(n3961) );
  NAND2_X1 U4673 ( .A1(n4537), .A2(n3961), .ZN(n3962) );
  NAND3_X1 U4674 ( .A1(n3964), .A2(n3963), .A3(n3962), .ZN(U3257) );
  INV_X1 U4675 ( .A(n4576), .ZN(n3966) );
  AOI22_X1 U4676 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3966), .B1(n4576), .B2(
        n3965), .ZN(n4544) );
  XNOR2_X1 U4677 ( .A(n4490), .B(REG1_REG_19__SCAN_IN), .ZN(n3968) );
  XNOR2_X1 U4678 ( .A(n3969), .B(n3968), .ZN(n3983) );
  NAND2_X1 U4679 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4576), .ZN(n3970) );
  OAI21_X1 U4680 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4576), .A(n3970), .ZN(n4543) );
  INV_X1 U4681 ( .A(n4491), .ZN(n3972) );
  NAND2_X1 U4682 ( .A1(n3972), .A2(n3971), .ZN(n3973) );
  MUX2_X1 U4683 ( .A(n4183), .B(REG2_REG_19__SCAN_IN), .S(n3979), .Z(n3975) );
  XNOR2_X1 U4684 ( .A(n3976), .B(n3975), .ZN(n3981) );
  NAND2_X1 U4685 ( .A1(n4527), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3977) );
  OAI211_X1 U4686 ( .C1(n4540), .C2(n3979), .A(n3978), .B(n3977), .ZN(n3980)
         );
  AOI21_X1 U4687 ( .B1(n3981), .B2(n4537), .A(n3980), .ZN(n3982) );
  OAI21_X1 U4688 ( .B1(n3983), .B2(n4546), .A(n3982), .ZN(U3259) );
  NAND2_X1 U4689 ( .A1(n4485), .A2(B_REG_SCAN_IN), .ZN(n3985) );
  AND2_X1 U4690 ( .A1(n4293), .A2(n3985), .ZN(n4011) );
  NAND2_X1 U4691 ( .A1(n3986), .A2(n4011), .ZN(n3995) );
  OAI21_X1 U4692 ( .B1(n3987), .B2(n4289), .A(n3995), .ZN(n4422) );
  NAND2_X1 U4693 ( .A1(n4570), .A2(n4422), .ZN(n3989) );
  NAND2_X1 U4694 ( .A1(n4276), .A2(REG2_REG_31__SCAN_IN), .ZN(n3988) );
  OAI211_X1 U4695 ( .C1(n4424), .C2(n4315), .A(n3989), .B(n3988), .ZN(U3260)
         );
  OAI21_X1 U4696 ( .B1(n4020), .B2(n3991), .A(n3990), .ZN(n3992) );
  INV_X1 U4697 ( .A(n3992), .ZN(n4426) );
  NAND2_X1 U4698 ( .A1(n4426), .A2(n4557), .ZN(n3997) );
  NAND2_X1 U4699 ( .A1(n4326), .A2(n3993), .ZN(n3994) );
  NAND2_X1 U4700 ( .A1(n3995), .A2(n3994), .ZN(n4427) );
  NAND2_X1 U4701 ( .A1(n4570), .A2(n4427), .ZN(n3996) );
  OAI211_X1 U4702 ( .C1(n4570), .C2(n3998), .A(n3997), .B(n3996), .ZN(U3261)
         );
  NAND2_X1 U4703 ( .A1(n2273), .A2(n4000), .ZN(n4345) );
  NAND2_X1 U4704 ( .A1(n4035), .A2(n4001), .ZN(n4343) );
  NAND2_X1 U4705 ( .A1(n4345), .A2(n4343), .ZN(n4003) );
  INV_X1 U4706 ( .A(n4344), .ZN(n4002) );
  XNOR2_X1 U4707 ( .A(n4003), .B(n4002), .ZN(n4004) );
  NAND2_X1 U4708 ( .A1(n4004), .A2(n4255), .ZN(n4027) );
  INV_X1 U4709 ( .A(n4005), .ZN(n4007) );
  XNOR2_X1 U4710 ( .A(n4009), .B(n4002), .ZN(n4010) );
  AOI22_X1 U4711 ( .A1(n4012), .A2(n4011), .B1(n4326), .B2(n4022), .ZN(n4013)
         );
  INV_X1 U4712 ( .A(n4342), .ZN(n4018) );
  OAI21_X1 U4713 ( .B1(n4019), .B2(n4313), .A(n4018), .ZN(n4025) );
  OAI22_X1 U4714 ( .A1(n2029), .A2(n4315), .B1(n4023), .B2(n4570), .ZN(n4024)
         );
  AOI21_X1 U4715 ( .B1(n4025), .B2(n4570), .A(n4024), .ZN(n4026) );
  NAND2_X1 U4716 ( .A1(n4027), .A2(n4026), .ZN(U3354) );
  XNOR2_X1 U4717 ( .A(n4029), .B(n4028), .ZN(n4349) );
  OAI22_X1 U4718 ( .A1(n4030), .A2(n4320), .B1(n4289), .B2(n4037), .ZN(n4034)
         );
  AOI21_X1 U4719 ( .B1(n4032), .B2(n4031), .A(n2027), .ZN(n4033) );
  NOR2_X1 U4720 ( .A1(n4350), .A2(n4276), .ZN(n4041) );
  OAI21_X1 U4721 ( .B1(n4053), .B2(n4037), .A(n4036), .ZN(n4352) );
  AOI22_X1 U4722 ( .A1(n4038), .A2(n4566), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4280), .ZN(n4039) );
  OAI21_X1 U4723 ( .B1(n4352), .B2(n4315), .A(n4039), .ZN(n4040) );
  INV_X1 U4724 ( .A(n4042), .ZN(U3263) );
  INV_X1 U4725 ( .A(n4354), .ZN(n4060) );
  INV_X1 U4726 ( .A(n4043), .ZN(n4044) );
  OR2_X1 U4727 ( .A1(n4045), .A2(n4044), .ZN(n4046) );
  XNOR2_X1 U4728 ( .A(n4046), .B(n2018), .ZN(n4047) );
  NAND2_X1 U4729 ( .A1(n4047), .A2(n4268), .ZN(n4052) );
  OAI22_X1 U4730 ( .A1(n4048), .A2(n4320), .B1(n4289), .B2(n4055), .ZN(n4049)
         );
  AOI21_X1 U4731 ( .B1(n4050), .B2(n4293), .A(n4049), .ZN(n4051) );
  NAND2_X1 U4732 ( .A1(n4052), .A2(n4051), .ZN(n4353) );
  INV_X1 U4733 ( .A(n4053), .ZN(n4054) );
  OAI21_X1 U4734 ( .B1(n4068), .B2(n4055), .A(n4054), .ZN(n4434) );
  AOI22_X1 U4735 ( .A1(n4056), .A2(n4566), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4280), .ZN(n4057) );
  OAI21_X1 U4736 ( .B1(n4434), .B2(n4315), .A(n4057), .ZN(n4058) );
  AOI21_X1 U4737 ( .B1(n4353), .B2(n4570), .A(n4058), .ZN(n4059) );
  OAI21_X1 U4738 ( .B1(n4060), .B2(n4143), .A(n4059), .ZN(U3264) );
  INV_X1 U4739 ( .A(n4356), .ZN(n4077) );
  XOR2_X1 U4740 ( .A(n4062), .B(n4061), .Z(n4067) );
  OAI22_X1 U4741 ( .A1(n4063), .A2(n4320), .B1(n4289), .B2(n4070), .ZN(n4064)
         );
  AOI21_X1 U4742 ( .B1(n4293), .B2(n4065), .A(n4064), .ZN(n4066) );
  OAI21_X1 U4743 ( .B1(n4067), .B2(n4330), .A(n4066), .ZN(n4355) );
  INV_X1 U4744 ( .A(n4086), .ZN(n4071) );
  INV_X1 U4745 ( .A(n4068), .ZN(n4069) );
  NOR2_X1 U4746 ( .A1(n4437), .A2(n4315), .ZN(n4075) );
  OAI22_X1 U4747 ( .A1(n4073), .A2(n4313), .B1(n4072), .B2(n4570), .ZN(n4074)
         );
  AOI211_X1 U4748 ( .C1(n4355), .C2(n4570), .A(n4075), .B(n4074), .ZN(n4076)
         );
  OAI21_X1 U4749 ( .B1(n4077), .B2(n4143), .A(n4076), .ZN(U3265) );
  XNOR2_X1 U4750 ( .A(n4078), .B(n4079), .ZN(n4360) );
  INV_X1 U4751 ( .A(n4360), .ZN(n4093) );
  XNOR2_X1 U4752 ( .A(n4080), .B(n4079), .ZN(n4084) );
  OAI22_X1 U4753 ( .A1(n4120), .A2(n4320), .B1(n4289), .B2(n4087), .ZN(n4081)
         );
  AOI21_X1 U4754 ( .B1(n4082), .B2(n4293), .A(n4081), .ZN(n4083) );
  OAI21_X1 U4755 ( .B1(n4084), .B2(n4330), .A(n4083), .ZN(n4359) );
  INV_X1 U4756 ( .A(n4085), .ZN(n4088) );
  OAI21_X1 U4757 ( .B1(n4088), .B2(n4087), .A(n4086), .ZN(n4440) );
  AOI22_X1 U4758 ( .A1(n4089), .A2(n4566), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4280), .ZN(n4090) );
  OAI21_X1 U4759 ( .B1(n4440), .B2(n4315), .A(n4090), .ZN(n4091) );
  AOI21_X1 U4760 ( .B1(n4359), .B2(n4570), .A(n4091), .ZN(n4092) );
  OAI21_X1 U4761 ( .B1(n4093), .B2(n4143), .A(n4092), .ZN(U3266) );
  XOR2_X1 U4762 ( .A(n4099), .B(n4094), .Z(n4364) );
  INV_X1 U4763 ( .A(n4364), .ZN(n4112) );
  OR2_X1 U4764 ( .A1(n4131), .A2(n4095), .ZN(n4097) );
  OAI21_X1 U4765 ( .B1(n4116), .B2(n4115), .A(n4098), .ZN(n4100) );
  XNOR2_X1 U4766 ( .A(n4100), .B(n4099), .ZN(n4104) );
  OAI22_X1 U4767 ( .A1(n4133), .A2(n4320), .B1(n4289), .B2(n4105), .ZN(n4101)
         );
  AOI21_X1 U4768 ( .B1(n4293), .B2(n4102), .A(n4101), .ZN(n4103) );
  OAI21_X1 U4769 ( .B1(n4104), .B2(n4330), .A(n4103), .ZN(n4363) );
  OR2_X1 U4770 ( .A1(n4368), .A2(n4105), .ZN(n4106) );
  NAND2_X1 U4771 ( .A1(n4085), .A2(n4106), .ZN(n4443) );
  INV_X1 U4772 ( .A(n4107), .ZN(n4108) );
  AOI22_X1 U4773 ( .A1(n4108), .A2(n4566), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4280), .ZN(n4109) );
  OAI21_X1 U4774 ( .B1(n4443), .B2(n4315), .A(n4109), .ZN(n4110) );
  AOI21_X1 U4775 ( .B1(n4363), .B2(n4570), .A(n4110), .ZN(n4111) );
  OAI21_X1 U4776 ( .B1(n4112), .B2(n4143), .A(n4111), .ZN(U3267) );
  OAI21_X1 U4777 ( .B1(n4114), .B2(n4115), .A(n4113), .ZN(n4371) );
  XNOR2_X1 U4778 ( .A(n4116), .B(n4115), .ZN(n4122) );
  NOR2_X1 U4779 ( .A1(n4289), .A2(n4125), .ZN(n4117) );
  AOI21_X1 U4780 ( .B1(n4118), .B2(n4223), .A(n4117), .ZN(n4119) );
  OAI21_X1 U4781 ( .B1(n4120), .B2(n4318), .A(n4119), .ZN(n4121) );
  AOI21_X1 U4782 ( .B1(n4122), .B2(n4268), .A(n4121), .ZN(n4370) );
  AOI22_X1 U4783 ( .A1(n4123), .A2(n4566), .B1(REG2_REG_22__SCAN_IN), .B2(
        n4280), .ZN(n4127) );
  NOR2_X1 U4784 ( .A1(n4124), .A2(n4125), .ZN(n4367) );
  OR3_X1 U4785 ( .A1(n4368), .A2(n4367), .A3(n4315), .ZN(n4126) );
  OAI211_X1 U4786 ( .C1(n4370), .C2(n4280), .A(n4127), .B(n4126), .ZN(n4128)
         );
  INV_X1 U4787 ( .A(n4128), .ZN(n4129) );
  OAI21_X1 U4788 ( .B1(n4371), .B2(n4143), .A(n4129), .ZN(U3268) );
  XOR2_X1 U4789 ( .A(n4130), .B(n4132), .Z(n4373) );
  INV_X1 U4790 ( .A(n4373), .ZN(n4144) );
  XOR2_X1 U4791 ( .A(n4132), .B(n4131), .Z(n4136) );
  OAI22_X1 U4792 ( .A1(n4133), .A2(n4318), .B1(n4289), .B2(n4138), .ZN(n4134)
         );
  AOI21_X1 U4793 ( .B1(n4223), .B2(n4177), .A(n4134), .ZN(n4135) );
  OAI21_X1 U4794 ( .B1(n4136), .B2(n4330), .A(n4135), .ZN(n4372) );
  INV_X1 U4795 ( .A(n4124), .ZN(n4137) );
  OAI21_X1 U4796 ( .B1(n3055), .B2(n4138), .A(n4137), .ZN(n4447) );
  AOI22_X1 U4797 ( .A1(n4139), .A2(n4566), .B1(n4276), .B2(
        REG2_REG_21__SCAN_IN), .ZN(n4140) );
  OAI21_X1 U4798 ( .B1(n4447), .B2(n4315), .A(n4140), .ZN(n4141) );
  AOI21_X1 U4799 ( .B1(n4372), .B2(n4570), .A(n4141), .ZN(n4142) );
  OAI21_X1 U4800 ( .B1(n4144), .B2(n4143), .A(n4142), .ZN(U3269) );
  XNOR2_X1 U4801 ( .A(n4145), .B(n4148), .ZN(n4157) );
  NAND2_X1 U4802 ( .A1(n4147), .A2(n4146), .ZN(n4149) );
  XNOR2_X1 U4803 ( .A(n4149), .B(n4148), .ZN(n4155) );
  AOI22_X1 U4804 ( .A1(n4151), .A2(n4223), .B1(n4326), .B2(n4150), .ZN(n4152)
         );
  OAI21_X1 U4805 ( .B1(n4153), .B2(n4318), .A(n4152), .ZN(n4154) );
  AOI21_X1 U4806 ( .B1(n4155), .B2(n4268), .A(n4154), .ZN(n4156) );
  OAI21_X1 U4807 ( .B1(n4157), .B2(n4322), .A(n4156), .ZN(n4376) );
  INV_X1 U4808 ( .A(n4376), .ZN(n4166) );
  INV_X1 U4809 ( .A(n4157), .ZN(n4377) );
  INV_X1 U4810 ( .A(n4158), .ZN(n4161) );
  OAI21_X1 U4811 ( .B1(n4161), .B2(n4160), .A(n4159), .ZN(n4451) );
  AOI22_X1 U4812 ( .A1(REG2_REG_20__SCAN_IN), .A2(n4276), .B1(n4162), .B2(
        n4566), .ZN(n4163) );
  OAI21_X1 U4813 ( .B1(n4451), .B2(n4315), .A(n4163), .ZN(n4164) );
  AOI21_X1 U4814 ( .B1(n4377), .B2(n4568), .A(n4164), .ZN(n4165) );
  OAI21_X1 U4815 ( .B1(n4166), .B2(n4280), .A(n4165), .ZN(U3270) );
  INV_X1 U4816 ( .A(n4167), .ZN(n4168) );
  OR2_X1 U4817 ( .A1(n4206), .A2(n4168), .ZN(n4170) );
  NAND2_X1 U4818 ( .A1(n4170), .A2(n4169), .ZN(n4188) );
  INV_X1 U4819 ( .A(n4171), .ZN(n4173) );
  OAI21_X1 U4820 ( .B1(n4188), .B2(n4173), .A(n4172), .ZN(n4174) );
  XNOR2_X1 U4821 ( .A(n4174), .B(n4180), .ZN(n4179) );
  OAI22_X1 U4822 ( .A1(n4175), .A2(n4320), .B1(n4289), .B2(n4181), .ZN(n4176)
         );
  AOI21_X1 U4823 ( .B1(n4293), .B2(n4177), .A(n4176), .ZN(n4178) );
  OAI21_X1 U4824 ( .B1(n4179), .B2(n4330), .A(n4178), .ZN(n4380) );
  INV_X1 U4825 ( .A(n4380), .ZN(n4187) );
  XNOR2_X1 U4826 ( .A(n2022), .B(n4180), .ZN(n4381) );
  OAI21_X1 U4827 ( .B1(n4196), .B2(n4181), .A(n4158), .ZN(n4455) );
  NOR2_X1 U4828 ( .A1(n4455), .A2(n4315), .ZN(n4185) );
  OAI22_X1 U4829 ( .A1(n4570), .A2(n4183), .B1(n4182), .B2(n4313), .ZN(n4184)
         );
  AOI211_X1 U4830 ( .C1(n4381), .C2(n4255), .A(n4185), .B(n4184), .ZN(n4186)
         );
  OAI21_X1 U4831 ( .B1(n4276), .B2(n4187), .A(n4186), .ZN(U3271) );
  XNOR2_X1 U4832 ( .A(n4188), .B(n2993), .ZN(n4192) );
  AOI22_X1 U4833 ( .A1(n4224), .A2(n4223), .B1(n4326), .B2(n4193), .ZN(n4189)
         );
  OAI21_X1 U4834 ( .B1(n4190), .B2(n4318), .A(n4189), .ZN(n4191) );
  AOI21_X1 U4835 ( .B1(n4192), .B2(n4268), .A(n4191), .ZN(n4386) );
  NAND2_X1 U4836 ( .A1(n4216), .A2(n4193), .ZN(n4194) );
  NAND2_X1 U4837 ( .A1(n4194), .A2(n4602), .ZN(n4195) );
  NOR2_X1 U4838 ( .A1(n4196), .A2(n4195), .ZN(n4384) );
  INV_X1 U4839 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4198) );
  OAI22_X1 U4840 ( .A1(n4570), .A2(n4198), .B1(n4197), .B2(n4313), .ZN(n4199)
         );
  AOI21_X1 U4841 ( .B1(n4384), .B2(n4200), .A(n4199), .ZN(n4205) );
  NOR2_X1 U4842 ( .A1(n2024), .A2(n4201), .ZN(n4202) );
  OR2_X1 U4843 ( .A1(n4203), .A2(n4202), .ZN(n4385) );
  NAND2_X1 U4844 ( .A1(n4385), .A2(n4255), .ZN(n4204) );
  OAI211_X1 U4845 ( .C1(n4386), .C2(n4276), .A(n4205), .B(n4204), .ZN(U3272)
         );
  XOR2_X1 U4846 ( .A(n4213), .B(n4206), .Z(n4212) );
  OAI22_X1 U4847 ( .A1(n4208), .A2(n4320), .B1(n4289), .B2(n4207), .ZN(n4209)
         );
  AOI21_X1 U4848 ( .B1(n4210), .B2(n4293), .A(n4209), .ZN(n4211) );
  OAI21_X1 U4849 ( .B1(n4212), .B2(n4330), .A(n4211), .ZN(n4388) );
  INV_X1 U4850 ( .A(n4388), .ZN(n4221) );
  XOR2_X1 U4851 ( .A(n4213), .B(n2300), .Z(n4389) );
  NAND2_X1 U4852 ( .A1(n4393), .A2(n4214), .ZN(n4215) );
  NAND2_X1 U4853 ( .A1(n4216), .A2(n4215), .ZN(n4460) );
  AOI22_X1 U4854 ( .A1(n4276), .A2(REG2_REG_17__SCAN_IN), .B1(n4217), .B2(
        n4566), .ZN(n4218) );
  OAI21_X1 U4855 ( .B1(n4460), .B2(n4315), .A(n4218), .ZN(n4219) );
  AOI21_X1 U4856 ( .B1(n4389), .B2(n4255), .A(n4219), .ZN(n4220) );
  OAI21_X1 U4857 ( .B1(n4221), .B2(n4276), .A(n4220), .ZN(U3273) );
  XNOR2_X1 U4858 ( .A(n4222), .B(n4231), .ZN(n4228) );
  AOI22_X1 U4859 ( .A1(n4224), .A2(n4293), .B1(n4223), .B2(n4264), .ZN(n4225)
         );
  OAI21_X1 U4860 ( .B1(n4289), .B2(n4226), .A(n4225), .ZN(n4227) );
  AOI21_X1 U4861 ( .B1(n4228), .B2(n4268), .A(n4227), .ZN(n4395) );
  OAI21_X1 U4862 ( .B1(n4232), .B2(n4231), .A(n4230), .ZN(n4396) );
  INV_X1 U4863 ( .A(n4396), .ZN(n4237) );
  NAND2_X1 U4864 ( .A1(n4251), .A2(n4233), .ZN(n4392) );
  AND3_X1 U4865 ( .A1(n4393), .A2(n4557), .A3(n4392), .ZN(n4236) );
  OAI22_X1 U4866 ( .A1(n4570), .A2(n4529), .B1(n4234), .B2(n4313), .ZN(n4235)
         );
  AOI211_X1 U4867 ( .C1(n4237), .C2(n4255), .A(n4236), .B(n4235), .ZN(n4238)
         );
  OAI21_X1 U4868 ( .B1(n4276), .B2(n4395), .A(n4238), .ZN(U3274) );
  NAND2_X1 U4869 ( .A1(n4265), .A2(n4239), .ZN(n4240) );
  XNOR2_X1 U4870 ( .A(n4240), .B(n4246), .ZN(n4245) );
  OAI22_X1 U4871 ( .A1(n4241), .A2(n4320), .B1(n4289), .B2(n4249), .ZN(n4242)
         );
  AOI21_X1 U4872 ( .B1(n4293), .B2(n4243), .A(n4242), .ZN(n4244) );
  OAI21_X1 U4873 ( .B1(n4245), .B2(n4330), .A(n4244), .ZN(n4397) );
  INV_X1 U4874 ( .A(n4397), .ZN(n4257) );
  XNOR2_X1 U4875 ( .A(n4247), .B(n4246), .ZN(n4398) );
  OR2_X1 U4876 ( .A1(n4248), .A2(n4249), .ZN(n4250) );
  NAND2_X1 U4877 ( .A1(n4251), .A2(n4250), .ZN(n4465) );
  AOI22_X1 U4878 ( .A1(n4276), .A2(REG2_REG_15__SCAN_IN), .B1(n4252), .B2(
        n4566), .ZN(n4253) );
  OAI21_X1 U4879 ( .B1(n4465), .B2(n4315), .A(n4253), .ZN(n4254) );
  AOI21_X1 U4880 ( .B1(n4398), .B2(n4255), .A(n4254), .ZN(n4256) );
  OAI21_X1 U4881 ( .B1(n4257), .B2(n4280), .A(n4256), .ZN(U3275) );
  INV_X1 U4882 ( .A(n4258), .ZN(n4259) );
  AOI21_X1 U4883 ( .B1(n4267), .B2(n4260), .A(n4259), .ZN(n4272) );
  INV_X1 U4884 ( .A(n4261), .ZN(n4262) );
  OAI22_X1 U4885 ( .A1(n4262), .A2(n4320), .B1(n4289), .B2(n4273), .ZN(n4263)
         );
  AOI21_X1 U4886 ( .B1(n4293), .B2(n4264), .A(n4263), .ZN(n4271) );
  OAI21_X1 U4887 ( .B1(n4267), .B2(n4266), .A(n4265), .ZN(n4269) );
  NAND2_X1 U4888 ( .A1(n4269), .A2(n4268), .ZN(n4270) );
  OAI211_X1 U4889 ( .C1(n4272), .C2(n4322), .A(n4271), .B(n4270), .ZN(n4401)
         );
  INV_X1 U4890 ( .A(n4401), .ZN(n4281) );
  INV_X1 U4891 ( .A(n4272), .ZN(n4402) );
  NOR2_X1 U4892 ( .A1(n4297), .A2(n4273), .ZN(n4274) );
  OR2_X1 U4893 ( .A1(n4248), .A2(n4274), .ZN(n4468) );
  AOI22_X1 U4894 ( .A1(n4276), .A2(REG2_REG_14__SCAN_IN), .B1(n4275), .B2(
        n4566), .ZN(n4277) );
  OAI21_X1 U4895 ( .B1(n4468), .B2(n4315), .A(n4277), .ZN(n4278) );
  AOI21_X1 U4896 ( .B1(n4402), .B2(n4568), .A(n4278), .ZN(n4279) );
  OAI21_X1 U4897 ( .B1(n4281), .B2(n4280), .A(n4279), .ZN(U3276) );
  XOR2_X1 U4898 ( .A(n4282), .B(n4287), .Z(n4405) );
  INV_X1 U4899 ( .A(n4283), .ZN(n4285) );
  OAI21_X1 U4900 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(n4288) );
  XOR2_X1 U4901 ( .A(n4288), .B(n4287), .Z(n4295) );
  OAI22_X1 U4902 ( .A1(n4319), .A2(n4320), .B1(n4289), .B2(n4298), .ZN(n4291)
         );
  NOR2_X1 U4903 ( .A1(n4405), .A2(n4322), .ZN(n4290) );
  AOI211_X1 U4904 ( .C1(n4293), .C2(n4292), .A(n4291), .B(n4290), .ZN(n4294)
         );
  OAI21_X1 U4905 ( .B1(n4330), .B2(n4295), .A(n4294), .ZN(n4406) );
  NAND2_X1 U4906 ( .A1(n4406), .A2(n4570), .ZN(n4305) );
  INV_X1 U4907 ( .A(n4296), .ZN(n4299) );
  OAI21_X1 U4908 ( .B1(n4299), .B2(n4298), .A(n2309), .ZN(n4472) );
  INV_X1 U4909 ( .A(n4472), .ZN(n4303) );
  OAI22_X1 U4910 ( .A1(n4570), .A2(n4301), .B1(n4300), .B2(n4313), .ZN(n4302)
         );
  AOI21_X1 U4911 ( .B1(n4303), .B2(n4557), .A(n4302), .ZN(n4304) );
  OAI211_X1 U4912 ( .C1(n4405), .C2(n4306), .A(n4305), .B(n4304), .ZN(U3277)
         );
  INV_X1 U4913 ( .A(n4307), .ZN(n4308) );
  AOI21_X1 U4914 ( .B1(n4316), .B2(n4309), .A(n4308), .ZN(n4323) );
  INV_X1 U4915 ( .A(n4323), .ZN(n4415) );
  OAI21_X1 U4916 ( .B1(n4312), .B2(n4311), .A(n4310), .ZN(n4481) );
  OAI22_X1 U4917 ( .A1(n4481), .A2(n4315), .B1(n4314), .B2(n4313), .ZN(n4332)
         );
  XOR2_X1 U4918 ( .A(n4317), .B(n4316), .Z(n4329) );
  OAI22_X1 U4919 ( .A1(n4321), .A2(n4320), .B1(n4319), .B2(n4318), .ZN(n4325)
         );
  NOR2_X1 U4920 ( .A1(n4323), .A2(n4322), .ZN(n4324) );
  AOI211_X1 U4921 ( .C1(n4327), .C2(n4326), .A(n4325), .B(n4324), .ZN(n4328)
         );
  OAI21_X1 U4922 ( .B1(n4330), .B2(n4329), .A(n4328), .ZN(n4414) );
  MUX2_X1 U4923 ( .A(REG2_REG_11__SCAN_IN), .B(n4414), .S(n4570), .Z(n4331) );
  AOI211_X1 U4924 ( .C1(n4568), .C2(n4415), .A(n4332), .B(n4331), .ZN(n4333)
         );
  INV_X1 U4925 ( .A(n4333), .ZN(U3279) );
  NAND2_X1 U4926 ( .A1(n4416), .A2(n4422), .ZN(n4336) );
  NAND2_X1 U4927 ( .A1(n4334), .A2(REG1_REG_31__SCAN_IN), .ZN(n4335) );
  OAI211_X1 U4928 ( .C1(n4424), .C2(n4419), .A(n4336), .B(n4335), .ZN(U3549)
         );
  INV_X1 U4929 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4340) );
  NAND2_X1 U4930 ( .A1(n4426), .A2(n4337), .ZN(n4339) );
  NAND2_X1 U4931 ( .A1(n4416), .A2(n4427), .ZN(n4338) );
  OAI211_X1 U4932 ( .C1(n4416), .C2(n4340), .A(n4339), .B(n4338), .ZN(U3548)
         );
  INV_X1 U4933 ( .A(n4411), .ZN(n4604) );
  NAND4_X1 U4934 ( .A1(n4345), .A2(n4411), .A3(n4344), .A4(n4343), .ZN(n4346)
         );
  NAND3_X1 U4935 ( .A1(n4348), .A2(n4347), .A3(n4346), .ZN(n4431) );
  MUX2_X1 U4936 ( .A(REG1_REG_29__SCAN_IN), .B(n4431), .S(n4416), .Z(U3547) );
  NAND2_X1 U4937 ( .A1(n4349), .A2(n4411), .ZN(n4351) );
  AOI21_X1 U4938 ( .B1(n4354), .B2(n4411), .A(n4353), .ZN(n4433) );
  INV_X1 U4939 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4357) );
  AOI21_X1 U4940 ( .B1(n4356), .B2(n4411), .A(n4355), .ZN(n4435) );
  INV_X1 U4941 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4361) );
  AOI21_X1 U4942 ( .B1(n4360), .B2(n4411), .A(n4359), .ZN(n4438) );
  OAI21_X1 U4943 ( .B1(n4419), .B2(n4440), .A(n4362), .ZN(U3542) );
  AOI21_X1 U4944 ( .B1(n4364), .B2(n4411), .A(n4363), .ZN(n4441) );
  MUX2_X1 U4945 ( .A(n4681), .B(n4441), .S(n4416), .Z(n4365) );
  OAI21_X1 U4946 ( .B1(n4419), .B2(n4443), .A(n4365), .ZN(U3541) );
  OR3_X1 U4947 ( .A1(n4368), .A2(n4367), .A3(n4366), .ZN(n4369) );
  OAI211_X1 U4948 ( .C1(n4371), .C2(n4604), .A(n4370), .B(n4369), .ZN(n4444)
         );
  MUX2_X1 U4949 ( .A(REG1_REG_22__SCAN_IN), .B(n4444), .S(n4416), .Z(U3540) );
  INV_X1 U4950 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4374) );
  AOI21_X1 U4951 ( .B1(n4373), .B2(n4411), .A(n4372), .ZN(n4445) );
  MUX2_X1 U4952 ( .A(n4374), .B(n4445), .S(n4416), .Z(n4375) );
  OAI21_X1 U4953 ( .B1(n4419), .B2(n4447), .A(n4375), .ZN(U3539) );
  INV_X1 U4954 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4378) );
  AOI21_X1 U4955 ( .B1(n4595), .B2(n4377), .A(n4376), .ZN(n4448) );
  MUX2_X1 U4956 ( .A(n4378), .B(n4448), .S(n4416), .Z(n4379) );
  OAI21_X1 U4957 ( .B1(n4419), .B2(n4451), .A(n4379), .ZN(U3538) );
  INV_X1 U4958 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4382) );
  AOI21_X1 U4959 ( .B1(n4381), .B2(n4411), .A(n4380), .ZN(n4452) );
  MUX2_X1 U4960 ( .A(n4382), .B(n4452), .S(n4416), .Z(n4383) );
  OAI21_X1 U4961 ( .B1(n4419), .B2(n4455), .A(n4383), .ZN(U3537) );
  AOI21_X1 U4962 ( .B1(n4385), .B2(n4411), .A(n4384), .ZN(n4387) );
  NAND2_X1 U4963 ( .A1(n4387), .A2(n4386), .ZN(n4456) );
  MUX2_X1 U4964 ( .A(REG1_REG_18__SCAN_IN), .B(n4456), .S(n4416), .Z(U3536) );
  INV_X1 U4965 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4390) );
  AOI21_X1 U4966 ( .B1(n4389), .B2(n4411), .A(n4388), .ZN(n4457) );
  MUX2_X1 U4967 ( .A(n4390), .B(n4457), .S(n4416), .Z(n4391) );
  OAI21_X1 U4968 ( .B1(n4419), .B2(n4460), .A(n4391), .ZN(U3535) );
  NAND3_X1 U4969 ( .A1(n4393), .A2(n4602), .A3(n4392), .ZN(n4394) );
  OAI211_X1 U4970 ( .C1(n4604), .C2(n4396), .A(n4395), .B(n4394), .ZN(n4461)
         );
  MUX2_X1 U4971 ( .A(REG1_REG_16__SCAN_IN), .B(n4461), .S(n4416), .Z(U3534) );
  AOI21_X1 U4972 ( .B1(n4411), .B2(n4398), .A(n4397), .ZN(n4462) );
  MUX2_X1 U4973 ( .A(n4399), .B(n4462), .S(n4416), .Z(n4400) );
  OAI21_X1 U4974 ( .B1(n4419), .B2(n4465), .A(n4400), .ZN(U3533) );
  AOI21_X1 U4975 ( .B1(n4595), .B2(n4402), .A(n4401), .ZN(n4466) );
  MUX2_X1 U4976 ( .A(n4403), .B(n4466), .S(n4416), .Z(n4404) );
  OAI21_X1 U4977 ( .B1(n4419), .B2(n4468), .A(n4404), .ZN(U3532) );
  INV_X1 U4978 ( .A(n4405), .ZN(n4407) );
  AOI21_X1 U4979 ( .B1(n4595), .B2(n4407), .A(n4406), .ZN(n4469) );
  MUX2_X1 U4980 ( .A(n4620), .B(n4469), .S(n4416), .Z(n4408) );
  OAI21_X1 U4981 ( .B1(n4419), .B2(n4472), .A(n4408), .ZN(U3531) );
  INV_X1 U4982 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4412) );
  AOI21_X1 U4983 ( .B1(n4411), .B2(n4410), .A(n4409), .ZN(n4473) );
  MUX2_X1 U4984 ( .A(n4412), .B(n4473), .S(n4416), .Z(n4413) );
  OAI21_X1 U4985 ( .B1(n4419), .B2(n4476), .A(n4413), .ZN(U3530) );
  AOI21_X1 U4986 ( .B1(n4595), .B2(n4415), .A(n4414), .ZN(n4477) );
  MUX2_X1 U4987 ( .A(n4417), .B(n4477), .S(n4416), .Z(n4418) );
  OAI21_X1 U4988 ( .B1(n4419), .B2(n4481), .A(n4418), .ZN(U3529) );
  NOR2_X1 U4989 ( .A1(n4612), .A2(n4420), .ZN(n4421) );
  AOI21_X1 U4990 ( .B1(n4612), .B2(n4422), .A(n4421), .ZN(n4423) );
  OAI21_X1 U4991 ( .B1(n4424), .B2(n4480), .A(n4423), .ZN(U3517) );
  NAND2_X1 U4992 ( .A1(n4426), .A2(n4425), .ZN(n4429) );
  NAND2_X1 U4993 ( .A1(n4612), .A2(n4427), .ZN(n4428) );
  OAI211_X1 U4994 ( .C1(n4612), .C2(n4430), .A(n4429), .B(n4428), .ZN(U3516)
         );
  MUX2_X1 U4995 ( .A(REG0_REG_29__SCAN_IN), .B(n4431), .S(n4612), .Z(U3515) );
  MUX2_X1 U4996 ( .A(REG0_REG_27__SCAN_IN), .B(n4432), .S(n4612), .Z(U3513) );
  INV_X1 U4997 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4436) );
  MUX2_X1 U4998 ( .A(n4758), .B(n4438), .S(n4612), .Z(n4439) );
  MUX2_X1 U4999 ( .A(n4759), .B(n4441), .S(n4612), .Z(n4442) );
  OAI21_X1 U5000 ( .B1(n4443), .B2(n4480), .A(n4442), .ZN(U3509) );
  MUX2_X1 U5001 ( .A(REG0_REG_22__SCAN_IN), .B(n4444), .S(n4612), .Z(U3508) );
  MUX2_X1 U5002 ( .A(n4718), .B(n4445), .S(n4612), .Z(n4446) );
  OAI21_X1 U5003 ( .B1(n4447), .B2(n4480), .A(n4446), .ZN(U3507) );
  INV_X1 U5004 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4449) );
  MUX2_X1 U5005 ( .A(n4449), .B(n4448), .S(n4612), .Z(n4450) );
  OAI21_X1 U5006 ( .B1(n4451), .B2(n4480), .A(n4450), .ZN(U3506) );
  INV_X1 U5007 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4453) );
  MUX2_X1 U5008 ( .A(n4453), .B(n4452), .S(n4612), .Z(n4454) );
  OAI21_X1 U5009 ( .B1(n4455), .B2(n4480), .A(n4454), .ZN(U3505) );
  MUX2_X1 U5010 ( .A(REG0_REG_18__SCAN_IN), .B(n4456), .S(n4612), .Z(U3503) );
  INV_X1 U5011 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4458) );
  MUX2_X1 U5012 ( .A(n4458), .B(n4457), .S(n4612), .Z(n4459) );
  OAI21_X1 U5013 ( .B1(n4460), .B2(n4480), .A(n4459), .ZN(U3501) );
  MUX2_X1 U5014 ( .A(REG0_REG_16__SCAN_IN), .B(n4461), .S(n4612), .Z(U3499) );
  MUX2_X1 U5015 ( .A(n4463), .B(n4462), .S(n4612), .Z(n4464) );
  OAI21_X1 U5016 ( .B1(n4465), .B2(n4480), .A(n4464), .ZN(U3497) );
  MUX2_X1 U5017 ( .A(n4640), .B(n4466), .S(n4612), .Z(n4467) );
  OAI21_X1 U5018 ( .B1(n4468), .B2(n4480), .A(n4467), .ZN(U3495) );
  INV_X1 U5019 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4470) );
  MUX2_X1 U5020 ( .A(n4470), .B(n4469), .S(n4612), .Z(n4471) );
  OAI21_X1 U5021 ( .B1(n4472), .B2(n4480), .A(n4471), .ZN(U3493) );
  MUX2_X1 U5022 ( .A(n4474), .B(n4473), .S(n4612), .Z(n4475) );
  OAI21_X1 U5023 ( .B1(n4476), .B2(n4480), .A(n4475), .ZN(U3491) );
  MUX2_X1 U5024 ( .A(n4478), .B(n4477), .S(n4612), .Z(n4479) );
  OAI21_X1 U5025 ( .B1(n4481), .B2(n4480), .A(n4479), .ZN(U3489) );
  MUX2_X1 U5026 ( .A(DATAI_30_), .B(n4482), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5027 ( .A(n4483), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5028 ( .A(DATAI_28_), .B(n4484), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5029 ( .A(n4485), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5030 ( .A(n2894), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5031 ( .A(n4486), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5032 ( .A(n4487), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5033 ( .A(n4488), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5034 ( .A(DATAI_20_), .B(n4489), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5035 ( .A(DATAI_19_), .B(n4490), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5036 ( .A(n4491), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5037 ( .A(DATAI_14_), .B(n2212), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5038 ( .A(DATAI_12_), .B(n4493), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5039 ( .A(DATAI_11_), .B(n4494), .S(STATE_REG_SCAN_IN), .Z(U3341)
         );
  MUX2_X1 U5040 ( .A(n4495), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5041 ( .A(n4496), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5042 ( .A(DATAI_8_), .B(n4497), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5043 ( .A(DATAI_7_), .B(n2208), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5044 ( .A(n4498), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5045 ( .A(n4499), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5046 ( .A(DATAI_4_), .B(n2479), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5047 ( .A(DATAI_3_), .B(n4500), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5048 ( .A(n4501), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5049 ( .A(n4503), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5050 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  AOI211_X1 U5051 ( .C1(n2015), .C2(n4505), .A(n4504), .B(n4546), .ZN(n4506)
         );
  AOI211_X1 U5052 ( .C1(n4527), .C2(ADDR_REG_13__SCAN_IN), .A(n4507), .B(n4506), .ZN(n4513) );
  AOI21_X1 U5053 ( .B1(n4301), .B2(n4514), .A(n4508), .ZN(n4511) );
  AOI21_X1 U5054 ( .B1(n4511), .B2(n4510), .A(n4541), .ZN(n4509) );
  OAI21_X1 U5055 ( .B1(n4511), .B2(n4510), .A(n4509), .ZN(n4512) );
  OAI211_X1 U5056 ( .C1(n4540), .C2(n4514), .A(n4513), .B(n4512), .ZN(U3253)
         );
  AOI211_X1 U5057 ( .C1(n2039), .C2(n4516), .A(n4515), .B(n4541), .ZN(n4517)
         );
  AOI211_X1 U5058 ( .C1(n4527), .C2(ADDR_REG_15__SCAN_IN), .A(n4518), .B(n4517), .ZN(n4524) );
  AOI21_X1 U5059 ( .B1(n4521), .B2(n4520), .A(n4519), .ZN(n4522) );
  NAND2_X1 U5060 ( .A1(n4535), .A2(n4522), .ZN(n4523) );
  OAI211_X1 U5061 ( .C1(n4540), .C2(n4581), .A(n4524), .B(n4523), .ZN(U3255)
         );
  INV_X1 U5062 ( .A(n4525), .ZN(n4526) );
  AOI21_X1 U5063 ( .B1(n4527), .B2(ADDR_REG_16__SCAN_IN), .A(n4526), .ZN(n4539) );
  OAI21_X1 U5064 ( .B1(n4530), .B2(n4529), .A(n4528), .ZN(n4536) );
  OAI21_X1 U5065 ( .B1(n4533), .B2(n4532), .A(n4531), .ZN(n4534) );
  AOI22_X1 U5066 ( .A1(n4537), .A2(n4536), .B1(n4535), .B2(n4534), .ZN(n4538)
         );
  OAI211_X1 U5067 ( .C1(n4579), .C2(n4540), .A(n4539), .B(n4538), .ZN(U3256)
         );
  INV_X1 U5068 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U5069 ( .A1(n4548), .A2(n4576), .ZN(n4549) );
  AOI22_X1 U5070 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4276), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4566), .ZN(n4560) );
  INV_X1 U5071 ( .A(n4555), .ZN(n4556) );
  AOI22_X1 U5072 ( .A1(n4558), .A2(n4568), .B1(n4557), .B2(n4556), .ZN(n4559)
         );
  OAI211_X1 U5073 ( .C1(n4280), .C2(n4561), .A(n4560), .B(n4559), .ZN(U3288)
         );
  INV_X1 U5074 ( .A(n4562), .ZN(n4564) );
  AOI21_X1 U5075 ( .B1(n4565), .B2(n4564), .A(n4563), .ZN(n4571) );
  AOI22_X1 U5076 ( .A1(n4568), .A2(n4567), .B1(REG3_REG_0__SCAN_IN), .B2(n4566), .ZN(n4569) );
  OAI221_X1 U5077 ( .B1(n4280), .B2(n4571), .C1(n4570), .C2(n2413), .A(n4569), 
        .ZN(U3290) );
  AND2_X1 U5078 ( .A1(D_REG_31__SCAN_IN), .A2(n4573), .ZN(U3291) );
  AND2_X1 U5079 ( .A1(D_REG_30__SCAN_IN), .A2(n4573), .ZN(U3292) );
  AND2_X1 U5080 ( .A1(D_REG_29__SCAN_IN), .A2(n4573), .ZN(U3293) );
  AND2_X1 U5081 ( .A1(D_REG_28__SCAN_IN), .A2(n4573), .ZN(U3294) );
  AND2_X1 U5082 ( .A1(D_REG_27__SCAN_IN), .A2(n4573), .ZN(U3295) );
  AND2_X1 U5083 ( .A1(D_REG_26__SCAN_IN), .A2(n4573), .ZN(U3296) );
  AND2_X1 U5084 ( .A1(D_REG_25__SCAN_IN), .A2(n4573), .ZN(U3297) );
  AND2_X1 U5085 ( .A1(D_REG_24__SCAN_IN), .A2(n4573), .ZN(U3298) );
  AND2_X1 U5086 ( .A1(D_REG_23__SCAN_IN), .A2(n4573), .ZN(U3299) );
  AND2_X1 U5087 ( .A1(D_REG_22__SCAN_IN), .A2(n4573), .ZN(U3300) );
  INV_X1 U5088 ( .A(n4573), .ZN(n4572) );
  INV_X1 U5089 ( .A(D_REG_21__SCAN_IN), .ZN(n4682) );
  NOR2_X1 U5090 ( .A1(n4572), .A2(n4682), .ZN(U3301) );
  AND2_X1 U5091 ( .A1(D_REG_20__SCAN_IN), .A2(n4573), .ZN(U3302) );
  AND2_X1 U5092 ( .A1(D_REG_19__SCAN_IN), .A2(n4573), .ZN(U3303) );
  AND2_X1 U5093 ( .A1(D_REG_18__SCAN_IN), .A2(n4573), .ZN(U3304) );
  AND2_X1 U5094 ( .A1(D_REG_17__SCAN_IN), .A2(n4573), .ZN(U3305) );
  AND2_X1 U5095 ( .A1(D_REG_16__SCAN_IN), .A2(n4573), .ZN(U3306) );
  INV_X1 U5096 ( .A(D_REG_15__SCAN_IN), .ZN(n4713) );
  NOR2_X1 U5097 ( .A1(n4572), .A2(n4713), .ZN(U3307) );
  AND2_X1 U5098 ( .A1(D_REG_14__SCAN_IN), .A2(n4573), .ZN(U3308) );
  AND2_X1 U5099 ( .A1(D_REG_13__SCAN_IN), .A2(n4573), .ZN(U3309) );
  AND2_X1 U5100 ( .A1(D_REG_12__SCAN_IN), .A2(n4573), .ZN(U3310) );
  AND2_X1 U5101 ( .A1(D_REG_11__SCAN_IN), .A2(n4573), .ZN(U3311) );
  AND2_X1 U5102 ( .A1(D_REG_10__SCAN_IN), .A2(n4573), .ZN(U3312) );
  AND2_X1 U5103 ( .A1(D_REG_9__SCAN_IN), .A2(n4573), .ZN(U3313) );
  AND2_X1 U5104 ( .A1(D_REG_8__SCAN_IN), .A2(n4573), .ZN(U3314) );
  AND2_X1 U5105 ( .A1(D_REG_7__SCAN_IN), .A2(n4573), .ZN(U3315) );
  INV_X1 U5106 ( .A(D_REG_6__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5107 ( .A1(n4572), .A2(n4714), .ZN(U3316) );
  AND2_X1 U5108 ( .A1(D_REG_5__SCAN_IN), .A2(n4573), .ZN(U3317) );
  INV_X1 U5109 ( .A(D_REG_4__SCAN_IN), .ZN(n4665) );
  NOR2_X1 U5110 ( .A1(n4572), .A2(n4665), .ZN(U3318) );
  AND2_X1 U5111 ( .A1(D_REG_3__SCAN_IN), .A2(n4573), .ZN(U3319) );
  AND2_X1 U5112 ( .A1(D_REG_2__SCAN_IN), .A2(n4573), .ZN(U3320) );
  OAI21_X1 U5113 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4574), .ZN(
        n4575) );
  INV_X1 U5114 ( .A(n4575), .ZN(U3329) );
  OAI22_X1 U5115 ( .A1(U3149), .A2(n4576), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4577) );
  INV_X1 U5116 ( .A(n4577), .ZN(U3334) );
  INV_X1 U5117 ( .A(DATAI_16_), .ZN(n4578) );
  AOI22_X1 U5118 ( .A1(STATE_REG_SCAN_IN), .A2(n4579), .B1(n4578), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5119 ( .A(DATAI_15_), .ZN(n4580) );
  AOI22_X1 U5120 ( .A1(STATE_REG_SCAN_IN), .A2(n4581), .B1(n4580), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5121 ( .A1(U3149), .A2(n4582), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4583) );
  INV_X1 U5122 ( .A(n4583), .ZN(U3339) );
  AOI22_X1 U5123 ( .A1(n4612), .A2(n4584), .B1(n2412), .B2(n4610), .ZN(U3467)
         );
  AOI22_X1 U5124 ( .A1(n4612), .A2(n4585), .B1(n2226), .B2(n4610), .ZN(U3469)
         );
  NOR2_X1 U5125 ( .A1(n4587), .A2(n4586), .ZN(n4589) );
  AOI211_X1 U5126 ( .C1(n4602), .C2(n4590), .A(n4589), .B(n4588), .ZN(n4614)
         );
  AOI22_X1 U5127 ( .A1(n4612), .A2(n4614), .B1(n2450), .B2(n4610), .ZN(U3473)
         );
  INV_X1 U5128 ( .A(n4591), .ZN(n4596) );
  INV_X1 U5129 ( .A(n4592), .ZN(n4594) );
  AOI211_X1 U5130 ( .C1(n4596), .C2(n4595), .A(n4594), .B(n4593), .ZN(n4616)
         );
  AOI22_X1 U5131 ( .A1(n4612), .A2(n4616), .B1(n2466), .B2(n4610), .ZN(U3475)
         );
  NOR2_X1 U5132 ( .A1(n4597), .A2(n4604), .ZN(n4600) );
  INV_X1 U5133 ( .A(n4598), .ZN(n4599) );
  AOI211_X1 U5134 ( .C1(n4602), .C2(n4601), .A(n4600), .B(n4599), .ZN(n4617)
         );
  INV_X1 U5135 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5136 ( .A1(n4612), .A2(n4617), .B1(n4603), .B2(n4610), .ZN(U3477)
         );
  NOR2_X1 U5137 ( .A1(n4605), .A2(n4604), .ZN(n4609) );
  AOI211_X1 U5138 ( .C1(n4609), .C2(n4608), .A(n4607), .B(n4606), .ZN(n4618)
         );
  INV_X1 U5139 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4611) );
  AOI22_X1 U5140 ( .A1(n4612), .A2(n4618), .B1(n4611), .B2(n4610), .ZN(U3481)
         );
  INV_X1 U5141 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4613) );
  AOI22_X1 U5142 ( .A1(n4619), .A2(n4614), .B1(n4613), .B2(n4334), .ZN(U3521)
         );
  INV_X1 U5143 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4615) );
  AOI22_X1 U5144 ( .A1(n4619), .A2(n4616), .B1(n4615), .B2(n4334), .ZN(U3522)
         );
  AOI22_X1 U5145 ( .A1(n4619), .A2(n4617), .B1(n2493), .B2(n4334), .ZN(U3523)
         );
  AOI22_X1 U5146 ( .A1(n4619), .A2(n4618), .B1(n2530), .B2(n4334), .ZN(U3525)
         );
  NOR4_X1 U5147 ( .A1(REG2_REG_12__SCAN_IN), .A2(REG2_REG_10__SCAN_IN), .A3(
        ADDR_REG_10__SCAN_IN), .A4(n3363), .ZN(n4623) );
  NOR4_X1 U5148 ( .A1(REG1_REG_1__SCAN_IN), .A2(n2493), .A3(n4620), .A4(n3091), 
        .ZN(n4622) );
  NOR3_X1 U5149 ( .A1(REG0_REG_21__SCAN_IN), .A2(REG1_REG_8__SCAN_IN), .A3(
        n4719), .ZN(n4621) );
  NAND4_X1 U5150 ( .A1(D_REG_6__SCAN_IN), .A2(n4623), .A3(n4622), .A4(n4621), 
        .ZN(n4631) );
  NOR4_X1 U5151 ( .A1(DATAI_9_), .A2(REG1_REG_23__SCAN_IN), .A3(
        REG2_REG_24__SCAN_IN), .A4(n4665), .ZN(n4626) );
  NOR3_X1 U5152 ( .A1(REG3_REG_4__SCAN_IN), .A2(DATAO_REG_1__SCAN_IN), .A3(
        DATAO_REG_10__SCAN_IN), .ZN(n4625) );
  NOR4_X1 U5153 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .A3(
        IR_REG_12__SCAN_IN), .A4(REG3_REG_27__SCAN_IN), .ZN(n4624) );
  NAND4_X1 U5154 ( .A1(n4626), .A2(DATAO_REG_28__SCAN_IN), .A3(n4625), .A4(
        n4624), .ZN(n4630) );
  NAND4_X1 U5155 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG2_REG_26__SCAN_IN), .A3(
        ADDR_REG_6__SCAN_IN), .A4(n4678), .ZN(n4629) );
  NAND4_X1 U5156 ( .A1(n4627), .A2(n4730), .A3(IR_REG_17__SCAN_IN), .A4(
        REG3_REG_12__SCAN_IN), .ZN(n4628) );
  NOR4_X1 U5157 ( .A1(n4631), .A2(n4630), .A3(n4629), .A4(n4628), .ZN(n4773)
         );
  INV_X1 U5158 ( .A(DATAI_12_), .ZN(n4632) );
  NAND3_X1 U5159 ( .A1(DATAO_REG_16__SCAN_IN), .A2(DATAO_REG_31__SCAN_IN), 
        .A3(n4632), .ZN(n4644) );
  NAND3_X1 U5160 ( .A1(REG3_REG_22__SCAN_IN), .A2(ADDR_REG_12__SCAN_IN), .A3(
        n3123), .ZN(n4643) );
  NOR4_X1 U5161 ( .A1(n4634), .A2(n4633), .A3(REG3_REG_3__SCAN_IN), .A4(
        DATAI_5_), .ZN(n4637) );
  NOR2_X1 U5162 ( .A1(n4635), .A2(n4669), .ZN(n4636) );
  NAND4_X1 U5163 ( .A1(n4637), .A2(IR_REG_1__SCAN_IN), .A3(n2662), .A4(n4636), 
        .ZN(n4642) );
  INV_X1 U5164 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4639) );
  NAND4_X1 U5165 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(REG0_REG_9__SCAN_IN), .ZN(n4641) );
  OR4_X1 U5166 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), .ZN(n4652) );
  NOR4_X1 U5167 ( .A1(IR_REG_25__SCAN_IN), .A2(REG0_REG_23__SCAN_IN), .A3(
        n4645), .A4(n4758), .ZN(n4648) );
  NOR4_X1 U5168 ( .A1(DATAO_REG_19__SCAN_IN), .A2(D_REG_1__SCAN_IN), .A3(
        DATAO_REG_24__SCAN_IN), .A4(n4753), .ZN(n4647) );
  NOR3_X1 U5169 ( .A1(IR_REG_21__SCAN_IN), .A2(DATAI_16_), .A3(
        ADDR_REG_18__SCAN_IN), .ZN(n4646) );
  NAND4_X1 U5170 ( .A1(DATAI_25_), .A2(n4648), .A3(n4647), .A4(n4646), .ZN(
        n4651) );
  INV_X1 U5171 ( .A(n4649), .ZN(n4650) );
  NOR3_X1 U5172 ( .A1(n4652), .A2(n4651), .A3(n4650), .ZN(n4772) );
  AOI22_X1 U5173 ( .A1(n4654), .A2(keyinput21), .B1(keyinput6), .B2(n3123), 
        .ZN(n4653) );
  OAI221_X1 U5174 ( .B1(n4654), .B2(keyinput21), .C1(n3123), .C2(keyinput6), 
        .A(n4653), .ZN(n4663) );
  INV_X1 U5175 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4656) );
  AOI22_X1 U5176 ( .A1(n4656), .A2(keyinput23), .B1(n4639), .B2(keyinput18), 
        .ZN(n4655) );
  OAI221_X1 U5177 ( .B1(n4656), .B2(keyinput23), .C1(n4639), .C2(keyinput18), 
        .A(n4655), .ZN(n4662) );
  XOR2_X1 U5178 ( .A(n4633), .B(keyinput7), .Z(n4660) );
  XOR2_X1 U5179 ( .A(n2662), .B(keyinput5), .Z(n4659) );
  XNOR2_X1 U5180 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput1), .ZN(n4658) );
  XNOR2_X1 U5181 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput39), .ZN(n4657) );
  NAND4_X1 U5182 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), .ZN(n4661)
         );
  NOR3_X1 U5183 ( .A1(n4663), .A2(n4662), .A3(n4661), .ZN(n4711) );
  INV_X1 U5184 ( .A(DATAI_9_), .ZN(n4666) );
  AOI22_X1 U5185 ( .A1(n4666), .A2(keyinput31), .B1(n4665), .B2(keyinput3), 
        .ZN(n4664) );
  OAI221_X1 U5186 ( .B1(n4666), .B2(keyinput31), .C1(n4665), .C2(keyinput3), 
        .A(n4664), .ZN(n4676) );
  AOI22_X1 U5187 ( .A1(n4634), .A2(keyinput55), .B1(keyinput19), .B2(n4668), 
        .ZN(n4667) );
  OAI221_X1 U5188 ( .B1(n4634), .B2(keyinput55), .C1(n4668), .C2(keyinput19), 
        .A(n4667), .ZN(n4675) );
  XNOR2_X1 U5189 ( .A(IR_REG_1__SCAN_IN), .B(keyinput47), .ZN(n4673) );
  XNOR2_X1 U5190 ( .A(REG0_REG_14__SCAN_IN), .B(keyinput27), .ZN(n4672) );
  XNOR2_X1 U5191 ( .A(n4669), .B(keyinput63), .ZN(n4671) );
  XNOR2_X1 U5192 ( .A(IR_REG_6__SCAN_IN), .B(keyinput16), .ZN(n4670) );
  NAND4_X1 U5193 ( .A1(n4673), .A2(n4672), .A3(n4671), .A4(n4670), .ZN(n4674)
         );
  NOR3_X1 U5194 ( .A1(n4676), .A2(n4675), .A3(n4674), .ZN(n4710) );
  AOI22_X1 U5195 ( .A1(n4679), .A2(keyinput17), .B1(n4678), .B2(keyinput12), 
        .ZN(n4677) );
  OAI221_X1 U5196 ( .B1(n4679), .B2(keyinput17), .C1(n4678), .C2(keyinput12), 
        .A(n4677), .ZN(n4691) );
  AOI22_X1 U5197 ( .A1(n4682), .A2(keyinput59), .B1(keyinput51), .B2(n4681), 
        .ZN(n4680) );
  OAI221_X1 U5198 ( .B1(n4682), .B2(keyinput59), .C1(n4681), .C2(keyinput51), 
        .A(n4680), .ZN(n4690) );
  AOI22_X1 U5199 ( .A1(n4685), .A2(keyinput11), .B1(n4684), .B2(keyinput15), 
        .ZN(n4683) );
  OAI221_X1 U5200 ( .B1(n4685), .B2(keyinput11), .C1(n4684), .C2(keyinput15), 
        .A(n4683), .ZN(n4689) );
  XNOR2_X1 U5201 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput10), .ZN(n4687) );
  XNOR2_X1 U5202 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput14), .ZN(n4686) );
  NAND2_X1 U5203 ( .A1(n4687), .A2(n4686), .ZN(n4688) );
  NOR4_X1 U5204 ( .A1(n4691), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4709)
         );
  XNOR2_X1 U5205 ( .A(n4692), .B(keyinput0), .ZN(n4697) );
  XNOR2_X1 U5206 ( .A(n4693), .B(keyinput4), .ZN(n4696) );
  XNOR2_X1 U5207 ( .A(n4694), .B(keyinput35), .ZN(n4695) );
  NOR3_X1 U5208 ( .A1(n4697), .A2(n4696), .A3(n4695), .ZN(n4700) );
  XNOR2_X1 U5209 ( .A(IR_REG_12__SCAN_IN), .B(keyinput43), .ZN(n4699) );
  XNOR2_X1 U5210 ( .A(IR_REG_26__SCAN_IN), .B(keyinput2), .ZN(n4698) );
  NAND3_X1 U5211 ( .A1(n4700), .A2(n4699), .A3(n4698), .ZN(n4707) );
  AOI22_X1 U5212 ( .A1(n4703), .A2(keyinput13), .B1(keyinput9), .B2(n4702), 
        .ZN(n4701) );
  OAI221_X1 U5213 ( .B1(n4703), .B2(keyinput13), .C1(n4702), .C2(keyinput9), 
        .A(n4701), .ZN(n4706) );
  XNOR2_X1 U5214 ( .A(n4704), .B(keyinput8), .ZN(n4705) );
  NOR3_X1 U5215 ( .A1(n4707), .A2(n4706), .A3(n4705), .ZN(n4708) );
  NAND4_X1 U5216 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4771)
         );
  AOI22_X1 U5217 ( .A1(n4714), .A2(keyinput40), .B1(n4713), .B2(keyinput62), 
        .ZN(n4712) );
  OAI221_X1 U5218 ( .B1(n4714), .B2(keyinput40), .C1(n4713), .C2(keyinput62), 
        .A(n4712), .ZN(n4725) );
  AOI22_X1 U5219 ( .A1(n2493), .A2(keyinput49), .B1(n4716), .B2(keyinput22), 
        .ZN(n4715) );
  OAI221_X1 U5220 ( .B1(n2493), .B2(keyinput49), .C1(n4716), .C2(keyinput22), 
        .A(n4715), .ZN(n4724) );
  AOI22_X1 U5221 ( .A1(n4719), .A2(keyinput50), .B1(keyinput41), .B2(n4718), 
        .ZN(n4717) );
  OAI221_X1 U5222 ( .B1(n4719), .B2(keyinput50), .C1(n4718), .C2(keyinput41), 
        .A(n4717), .ZN(n4723) );
  XNOR2_X1 U5223 ( .A(REG1_REG_13__SCAN_IN), .B(keyinput48), .ZN(n4721) );
  XNOR2_X1 U5224 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput32), .ZN(n4720) );
  NAND2_X1 U5225 ( .A1(n4721), .A2(n4720), .ZN(n4722) );
  NOR4_X1 U5226 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .ZN(n4769)
         );
  AOI22_X1 U5227 ( .A1(n3935), .A2(keyinput53), .B1(keyinput57), .B2(n3091), 
        .ZN(n4726) );
  OAI221_X1 U5228 ( .B1(n3935), .B2(keyinput53), .C1(n3091), .C2(keyinput57), 
        .A(n4726), .ZN(n4737) );
  INV_X1 U5229 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4728) );
  AOI22_X1 U5230 ( .A1(n3409), .A2(keyinput28), .B1(keyinput26), .B2(n4728), 
        .ZN(n4727) );
  OAI221_X1 U5231 ( .B1(n3409), .B2(keyinput28), .C1(n4728), .C2(keyinput26), 
        .A(n4727), .ZN(n4736) );
  AOI22_X1 U5232 ( .A1(n4731), .A2(keyinput24), .B1(keyinput60), .B2(n4730), 
        .ZN(n4729) );
  OAI221_X1 U5233 ( .B1(n4731), .B2(keyinput24), .C1(n4730), .C2(keyinput60), 
        .A(n4729), .ZN(n4735) );
  XOR2_X1 U5234 ( .A(n3363), .B(keyinput56), .Z(n4733) );
  XNOR2_X1 U5235 ( .A(IR_REG_0__SCAN_IN), .B(keyinput54), .ZN(n4732) );
  NAND2_X1 U5236 ( .A1(n4733), .A2(n4732), .ZN(n4734) );
  NOR4_X1 U5237 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(n4768)
         );
  AOI22_X1 U5238 ( .A1(n4740), .A2(keyinput52), .B1(keyinput29), .B2(n4739), 
        .ZN(n4738) );
  OAI221_X1 U5239 ( .B1(n4740), .B2(keyinput52), .C1(n4739), .C2(keyinput29), 
        .A(n4738), .ZN(n4750) );
  INV_X1 U5240 ( .A(DATAI_25_), .ZN(n4742) );
  AOI22_X1 U5241 ( .A1(n4743), .A2(keyinput34), .B1(n4742), .B2(keyinput37), 
        .ZN(n4741) );
  OAI221_X1 U5242 ( .B1(n4743), .B2(keyinput34), .C1(n4742), .C2(keyinput37), 
        .A(n4741), .ZN(n4749) );
  XNOR2_X1 U5243 ( .A(DATAI_5_), .B(keyinput30), .ZN(n4747) );
  XNOR2_X1 U5244 ( .A(DATAI_16_), .B(keyinput33), .ZN(n4746) );
  XNOR2_X1 U5245 ( .A(IR_REG_21__SCAN_IN), .B(keyinput38), .ZN(n4745) );
  XNOR2_X1 U5246 ( .A(keyinput25), .B(DATAI_12_), .ZN(n4744) );
  NAND4_X1 U5247 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4748)
         );
  NOR3_X1 U5248 ( .A1(n4750), .A2(n4749), .A3(n4748), .ZN(n4767) );
  AOI22_X1 U5249 ( .A1(n4753), .A2(keyinput58), .B1(keyinput61), .B2(n4752), 
        .ZN(n4751) );
  OAI221_X1 U5250 ( .B1(n4753), .B2(keyinput58), .C1(n4752), .C2(keyinput61), 
        .A(n4751), .ZN(n4765) );
  AOI22_X1 U5251 ( .A1(n4756), .A2(keyinput45), .B1(n4755), .B2(keyinput46), 
        .ZN(n4754) );
  OAI221_X1 U5252 ( .B1(n4756), .B2(keyinput45), .C1(n4755), .C2(keyinput46), 
        .A(n4754), .ZN(n4764) );
  AOI22_X1 U5253 ( .A1(n4759), .A2(keyinput44), .B1(keyinput20), .B2(n4758), 
        .ZN(n4757) );
  OAI221_X1 U5254 ( .B1(n4759), .B2(keyinput44), .C1(n4758), .C2(keyinput20), 
        .A(n4757), .ZN(n4763) );
  XNOR2_X1 U5255 ( .A(REG0_REG_26__SCAN_IN), .B(keyinput36), .ZN(n4761) );
  XNOR2_X1 U5256 ( .A(IR_REG_25__SCAN_IN), .B(keyinput42), .ZN(n4760) );
  NAND2_X1 U5257 ( .A1(n4761), .A2(n4760), .ZN(n4762) );
  NOR4_X1 U5258 ( .A1(n4765), .A2(n4764), .A3(n4763), .A4(n4762), .ZN(n4766)
         );
  NAND4_X1 U5259 ( .A1(n4769), .A2(n4768), .A3(n4767), .A4(n4766), .ZN(n4770)
         );
  AOI211_X1 U5260 ( .C1(n4773), .C2(n4772), .A(n4771), .B(n4770), .ZN(n4778)
         );
  INV_X1 U5261 ( .A(n4774), .ZN(n4775) );
  NAND2_X1 U5262 ( .A1(n4775), .A2(U4043), .ZN(n4776) );
  OAI21_X1 U5263 ( .B1(U4043), .B2(DATAO_REG_29__SCAN_IN), .A(n4776), .ZN(
        n4777) );
  XNOR2_X1 U5264 ( .A(n4778), .B(n4777), .ZN(U3579) );
  INV_X1 U2251 ( .A(n3751), .ZN(n2936) );
  AND2_X1 U3145 ( .A1(n2500), .A2(n2372), .ZN(n2668) );
endmodule

