

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11149, n11150, n11151, n11152, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
         n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
         n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
         n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
         n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
         n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
         n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
         n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
         n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
         n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
         n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
         n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746,
         n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
         n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
         n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
         n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
         n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
         n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818,
         n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
         n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
         n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
         n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855;

  AND2_X1 U11257 ( .A1(n22255), .A2(n14315), .ZN(n22353) );
  NAND2_X1 U11258 ( .A1(n16549), .A2(n16550), .ZN(n16537) );
  NAND2_X1 U11259 ( .A1(n12641), .A2(n17636), .ZN(n17618) );
  INV_X2 U11260 ( .A(n11252), .ZN(n19396) );
  CLKBUF_X2 U11261 ( .A(n16494), .Z(n11155) );
  CLKBUF_X2 U11262 ( .A(n12159), .Z(n12196) );
  CLKBUF_X2 U11263 ( .A(n14404), .Z(n11164) );
  INV_X1 U11264 ( .A(n18616), .ZN(n18496) );
  CLKBUF_X2 U11265 ( .A(n14419), .Z(n18663) );
  CLKBUF_X1 U11266 ( .A(n18617), .Z(n11156) );
  CLKBUF_X3 U11267 ( .A(n18627), .Z(n18679) );
  AND2_X1 U11268 ( .A1(n11996), .A2(n15297), .ZN(n13950) );
  AND2_X1 U11269 ( .A1(n11996), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13948) );
  AND2_X1 U11270 ( .A1(n14175), .A2(n15297), .ZN(n13949) );
  AND2_X1 U11271 ( .A1(n13925), .A2(n11783), .ZN(n13963) );
  NOR2_X1 U11272 ( .A1(n14522), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n21625) );
  NAND2_X2 U11273 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14522) );
  NOR2_X1 U11274 ( .A1(n12064), .A2(n12772), .ZN(n12054) );
  NAND2_X2 U11275 ( .A1(n11588), .A2(n12046), .ZN(n12064) );
  INV_X1 U11277 ( .A(n12928), .ZN(n12981) );
  BUF_X1 U11278 ( .A(n12772), .Z(n11245) );
  BUF_X2 U11279 ( .A(n12931), .Z(n13694) );
  CLKBUF_X2 U11280 ( .A(n12956), .Z(n13651) );
  BUF_X1 U11281 ( .A(n13127), .Z(n13754) );
  INV_X2 U11282 ( .A(n12045), .ZN(n11590) );
  AND2_X1 U11283 ( .A1(n14826), .A2(n14822), .ZN(n13069) );
  AND2_X1 U11284 ( .A1(n12887), .A2(n14660), .ZN(n13027) );
  CLKBUF_X2 U11285 ( .A(n12956), .Z(n13584) );
  AND2_X2 U11286 ( .A1(n12887), .A2(n14826), .ZN(n12942) );
  CLKBUF_X1 U11287 ( .A(n22673), .Z(n11149) );
  CLKBUF_X1 U11288 ( .A(n22770), .Z(n11150) );
  AND4_X1 U11289 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12510) );
  AND2_X1 U11290 ( .A1(n12886), .A2(n14660), .ZN(n12966) );
  NAND2_X1 U11291 ( .A1(n16494), .A2(n14293), .ZN(n14286) );
  AND2_X1 U11292 ( .A1(n14822), .A2(n14660), .ZN(n13034) );
  NAND2_X1 U11293 ( .A1(n11273), .A2(n11774), .ZN(n14096) );
  AND2_X1 U11294 ( .A1(n13925), .A2(n11781), .ZN(n13957) );
  NAND2_X1 U11295 ( .A1(n12501), .A2(n12463), .ZN(n20128) );
  NOR2_X1 U11296 ( .A1(n21638), .A2(n14459), .ZN(n18627) );
  AND3_X1 U11297 ( .A1(n14686), .A2(n14931), .A3(n12975), .ZN(n14696) );
  AND2_X1 U11298 ( .A1(n14163), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12219) );
  AND2_X1 U11299 ( .A1(n14175), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13962) );
  NAND2_X1 U11300 ( .A1(n11743), .A2(n11343), .ZN(n11735) );
  INV_X1 U11301 ( .A(n15973), .ZN(n11159) );
  NAND2_X1 U11302 ( .A1(n12604), .A2(n15665), .ZN(n12605) );
  INV_X1 U11303 ( .A(n12529), .ZN(n20166) );
  OR2_X1 U11304 ( .A1(n12500), .A2(n12463), .ZN(n20111) );
  AND2_X1 U11305 ( .A1(n11992), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13956) );
  NAND2_X1 U11306 ( .A1(n15007), .A2(n11243), .ZN(n14295) );
  AND4_X1 U11307 ( .A1(n12960), .A2(n12959), .A3(n12958), .A4(n12957), .ZN(
        n12961) );
  NAND2_X2 U11308 ( .A1(n11299), .A2(n11723), .ZN(n14784) );
  NAND2_X1 U11309 ( .A1(n11734), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11732) );
  INV_X1 U11310 ( .A(n11683), .ZN(n12708) );
  NAND2_X1 U11311 ( .A1(n17826), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17783) );
  INV_X1 U11312 ( .A(n21341), .ZN(n21419) );
  INV_X1 U11313 ( .A(n21964), .ZN(n21985) );
  INV_X1 U11314 ( .A(n14777), .ZN(n16741) );
  XNOR2_X1 U11315 ( .A(n15986), .B(n15985), .ZN(n19449) );
  AND2_X2 U11316 ( .A1(n17567), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17826) );
  XNOR2_X1 U11317 ( .A(n12708), .B(n12707), .ZN(n17503) );
  CLKBUF_X3 U11318 ( .A(n13810), .Z(n19551) );
  INV_X1 U11319 ( .A(n21327), .ZN(n21341) );
  INV_X1 U11320 ( .A(n21533), .ZN(n21435) );
  INV_X1 U11321 ( .A(n22353), .ZN(n22383) );
  BUF_X1 U11323 ( .A(n18617), .Z(n11158) );
  AND2_X1 U11325 ( .A1(n12923), .A2(n12924), .ZN(n11151) );
  NAND4_X1 U11326 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n11244) );
  AND2_X2 U11327 ( .A1(n12831), .A2(n11368), .ZN(n12077) );
  NOR2_X4 U11328 ( .A1(n16904), .A2(n22205), .ZN(n11421) );
  AND2_X2 U11329 ( .A1(n11219), .A2(n11194), .ZN(n16904) );
  XNOR2_X2 U11330 ( .A(n13196), .B(n13205), .ZN(n13359) );
  NAND2_X1 U11331 ( .A1(n12456), .A2(n12472), .ZN(n12460) );
  NAND2_X2 U11333 ( .A1(n21618), .A2(n21624), .ZN(n14523) );
  XNOR2_X2 U11334 ( .A(n13200), .B(n15786), .ZN(n15571) );
  NAND2_X1 U11335 ( .A1(n15963), .A2(n11719), .ZN(n15973) );
  CLKBUF_X3 U11336 ( .A(n12032), .Z(n11242) );
  AND2_X1 U11337 ( .A1(n15300), .A2(n13925), .ZN(n13964) );
  BUF_X2 U11338 ( .A(n12792), .Z(n12800) );
  XNOR2_X2 U11339 ( .A(n11418), .B(n12608), .ZN(n12792) );
  OAI21_X2 U11340 ( .B1(n11159), .B2(n11488), .A(n11486), .ZN(n17451) );
  OAI21_X2 U11341 ( .B1(n13344), .B2(n13258), .A(n13191), .ZN(n13192) );
  AND2_X1 U11344 ( .A1(n14784), .A2(n11244), .ZN(n16494) );
  XNOR2_X2 U11345 ( .A(n12094), .B(n12095), .ZN(n12457) );
  NOR2_X1 U11347 ( .A1(n14523), .A2(n14515), .ZN(n18617) );
  OAI211_X2 U11348 ( .C1(n11199), .C2(n11203), .A(n11197), .B(n11196), .ZN(
        n13313) );
  NAND2_X1 U11349 ( .A1(n11420), .A2(n11160), .ZN(n11645) );
  AOI21_X1 U11350 ( .B1(n13232), .B2(n13231), .A(n11160), .ZN(n16905) );
  NOR2_X2 U11351 ( .A1(n16563), .A2(n16565), .ZN(n16549) );
  NAND2_X1 U11352 ( .A1(n12797), .A2(n12796), .ZN(n11586) );
  NOR3_X1 U11353 ( .A1(n17262), .A2(n11345), .A3(n17182), .ZN(n12202) );
  OR2_X1 U11354 ( .A1(n12633), .A2(n12798), .ZN(n11382) );
  AOI211_X1 U11355 ( .C1(n21964), .C2(n22008), .A(n21819), .B(n21947), .ZN(
        n22037) );
  OAI21_X1 U11356 ( .B1(n11636), .B2(n13230), .A(n11160), .ZN(n11220) );
  INV_X1 U11357 ( .A(n12575), .ZN(n20121) );
  NAND2_X1 U11358 ( .A1(n14974), .A2(n14973), .ZN(n14972) );
  INV_X1 U11359 ( .A(n12622), .ZN(n20154) );
  NAND2_X1 U11360 ( .A1(n12494), .A2(n12493), .ZN(n12568) );
  NOR2_X1 U11361 ( .A1(n18879), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18878) );
  AND2_X1 U11362 ( .A1(n13831), .A2(n13809), .ZN(n14899) );
  NOR2_X1 U11363 ( .A1(n22562), .A2(n15198), .ZN(n22776) );
  NOR2_X1 U11364 ( .A1(n15050), .A2(n15392), .ZN(n22834) );
  AND2_X1 U11365 ( .A1(n12695), .A2(n12696), .ZN(n12702) );
  OAI21_X1 U11366 ( .B1(n17159), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13080), 
        .ZN(n13151) );
  NAND2_X1 U11367 ( .A1(n13066), .A2(n13067), .ZN(n17974) );
  NAND2_X1 U11368 ( .A1(n11162), .A2(n11180), .ZN(n13065) );
  AOI21_X1 U11369 ( .B1(n12098), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n12090), .ZN(n12094) );
  INV_X1 U11370 ( .A(n11251), .ZN(n11253) );
  INV_X1 U11371 ( .A(n11737), .ZN(n11251) );
  AND2_X1 U11372 ( .A1(n11235), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U11373 ( .A1(n13055), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11203) );
  NAND2_X1 U11374 ( .A1(n14685), .A2(n11208), .ZN(n17167) );
  NAND2_X1 U11375 ( .A1(n12855), .A2(n14653), .ZN(n12079) );
  INV_X4 U11376 ( .A(n12192), .ZN(n16023) );
  NAND2_X1 U11377 ( .A1(n12029), .A2(n12028), .ZN(n12053) );
  AND2_X1 U11378 ( .A1(n11736), .A2(n11499), .ZN(n11734) );
  CLKBUF_X2 U11379 ( .A(n12255), .Z(n16040) );
  NOR2_X2 U11380 ( .A1(n19739), .A2(n19698), .ZN(n21439) );
  NOR2_X2 U11381 ( .A1(n11735), .A2(n19375), .ZN(n11736) );
  NAND2_X1 U11382 ( .A1(n12045), .A2(n12041), .ZN(n12772) );
  INV_X2 U11383 ( .A(n15778), .ZN(n11588) );
  INV_X1 U11384 ( .A(n14784), .ZN(n14986) );
  NOR2_X1 U11385 ( .A1(n11757), .A2(n11518), .ZN(n11744) );
  NAND3_X2 U11386 ( .A1(n12899), .A2(n12898), .A3(n11722), .ZN(n14770) );
  AND4_X1 U11387 ( .A1(n12946), .A2(n12945), .A3(n12944), .A4(n12943), .ZN(
        n12964) );
  AND4_X1 U11388 ( .A1(n12894), .A2(n12893), .A3(n12892), .A4(n12891), .ZN(
        n12899) );
  CLKBUF_X2 U11389 ( .A(n11968), .Z(n14176) );
  BUF_X2 U11390 ( .A(n13069), .Z(n13756) );
  CLKBUF_X2 U11391 ( .A(n13523), .Z(n13765) );
  CLKBUF_X3 U11392 ( .A(n14372), .Z(n11163) );
  BUF_X2 U11393 ( .A(n13376), .Z(n13764) );
  BUF_X2 U11394 ( .A(n13604), .Z(n13766) );
  CLKBUF_X2 U11395 ( .A(n12900), .Z(n13755) );
  CLKBUF_X2 U11396 ( .A(n13028), .Z(n13757) );
  CLKBUF_X2 U11397 ( .A(n13027), .Z(n13767) );
  INV_X1 U11398 ( .A(n21625), .ZN(n14459) );
  CLKBUF_X2 U11399 ( .A(n13034), .Z(n13739) );
  BUF_X2 U11400 ( .A(n12966), .Z(n13619) );
  BUF_X1 U11401 ( .A(n12886), .Z(n17162) );
  NAND2_X1 U11402 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14340) );
  INV_X1 U11403 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11416) );
  AND2_X1 U11404 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14660) );
  INV_X4 U11405 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11476) );
  BUF_X1 U11406 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11237) );
  AOI21_X1 U11407 ( .B1(n17416), .B2(n19537), .A(n16047), .ZN(n16048) );
  AND2_X1 U11408 ( .A1(n16021), .A2(n16020), .ZN(n17416) );
  AOI211_X1 U11409 ( .C1(n18088), .C2(n19450), .A(n17461), .B(n17460), .ZN(
        n17462) );
  OAI21_X1 U11410 ( .B1(n12879), .B2(n18063), .A(n12878), .ZN(n12880) );
  OAI21_X1 U11411 ( .B1(n12879), .B2(n17944), .A(n12864), .ZN(n12865) );
  NOR2_X1 U11412 ( .A1(n17436), .A2(n17435), .ZN(n17669) );
  OAI21_X1 U11413 ( .B1(n17419), .B2(n17422), .A(n11309), .ZN(n16017) );
  AND2_X1 U11414 ( .A1(n16057), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17444) );
  AND2_X1 U11415 ( .A1(n17458), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16057) );
  OAI211_X1 U11416 ( .C1(n16841), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16850), .B(n16840), .ZN(n16842) );
  AND2_X1 U11417 ( .A1(n17477), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17458) );
  NOR2_X1 U11418 ( .A1(n17902), .A2(n17894), .ZN(n17893) );
  XNOR2_X1 U11419 ( .A(n11172), .B(n17016), .ZN(n17021) );
  OAI21_X1 U11420 ( .B1(n16861), .B2(n20853), .A(n11407), .ZN(n11406) );
  NAND2_X1 U11421 ( .A1(n16525), .A2(n16526), .ZN(n16861) );
  OAI211_X1 U11422 ( .C1(n11176), .C2(n11175), .A(n11174), .B(n11173), .ZN(
        n11172) );
  NAND2_X1 U11423 ( .A1(n11439), .A2(n11294), .ZN(n16839) );
  AND2_X1 U11424 ( .A1(n14094), .A2(n14093), .ZN(n14116) );
  XNOR2_X1 U11425 ( .A(n11296), .B(n13788), .ZN(n16743) );
  NAND2_X1 U11426 ( .A1(n11176), .A2(n17024), .ZN(n11174) );
  NOR2_X1 U11427 ( .A1(n16897), .A2(n16856), .ZN(n11176) );
  XNOR2_X1 U11428 ( .A(n11411), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20848) );
  NOR2_X1 U11429 ( .A1(n16537), .A2(n16538), .ZN(n16536) );
  AOI21_X1 U11430 ( .B1(n11267), .B2(n11579), .A(n11314), .ZN(n11574) );
  CLKBUF_X1 U11431 ( .A(n16563), .Z(n16564) );
  AND2_X1 U11432 ( .A1(n16925), .A2(n16916), .ZN(n17083) );
  AND2_X1 U11433 ( .A1(n11577), .A2(n17622), .ZN(n11267) );
  NAND2_X1 U11434 ( .A1(n16027), .A2(n12205), .ZN(n17651) );
  NAND2_X1 U11435 ( .A1(n11183), .A2(n11636), .ZN(n16914) );
  XNOR2_X1 U11436 ( .A(n16027), .B(n16026), .ZN(n17241) );
  OR2_X1 U11437 ( .A1(n11584), .A2(n12794), .ZN(n11583) );
  INV_X1 U11438 ( .A(n11586), .ZN(n11584) );
  OR2_X1 U11439 ( .A1(n12806), .A2(n17935), .ZN(n17632) );
  CLKBUF_X1 U11440 ( .A(n16942), .Z(n17137) );
  NAND2_X1 U11441 ( .A1(n12202), .A2(n12201), .ZN(n16027) );
  NAND2_X1 U11442 ( .A1(n16942), .A2(n11635), .ZN(n11183) );
  NAND2_X1 U11443 ( .A1(n17135), .A2(n13220), .ZN(n16942) );
  OR2_X1 U11444 ( .A1(n12804), .A2(n16007), .ZN(n12807) );
  OR2_X1 U11445 ( .A1(n11222), .A2(n15785), .ZN(n11221) );
  NAND2_X1 U11446 ( .A1(n17295), .A2(n17296), .ZN(n17286) );
  NAND2_X1 U11447 ( .A1(n12633), .A2(n12798), .ZN(n12804) );
  OAI21_X1 U11448 ( .B1(n11628), .B2(n11430), .A(n11410), .ZN(n11222) );
  NAND2_X1 U11449 ( .A1(n15670), .A2(n15671), .ZN(n11628) );
  NAND2_X1 U11450 ( .A1(n11177), .A2(n11223), .ZN(n15670) );
  NAND2_X1 U11451 ( .A1(n11226), .A2(n13193), .ZN(n15572) );
  NAND2_X1 U11452 ( .A1(n15474), .A2(n11178), .ZN(n11177) );
  AOI211_X1 U11453 ( .C1(n21964), .C2(n21963), .A(n21962), .B(n21961), .ZN(
        n21965) );
  NAND2_X1 U11454 ( .A1(n15474), .A2(n15473), .ZN(n11226) );
  NOR2_X1 U11455 ( .A1(n17312), .A2(n17311), .ZN(n12164) );
  NAND2_X1 U11456 ( .A1(n13182), .A2(n13181), .ZN(n15474) );
  AOI21_X1 U11457 ( .B1(n11487), .B2(n11495), .A(n11330), .ZN(n11486) );
  INV_X1 U11458 ( .A(n11220), .ZN(n11219) );
  NAND2_X1 U11459 ( .A1(n11216), .A2(n13174), .ZN(n15360) );
  NAND2_X1 U11460 ( .A1(n18944), .A2(n18943), .ZN(n21933) );
  XNOR2_X1 U11461 ( .A(n16002), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16055) );
  OAI211_X1 U11462 ( .C1(n11627), .C2(n11423), .A(n11217), .B(n15379), .ZN(
        n11216) );
  AND2_X1 U11463 ( .A1(n12599), .A2(n12598), .ZN(n12608) );
  INV_X1 U11464 ( .A(n11649), .ZN(n18944) );
  NOR2_X1 U11465 ( .A1(n16932), .A2(n13228), .ZN(n11636) );
  AND4_X1 U11466 ( .A1(n12619), .A2(n12618), .A3(n12617), .A4(n12616), .ZN(
        n12628) );
  NAND2_X1 U11467 ( .A1(n11218), .A2(n11627), .ZN(n11217) );
  INV_X1 U11468 ( .A(n16859), .ZN(n11173) );
  NOR2_X1 U11469 ( .A1(n11225), .A2(n11179), .ZN(n11178) );
  AOI21_X1 U11470 ( .B1(n15571), .B2(n11224), .A(n13201), .ZN(n11223) );
  AOI211_X1 U11471 ( .C1(n21964), .C2(n21785), .A(n21813), .B(n21784), .ZN(
        n21787) );
  OR2_X1 U11472 ( .A1(n16943), .A2(n17093), .ZN(n16932) );
  INV_X1 U11473 ( .A(n15571), .ZN(n11225) );
  AOI211_X1 U11474 ( .C1(n20154), .C2(n20253), .A(n20184), .B(n20601), .ZN(
        n20151) );
  AND4_X1 U11475 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        n12595) );
  AND2_X1 U11476 ( .A1(n11427), .A2(n11426), .ZN(n11218) );
  NOR2_X1 U11477 ( .A1(n15971), .A2(n15970), .ZN(n15972) );
  NOR3_X1 U11478 ( .A1(n18878), .A2(n21958), .A3(n18874), .ZN(n18927) );
  INV_X1 U11479 ( .A(n15473), .ZN(n11179) );
  AND2_X1 U11480 ( .A1(n13200), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13201) );
  INV_X1 U11481 ( .A(n13193), .ZN(n11224) );
  NAND2_X1 U11482 ( .A1(n13221), .A2(n16945), .ZN(n16960) );
  NAND2_X1 U11483 ( .A1(n15255), .A2(n15589), .ZN(n15588) );
  INV_X1 U11484 ( .A(n12621), .ZN(n20088) );
  NAND2_X1 U11485 ( .A1(n14888), .A2(n14887), .ZN(n11627) );
  OR2_X1 U11486 ( .A1(n13229), .A2(n22138), .ZN(n16945) );
  INV_X4 U11487 ( .A(n17134), .ZN(n11160) );
  NOR2_X1 U11488 ( .A1(n21539), .A2(n21540), .ZN(n21564) );
  NAND2_X1 U11489 ( .A1(n12459), .A2(n12463), .ZN(n12622) );
  NAND2_X1 U11490 ( .A1(n18873), .A2(n18753), .ZN(n18813) );
  NOR2_X1 U11491 ( .A1(n14906), .A2(n14966), .ZN(n14967) );
  NOR2_X1 U11492 ( .A1(n15050), .A2(n15197), .ZN(n22819) );
  OAI21_X1 U11493 ( .B1(n13328), .B2(n13258), .A(n13178), .ZN(n13180) );
  NAND2_X1 U11494 ( .A1(n13327), .A2(n13326), .ZN(n14973) );
  OAI21_X1 U11495 ( .B1(n13344), .B2(n13404), .A(n13343), .ZN(n15367) );
  CLKBUF_X1 U11496 ( .A(n12574), .Z(n20226) );
  XNOR2_X1 U11497 ( .A(n13165), .B(n22148), .ZN(n14888) );
  NAND2_X1 U11498 ( .A1(n18979), .A2(n19019), .ZN(n18873) );
  NAND2_X1 U11499 ( .A1(n11182), .A2(n13184), .ZN(n13328) );
  NAND2_X1 U11500 ( .A1(n13150), .A2(n13149), .ZN(n13165) );
  NOR2_X1 U11501 ( .A1(n15118), .A2(n22548), .ZN(n22803) );
  OR2_X1 U11502 ( .A1(n15196), .A2(n13404), .ZN(n13327) );
  NAND2_X1 U11503 ( .A1(n11417), .A2(n13134), .ZN(n13196) );
  NAND2_X1 U11504 ( .A1(n14768), .A2(n14767), .ZN(n14910) );
  NAND2_X1 U11505 ( .A1(n13176), .A2(n13175), .ZN(n11182) );
  AND2_X1 U11506 ( .A1(n14883), .A2(n14882), .ZN(n14905) );
  NAND2_X1 U11507 ( .A1(n13176), .A2(n13168), .ZN(n15196) );
  NAND2_X1 U11508 ( .A1(n18980), .A2(n22028), .ZN(n18979) );
  NAND2_X1 U11509 ( .A1(n14799), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13150) );
  INV_X1 U11510 ( .A(n13112), .ZN(n13176) );
  NAND2_X1 U11511 ( .A1(n13310), .A2(n13309), .ZN(n14768) );
  NOR3_X2 U11512 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n19112), .A3(n21619), 
        .ZN(n18964) );
  OAI21_X1 U11513 ( .B1(n13301), .B2(n13258), .A(n13164), .ZN(n14887) );
  NAND2_X1 U11514 ( .A1(n13112), .A2(n13111), .ZN(n13184) );
  NAND2_X1 U11515 ( .A1(n11212), .A2(n11209), .ZN(n14799) );
  AOI211_X1 U11516 ( .C1(n19551), .C2(n19550), .A(n19549), .B(n19548), .ZN(
        n19552) );
  AOI222_X2 U11517 ( .A1(n15040), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(n15433), 
        .B2(n15061), .C1(n17151), .C2(n22825), .ZN(n22824) );
  NAND2_X1 U11518 ( .A1(n11626), .A2(n12097), .ZN(n11587) );
  OAI21_X1 U11519 ( .B1(n11211), .B2(n11210), .A(n13148), .ZN(n11209) );
  NAND2_X1 U11520 ( .A1(n12476), .A2(n12475), .ZN(n17238) );
  CLKBUF_X1 U11521 ( .A(n14936), .Z(n11254) );
  INV_X1 U11522 ( .A(n14935), .ZN(n13100) );
  NOR2_X1 U11523 ( .A1(n22266), .A2(n11208), .ZN(n11207) );
  AOI222_X2 U11524 ( .A1(n15062), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(n22585), 
        .B2(n15061), .C1(n17151), .C2(n22597), .ZN(n22596) );
  NOR2_X2 U11525 ( .A1(n20959), .A2(n22101), .ZN(n19137) );
  NAND2_X1 U11526 ( .A1(n11184), .A2(n13054), .ZN(n13153) );
  INV_X1 U11527 ( .A(n13148), .ZN(n11161) );
  NAND2_X2 U11528 ( .A1(n16834), .A2(n14930), .ZN(n16837) );
  AOI221_X1 U11529 ( .B1(n22016), .B2(n21654), .C1(n21964), .C2(n21654), .A(
        n14492), .ZN(n22100) );
  CLKBUF_X1 U11530 ( .A(n14817), .Z(n22237) );
  INV_X1 U11531 ( .A(n11215), .ZN(n11211) );
  NAND2_X1 U11532 ( .A1(n11215), .A2(n11213), .ZN(n14857) );
  NAND2_X1 U11533 ( .A1(n13302), .A2(n13303), .ZN(n11184) );
  NAND2_X1 U11534 ( .A1(n13311), .A2(n13147), .ZN(n11215) );
  OAI21_X1 U11535 ( .B1(n13311), .B2(n13258), .A(n13147), .ZN(n14855) );
  NOR2_X1 U11536 ( .A1(n15187), .A2(n14986), .ZN(n22671) );
  NOR2_X1 U11537 ( .A1(n15187), .A2(n15025), .ZN(n22687) );
  OAI21_X1 U11538 ( .B1(n15394), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13012), 
        .ZN(n13051) );
  CLKBUF_X1 U11539 ( .A(n15394), .Z(n22611) );
  NOR2_X1 U11540 ( .A1(n19067), .A2(n21755), .ZN(n19066) );
  INV_X2 U11541 ( .A(n17309), .ZN(n15680) );
  INV_X2 U11542 ( .A(n21591), .ZN(n21600) );
  NAND2_X1 U11543 ( .A1(n13065), .A2(n13064), .ZN(n13066) );
  NAND2_X1 U11544 ( .A1(n13043), .A2(n13042), .ZN(n13145) );
  NAND2_X1 U11545 ( .A1(n13065), .A2(n15046), .ZN(n15394) );
  NOR2_X2 U11546 ( .A1(n20085), .A2(n20558), .ZN(n20086) );
  NOR2_X2 U11547 ( .A1(n20271), .A2(n20558), .ZN(n20272) );
  NAND2_X1 U11548 ( .A1(n13313), .A2(n22392), .ZN(n13043) );
  NOR2_X2 U11549 ( .A1(n20320), .A2(n20558), .ZN(n20321) );
  NOR2_X2 U11550 ( .A1(n20361), .A2(n20558), .ZN(n20362) );
  NOR2_X2 U11551 ( .A1(n20452), .A2(n20558), .ZN(n20453) );
  NOR2_X2 U11552 ( .A1(n20409), .A2(n20558), .ZN(n15775) );
  NAND2_X1 U11553 ( .A1(n12085), .A2(n12084), .ZN(n12454) );
  INV_X1 U11554 ( .A(n13001), .ZN(n11180) );
  OR2_X1 U11555 ( .A1(n19087), .A2(n11653), .ZN(n11652) );
  CLKBUF_X2 U11556 ( .A(n22067), .Z(n11250) );
  INV_X1 U11557 ( .A(n14987), .ZN(n11162) );
  NAND2_X1 U11558 ( .A1(n11203), .A2(n12992), .ZN(n11422) );
  CLKBUF_X3 U11559 ( .A(n12098), .Z(n16025) );
  NAND2_X1 U11560 ( .A1(n11200), .A2(n11198), .ZN(n11197) );
  INV_X1 U11561 ( .A(n11200), .ZN(n11199) );
  NOR2_X2 U11562 ( .A1(n14551), .A2(n19264), .ZN(n14552) );
  INV_X1 U11563 ( .A(n12991), .ZN(n13062) );
  INV_X1 U11564 ( .A(n13026), .ZN(n11200) );
  NAND2_X1 U11565 ( .A1(n12999), .A2(n11201), .ZN(n13026) );
  OAI21_X1 U11566 ( .B1(n11167), .B2(n11166), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11165) );
  INV_X1 U11567 ( .A(n11202), .ZN(n11201) );
  OAI211_X1 U11568 ( .C1(n16023), .C2(n12089), .A(n12088), .B(n12087), .ZN(
        n12090) );
  NAND2_X1 U11569 ( .A1(n11208), .A2(n12976), .ZN(n14795) );
  NAND2_X1 U11570 ( .A1(n12820), .A2(n12057), .ZN(n12067) );
  AND2_X1 U11571 ( .A1(n11549), .A2(n12642), .ZN(n11548) );
  NAND2_X1 U11572 ( .A1(n14198), .A2(n14986), .ZN(n11208) );
  CLKBUF_X1 U11573 ( .A(n14198), .Z(n16097) );
  AND2_X1 U11574 ( .A1(n11391), .A2(n11390), .ZN(n12820) );
  INV_X1 U11575 ( .A(n11213), .ZN(n11210) );
  NAND3_X1 U11576 ( .A1(n12053), .A2(n11589), .A3(n12030), .ZN(n12075) );
  NAND2_X1 U11577 ( .A1(n12998), .A2(n13044), .ZN(n11168) );
  NAND2_X1 U11578 ( .A1(n12024), .A2(n11311), .ZN(n12026) );
  INV_X1 U11579 ( .A(n12053), .ZN(n12833) );
  AOI21_X1 U11580 ( .B1(n13147), .B2(n13258), .A(n11214), .ZN(n11213) );
  INV_X1 U11581 ( .A(n12042), .ZN(n12058) );
  NAND2_X1 U11582 ( .A1(n12984), .A2(n12983), .ZN(n11166) );
  AND2_X1 U11583 ( .A1(n12551), .A2(n12550), .ZN(n12538) );
  AND2_X1 U11584 ( .A1(n14801), .A2(n16690), .ZN(n12983) );
  AND2_X1 U11585 ( .A1(n12829), .A2(n12055), .ZN(n11390) );
  OR2_X1 U11586 ( .A1(n19133), .A2(n19142), .ZN(n11658) );
  NAND2_X1 U11587 ( .A1(n14696), .A2(n11243), .ZN(n14722) );
  NAND2_X1 U11588 ( .A1(n12728), .A2(n12772), .ZN(n12829) );
  OR2_X1 U11589 ( .A1(n13293), .A2(n12987), .ZN(n14758) );
  INV_X1 U11590 ( .A(n11245), .ZN(n12721) );
  AND2_X2 U11591 ( .A1(n12239), .A2(n14139), .ZN(n16041) );
  OR2_X1 U11592 ( .A1(n12776), .A2(n20322), .ZN(n12247) );
  AOI21_X1 U11593 ( .B1(n12988), .B2(n11244), .A(n14819), .ZN(n11169) );
  NAND2_X1 U11594 ( .A1(n12981), .A2(n14770), .ZN(n14674) );
  AND3_X2 U11595 ( .A1(n11922), .A2(n11921), .A3(n11920), .ZN(n16007) );
  CLKBUF_X2 U11596 ( .A(n12928), .Z(n14771) );
  NAND2_X1 U11597 ( .A1(n13800), .A2(n12218), .ZN(n12030) );
  CLKBUF_X1 U11598 ( .A(n12032), .Z(n11241) );
  CLKBUF_X1 U11599 ( .A(n11589), .Z(n19264) );
  AND4_X1 U11600 ( .A1(n11866), .A2(n11865), .A3(n11864), .A4(n11863), .ZN(
        n11873) );
  INV_X1 U11601 ( .A(n12982), .ZN(n13044) );
  AND2_X1 U11602 ( .A1(n15016), .A2(n14777), .ZN(n14931) );
  INV_X1 U11603 ( .A(n15033), .ZN(n14772) );
  INV_X1 U11604 ( .A(n12041), .ZN(n11589) );
  OR2_X1 U11605 ( .A1(n14770), .A2(n15033), .ZN(n12980) );
  INV_X1 U11606 ( .A(n14786), .ZN(n15025) );
  NAND2_X2 U11607 ( .A1(n11981), .A2(n11980), .ZN(n12737) );
  AND4_X1 U11608 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11921) );
  NAND2_X1 U11609 ( .A1(n14770), .A2(n15033), .ZN(n13293) );
  OR2_X2 U11610 ( .A1(n20947), .A2(n20884), .ZN(n20933) );
  OR2_X2 U11611 ( .A1(n12919), .A2(n12918), .ZN(n14777) );
  MUX2_X1 U11612 ( .A(n11842), .B(n11841), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12041) );
  AND3_X2 U11613 ( .A1(n11204), .A2(n12922), .A3(n11151), .ZN(n15033) );
  NOR2_X1 U11614 ( .A1(n11192), .A2(n11190), .ZN(n11189) );
  OAI21_X1 U11615 ( .B1(n11953), .B2(n11952), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11954) );
  MUX2_X1 U11616 ( .A(n11941), .B(n11940), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15778) );
  NAND4_X1 U11617 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n12982) );
  NOR2_X1 U11618 ( .A1(n11186), .A2(n11185), .ZN(n11188) );
  AND4_X1 U11619 ( .A1(n12904), .A2(n12903), .A3(n12902), .A4(n12901), .ZN(
        n12909) );
  AND2_X2 U11620 ( .A1(n14176), .A2(n15297), .ZN(n13946) );
  NAND2_X1 U11621 ( .A1(n14160), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12404) );
  NOR2_X1 U11622 ( .A1(n11206), .A2(n11205), .ZN(n11204) );
  AND2_X1 U11623 ( .A1(n11987), .A2(n11986), .ZN(n11991) );
  AND4_X1 U11624 ( .A1(n12950), .A2(n12949), .A3(n12948), .A4(n12947), .ZN(
        n12963) );
  AND4_X1 U11625 ( .A1(n12955), .A2(n12954), .A3(n12953), .A4(n12952), .ZN(
        n12962) );
  INV_X2 U11626 ( .A(U214), .ZN(n20947) );
  AOI21_X1 U11627 ( .B1(n11968), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n11848), .ZN(n11852) );
  NAND2_X1 U11628 ( .A1(n11951), .A2(n11950), .ZN(n11952) );
  AND2_X1 U11629 ( .A1(n11631), .A2(n11634), .ZN(n11191) );
  INV_X1 U11630 ( .A(n12883), .ZN(n11192) );
  NAND2_X1 U11631 ( .A1(n12890), .A2(n11630), .ZN(n11185) );
  NAND2_X1 U11632 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11187) );
  INV_X2 U11633 ( .A(n14336), .ZN(n18644) );
  AND2_X2 U11634 ( .A1(n11784), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12300) );
  NAND2_X1 U11635 ( .A1(n12921), .A2(n12920), .ZN(n11206) );
  INV_X1 U11636 ( .A(n12992), .ZN(n11198) );
  CLKBUF_X3 U11637 ( .A(n18633), .Z(n18659) );
  CLKBUF_X3 U11638 ( .A(n18634), .Z(n18664) );
  CLKBUF_X3 U11639 ( .A(n18632), .Z(n18648) );
  AND2_X1 U11640 ( .A1(n11248), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11717) );
  CLKBUF_X2 U11641 ( .A(n14419), .Z(n18615) );
  AND2_X1 U11642 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11848) );
  CLKBUF_X2 U11643 ( .A(n11995), .Z(n11968) );
  INV_X1 U11644 ( .A(n13230), .ZN(n11195) );
  NAND2_X2 U11645 ( .A1(n22855), .A2(n22433), .ZN(n20780) );
  BUF_X2 U11646 ( .A(n13999), .Z(n14175) );
  AND2_X2 U11647 ( .A1(n11992), .A2(n15297), .ZN(n13947) );
  NOR2_X1 U11648 ( .A1(n20247), .A2(n20159), .ZN(n20601) );
  CLKBUF_X2 U11649 ( .A(n12931), .Z(n13656) );
  AND2_X2 U11651 ( .A1(n17162), .A2(n14826), .ZN(n13604) );
  NOR2_X1 U11652 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20137), .ZN(
        n20594) );
  AND2_X2 U11653 ( .A1(n12885), .A2(n14826), .ZN(n13376) );
  NOR2_X1 U11654 ( .A1(n14339), .A2(n14340), .ZN(n18630) );
  AND2_X2 U11656 ( .A1(n15264), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11249) );
  INV_X2 U11657 ( .A(n20674), .ZN(n20700) );
  NOR3_X1 U11658 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n14523), .ZN(n18677) );
  NAND2_X1 U11659 ( .A1(n21618), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14339) );
  OR2_X1 U11660 ( .A1(n16975), .A2(n16915), .ZN(n13230) );
  CLKBUF_X1 U11661 ( .A(n13626), .Z(n13782) );
  AND2_X1 U11662 ( .A1(n11553), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12887) );
  AND2_X1 U11663 ( .A1(n14818), .A2(n12886), .ZN(n12931) );
  NAND2_X2 U11664 ( .A1(n12212), .A2(n20222), .ZN(n19301) );
  AND2_X2 U11665 ( .A1(n11431), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14823) );
  AND2_X1 U11666 ( .A1(n16858), .A2(n17034), .ZN(n11175) );
  AND2_X2 U11667 ( .A1(n11416), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14826) );
  AND2_X2 U11668 ( .A1(n14818), .A2(n14822), .ZN(n13033) );
  INV_X1 U11669 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n11214) );
  AND4_X1 U11670 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11517) );
  NOR2_X2 U11671 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12886) );
  INV_X1 U11673 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11431) );
  AND2_X2 U11674 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14822) );
  INV_X1 U11675 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11782) );
  INV_X1 U11676 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15306) );
  NAND2_X2 U11677 ( .A1(n12991), .A2(n11165), .ZN(n13055) );
  NAND3_X1 U11678 ( .A1(n13000), .A2(n11169), .A3(n11168), .ZN(n11167) );
  NAND3_X1 U11679 ( .A1(n12941), .A2(n12993), .A3(n12940), .ZN(n12998) );
  OAI21_X2 U11680 ( .B1(n14795), .B2(n11170), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12991) );
  OAI21_X2 U11681 ( .B1(n14722), .B2(n14305), .A(n14806), .ZN(n11170) );
  NAND2_X1 U11682 ( .A1(n14987), .A2(n13001), .ZN(n15046) );
  XNOR2_X2 U11683 ( .A(n11181), .B(n13062), .ZN(n14987) );
  NAND2_X1 U11684 ( .A1(n11409), .A2(n12990), .ZN(n11181) );
  NAND2_X1 U11685 ( .A1(n11222), .A2(n15785), .ZN(n17135) );
  NAND3_X1 U11686 ( .A1(n11184), .A2(n13054), .A3(n13151), .ZN(n13167) );
  NAND3_X1 U11687 ( .A1(n12889), .A2(n11632), .A3(n11187), .ZN(n11186) );
  NAND3_X1 U11688 ( .A1(n11189), .A2(n11188), .A3(n12884), .ZN(n12928) );
  NAND3_X1 U11689 ( .A1(n12888), .A2(n11633), .A3(n11191), .ZN(n11190) );
  NAND2_X2 U11690 ( .A1(n13196), .A2(n13137), .ZN(n13229) );
  NAND2_X1 U11691 ( .A1(n13112), .A2(n11408), .ZN(n13195) );
  NOR2_X2 U11692 ( .A1(n13100), .A2(n13167), .ZN(n13112) );
  NOR2_X4 U11693 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14818) );
  OAI21_X2 U11694 ( .B1(n16871), .B2(n17004), .A(n11160), .ZN(n16840) );
  NAND4_X2 U11695 ( .A1(n11645), .A2(n11638), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(n11637), .ZN(n16871) );
  NAND3_X1 U11696 ( .A1(n11635), .A2(n16942), .A3(n11195), .ZN(n11194) );
  NAND3_X1 U11697 ( .A1(n11199), .A2(n11203), .A3(n12992), .ZN(n11196) );
  OAI21_X1 U11698 ( .B1(n13000), .B2(n14986), .A(n14680), .ZN(n11202) );
  NAND3_X1 U11699 ( .A1(n12925), .A2(n12926), .A3(n12927), .ZN(n11205) );
  NAND3_X1 U11700 ( .A1(n11161), .A2(n11215), .A3(n11213), .ZN(n11212) );
  NAND2_X1 U11701 ( .A1(n17135), .A2(n11221), .ZN(n15880) );
  OR2_X2 U11702 ( .A1(n12673), .A2(n11541), .ZN(n11291) );
  CLKBUF_X1 U11703 ( .A(n11401), .Z(n11227) );
  AND2_X1 U11704 ( .A1(n12506), .A2(n19551), .ZN(n11228) );
  NAND2_X1 U11705 ( .A1(n17826), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11229) );
  AOI21_X1 U11706 ( .B1(n13145), .B2(n13144), .A(n13135), .ZN(n13303) );
  OR2_X1 U11707 ( .A1(n14674), .A2(n14215), .ZN(n14801) );
  NAND2_X2 U11708 ( .A1(n14879), .A2(n11278), .ZN(n15374) );
  NAND2_X2 U11709 ( .A1(n14901), .A2(n13832), .ZN(n14879) );
  NAND2_X2 U11710 ( .A1(n12040), .A2(n12039), .ZN(n12773) );
  NAND2_X2 U11711 ( .A1(n17618), .A2(n17620), .ZN(n12648) );
  NAND2_X1 U11712 ( .A1(n13167), .A2(n13154), .ZN(n13301) );
  AND2_X1 U11713 ( .A1(n12506), .A2(n19551), .ZN(n12567) );
  OR2_X1 U11714 ( .A1(n19551), .A2(n12482), .ZN(n12483) );
  XNOR2_X1 U11715 ( .A(n13180), .B(n13179), .ZN(n15359) );
  XNOR2_X1 U11716 ( .A(n13051), .B(n13052), .ZN(n13302) );
  NAND2_X2 U11717 ( .A1(n11781), .A2(n11232), .ZN(n14024) );
  OR2_X1 U11718 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  NOR2_X2 U11719 ( .A1(n14972), .A2(n15113), .ZN(n15112) );
  INV_X2 U11720 ( .A(n15537), .ZN(n13361) );
  AOI21_X2 U11721 ( .B1(n14190), .B2(n16526), .A(n16517), .ZN(n16854) );
  OR2_X2 U11722 ( .A1(n16537), .A2(n11710), .ZN(n16526) );
  NOR2_X2 U11723 ( .A1(n16584), .A2(n16586), .ZN(n16573) );
  AND2_X1 U11725 ( .A1(n17580), .A2(n11231), .ZN(n17477) );
  AND2_X1 U11726 ( .A1(n11402), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11231) );
  INV_X2 U11727 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11232) );
  AND2_X1 U11728 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11233) );
  AND2_X1 U11729 ( .A1(n11995), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11234) );
  NOR2_X1 U11730 ( .A1(n11233), .A2(n11234), .ZN(n11963) );
  NAND2_X1 U11731 ( .A1(n11400), .A2(n12803), .ZN(n17633) );
  NOR2_X1 U11732 ( .A1(n19515), .A2(n12456), .ZN(n12478) );
  CLKBUF_X3 U11733 ( .A(n12489), .Z(n11261) );
  AND2_X1 U11734 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11273) );
  NAND3_X1 U11735 ( .A1(n12067), .A2(n12060), .A3(n12059), .ZN(n11235) );
  AND2_X1 U11736 ( .A1(n11391), .A2(n11390), .ZN(n11236) );
  NAND3_X1 U11737 ( .A1(n12067), .A2(n12060), .A3(n12059), .ZN(n11397) );
  AND2_X2 U11738 ( .A1(n14823), .A2(n14822), .ZN(n12956) );
  NAND2_X1 U11739 ( .A1(n12460), .A2(n12086), .ZN(n11238) );
  NAND2_X1 U11740 ( .A1(n12460), .A2(n12086), .ZN(n12458) );
  NOR2_X4 U11741 ( .A1(n15374), .A2(n15375), .ZN(n15251) );
  NAND2_X1 U11742 ( .A1(n11227), .A2(n11580), .ZN(n11239) );
  BUF_X1 U11743 ( .A(n12788), .Z(n11240) );
  NAND2_X1 U11744 ( .A1(n11401), .A2(n11580), .ZN(n18073) );
  NAND2_X1 U11745 ( .A1(n11573), .A2(n12784), .ZN(n12788) );
  AND2_X1 U11746 ( .A1(n12045), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14653) );
  NOR2_X1 U11747 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11775) );
  BUF_X1 U11748 ( .A(n12062), .Z(n12102) );
  INV_X1 U11749 ( .A(n12519), .ZN(n12586) );
  NOR2_X1 U11750 ( .A1(n12505), .A2(n12495), .ZN(n12519) );
  NAND2_X1 U11751 ( .A1(n11955), .A2(n11954), .ZN(n12032) );
  AND2_X2 U11752 ( .A1(n14176), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12228) );
  NAND2_X1 U11753 ( .A1(n12014), .A2(n12013), .ZN(n12027) );
  AOI21_X2 U11754 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12101), .ZN(n12106) );
  NAND4_X1 U11755 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n11243) );
  NOR2_X2 U11756 ( .A1(n12505), .A2(n17238), .ZN(n12506) );
  INV_X2 U11757 ( .A(n12737), .ZN(n12046) );
  INV_X1 U11758 ( .A(n14170), .ZN(n11246) );
  INV_X1 U11759 ( .A(n14160), .ZN(n11247) );
  INV_X2 U11760 ( .A(n12017), .ZN(n12014) );
  AND2_X1 U11761 ( .A1(n15264), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11248) );
  XNOR2_X1 U11762 ( .A(n11238), .B(n12457), .ZN(n13810) );
  NAND2_X1 U11763 ( .A1(n12458), .A2(n12457), .ZN(n11626) );
  OR2_X1 U11764 ( .A1(n11260), .A2(n12468), .ZN(n12577) );
  INV_X1 U11766 ( .A(n11251), .ZN(n11252) );
  NOR2_X2 U11767 ( .A1(n17267), .A2(n14023), .ZN(n14045) );
  AND2_X2 U11768 ( .A1(n12496), .A2(n14646), .ZN(n12488) );
  OR2_X2 U11769 ( .A1(n11260), .A2(n15700), .ZN(n12505) );
  OR2_X1 U11770 ( .A1(n12455), .A2(n12454), .ZN(n12461) );
  AND2_X2 U11771 ( .A1(n12052), .A2(n12051), .ZN(n11374) );
  NOR2_X2 U11772 ( .A1(n17300), .A2(n17302), .ZN(n17295) );
  INV_X1 U11773 ( .A(n12030), .ZN(n14125) );
  NAND2_X2 U11774 ( .A1(n12455), .A2(n12454), .ZN(n12472) );
  INV_X2 U11775 ( .A(n14170), .ZN(n11985) );
  NOR2_X2 U11776 ( .A1(n11261), .A2(n12480), .ZN(n12573) );
  NAND2_X1 U11777 ( .A1(n11780), .A2(n11232), .ZN(n14170) );
  NAND2_X2 U11778 ( .A1(n12536), .A2(n12535), .ZN(n12563) );
  NOR2_X4 U11779 ( .A1(n17783), .A2(n17544), .ZN(n17543) );
  AOI211_X2 U11780 ( .C1(n18088), .C2(n17790), .A(n17546), .B(n17545), .ZN(
        n17547) );
  NOR2_X4 U11781 ( .A1(n11295), .A2(n15919), .ZN(n15918) );
  OR2_X2 U11782 ( .A1(n15634), .A2(n11670), .ZN(n11295) );
  INV_X1 U11783 ( .A(n19551), .ZN(n12463) );
  INV_X2 U11784 ( .A(n14024), .ZN(n11255) );
  INV_X1 U11785 ( .A(n11255), .ZN(n11256) );
  INV_X1 U11786 ( .A(n14177), .ZN(n11257) );
  INV_X1 U11787 ( .A(n11994), .ZN(n11258) );
  NOR2_X4 U11788 ( .A1(n11773), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15264) );
  BUF_X2 U11789 ( .A(n12489), .Z(n11260) );
  NAND2_X1 U11790 ( .A1(n11803), .A2(n11802), .ZN(n12018) );
  INV_X4 U11791 ( .A(n12218), .ZN(n20322) );
  INV_X2 U11792 ( .A(n12018), .ZN(n12218) );
  CLKBUF_X1 U11793 ( .A(n21342), .Z(n11262) );
  NOR4_X1 U11794 ( .A1(n21869), .A2(n14455), .A3(n11533), .A4(n22090), .ZN(
        n21342) );
  NAND2_X1 U11795 ( .A1(n12075), .A2(n11590), .ZN(n11368) );
  NAND2_X1 U11796 ( .A1(n16524), .A2(n11711), .ZN(n11710) );
  INV_X1 U11797 ( .A(n16538), .ZN(n11711) );
  NAND2_X1 U11798 ( .A1(n16598), .A2(n16600), .ZN(n16584) );
  NOR2_X1 U11799 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13626) );
  NAND2_X1 U11800 ( .A1(n15909), .A2(n11403), .ZN(n15935) );
  AND2_X1 U11801 ( .A1(n11404), .A2(n13449), .ZN(n11403) );
  OR2_X1 U11802 ( .A1(n15908), .A2(n16660), .ZN(n11404) );
  NAND2_X1 U11803 ( .A1(n15033), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13404) );
  NAND2_X1 U11804 ( .A1(n11339), .A2(n16979), .ZN(n11629) );
  INV_X1 U11805 ( .A(n11155), .ZN(n16498) );
  INV_X1 U11806 ( .A(n15855), .ZN(n11565) );
  NAND2_X1 U11807 ( .A1(n11427), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11423) );
  NOR2_X1 U11808 ( .A1(n13068), .A2(n22392), .ZN(n13283) );
  AOI21_X1 U11809 ( .B1(n12816), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12050), 
        .ZN(n12051) );
  AND2_X1 U11810 ( .A1(n12212), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12050) );
  NAND2_X1 U11811 ( .A1(n12159), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11395) );
  AOI21_X1 U11812 ( .B1(n12192), .B2(P2_EBX_REG_1__SCAN_IN), .A(n11338), .ZN(
        n11396) );
  NAND2_X1 U11813 ( .A1(n11397), .A2(n11335), .ZN(n12061) );
  AND2_X1 U11814 ( .A1(n17275), .A2(n14019), .ZN(n14023) );
  AND2_X1 U11815 ( .A1(n12814), .A2(n11625), .ZN(n11624) );
  INV_X1 U11816 ( .A(n17289), .ZN(n11625) );
  NOR2_X1 U11817 ( .A1(n11259), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12239) );
  AND2_X1 U11818 ( .A1(n20322), .A2(n11242), .ZN(n14139) );
  NOR2_X1 U11819 ( .A1(n17889), .A2(n11681), .ZN(n11680) );
  INV_X1 U11820 ( .A(n11682), .ZN(n11681) );
  AND4_X1 U11821 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11920) );
  AOI21_X1 U11822 ( .B1(n12556), .B2(n11379), .A(n11378), .ZN(n11377) );
  INV_X1 U11823 ( .A(n15619), .ZN(n11378) );
  INV_X1 U11824 ( .A(n15547), .ZN(n11379) );
  AND2_X1 U11825 ( .A1(n12054), .A2(n12833), .ZN(n14148) );
  NAND2_X1 U11826 ( .A1(n11991), .A2(n11990), .ZN(n12002) );
  AOI21_X1 U11827 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20140), .A(
        n11859), .ZN(n12005) );
  NOR2_X1 U11828 ( .A1(n11858), .A2(n11857), .ZN(n11859) );
  INV_X1 U11829 ( .A(n11856), .ZN(n11858) );
  AND3_X1 U11830 ( .A1(n11652), .A2(n11310), .A3(n11650), .ZN(n18767) );
  NOR2_X1 U11831 ( .A1(n18695), .A2(n19100), .ZN(n18697) );
  AOI21_X1 U11832 ( .B1(n21622), .B2(n11459), .A(n11458), .ZN(n14526) );
  INV_X1 U11833 ( .A(n22402), .ZN(n14927) );
  AND2_X1 U11834 ( .A1(n22556), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13786) );
  NOR2_X1 U11835 ( .A1(n16108), .A2(n22402), .ZN(n14783) );
  CLKBUF_X1 U11836 ( .A(n12049), .Z(n12019) );
  NOR2_X1 U11837 ( .A1(n15339), .A2(n19580), .ZN(n12021) );
  XNOR2_X1 U11838 ( .A(n11728), .B(n11727), .ZN(n17411) );
  NAND2_X1 U11839 ( .A1(n11726), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11728) );
  INV_X1 U11840 ( .A(n11610), .ZN(n11607) );
  INV_X1 U11841 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20162) );
  AOI21_X1 U11842 ( .B1(n18202), .B2(n18201), .A(n21653), .ZN(n21431) );
  OAI211_X1 U11843 ( .C1(n14490), .C2(n14480), .A(n14479), .B(n14491), .ZN(
        n21654) );
  OAI211_X1 U11844 ( .C1(n14484), .C2(n14483), .A(n14482), .B(n18202), .ZN(
        n17969) );
  NAND2_X1 U11845 ( .A1(n15345), .A2(n19570), .ZN(n19583) );
  NOR2_X1 U11846 ( .A1(n22082), .A2(n11365), .ZN(n22094) );
  INV_X1 U11847 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11553) );
  OAI22_X1 U11848 ( .A1(n15294), .A2(n11861), .B1(n14058), .B2(n12404), .ZN(
        n11547) );
  NAND2_X1 U11849 ( .A1(n20197), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12524) );
  BUF_X1 U11850 ( .A(n13754), .Z(n13709) );
  NOR2_X1 U11851 ( .A1(n13183), .A2(n13175), .ZN(n11408) );
  INV_X1 U11852 ( .A(n12027), .ZN(n12029) );
  NAND2_X1 U11853 ( .A1(n11540), .A2(n11539), .ZN(n12558) );
  NAND2_X1 U11854 ( .A1(n20322), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11539) );
  OR2_X1 U11855 ( .A1(n12718), .A2(n20322), .ZN(n11540) );
  NOR2_X1 U11856 ( .A1(n12017), .A2(n12737), .ZN(n11982) );
  AND2_X1 U11857 ( .A1(n15778), .A2(n11242), .ZN(n11983) );
  NAND2_X1 U11858 ( .A1(n12030), .A2(n12017), .ZN(n12825) );
  AOI22_X1 U11859 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11255), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U11860 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11987) );
  NOR2_X1 U11861 ( .A1(n21479), .A2(n18715), .ZN(n18676) );
  NOR2_X1 U11862 ( .A1(n16558), .A2(n11571), .ZN(n11570) );
  OR2_X1 U11863 ( .A1(n16540), .A2(n11572), .ZN(n11571) );
  INV_X1 U11864 ( .A(n16528), .ZN(n11572) );
  NOR2_X1 U11865 ( .A1(n11563), .A2(n16734), .ZN(n11562) );
  NOR2_X1 U11866 ( .A1(n11710), .A2(n14190), .ZN(n11709) );
  INV_X1 U11867 ( .A(n16721), .ZN(n11703) );
  INV_X1 U11868 ( .A(n13748), .ZN(n13778) );
  NAND2_X1 U11869 ( .A1(n17163), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13748) );
  INV_X1 U11870 ( .A(n16620), .ZN(n13537) );
  INV_X1 U11871 ( .A(n13626), .ZN(n13751) );
  NOR2_X1 U11872 ( .A1(n14777), .A2(n22556), .ZN(n13345) );
  INV_X1 U11873 ( .A(n15689), .ZN(n11566) );
  INV_X1 U11874 ( .A(n13214), .ZN(n11429) );
  NAND2_X1 U11875 ( .A1(n16496), .A2(n11155), .ZN(n14301) );
  AND2_X1 U11876 ( .A1(n13025), .A2(n13024), .ZN(n13052) );
  NAND2_X1 U11877 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11793) );
  INV_X1 U11878 ( .A(n11544), .ZN(n11543) );
  NAND2_X1 U11879 ( .A1(n12683), .A2(n11545), .ZN(n11544) );
  INV_X1 U11880 ( .A(n11348), .ZN(n11545) );
  NAND2_X1 U11881 ( .A1(n15342), .A2(n11590), .ZN(n12049) );
  INV_X1 U11882 ( .A(n11372), .ZN(n11370) );
  AOI22_X1 U11883 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11947) );
  NAND2_X1 U11884 ( .A1(n11995), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11951) );
  AOI211_X1 U11885 ( .C1(n14091), .C2(n14070), .A(n14069), .B(n17245), .ZN(
        n14089) );
  NAND2_X1 U11886 ( .A1(n11667), .A2(n11666), .ZN(n11665) );
  INV_X1 U11887 ( .A(n11714), .ZN(n11664) );
  NAND2_X1 U11888 ( .A1(n11671), .A2(n15888), .ZN(n11670) );
  INV_X1 U11889 ( .A(n11672), .ZN(n11671) );
  INV_X1 U11890 ( .A(n13962), .ZN(n13919) );
  INV_X1 U11891 ( .A(n13956), .ZN(n13915) );
  AND4_X1 U11892 ( .A1(n11588), .A2(n11589), .A3(n11590), .A4(n12046), .ZN(
        n12832) );
  NOR2_X1 U11893 ( .A1(n11245), .A2(n17995), .ZN(n12063) );
  NOR2_X1 U11894 ( .A1(n12874), .A2(n11501), .ZN(n11500) );
  AND2_X1 U11895 ( .A1(n11621), .A2(n15845), .ZN(n11620) );
  AND2_X1 U11896 ( .A1(n15638), .A2(n12140), .ZN(n11621) );
  OR2_X1 U11897 ( .A1(n11521), .A2(n19313), .ZN(n11520) );
  NOR2_X1 U11898 ( .A1(n11615), .A2(n15370), .ZN(n11614) );
  INV_X1 U11899 ( .A(n14960), .ZN(n11615) );
  NOR2_X1 U11900 ( .A1(n17485), .A2(n11331), .ZN(n11496) );
  NAND2_X1 U11901 ( .A1(n11498), .A2(n15972), .ZN(n11497) );
  INV_X1 U11902 ( .A(n12852), .ZN(n11604) );
  NAND2_X1 U11903 ( .A1(n11387), .A2(n11481), .ZN(n15963) );
  NOR2_X1 U11904 ( .A1(n11483), .A2(n11482), .ZN(n11481) );
  OAI21_X1 U11905 ( .B1(n12648), .B2(n11386), .A(n11384), .ZN(n11387) );
  AND2_X1 U11906 ( .A1(n11485), .A2(n11484), .ZN(n11483) );
  INV_X1 U11907 ( .A(n11688), .ZN(n11685) );
  INV_X1 U11908 ( .A(n11689), .ZN(n11687) );
  OR2_X1 U11909 ( .A1(n19394), .A2(n16007), .ZN(n15967) );
  AND2_X1 U11910 ( .A1(n12698), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15968) );
  NAND2_X1 U11911 ( .A1(n11692), .A2(n17527), .ZN(n11688) );
  NAND2_X1 U11912 ( .A1(n11690), .A2(n17527), .ZN(n11689) );
  INV_X1 U11913 ( .A(n15965), .ZN(n11690) );
  AND2_X1 U11914 ( .A1(n12415), .A2(n11603), .ZN(n11602) );
  INV_X1 U11915 ( .A(n15868), .ZN(n11603) );
  AND2_X1 U11916 ( .A1(n12687), .A2(n17536), .ZN(n17550) );
  INV_X1 U11917 ( .A(n17815), .ZN(n12416) );
  NAND2_X1 U11918 ( .A1(n11363), .A2(n11598), .ZN(n11597) );
  INV_X1 U11919 ( .A(n15806), .ZN(n11598) );
  NAND2_X1 U11920 ( .A1(n12541), .A2(n16090), .ZN(n12555) );
  AND2_X1 U11921 ( .A1(n11255), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13961) );
  NAND2_X1 U11922 ( .A1(n12497), .A2(n12496), .ZN(n20138) );
  AOI22_X1 U11923 ( .A1(n11995), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13935), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11840) );
  AND2_X1 U11924 ( .A1(n17995), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13824) );
  NOR2_X1 U11925 ( .A1(n14515), .A2(n14339), .ZN(n14372) );
  NOR2_X1 U11926 ( .A1(n11454), .A2(n14515), .ZN(n14419) );
  NOR2_X1 U11927 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14459), .ZN(
        n18612) );
  AND2_X1 U11928 ( .A1(n19019), .A2(n11302), .ZN(n18769) );
  NAND2_X1 U11929 ( .A1(n18813), .A2(n11361), .ZN(n18874) );
  AOI21_X1 U11930 ( .B1(n18742), .B2(n18741), .A(n21946), .ZN(n18746) );
  OAI21_X1 U11931 ( .B1(n19066), .B2(n11661), .A(n11346), .ZN(n18742) );
  OR2_X1 U11932 ( .A1(n18704), .A2(n11662), .ZN(n11661) );
  INV_X1 U11933 ( .A(n18800), .ZN(n11662) );
  NOR2_X1 U11934 ( .A1(n19068), .A2(n21755), .ZN(n18729) );
  NAND2_X1 U11935 ( .A1(n19090), .A2(n18725), .ZN(n18727) );
  NAND2_X1 U11936 ( .A1(n19115), .A2(n18721), .ZN(n18722) );
  XNOR2_X1 U11937 ( .A(n18719), .B(n21484), .ZN(n18690) );
  INV_X1 U11938 ( .A(n21652), .ZN(n14440) );
  NAND2_X1 U11939 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19653), .ZN(
        n14475) );
  AOI22_X1 U11940 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n19636), .B2(n21624), .ZN(
        n14476) );
  INV_X1 U11941 ( .A(n14367), .ZN(n14491) );
  AOI21_X1 U11942 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17987), .A(
        n14370), .ZN(n14479) );
  NOR2_X1 U11943 ( .A1(n21435), .A2(n19819), .ZN(n14489) );
  NOR2_X1 U11944 ( .A1(n14515), .A2(n14522), .ZN(n18238) );
  NAND2_X1 U11945 ( .A1(n22255), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16691) );
  INV_X1 U11946 ( .A(n15793), .ZN(n16757) );
  NAND2_X1 U11947 ( .A1(n11709), .A2(n16515), .ZN(n11708) );
  AND2_X1 U11948 ( .A1(n13727), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13728) );
  NAND2_X1 U11949 ( .A1(n13728), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13791) );
  INV_X1 U11950 ( .A(n15938), .ZN(n13466) );
  INV_X1 U11951 ( .A(n15538), .ZN(n13351) );
  NAND2_X1 U11952 ( .A1(n13329), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13337) );
  NAND2_X1 U11953 ( .A1(n14913), .A2(n13320), .ZN(n14974) );
  AOI21_X1 U11954 ( .B1(n13300), .B2(n13404), .A(n11696), .ZN(n11695) );
  INV_X1 U11955 ( .A(n13320), .ZN(n11696) );
  AOI21_X1 U11956 ( .B1(n16905), .B2(n17134), .A(n11641), .ZN(n11637) );
  NAND2_X1 U11957 ( .A1(n11644), .A2(n11642), .ZN(n11641) );
  NAND2_X1 U11958 ( .A1(n17134), .A2(n11643), .ZN(n11642) );
  INV_X1 U11959 ( .A(n16856), .ZN(n11644) );
  INV_X1 U11960 ( .A(n13166), .ZN(n11428) );
  NAND2_X1 U11961 ( .A1(n13166), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11426) );
  AND2_X1 U11962 ( .A1(n14792), .A2(n14791), .ZN(n14811) );
  NAND2_X1 U11963 ( .A1(n13049), .A2(n13048), .ZN(n13144) );
  INV_X1 U11964 ( .A(n14758), .ZN(n17163) );
  NOR2_X1 U11965 ( .A1(n13301), .A2(n13100), .ZN(n15149) );
  NAND2_X1 U11966 ( .A1(n13291), .A2(n13290), .ZN(n16108) );
  OAI21_X1 U11967 ( .B1(n14197), .B2(n13287), .A(n13286), .ZN(n13291) );
  INV_X1 U11968 ( .A(n11510), .ZN(n11509) );
  OAI21_X1 U11969 ( .B1(n11252), .B2(n11511), .A(n19484), .ZN(n11510) );
  NAND2_X1 U11970 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19386), .ZN(n19462) );
  NAND2_X1 U11971 ( .A1(n11669), .A2(n17280), .ZN(n11668) );
  INV_X1 U11972 ( .A(n17288), .ZN(n11669) );
  BUF_X1 U11973 ( .A(n14021), .Z(n17275) );
  AND2_X1 U11974 ( .A1(n20546), .A2(n14128), .ZN(n15614) );
  NAND2_X1 U11975 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11512) );
  INV_X1 U11976 ( .A(n15881), .ZN(n12153) );
  NAND2_X1 U11977 ( .A1(n17602), .A2(n12661), .ZN(n11484) );
  NOR2_X1 U11978 ( .A1(n17602), .A2(n12661), .ZN(n11485) );
  NAND2_X1 U11979 ( .A1(n11610), .A2(n11609), .ZN(n11608) );
  NOR2_X1 U11980 ( .A1(n17177), .A2(n16038), .ZN(n11609) );
  NAND2_X1 U11981 ( .A1(n15991), .A2(n11308), .ZN(n11389) );
  INV_X1 U11982 ( .A(n16049), .ZN(n11478) );
  AND2_X1 U11983 ( .A1(n11328), .A2(n17271), .ZN(n11622) );
  AOI21_X1 U11984 ( .B1(n11496), .B2(n11497), .A(n11327), .ZN(n11494) );
  INV_X1 U11985 ( .A(n11497), .ZN(n11493) );
  OAI21_X1 U11986 ( .B1(n17551), .B2(n11689), .A(n11688), .ZN(n17512) );
  NOR2_X1 U11987 ( .A1(n17922), .A2(n11322), .ZN(n17874) );
  NAND2_X1 U11988 ( .A1(n12648), .A2(n11680), .ZN(n11383) );
  INV_X1 U11989 ( .A(n12800), .ZN(n12796) );
  NAND2_X1 U11990 ( .A1(n15627), .A2(n15834), .ZN(n15629) );
  AND3_X1 U11991 ( .A1(n12268), .A2(n12267), .A3(n12266), .ZN(n15556) );
  AND2_X1 U11992 ( .A1(n20132), .A2(n20447), .ZN(n20249) );
  INV_X1 U11993 ( .A(n15767), .ZN(n15766) );
  NOR2_X1 U11994 ( .A1(n20108), .A2(n20554), .ZN(n20218) );
  CLKBUF_X1 U11995 ( .A(n13800), .Z(n13801) );
  OR2_X1 U11996 ( .A1(n20132), .A2(n20447), .ZN(n20109) );
  OR2_X1 U11997 ( .A1(n12762), .A2(n12011), .ZN(n15339) );
  INV_X1 U11998 ( .A(n21647), .ZN(n14494) );
  NOR2_X1 U11999 ( .A1(n11454), .A2(n11453), .ZN(n14404) );
  NAND2_X1 U12000 ( .A1(n21638), .A2(n14501), .ZN(n11453) );
  AOI22_X1 U12001 ( .A1(n21432), .A2(n21431), .B1(n21430), .B2(n21429), .ZN(
        n21605) );
  NOR3_X1 U12002 ( .A1(n22418), .A2(n21647), .A3(n21653), .ZN(n21430) );
  OR2_X1 U12003 ( .A1(n18901), .A2(n21874), .ZN(n11649) );
  AND2_X1 U12004 ( .A1(n18816), .A2(n11288), .ZN(n18890) );
  INV_X1 U12005 ( .A(n21661), .ZN(n21935) );
  NOR2_X1 U12006 ( .A1(n19070), .A2(n19069), .ZN(n19068) );
  OR2_X1 U12007 ( .A1(n19081), .A2(n21730), .ZN(n11653) );
  NAND2_X1 U12008 ( .A1(n18699), .A2(n11651), .ZN(n11650) );
  INV_X1 U12009 ( .A(n19081), .ZN(n11651) );
  OR2_X1 U12010 ( .A1(n19087), .A2(n21730), .ZN(n11655) );
  NOR2_X1 U12011 ( .A1(n19739), .A2(n14440), .ZN(n21648) );
  INV_X1 U12012 ( .A(n21894), .ZN(n22016) );
  OAI21_X1 U12013 ( .B1(n14528), .B2(n14529), .A(n11470), .ZN(n11469) );
  AOI21_X1 U12014 ( .B1(n14531), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11470) );
  AOI21_X1 U12015 ( .B1(n14528), .B2(n14529), .A(n19609), .ZN(n11467) );
  OAI21_X1 U12016 ( .B1(n14530), .B2(n14531), .A(n11334), .ZN(n11464) );
  OR2_X1 U12017 ( .A1(n17970), .A2(n14532), .ZN(n11465) );
  NOR2_X1 U12018 ( .A1(n14314), .A2(n22388), .ZN(n14205) );
  NAND2_X1 U12019 ( .A1(n11558), .A2(n11557), .ZN(n16967) );
  NAND2_X1 U12020 ( .A1(n16501), .A2(n16500), .ZN(n11557) );
  NAND2_X1 U12021 ( .A1(n16502), .A2(n11559), .ZN(n11558) );
  OR2_X1 U12022 ( .A1(n16536), .A2(n16524), .ZN(n16525) );
  NAND2_X1 U12023 ( .A1(n22385), .A2(n13790), .ZN(n20842) );
  AND2_X1 U12024 ( .A1(n20842), .A2(n14858), .ZN(n20862) );
  NAND2_X2 U12025 ( .A1(n14783), .A2(n18031), .ZN(n22385) );
  INV_X1 U12026 ( .A(n16967), .ZN(n11556) );
  AND2_X1 U12027 ( .A1(n11340), .A2(n11285), .ZN(n11436) );
  OR2_X1 U12028 ( .A1(n15196), .A2(n14937), .ZN(n15050) );
  NAND2_X1 U12029 ( .A1(n14547), .A2(n17240), .ZN(n19275) );
  NAND2_X1 U12030 ( .A1(n19483), .A2(n11252), .ZN(n19499) );
  NOR2_X1 U12031 ( .A1(n11508), .A2(n17439), .ZN(n11504) );
  NAND2_X1 U12032 ( .A1(n11509), .A2(n11511), .ZN(n11508) );
  AND2_X1 U12033 ( .A1(n11253), .A2(n11515), .ZN(n19353) );
  NAND2_X1 U12034 ( .A1(n19336), .A2(n17566), .ZN(n11515) );
  INV_X1 U12035 ( .A(n19464), .ZN(n19491) );
  OR2_X1 U12036 ( .A1(n17651), .A2(n15680), .ZN(n14187) );
  AND2_X1 U12037 ( .A1(n17309), .A2(n11242), .ZN(n17303) );
  AND2_X1 U12038 ( .A1(n14149), .A2(n19570), .ZN(n17309) );
  AND2_X1 U12039 ( .A1(n20546), .A2(n14125), .ZN(n20551) );
  NAND2_X1 U12040 ( .A1(n19583), .A2(n12871), .ZN(n18093) );
  AND2_X1 U12041 ( .A1(n18093), .A2(n14544), .ZN(n18083) );
  INV_X1 U12042 ( .A(n18083), .ZN(n17638) );
  INV_X1 U12043 ( .A(n18088), .ZN(n17641) );
  INV_X1 U12044 ( .A(n18063), .ZN(n18086) );
  XNOR2_X1 U12045 ( .A(n16039), .B(n16038), .ZN(n17652) );
  AND2_X1 U12046 ( .A1(n11617), .A2(n11616), .ZN(n14152) );
  AND2_X1 U12047 ( .A1(n16063), .A2(n16064), .ZN(n14127) );
  NAND2_X1 U12048 ( .A1(n12860), .A2(n12859), .ZN(n19542) );
  NAND2_X1 U12049 ( .A1(n12860), .A2(n12819), .ZN(n19514) );
  AND2_X1 U12050 ( .A1(n12860), .A2(n15326), .ZN(n19537) );
  INV_X1 U12051 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20247) );
  INV_X1 U12052 ( .A(n20554), .ZN(n18098) );
  INV_X1 U12053 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20245) );
  NAND2_X1 U12054 ( .A1(n11531), .A2(n11530), .ZN(n11529) );
  OR2_X1 U12055 ( .A1(n21401), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n11530) );
  NAND2_X1 U12056 ( .A1(n11532), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n11531) );
  OR2_X1 U12057 ( .A1(n21406), .A2(n21424), .ZN(n11532) );
  NOR2_X2 U12058 ( .A1(n11262), .A2(n22084), .ZN(n21404) );
  INV_X1 U12059 ( .A(n18958), .ZN(n11451) );
  NAND2_X1 U12060 ( .A1(n18964), .A2(n18959), .ZN(n11450) );
  AOI21_X1 U12061 ( .B1(n21886), .B2(n19072), .A(n18974), .ZN(n18978) );
  INV_X1 U12062 ( .A(n19054), .ZN(n18961) );
  INV_X1 U12063 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19609) );
  NAND2_X1 U12064 ( .A1(n11463), .A2(n11462), .ZN(n11461) );
  AOI211_X1 U12065 ( .C1(n22097), .C2(n17969), .A(n19613), .B(n17968), .ZN(
        n21639) );
  NOR2_X1 U12066 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n22095), .ZN(n14535) );
  NOR3_X1 U12067 ( .A1(n22091), .A2(n21653), .A3(n11362), .ZN(n22082) );
  NAND2_X1 U12068 ( .A1(n15033), .A2(n14771), .ZN(n12929) );
  AND2_X1 U12069 ( .A1(n13247), .A2(n13246), .ZN(n13249) );
  AOI21_X1 U12070 ( .B1(n20171), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n19264), .ZN(n12516) );
  AND2_X1 U12071 ( .A1(n14163), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11974) );
  OR2_X1 U12072 ( .A1(n14365), .A2(n14366), .ZN(n14361) );
  NOR2_X1 U12073 ( .A1(n11160), .A2(n13226), .ZN(n16943) );
  OR2_X1 U12074 ( .A1(n13022), .A2(n13021), .ZN(n13216) );
  OR2_X1 U12075 ( .A1(n13011), .A2(n13010), .ZN(n13158) );
  NAND2_X1 U12076 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11630) );
  NAND2_X1 U12077 ( .A1(n13028), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11632) );
  NAND2_X1 U12078 ( .A1(n13376), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U12079 ( .A1(n13127), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11633) );
  NAND2_X1 U12080 ( .A1(n12900), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11634) );
  AOI21_X1 U12081 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n22553), .A(
        n13249), .ZN(n13244) );
  AND2_X1 U12082 ( .A1(n20247), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12009) );
  INV_X1 U12083 ( .A(n17276), .ZN(n11666) );
  INV_X1 U12084 ( .A(n11668), .ZN(n11667) );
  INV_X1 U12085 ( .A(n17474), .ZN(n11489) );
  AND2_X1 U12086 ( .A1(n11385), .A2(n11484), .ZN(n11384) );
  OR2_X1 U12087 ( .A1(n11680), .A2(n11386), .ZN(n11385) );
  INV_X1 U12088 ( .A(n12658), .ZN(n11386) );
  INV_X1 U12089 ( .A(n17594), .ZN(n11482) );
  NOR2_X1 U12090 ( .A1(n11862), .A2(n11547), .ZN(n11874) );
  NOR2_X1 U12091 ( .A1(n12031), .A2(n15778), .ZN(n12056) );
  NAND2_X1 U12092 ( .A1(n11588), .A2(n12053), .ZN(n12036) );
  AND3_X1 U12093 ( .A1(n11989), .A2(n15297), .A3(n11988), .ZN(n11990) );
  AOI22_X1 U12094 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U12095 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U12096 ( .A1(n11832), .A2(n11831), .ZN(n11856) );
  XNOR2_X1 U12097 ( .A(n15297), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U12098 ( .A1(n12040), .A2(n12003), .ZN(n12042) );
  INV_X1 U12099 ( .A(n12031), .ZN(n12003) );
  NAND2_X1 U12100 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14501), .ZN(
        n14337) );
  NOR2_X1 U12101 ( .A1(n18718), .A2(n18706), .ZN(n18714) );
  AOI21_X1 U12102 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19636), .A(
        n14360), .ZN(n14366) );
  NOR2_X1 U12103 ( .A1(n14475), .A2(n14476), .ZN(n14360) );
  AND2_X1 U12104 ( .A1(n11705), .A2(n16612), .ZN(n11704) );
  NOR2_X1 U12105 ( .A1(n16726), .A2(n16624), .ZN(n11705) );
  NOR2_X1 U12106 ( .A1(n13517), .A2(n16639), .ZN(n13552) );
  AND2_X1 U12107 ( .A1(n17089), .A2(n11318), .ZN(n11635) );
  NAND2_X1 U12108 ( .A1(n11699), .A2(n11697), .ZN(n16620) );
  NOR2_X1 U12109 ( .A1(n11701), .A2(n11698), .ZN(n11697) );
  INV_X1 U12110 ( .A(n16635), .ZN(n11698) );
  NAND2_X1 U12111 ( .A1(n11702), .A2(n13485), .ZN(n11701) );
  INV_X1 U12112 ( .A(n16646), .ZN(n11702) );
  OR2_X1 U12113 ( .A1(n16960), .A2(n16958), .ZN(n16944) );
  NAND2_X1 U12114 ( .A1(n13400), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13406) );
  INV_X1 U12115 ( .A(n16858), .ZN(n11643) );
  NAND2_X1 U12116 ( .A1(n14271), .A2(n11562), .ZN(n11561) );
  INV_X1 U12117 ( .A(n13195), .ZN(n11417) );
  INV_X1 U12118 ( .A(n16495), .ZN(n16499) );
  AND2_X1 U12119 ( .A1(n14702), .A2(n14701), .ZN(n14788) );
  OR2_X1 U12120 ( .A1(n13040), .A2(n13039), .ZN(n13157) );
  NOR2_X1 U12121 ( .A1(n14771), .A2(n22392), .ZN(n13050) );
  OR2_X1 U12122 ( .A1(n13079), .A2(n13078), .ZN(n13159) );
  OR2_X1 U12123 ( .A1(n22237), .A2(n22224), .ZN(n22566) );
  NAND2_X1 U12124 ( .A1(n14817), .A2(n22392), .ZN(n13099) );
  INV_X1 U12125 ( .A(n13311), .ZN(n15044) );
  AND2_X1 U12126 ( .A1(n22840), .A2(n13082), .ZN(n15437) );
  AOI21_X1 U12127 ( .B1(n18051), .B2(n22391), .A(n22396), .ZN(n14985) );
  INV_X1 U12128 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22552) );
  AND2_X1 U12129 ( .A1(n13068), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13288) );
  AOI21_X1 U12130 ( .B1(n11996), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n15297), .ZN(n11792) );
  NAND2_X1 U12131 ( .A1(n14163), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11796) );
  AND2_X1 U12132 ( .A1(n11930), .A2(n15996), .ZN(n16006) );
  NAND2_X1 U12133 ( .A1(n11875), .A2(n11538), .ZN(n12602) );
  INV_X1 U12134 ( .A(n12558), .ZN(n11538) );
  INV_X1 U12135 ( .A(n13949), .ZN(n12401) );
  INV_X1 U12136 ( .A(n13948), .ZN(n12399) );
  NOR2_X1 U12137 ( .A1(n17957), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13925) );
  NAND2_X1 U12138 ( .A1(n17244), .A2(n17252), .ZN(n14093) );
  AND2_X1 U12139 ( .A1(n14114), .A2(n14113), .ZN(n14115) );
  NAND2_X1 U12140 ( .A1(n11674), .A2(n11673), .ZN(n11672) );
  INV_X1 U12141 ( .A(n15867), .ZN(n11673) );
  INV_X1 U12142 ( .A(n11675), .ZN(n11674) );
  AND2_X1 U12143 ( .A1(n11259), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13802) );
  NAND2_X1 U12144 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11513) );
  NAND2_X1 U12145 ( .A1(n11519), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11518) );
  INV_X1 U12146 ( .A(n11520), .ZN(n11519) );
  INV_X1 U12147 ( .A(n15679), .ZN(n12140) );
  NAND2_X1 U12148 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11521) );
  NOR2_X1 U12149 ( .A1(n11611), .A2(n11612), .ZN(n11610) );
  INV_X1 U12150 ( .A(n14126), .ZN(n11611) );
  NAND2_X1 U12151 ( .A1(n16050), .A2(n15995), .ZN(n15998) );
  INV_X1 U12152 ( .A(n16025), .ZN(n12195) );
  INV_X1 U12153 ( .A(n17281), .ZN(n11623) );
  AND2_X1 U12154 ( .A1(n12843), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11592) );
  AND2_X1 U12155 ( .A1(n12424), .A2(n11606), .ZN(n11605) );
  INV_X1 U12156 ( .A(n17389), .ZN(n11606) );
  INV_X1 U12157 ( .A(n17400), .ZN(n12425) );
  AND2_X1 U12158 ( .A1(n12651), .A2(n17619), .ZN(n11682) );
  AOI21_X1 U12159 ( .B1(n12794), .B2(n15837), .A(n11584), .ZN(n12802) );
  NOR2_X1 U12160 ( .A1(n12800), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11419) );
  NAND2_X1 U12161 ( .A1(n11381), .A2(n15722), .ZN(n12637) );
  NAND2_X1 U12162 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  NAND2_X1 U12163 ( .A1(n15598), .A2(n11599), .ZN(n15610) );
  AND2_X1 U12164 ( .A1(n12261), .A2(n11319), .ZN(n11599) );
  OAI22_X1 U12165 ( .A1(n12062), .A2(n12066), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12192), .ZN(n12071) );
  OAI211_X1 U12166 ( .C1(n12390), .C2(n12544), .A(n12238), .B(n12253), .ZN(
        n15601) );
  INV_X1 U12167 ( .A(n15556), .ZN(n11600) );
  INV_X1 U12168 ( .A(n12500), .ZN(n12459) );
  AOI22_X1 U12169 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U12170 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U12171 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11936) );
  NAND2_X1 U12172 ( .A1(n12501), .A2(n19551), .ZN(n12621) );
  AND2_X1 U12173 ( .A1(n12755), .A2(n12754), .ZN(n15280) );
  AOI221_X1 U12174 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12005), 
        .C1(n19509), .C2(n12005), .A(n12004), .ZN(n12762) );
  INV_X1 U12175 ( .A(n18631), .ZN(n18433) );
  NOR2_X1 U12176 ( .A1(n14523), .A2(n14337), .ZN(n18634) );
  NOR2_X1 U12177 ( .A1(n11454), .A2(n14337), .ZN(n18633) );
  NOR2_X1 U12178 ( .A1(n14337), .A2(n14339), .ZN(n18632) );
  NOR2_X1 U12179 ( .A1(n14523), .A2(n14340), .ZN(n18631) );
  NAND2_X1 U12180 ( .A1(n21624), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11454) );
  NAND2_X1 U12181 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11445) );
  AOI21_X1 U12182 ( .B1(n18630), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n11447), .ZN(n11446) );
  NOR2_X1 U12183 ( .A1(n18433), .A2(n11448), .ZN(n11447) );
  INV_X1 U12184 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11448) );
  NOR2_X1 U12185 ( .A1(n14456), .A2(n11524), .ZN(n11523) );
  NOR2_X1 U12186 ( .A1(n21229), .A2(n11537), .ZN(n11536) );
  NAND2_X1 U12187 ( .A1(n18868), .A2(n21658), .ZN(n18753) );
  NAND2_X1 U12188 ( .A1(n14449), .A2(n11307), .ZN(n14497) );
  AND2_X1 U12189 ( .A1(n18700), .A2(n18708), .ZN(n18702) );
  NAND2_X1 U12190 ( .A1(n14509), .A2(n14507), .ZN(n14498) );
  NAND2_X1 U12191 ( .A1(n11443), .A2(n11442), .ZN(n18716) );
  OR2_X1 U12192 ( .A1(n18717), .A2(n18715), .ZN(n11442) );
  INV_X1 U12193 ( .A(n18714), .ZN(n11443) );
  NAND2_X1 U12194 ( .A1(n11657), .A2(n11656), .ZN(n18691) );
  NOR2_X1 U12195 ( .A1(n14516), .A2(n14497), .ZN(n14506) );
  OAI21_X1 U12196 ( .B1(n22088), .B2(n18578), .A(n17965), .ZN(n19612) );
  NAND2_X1 U12197 ( .A1(n20969), .A2(n14495), .ZN(n21429) );
  INV_X1 U12198 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16639) );
  AND2_X1 U12199 ( .A1(n13477), .A2(n13420), .ZN(n16660) );
  INV_X1 U12200 ( .A(n16500), .ZN(n11559) );
  OR2_X1 U12201 ( .A1(n16561), .A2(n11569), .ZN(n16497) );
  NAND2_X1 U12202 ( .A1(n14302), .A2(n11570), .ZN(n11569) );
  INV_X1 U12203 ( .A(n11570), .ZN(n11568) );
  AND2_X1 U12204 ( .A1(n14264), .A2(n14263), .ZN(n16647) );
  NOR2_X1 U12205 ( .A1(n16735), .A2(n11560), .ZN(n16649) );
  INV_X1 U12206 ( .A(n11562), .ZN(n11560) );
  AND2_X1 U12207 ( .A1(n14260), .A2(n14259), .ZN(n16734) );
  NOR2_X1 U12208 ( .A1(n16735), .A2(n16734), .ZN(n16736) );
  AND2_X1 U12209 ( .A1(n14295), .A2(n14293), .ZN(n16495) );
  NAND2_X1 U12210 ( .A1(n16834), .A2(n12978), .ZN(n16744) );
  AND2_X1 U12211 ( .A1(n14749), .A2(n18044), .ZN(n20709) );
  INV_X1 U12212 ( .A(n11709), .ZN(n11707) );
  AOI21_X1 U12213 ( .B1(n13782), .B2(n16863), .A(n13725), .ZN(n16524) );
  AND2_X1 U12214 ( .A1(n13688), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13689) );
  NAND2_X1 U12215 ( .A1(n13648), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13687) );
  AND2_X1 U12216 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n13602), .ZN(
        n13603) );
  INV_X1 U12217 ( .A(n13601), .ZN(n13602) );
  NAND2_X1 U12218 ( .A1(n13603), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13647) );
  CLKBUF_X1 U12219 ( .A(n16584), .Z(n16585) );
  CLKBUF_X1 U12220 ( .A(n16598), .Z(n16599) );
  AND2_X1 U12221 ( .A1(n13552), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13553) );
  NAND2_X1 U12222 ( .A1(n13553), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13569) );
  CLKBUF_X1 U12223 ( .A(n16620), .Z(n16621) );
  NAND2_X1 U12224 ( .A1(n13504), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13517) );
  OR2_X1 U12225 ( .A1(n13468), .A2(n13451), .ZN(n13486) );
  INV_X1 U12226 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13421) );
  CLKBUF_X1 U12227 ( .A(n15935), .Z(n15936) );
  NOR2_X1 U12228 ( .A1(n13406), .A2(n13401), .ZN(n13407) );
  AND2_X1 U12229 ( .A1(n13375), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13400) );
  AND3_X1 U12230 ( .A1(n13374), .A2(n13373), .A3(n13372), .ZN(n15756) );
  NOR2_X1 U12231 ( .A1(n13353), .A2(n22291), .ZN(n13375) );
  NAND2_X1 U12232 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13353) );
  NOR2_X1 U12233 ( .A1(n13337), .A2(n22270), .ZN(n13346) );
  AOI21_X1 U12234 ( .B1(n13336), .B2(n13477), .A(n13335), .ZN(n15113) );
  INV_X1 U12235 ( .A(n13334), .ZN(n13335) );
  NOR2_X1 U12236 ( .A1(n13322), .A2(n15381), .ZN(n13329) );
  INV_X1 U12237 ( .A(n14910), .ZN(n13319) );
  AND2_X1 U12238 ( .A1(n11629), .A2(n11285), .ZN(n11435) );
  NAND2_X1 U12239 ( .A1(n11629), .A2(n11332), .ZN(n11434) );
  AND2_X1 U12240 ( .A1(n14291), .A2(n14290), .ZN(n16540) );
  NOR2_X1 U12241 ( .A1(n16557), .A2(n16540), .ZN(n16539) );
  NOR2_X1 U12242 ( .A1(n16593), .A2(n16581), .ZN(n16580) );
  AND2_X1 U12243 ( .A1(n16983), .A2(n16982), .ZN(n17053) );
  OR2_X1 U12244 ( .A1(n16718), .A2(n16601), .ZN(n16603) );
  OR2_X1 U12245 ( .A1(n16603), .A2(n16595), .ZN(n16593) );
  NOR2_X1 U12246 ( .A1(n11292), .A2(n16614), .ZN(n16720) );
  AND3_X1 U12247 ( .A1(n14274), .A2(n14273), .A3(n14272), .ZN(n16724) );
  OR2_X1 U12248 ( .A1(n16666), .A2(n15944), .ZN(n16735) );
  AND2_X1 U12249 ( .A1(n13229), .A2(n16970), .ZN(n16958) );
  AND2_X1 U12250 ( .A1(n15650), .A2(n11564), .ZN(n17119) );
  AND2_X1 U12251 ( .A1(n11282), .A2(n11341), .ZN(n11564) );
  NAND2_X1 U12252 ( .A1(n11414), .A2(n17134), .ZN(n11413) );
  NAND2_X1 U12253 ( .A1(n15650), .A2(n11282), .ZN(n17115) );
  AND2_X1 U12254 ( .A1(n14240), .A2(n14239), .ZN(n15689) );
  NAND2_X1 U12255 ( .A1(n15650), .A2(n11323), .ZN(n15856) );
  AOI21_X1 U12256 ( .B1(n15643), .B2(n11429), .A(n11300), .ZN(n11410) );
  AND2_X1 U12257 ( .A1(n15595), .A2(n15594), .ZN(n15650) );
  NAND2_X1 U12258 ( .A1(n15650), .A2(n14236), .ZN(n15690) );
  INV_X1 U12259 ( .A(n22147), .ZN(n17122) );
  OR2_X1 U12260 ( .A1(n15115), .A2(n15114), .ZN(n15542) );
  NAND2_X1 U12261 ( .A1(n11627), .A2(n13166), .ZN(n13173) );
  AND2_X1 U12262 ( .A1(n14893), .A2(n14892), .ZN(n14976) );
  OR2_X1 U12263 ( .A1(n14811), .A2(n16105), .ZN(n22119) );
  NOR2_X1 U12264 ( .A1(n14811), .A2(n14804), .ZN(n22123) );
  INV_X1 U12265 ( .A(n22119), .ZN(n17125) );
  INV_X1 U12266 ( .A(n14682), .ZN(n12979) );
  NAND2_X1 U12267 ( .A1(n13060), .A2(n13059), .ZN(n13067) );
  NAND2_X1 U12268 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  XNOR2_X1 U12269 ( .A(n17974), .B(n15059), .ZN(n14817) );
  INV_X1 U12270 ( .A(n18037), .ZN(n18017) );
  NAND2_X1 U12271 ( .A1(n11254), .A2(n13311), .ZN(n22548) );
  NOR2_X1 U12272 ( .A1(n13301), .A2(n14935), .ZN(n15120) );
  INV_X1 U12273 ( .A(n15050), .ZN(n15045) );
  NAND2_X1 U12274 ( .A1(n11254), .A2(n15044), .ZN(n15392) );
  INV_X1 U12275 ( .A(n15198), .ZN(n15148) );
  INV_X1 U12276 ( .A(n15197), .ZN(n15147) );
  NAND2_X1 U12277 ( .A1(n16757), .A2(n20873), .ZN(n15184) );
  OR2_X1 U12278 ( .A1(n16757), .A2(n20853), .ZN(n15186) );
  AND2_X1 U12279 ( .A1(n22388), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U12280 ( .A1(n11903), .A2(n12634), .ZN(n16013) );
  INV_X1 U12281 ( .A(n19500), .ZN(n11511) );
  NOR2_X1 U12282 ( .A1(n15988), .A2(n11552), .ZN(n11551) );
  INV_X1 U12283 ( .A(n15982), .ZN(n11552) );
  NAND2_X1 U12284 ( .A1(n12702), .A2(n12703), .ZN(n12711) );
  INV_X1 U12285 ( .A(n12688), .ZN(n11546) );
  INV_X1 U12286 ( .A(n12667), .ZN(n11542) );
  NAND2_X1 U12287 ( .A1(n11903), .A2(n11548), .ZN(n12650) );
  NAND2_X1 U12288 ( .A1(n15656), .A2(n12273), .ZN(n15718) );
  NAND2_X1 U12289 ( .A1(n15798), .A2(n11676), .ZN(n11675) );
  INV_X1 U12290 ( .A(n15849), .ZN(n11676) );
  INV_X1 U12291 ( .A(n15683), .ZN(n11677) );
  AND2_X1 U12292 ( .A1(n15254), .A2(n11679), .ZN(n11678) );
  INV_X1 U12293 ( .A(n15590), .ZN(n11679) );
  INV_X1 U12294 ( .A(n11374), .ZN(n11373) );
  INV_X1 U12295 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11774) );
  AND2_X1 U12296 ( .A1(n12429), .A2(n12428), .ZN(n12852) );
  OR3_X1 U12297 ( .A1(n13907), .A2(n13906), .A3(n13905), .ZN(n17296) );
  CLKBUF_X1 U12298 ( .A(n17286), .Z(n17287) );
  CLKBUF_X1 U12299 ( .A(n17300), .Z(n17301) );
  CLKBUF_X1 U12300 ( .A(n11295), .Z(n15887) );
  AND2_X1 U12301 ( .A1(n12418), .A2(n12417), .ZN(n15868) );
  AND3_X1 U12302 ( .A1(n12375), .A2(n12374), .A3(n12373), .ZN(n15806) );
  AND2_X1 U12303 ( .A1(n13831), .A2(n11720), .ZN(n13832) );
  AND2_X1 U12304 ( .A1(n14652), .A2(n19266), .ZN(n18127) );
  INV_X1 U12305 ( .A(n14138), .ZN(n15777) );
  OAI21_X1 U12306 ( .B1(n14137), .B2(n14136), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14138) );
  INV_X1 U12307 ( .A(n11617), .ZN(n17184) );
  AND2_X1 U12308 ( .A1(n11271), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U12309 ( .A1(n17305), .A2(n12814), .ZN(n17290) );
  NAND2_X1 U12310 ( .A1(n17305), .A2(n11624), .ZN(n17292) );
  INV_X1 U12311 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12874) );
  INV_X1 U12312 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19375) );
  AND2_X1 U12313 ( .A1(n11620), .A2(n11619), .ZN(n11618) );
  INV_X1 U12314 ( .A(n15801), .ZN(n11619) );
  AND2_X1 U12315 ( .A1(n15387), .A2(n11621), .ZN(n15846) );
  AND2_X1 U12316 ( .A1(n15387), .A2(n12140), .ZN(n15677) );
  NOR2_X1 U12317 ( .A1(n11757), .A2(n18094), .ZN(n11759) );
  INV_X1 U12318 ( .A(n15256), .ZN(n11613) );
  NAND2_X1 U12319 ( .A1(n14967), .A2(n11614), .ZN(n15373) );
  INV_X1 U12320 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U12321 ( .A1(n17433), .A2(n17431), .ZN(n17419) );
  INV_X1 U12322 ( .A(n16058), .ZN(n11616) );
  AND2_X1 U12323 ( .A1(n12440), .A2(n12439), .ZN(n17177) );
  NOR2_X1 U12324 ( .A1(n11265), .A2(n17351), .ZN(n17341) );
  AND2_X1 U12325 ( .A1(n17305), .A2(n11328), .ZN(n17282) );
  AND2_X1 U12326 ( .A1(n11591), .A2(n12810), .ZN(n11402) );
  AND2_X1 U12327 ( .A1(n11592), .A2(n16031), .ZN(n11591) );
  AND2_X1 U12328 ( .A1(n12425), .A2(n11347), .ZN(n17372) );
  OR2_X1 U12329 ( .A1(n15969), .A2(n15968), .ZN(n15971) );
  NAND2_X1 U12330 ( .A1(n17572), .A2(n11592), .ZN(n17500) );
  NAND2_X1 U12331 ( .A1(n17511), .A2(n11687), .ZN(n11686) );
  AOI21_X1 U12332 ( .B1(n11685), .B2(n17511), .A(n15959), .ZN(n11684) );
  NAND2_X1 U12333 ( .A1(n12425), .A2(n11605), .ZN(n17391) );
  NAND2_X1 U12334 ( .A1(n12425), .A2(n12424), .ZN(n17402) );
  NAND2_X1 U12335 ( .A1(n12416), .A2(n11601), .ZN(n17400) );
  AND2_X1 U12336 ( .A1(n11329), .A2(n15920), .ZN(n11601) );
  AND2_X1 U12337 ( .A1(n12416), .A2(n11329), .ZN(n15921) );
  NAND2_X1 U12338 ( .A1(n12416), .A2(n12415), .ZN(n17816) );
  NOR2_X1 U12339 ( .A1(n11597), .A2(n11596), .ZN(n11595) );
  INV_X1 U12340 ( .A(n17841), .ZN(n11596) );
  INV_X1 U12341 ( .A(n17567), .ZN(n17795) );
  NAND2_X1 U12342 ( .A1(n12648), .A2(n11682), .ZN(n17887) );
  AND2_X1 U12343 ( .A1(n12655), .A2(n17894), .ZN(n17889) );
  AND3_X1 U12344 ( .A1(n12327), .A2(n12326), .A3(n12325), .ZN(n15732) );
  NAND2_X1 U12345 ( .A1(n11578), .A2(n17632), .ZN(n11577) );
  INV_X1 U12346 ( .A(n17631), .ZN(n11578) );
  INV_X1 U12347 ( .A(n17632), .ZN(n11579) );
  NAND2_X1 U12348 ( .A1(n14967), .A2(n14960), .ZN(n15371) );
  INV_X1 U12349 ( .A(n15610), .ZN(n15658) );
  OAI21_X1 U12350 ( .B1(n15546), .B2(n11380), .A(n11377), .ZN(n12562) );
  NAND4_X1 U12351 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n14542) );
  BUF_X1 U12352 ( .A(n12067), .Z(n15261) );
  AND2_X1 U12353 ( .A1(n12860), .A2(n12839), .ZN(n17919) );
  NOR2_X1 U12354 ( .A1(n12823), .A2(n15333), .ZN(n19539) );
  MUX2_X1 U12355 ( .A(n12249), .B(n20245), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n14840) );
  NAND2_X1 U12356 ( .A1(n14839), .A2(n14840), .ZN(n14838) );
  NOR2_X2 U12357 ( .A1(n11782), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15300) );
  AOI21_X1 U12358 ( .B1(n17238), .B2(n13824), .A(n13823), .ZN(n14714) );
  CLKBUF_X1 U12359 ( .A(n12816), .Z(n12817) );
  INV_X1 U12360 ( .A(n12577), .ZN(n20171) );
  AND2_X1 U12361 ( .A1(n20108), .A2(n18098), .ZN(n20191) );
  INV_X1 U12362 ( .A(n20100), .ZN(n20096) );
  NAND2_X2 U12363 ( .A1(n11855), .A2(n11854), .ZN(n12045) );
  NAND2_X1 U12364 ( .A1(n11847), .A2(n15297), .ZN(n11855) );
  NAND3_X1 U12365 ( .A1(n15776), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20184), 
        .ZN(n20456) );
  NAND3_X1 U12366 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15777), .A3(n20184), 
        .ZN(n20455) );
  INV_X1 U12367 ( .A(n20456), .ZN(n20564) );
  INV_X1 U12368 ( .A(n20455), .ZN(n20563) );
  NOR2_X1 U12369 ( .A1(n20108), .A2(n18098), .ZN(n20203) );
  INV_X1 U12370 ( .A(n20109), .ZN(n20114) );
  INV_X1 U12371 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n22444) );
  INV_X1 U12372 ( .A(n21932), .ZN(n21657) );
  OAI22_X1 U12373 ( .A1(n21654), .A2(n21985), .B1(n14496), .B2(n21657), .ZN(
        n18705) );
  NAND2_X1 U12374 ( .A1(n18894), .A2(n11289), .ZN(n18965) );
  NOR2_X1 U12375 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n21128), .ZN(n21146) );
  NOR2_X1 U12376 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n21100), .ZN(n21118) );
  NAND2_X1 U12377 ( .A1(n21638), .A2(n14501), .ZN(n11646) );
  INV_X1 U12378 ( .A(n19198), .ZN(n19199) );
  AOI211_X1 U12379 ( .C1(n22463), .C2(n17980), .A(n19254), .B(
        P3_STATE_REG_0__SCAN_IN), .ZN(n17989) );
  OR2_X1 U12380 ( .A1(n20959), .A2(n14439), .ZN(n20969) );
  INV_X1 U12381 ( .A(n18574), .ZN(n20966) );
  AND2_X1 U12382 ( .A1(n18894), .A2(n11522), .ZN(n14457) );
  AND2_X1 U12383 ( .A1(n11289), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11522) );
  NAND2_X1 U12384 ( .A1(n18894), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18968) );
  NOR2_X1 U12385 ( .A1(n18909), .A2(n21358), .ZN(n18894) );
  NOR2_X1 U12386 ( .A1(n11527), .A2(n11526), .ZN(n11525) );
  NAND2_X1 U12387 ( .A1(n18816), .A2(n11280), .ZN(n18848) );
  NOR2_X1 U12388 ( .A1(n18836), .A2(n18835), .ZN(n18816) );
  AND2_X1 U12389 ( .A1(n21167), .A2(n11535), .ZN(n18737) );
  AND2_X1 U12390 ( .A1(n11281), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11535) );
  NAND2_X1 U12391 ( .A1(n21167), .A2(n11281), .ZN(n18736) );
  AND2_X1 U12392 ( .A1(n21167), .A2(n11536), .ZN(n18984) );
  OAI21_X1 U12393 ( .B1(n18937), .B2(n21027), .A(n19862), .ZN(n18936) );
  AND2_X1 U12394 ( .A1(n19001), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18812) );
  NAND2_X1 U12395 ( .A1(n21167), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18772) );
  NOR2_X1 U12396 ( .A1(n21154), .A2(n18995), .ZN(n21167) );
  INV_X1 U12397 ( .A(n18936), .ZN(n18889) );
  NAND2_X1 U12398 ( .A1(n18993), .A2(n19055), .ZN(n21154) );
  NOR2_X1 U12399 ( .A1(n18769), .A2(n21756), .ZN(n21766) );
  AOI22_X1 U12400 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18664), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14348) );
  AOI22_X1 U12401 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14349) );
  AOI211_X1 U12402 ( .C1(n11163), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n14346), .B(n14345), .ZN(n14347) );
  NOR2_X1 U12403 ( .A1(n19079), .A2(n21078), .ZN(n19055) );
  NAND2_X1 U12404 ( .A1(n19097), .A2(n18724), .ZN(n19091) );
  INV_X1 U12405 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21051) );
  XNOR2_X1 U12406 ( .A(n18716), .B(n21699), .ZN(n19126) );
  INV_X1 U12407 ( .A(n19144), .ZN(n19112) );
  AOI211_X1 U12408 ( .C1(n11152), .C2(n18900), .A(n18899), .B(n18898), .ZN(
        n18901) );
  AND2_X1 U12409 ( .A1(n21931), .A2(n21932), .ZN(n21945) );
  INV_X1 U12410 ( .A(n21952), .ZN(n18942) );
  NAND2_X1 U12411 ( .A1(n18873), .A2(n18872), .ZN(n18879) );
  INV_X1 U12412 ( .A(n22022), .ZN(n22013) );
  NOR2_X1 U12413 ( .A1(n18746), .A2(n18745), .ZN(n18980) );
  NAND2_X1 U12414 ( .A1(n18747), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18744) );
  INV_X1 U12415 ( .A(n18812), .ZN(n22008) );
  INV_X1 U12416 ( .A(n19019), .ZN(n21946) );
  INV_X1 U12417 ( .A(n18755), .ZN(n21812) );
  NOR2_X1 U12418 ( .A1(n21811), .A2(n19002), .ZN(n19001) );
  OAI21_X1 U12419 ( .B1(n14497), .B2(n11475), .A(n11474), .ZN(n21892) );
  INV_X1 U12420 ( .A(n14498), .ZN(n11475) );
  INV_X1 U12421 ( .A(n14516), .ZN(n11474) );
  INV_X1 U12422 ( .A(n18742), .ZN(n19021) );
  NOR2_X1 U12423 ( .A1(n17988), .A2(n21429), .ZN(n14500) );
  NAND2_X1 U12424 ( .A1(n18734), .A2(n19050), .ZN(n21769) );
  NOR2_X1 U12425 ( .A1(n21657), .A2(n21935), .ZN(n22011) );
  INV_X1 U12426 ( .A(n18704), .ZN(n11659) );
  INV_X1 U12427 ( .A(n19066), .ZN(n11660) );
  NAND2_X1 U12428 ( .A1(n19075), .A2(n18728), .ZN(n19069) );
  XNOR2_X1 U12429 ( .A(n18727), .B(n11441), .ZN(n19076) );
  INV_X1 U12430 ( .A(n18726), .ZN(n11441) );
  NAND2_X1 U12431 ( .A1(n19076), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19075) );
  NOR2_X1 U12432 ( .A1(n14518), .A2(n14498), .ZN(n22067) );
  XNOR2_X1 U12433 ( .A(n18722), .B(n11440), .ZN(n19099) );
  INV_X1 U12434 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U12435 ( .A1(n19099), .A2(n19098), .ZN(n19097) );
  AND3_X1 U12436 ( .A1(n14489), .A2(n21648), .A3(n14505), .ZN(n14487) );
  OAI21_X1 U12437 ( .B1(n14371), .B2(n14491), .A(n14479), .ZN(n21647) );
  NAND2_X1 U12438 ( .A1(n14506), .A2(n14488), .ZN(n14518) );
  NAND2_X1 U12439 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21638), .ZN(
        n14515) );
  OR2_X1 U12440 ( .A1(n21624), .A2(n14340), .ZN(n17963) );
  NOR2_X1 U12441 ( .A1(n14414), .A2(n14413), .ZN(n21652) );
  NOR2_X1 U12442 ( .A1(n14403), .A2(n14402), .ZN(n19819) );
  NOR2_X1 U12443 ( .A1(n14425), .A2(n14424), .ZN(n21656) );
  NOR2_X1 U12444 ( .A1(n14383), .A2(n14382), .ZN(n19739) );
  INV_X1 U12445 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19653) );
  NAND2_X1 U12446 ( .A1(n22095), .A2(n19612), .ZN(n19863) );
  NOR2_X1 U12447 ( .A1(n21641), .A2(n14439), .ZN(n20967) );
  AOI211_X1 U12448 ( .C1(n20959), .C2(n20958), .A(n22418), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n14534) );
  INV_X1 U12449 ( .A(n22470), .ZN(n22418) );
  OR2_X1 U12450 ( .A1(n16578), .A2(n14309), .ZN(n16569) );
  OR2_X1 U12451 ( .A1(n22104), .A2(n14204), .ZN(n22255) );
  INV_X1 U12452 ( .A(n22358), .ZN(n22374) );
  INV_X1 U12453 ( .A(n22371), .ZN(n22337) );
  INV_X1 U12454 ( .A(n22248), .ZN(n22323) );
  NOR2_X2 U12455 ( .A1(n14313), .A2(n14304), .ZN(n22327) );
  OR2_X1 U12456 ( .A1(n22248), .A2(n22238), .ZN(n22339) );
  INV_X1 U12457 ( .A(n22275), .ZN(n22259) );
  INV_X1 U12458 ( .A(n20833), .ZN(n16714) );
  AND2_X2 U12459 ( .A1(n14776), .A2(n14775), .ZN(n20833) );
  AND2_X1 U12460 ( .A1(n11155), .A2(n14927), .ZN(n14775) );
  INV_X1 U12461 ( .A(n16854), .ZN(n16756) );
  NAND2_X1 U12462 ( .A1(n16834), .A2(n14931), .ZN(n16792) );
  INV_X1 U12463 ( .A(n16823), .ZN(n16794) );
  NOR2_X2 U12464 ( .A1(n16744), .A2(n16757), .ZN(n16825) );
  AND2_X1 U12465 ( .A1(n16792), .A2(n16744), .ZN(n16836) );
  NOR2_X1 U12466 ( .A1(n20709), .A2(n22106), .ZN(n20722) );
  BUF_X1 U12468 ( .A(n20725), .Z(n22106) );
  OAI21_X1 U12469 ( .B1(n14721), .B2(n22424), .A(n14720), .ZN(n22528) );
  INV_X1 U12471 ( .A(n22525), .ZN(n22527) );
  XNOR2_X1 U12472 ( .A(n13793), .B(n13792), .ZN(n14314) );
  INV_X1 U12473 ( .A(n13787), .ZN(n13788) );
  INV_X1 U12474 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15381) );
  NAND2_X1 U12475 ( .A1(n16839), .A2(n16840), .ZN(n16849) );
  AND3_X1 U12476 ( .A1(n11645), .A2(n11637), .A3(n11638), .ZN(n16872) );
  INV_X1 U12477 ( .A(n11645), .ZN(n16879) );
  NOR2_X1 U12478 ( .A1(n20881), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22190) );
  INV_X1 U12479 ( .A(n22223), .ZN(n22188) );
  NAND2_X1 U12480 ( .A1(n11627), .A2(n11425), .ZN(n11424) );
  INV_X1 U12481 ( .A(n11426), .ZN(n11425) );
  INV_X1 U12482 ( .A(n15120), .ZN(n15118) );
  INV_X1 U12483 ( .A(n22609), .ZN(n17151) );
  INV_X1 U12484 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14761) );
  NOR2_X1 U12485 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17977) );
  INV_X1 U12486 ( .A(n22782), .ZN(n22696) );
  OR2_X1 U12487 ( .A1(n22562), .A2(n15197), .ZN(n22782) );
  NOR2_X2 U12488 ( .A1(n22562), .A2(n22548), .ZN(n22789) );
  NAND2_X1 U12489 ( .A1(n15120), .A2(n15057), .ZN(n22602) );
  NAND2_X1 U12490 ( .A1(n15045), .A2(n15148), .ZN(n22814) );
  OAI211_X1 U12491 ( .C1(n17151), .C2(n15052), .A(n15051), .B(n15205), .ZN(
        n22811) );
  NOR2_X1 U12492 ( .A1(n15187), .A2(n15007), .ZN(n22708) );
  NOR2_X1 U12493 ( .A1(n15187), .A2(n15033), .ZN(n22769) );
  AND2_X1 U12494 ( .A1(n15149), .A2(n15148), .ZN(n22832) );
  NAND2_X1 U12495 ( .A1(n15149), .A2(n15147), .ZN(n22650) );
  OAI21_X1 U12496 ( .B1(n14983), .B2(n14982), .A(n15205), .ZN(n22847) );
  INV_X1 U12497 ( .A(n22838), .ZN(n22844) );
  NAND2_X1 U12498 ( .A1(n13292), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22402) );
  NOR2_X1 U12499 ( .A1(n16108), .A2(n22393), .ZN(n22396) );
  INV_X1 U12500 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22556) );
  INV_X1 U12501 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n22388) );
  INV_X1 U12502 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22392) );
  INV_X1 U12503 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22393) );
  OR2_X1 U12504 ( .A1(n17193), .A2(n17194), .ZN(n17196) );
  NOR2_X1 U12505 ( .A1(n19361), .A2(n19360), .ZN(n19359) );
  AND2_X1 U12506 ( .A1(n11729), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11516) );
  OR3_X1 U12507 ( .A1(n19275), .A2(n12214), .A3(n12213), .ZN(n19386) );
  INV_X1 U12508 ( .A(n19386), .ZN(n19494) );
  INV_X1 U12509 ( .A(n19393), .ZN(n19492) );
  NAND2_X1 U12510 ( .A1(n19275), .A2(n12206), .ZN(n19467) );
  INV_X1 U12511 ( .A(n19563), .ZN(n19484) );
  NAND2_X1 U12512 ( .A1(n12021), .A2(n12020), .ZN(n17240) );
  OR3_X1 U12513 ( .A1(n14547), .A2(n12448), .A3(n12211), .ZN(n19464) );
  INV_X1 U12514 ( .A(n19467), .ZN(n19498) );
  CLKBUF_X1 U12515 ( .A(n15634), .Z(n15635) );
  CLKBUF_X1 U12516 ( .A(n15632), .Z(n15633) );
  CLKBUF_X1 U12517 ( .A(n15251), .Z(n15252) );
  INV_X1 U12518 ( .A(n17303), .ZN(n17316) );
  NOR2_X1 U12519 ( .A1(n17286), .A2(n11668), .ZN(n11663) );
  AND2_X1 U12520 ( .A1(n15614), .A2(n15776), .ZN(n20048) );
  OR2_X1 U12521 ( .A1(n15614), .A2(n17344), .ZN(n20072) );
  AND2_X1 U12522 ( .A1(n20405), .A2(n20548), .ZN(n20081) );
  INV_X1 U12523 ( .A(n20548), .ZN(n20497) );
  INV_X2 U12525 ( .A(n14650), .ZN(n14607) );
  OR2_X1 U12526 ( .A1(n17601), .A2(n11485), .ZN(n11480) );
  INV_X1 U12527 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17626) );
  AND2_X1 U12528 ( .A1(n18093), .A2(n12875), .ZN(n18088) );
  OR2_X1 U12529 ( .A1(n19583), .A2(n11259), .ZN(n18063) );
  INV_X1 U12530 ( .A(n18093), .ZN(n17612) );
  NOR2_X1 U12531 ( .A1(n11264), .A2(n11608), .ZN(n16044) );
  NAND2_X1 U12532 ( .A1(n16019), .A2(n11729), .ZN(n16021) );
  NAND2_X1 U12533 ( .A1(n16051), .A2(n16052), .ZN(n16053) );
  AND2_X1 U12534 ( .A1(n17262), .A2(n17261), .ZN(n19450) );
  NAND2_X1 U12535 ( .A1(n11159), .A2(n11491), .ZN(n11490) );
  AOI21_X1 U12536 ( .B1(n15973), .B2(n11493), .A(n11331), .ZN(n11492) );
  OAI21_X1 U12537 ( .B1(n17551), .B2(n15965), .A(n11691), .ZN(n17526) );
  NAND2_X1 U12538 ( .A1(n11576), .A2(n17632), .ZN(n17623) );
  NAND2_X1 U12539 ( .A1(n11230), .A2(n17631), .ZN(n11576) );
  NAND2_X1 U12540 ( .A1(n11585), .A2(n11586), .ZN(n15824) );
  OR2_X1 U12541 ( .A1(n12796), .A2(n12797), .ZN(n11585) );
  NAND2_X1 U12542 ( .A1(n15546), .A2(n15547), .ZN(n11376) );
  INV_X1 U12543 ( .A(n19514), .ZN(n19550) );
  INV_X1 U12544 ( .A(n19542), .ZN(n19527) );
  NAND2_X1 U12545 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18096) );
  INV_X1 U12546 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20161) );
  INV_X1 U12547 ( .A(n20222), .ZN(n20254) );
  INV_X1 U12548 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20140) );
  NAND2_X1 U12549 ( .A1(n15598), .A2(n12261), .ZN(n15555) );
  NOR2_X1 U12550 ( .A1(n14658), .A2(n14657), .ZN(n20554) );
  BUF_X1 U12551 ( .A(n11237), .Z(n17957) );
  INV_X1 U12552 ( .A(n20447), .ZN(n18109) );
  CLKBUF_X1 U12553 ( .A(n14901), .Z(n14902) );
  INV_X1 U12554 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15784) );
  INV_X1 U12555 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20400) );
  AOI21_X1 U12556 ( .B1(n15769), .B2(n15779), .A(n20558), .ZN(n20672) );
  AND2_X1 U12557 ( .A1(n20249), .A2(n20191), .ZN(n20668) );
  AND2_X1 U12558 ( .A1(n20249), .A2(n20218), .ZN(n20649) );
  INV_X1 U12559 ( .A(n20632), .ZN(n20634) );
  OAI21_X1 U12560 ( .B1(n20200), .B2(n20196), .A(n20195), .ZN(n20629) );
  INV_X1 U12561 ( .A(n20625), .ZN(n20615) );
  NAND2_X1 U12562 ( .A1(n20149), .A2(n20232), .ZN(n20606) );
  OR3_X1 U12563 ( .A1(n20142), .A2(n20558), .A3(n20141), .ZN(n20597) );
  OAI21_X1 U12564 ( .B1(n20146), .B2(n20145), .A(n20144), .ZN(n20596) );
  INV_X1 U12565 ( .A(n20600), .ZN(n20589) );
  OAI22_X1 U12566 ( .A1(n20926), .A2(n20455), .B1(n21504), .B2(n20456), .ZN(
        n20397) );
  AOI22_X1 U12567 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n20564), .B1(
        BUF1_REG_16__SCAN_IN), .B2(n20563), .ZN(n20660) );
  INV_X1 U12568 ( .A(n20653), .ZN(n20664) );
  INV_X1 U12569 ( .A(n20351), .ZN(n20356) );
  INV_X1 U12570 ( .A(n20510), .ZN(n20583) );
  AOI22_X1 U12571 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n20564), .B1(
        BUF1_REG_17__SCAN_IN), .B2(n20563), .ZN(n20538) );
  INV_X1 U12572 ( .A(n20485), .ZN(n20490) );
  INV_X1 U12573 ( .A(n20445), .ZN(n20437) );
  INV_X1 U12574 ( .A(n20580), .ZN(n20507) );
  NAND2_X1 U12575 ( .A1(n20114), .A2(n20232), .ZN(n20580) );
  AOI22_X1 U12576 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20563), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20564), .ZN(n20244) );
  OAI21_X1 U12577 ( .B1(n20103), .B2(n20102), .A(n20101), .ZN(n20571) );
  INV_X1 U12578 ( .A(n20660), .ZN(n20667) );
  AOI22_X1 U12579 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20563), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20564), .ZN(n20653) );
  INV_X1 U12580 ( .A(n20538), .ZN(n20542) );
  AND2_X1 U12581 ( .A1(n11259), .A2(n20560), .ZN(n20539) );
  OAI22_X1 U12582 ( .A1(n21520), .A2(n20456), .B1(n20922), .B2(n20455), .ZN(
        n20491) );
  AOI22_X1 U12583 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20564), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n20563), .ZN(n20485) );
  AND2_X1 U12584 ( .A1(n15778), .A2(n20560), .ZN(n20441) );
  AOI22_X1 U12585 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n20564), .B1(
        BUF1_REG_19__SCAN_IN), .B2(n20563), .ZN(n20445) );
  INV_X1 U12586 ( .A(n20391), .ZN(n20396) );
  INV_X1 U12587 ( .A(n20397), .ZN(n20394) );
  OAI22_X1 U12588 ( .A1(n20928), .A2(n20455), .B1(n21498), .B2(n20456), .ZN(
        n20357) );
  AOI22_X1 U12589 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20563), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20564), .ZN(n20351) );
  INV_X1 U12590 ( .A(n20412), .ZN(n20663) );
  INV_X1 U12591 ( .A(n20305), .ZN(n20308) );
  AOI22_X1 U12592 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20563), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20564), .ZN(n20302) );
  INV_X1 U12593 ( .A(n20568), .ZN(n20570) );
  AND3_X1 U12594 ( .A1(n17948), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n19570) );
  AND2_X1 U12595 ( .A1(n15356), .A2(n15355), .ZN(n19571) );
  NOR2_X1 U12596 ( .A1(n18186), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n18184) );
  NOR2_X1 U12598 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n22444), .ZN(n22449) );
  INV_X1 U12599 ( .A(n14455), .ZN(n20954) );
  NOR2_X1 U12600 ( .A1(n14486), .A2(n14485), .ZN(n20961) );
  NAND2_X1 U12601 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n14535), .ZN(n21653) );
  NAND2_X1 U12602 ( .A1(n22097), .A2(n18705), .ZN(n22101) );
  NAND2_X1 U12603 ( .A1(n21242), .A2(n21399), .ZN(n21243) );
  NOR2_X1 U12604 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n21209), .ZN(n21233) );
  NAND2_X1 U12605 ( .A1(n21230), .A2(n21231), .ZN(n21242) );
  OR2_X1 U12606 ( .A1(n21214), .A2(n11528), .ZN(n21230) );
  NOR2_X1 U12607 ( .A1(n21228), .A2(n21229), .ZN(n11528) );
  INV_X1 U12608 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n21149) );
  INV_X1 U12609 ( .A(n21404), .ZN(n21357) );
  INV_X1 U12610 ( .A(n21397), .ZN(n21423) );
  AND2_X1 U12611 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18483), .ZN(n18478) );
  AND2_X1 U12612 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n18508), .ZN(n18493) );
  AND2_X1 U12613 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18494), .ZN(n18508) );
  NAND3_X1 U12614 ( .A1(n14393), .A2(n14392), .A3(n14391), .ZN(n21533) );
  INV_X1 U12615 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18662) );
  INV_X1 U12616 ( .A(n18562), .ZN(n18572) );
  NOR2_X1 U12617 ( .A1(n21563), .A2(n21558), .ZN(n21557) );
  INV_X1 U12618 ( .A(n21569), .ZN(n21534) );
  NOR2_X1 U12619 ( .A1(n21533), .A2(n21574), .ZN(n21570) );
  NOR3_X1 U12620 ( .A1(n21581), .A2(n21532), .A3(n21531), .ZN(n21575) );
  NOR2_X1 U12621 ( .A1(n21533), .A2(n21581), .ZN(n21527) );
  NOR2_X1 U12622 ( .A1(n21645), .A2(n21600), .ZN(n21579) );
  NOR2_X2 U12623 ( .A1(n21497), .A2(n21600), .ZN(n21580) );
  NOR2_X1 U12624 ( .A1(n21593), .A2(n21592), .ZN(n21590) );
  NOR2_X1 U12625 ( .A1(n21435), .A2(n21605), .ZN(n21591) );
  AND2_X1 U12626 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n21468), .ZN(n21598) );
  NOR2_X1 U12627 ( .A1(n18591), .A2(n18590), .ZN(n21661) );
  NOR2_X1 U12628 ( .A1(n18601), .A2(n18600), .ZN(n21470) );
  NOR2_X1 U12629 ( .A1(n18611), .A2(n18610), .ZN(n21479) );
  NOR2_X1 U12630 ( .A1(n21490), .A2(n21614), .ZN(n21486) );
  INV_X1 U12631 ( .A(n21611), .ZN(n21603) );
  INV_X1 U12632 ( .A(n21612), .ZN(n21487) );
  NOR2_X1 U12633 ( .A1(n18686), .A2(n11444), .ZN(n18687) );
  NOR2_X1 U12634 ( .A1(n19216), .A2(n19199), .ZN(n19208) );
  NOR2_X1 U12637 ( .A1(n21888), .A2(n21957), .ZN(n21885) );
  NOR2_X1 U12638 ( .A1(n18947), .A2(n21888), .ZN(n18962) );
  NAND2_X1 U12639 ( .A1(n18903), .A2(n21951), .ZN(n21931) );
  NAND2_X1 U12640 ( .A1(n18816), .A2(n11263), .ZN(n18923) );
  NAND2_X1 U12641 ( .A1(n18812), .A2(n18866), .ZN(n18947) );
  NAND2_X1 U12642 ( .A1(n18866), .A2(n21812), .ZN(n21957) );
  NAND2_X1 U12643 ( .A1(n18737), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18836) );
  AND3_X1 U12644 ( .A1(n21658), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18988), .ZN(n18885) );
  NOR2_X1 U12645 ( .A1(n19104), .A2(n21051), .ZN(n19088) );
  INV_X1 U12646 ( .A(n19140), .ZN(n19107) );
  INV_X1 U12647 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21619) );
  INV_X1 U12648 ( .A(n19072), .ZN(n19148) );
  INV_X1 U12649 ( .A(n22011), .ZN(n21987) );
  NAND2_X1 U12650 ( .A1(n18901), .A2(n21874), .ZN(n21952) );
  AOI21_X1 U12651 ( .B1(n11648), .B2(n11647), .A(n21947), .ZN(n21948) );
  NAND2_X1 U12652 ( .A1(n21944), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11647) );
  NAND2_X1 U12653 ( .A1(n21945), .A2(n21946), .ZN(n11648) );
  NOR2_X1 U12654 ( .A1(n21811), .A2(n18992), .ZN(n21820) );
  INV_X1 U12655 ( .A(n21892), .ZN(n22068) );
  INV_X1 U12656 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21755) );
  NAND2_X1 U12657 ( .A1(n11652), .A2(n11650), .ZN(n19080) );
  NAND2_X1 U12658 ( .A1(n20961), .A2(n14487), .ZN(n21894) );
  NOR2_X1 U12659 ( .A1(n19123), .A2(n19122), .ZN(n19121) );
  AND2_X1 U12660 ( .A1(n11658), .A2(n11272), .ZN(n19123) );
  NOR2_X1 U12661 ( .A1(n21869), .A2(n22048), .ZN(n21962) );
  AOI22_X1 U12662 ( .A1(n22087), .A2(n21618), .B1(P3_STATE2_REG_1__SCAN_IN), 
        .B2(n21834), .ZN(n11456) );
  INV_X1 U12663 ( .A(n21653), .ZN(n22097) );
  AOI21_X1 U12664 ( .B1(n11468), .B2(n11466), .A(n11464), .ZN(n14533) );
  INV_X1 U12665 ( .A(n11467), .ZN(n11466) );
  INV_X1 U12666 ( .A(n11469), .ZN(n11468) );
  INV_X1 U12667 ( .A(n14332), .ZN(n15793) );
  OAI21_X1 U12668 ( .B1(n14331), .B2(n14330), .A(P1_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14332) );
  CLKBUF_X1 U12669 ( .A(n19738), .Z(n19945) );
  INV_X1 U12670 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20675) );
  OAI21_X1 U12671 ( .B1(n17021), .B2(n22385), .A(n11405), .ZN(P1_U2971) );
  INV_X1 U12672 ( .A(n11406), .ZN(n11405) );
  AOI21_X1 U12673 ( .B1(n16863), .B2(n20862), .A(n16862), .ZN(n11407) );
  OAI211_X1 U12674 ( .C1(n16991), .C2(n22218), .A(n11555), .B(n11554), .ZN(
        P1_U3000) );
  NOR3_X1 U12675 ( .A1(n16990), .A2(n16989), .A3(n16988), .ZN(n11554) );
  NAND2_X1 U12676 ( .A1(n11556), .A2(n22199), .ZN(n11555) );
  NAND2_X1 U12677 ( .A1(n11506), .A2(n17439), .ZN(n11505) );
  AND2_X1 U12678 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  AND2_X1 U12679 ( .A1(n14154), .A2(n14153), .ZN(n14155) );
  AND2_X1 U12680 ( .A1(n14144), .A2(n14143), .ZN(n14145) );
  NAND2_X1 U12681 ( .A1(n11301), .A2(n18089), .ZN(n11399) );
  NAND2_X1 U12682 ( .A1(n11301), .A2(n19530), .ZN(n11398) );
  AOI211_X1 U12683 ( .C1(n17669), .C2(n19537), .A(n17668), .B(n17667), .ZN(
        n17670) );
  AOI21_X1 U12684 ( .B1(n11534), .B2(n11533), .A(n11529), .ZN(n21402) );
  XNOR2_X1 U12685 ( .A(n21408), .B(n18959), .ZN(n11534) );
  AOI21_X1 U12686 ( .B1(n18957), .B2(n11452), .A(n11449), .ZN(n18960) );
  OAI211_X1 U12687 ( .C1(n18978), .C2(n11452), .A(n11451), .B(n11450), .ZN(
        n11449) );
  INV_X1 U12688 ( .A(n11455), .ZN(n21617) );
  INV_X1 U12689 ( .A(n21634), .ZN(n11457) );
  NAND2_X1 U12690 ( .A1(n11473), .A2(n11471), .ZN(P3_U2997) );
  NOR2_X1 U12691 ( .A1(n11533), .A2(n11472), .ZN(n11471) );
  OR2_X1 U12692 ( .A1(n22086), .A2(n17984), .ZN(n11472) );
  AND2_X1 U12693 ( .A1(n11284), .A2(n11525), .ZN(n11263) );
  NAND2_X1 U12694 ( .A1(n11594), .A2(n11363), .ZN(n15804) );
  OR2_X2 U12695 ( .A1(n21618), .A2(n17963), .ZN(n11293) );
  OR2_X1 U12696 ( .A1(n17330), .A2(n17331), .ZN(n11264) );
  OR2_X1 U12697 ( .A1(n17364), .A2(n17365), .ZN(n11265) );
  AND2_X1 U12698 ( .A1(n13537), .A2(n11705), .ZN(n16610) );
  NAND2_X1 U12699 ( .A1(n11700), .A2(n13485), .ZN(n16645) );
  OR2_X1 U12700 ( .A1(n11757), .A2(n11521), .ZN(n11266) );
  NOR2_X1 U12701 ( .A1(n11753), .A2(n18071), .ZN(n11754) );
  AND2_X1 U12702 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11755) );
  OR3_X1 U12703 ( .A1(n12673), .A2(n12667), .A3(n11348), .ZN(n11268) );
  AND2_X1 U12704 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11269) );
  AND2_X1 U12705 ( .A1(n14881), .A2(n11351), .ZN(n11270) );
  AND2_X1 U12706 ( .A1(n11500), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11271) );
  INV_X1 U12707 ( .A(n11492), .ZN(n17484) );
  OR2_X1 U12708 ( .A1(n21606), .A2(n21691), .ZN(n11272) );
  INV_X1 U12709 ( .A(n11495), .ZN(n11491) );
  INV_X1 U12710 ( .A(n11496), .ZN(n11495) );
  INV_X1 U12711 ( .A(n12064), .ZN(n12057) );
  AND3_X1 U12712 ( .A1(n12800), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n12799), .ZN(n11274) );
  AND2_X1 U12713 ( .A1(n11269), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11275) );
  AND2_X1 U12714 ( .A1(n12638), .A2(n11352), .ZN(n11276) );
  AND2_X1 U12715 ( .A1(n11312), .A2(n11505), .ZN(n11277) );
  AND2_X1 U12716 ( .A1(n11270), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11278) );
  NAND2_X1 U12717 ( .A1(n14879), .A2(n14881), .ZN(n14880) );
  NAND2_X1 U12718 ( .A1(n15600), .A2(n15599), .ZN(n15598) );
  AND2_X1 U12719 ( .A1(n15251), .A2(n11678), .ZN(n15385) );
  OR2_X1 U12720 ( .A1(n15634), .A2(n11675), .ZN(n11279) );
  AND2_X1 U12721 ( .A1(n11356), .A2(n15598), .ZN(n15554) );
  AND2_X1 U12722 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11280) );
  AND3_X1 U12723 ( .A1(n12292), .A2(n12291), .A3(n12290), .ZN(n17921) );
  NAND2_X1 U12724 ( .A1(n15387), .A2(n11620), .ZN(n15799) );
  AND2_X1 U12725 ( .A1(n11536), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11281) );
  AND2_X1 U12726 ( .A1(n11323), .A2(n11565), .ZN(n11282) );
  AND2_X1 U12727 ( .A1(n11706), .A2(n15687), .ZN(n11283) );
  AND2_X1 U12728 ( .A1(n11280), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11284) );
  NAND2_X1 U12729 ( .A1(n11743), .A2(n11269), .ZN(n11738) );
  NAND2_X1 U12730 ( .A1(n11160), .A2(n16987), .ZN(n11285) );
  OR2_X1 U12731 ( .A1(n17921), .A2(n17223), .ZN(n11286) );
  AND2_X1 U12732 ( .A1(n11283), .A2(n15853), .ZN(n11287) );
  AND2_X1 U12733 ( .A1(n11263), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11288) );
  AND2_X1 U12734 ( .A1(n14879), .A2(n11270), .ZN(n14959) );
  NOR3_X1 U12735 ( .A1(n11732), .A2(n11514), .A3(n17468), .ZN(n11768) );
  NAND2_X1 U12736 ( .A1(n11736), .A2(n11271), .ZN(n11767) );
  NAND2_X1 U12737 ( .A1(n11736), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11765) );
  AND2_X1 U12738 ( .A1(n11523), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11289) );
  AND2_X1 U12739 ( .A1(n11551), .A2(n15985), .ZN(n11290) );
  OR3_X1 U12740 ( .A1(n16735), .A2(n11561), .A3(n16724), .ZN(n11292) );
  NAND2_X1 U12741 ( .A1(n11639), .A2(n17134), .ZN(n11294) );
  NAND3_X1 U12742 ( .A1(n14349), .A2(n14348), .A3(n14347), .ZN(n21641) );
  INV_X2 U12743 ( .A(n21641), .ZN(n20959) );
  OR2_X1 U12744 ( .A1(n16537), .A2(n11708), .ZN(n11296) );
  NAND2_X1 U12745 ( .A1(n13537), .A2(n11704), .ZN(n16611) );
  AND4_X1 U12746 ( .A1(n12908), .A2(n12907), .A3(n12906), .A4(n12905), .ZN(
        n11297) );
  OR2_X1 U12747 ( .A1(n12673), .A2(n12667), .ZN(n11298) );
  AND4_X1 U12748 ( .A1(n12970), .A2(n12969), .A3(n12968), .A4(n12967), .ZN(
        n11299) );
  NAND2_X1 U12749 ( .A1(n15909), .A2(n15908), .ZN(n15910) );
  NAND2_X1 U12750 ( .A1(n13537), .A2(n13536), .ZN(n16622) );
  AND2_X1 U12751 ( .A1(n13219), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11300) );
  XOR2_X1 U12752 ( .A(n17424), .B(n17423), .Z(n11301) );
  AND2_X1 U12753 ( .A1(n11660), .A2(n11659), .ZN(n11302) );
  NAND2_X1 U12754 ( .A1(n12648), .A2(n17619), .ZN(n17610) );
  NAND2_X1 U12755 ( .A1(n11490), .A2(n11494), .ZN(n17473) );
  NAND2_X1 U12756 ( .A1(n11383), .A2(n12658), .ZN(n17601) );
  AND2_X1 U12757 ( .A1(n13816), .A2(n13828), .ZN(n14764) );
  AND2_X1 U12758 ( .A1(n17551), .A2(n17550), .ZN(n17535) );
  OR2_X1 U12759 ( .A1(n16756), .A2(n22377), .ZN(n11303) );
  INV_X1 U12760 ( .A(n14770), .ZN(n15016) );
  OR3_X1 U12761 ( .A1(n12673), .A2(n11544), .A3(n12667), .ZN(n11304) );
  AND2_X1 U12762 ( .A1(n16942), .A2(n17089), .ZN(n11305) );
  NAND2_X1 U12763 ( .A1(n13099), .A2(n13098), .ZN(n14935) );
  OR2_X1 U12764 ( .A1(n21699), .A2(n18690), .ZN(n11306) );
  AND2_X1 U12765 ( .A1(n20969), .A2(n14499), .ZN(n11307) );
  AND2_X1 U12766 ( .A1(n15998), .A2(n16055), .ZN(n11308) );
  INV_X1 U12767 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14501) );
  NAND2_X1 U12768 ( .A1(n17580), .A2(n12810), .ZN(n17571) );
  AND2_X1 U12769 ( .A1(n17420), .A2(n17432), .ZN(n11309) );
  NAND2_X1 U12770 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18701), .ZN(
        n11310) );
  AND4_X1 U12771 ( .A1(n11242), .A2(n12737), .A3(n12014), .A4(n12218), .ZN(
        n11311) );
  AND2_X1 U12772 ( .A1(n12452), .A2(n12451), .ZN(n11312) );
  NAND2_X1 U12773 ( .A1(n11929), .A2(n11290), .ZN(n11313) );
  AND2_X1 U12774 ( .A1(n12808), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11314) );
  INV_X1 U12775 ( .A(n11692), .ZN(n11691) );
  OAI21_X1 U12776 ( .B1(n15965), .B2(n17550), .A(n17534), .ZN(n11692) );
  NAND2_X1 U12777 ( .A1(n17580), .A2(n11402), .ZN(n17478) );
  INV_X1 U12778 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21638) );
  AND3_X1 U12779 ( .A1(n18684), .A2(n11446), .A3(n11445), .ZN(n11315) );
  NAND2_X1 U12780 ( .A1(n11480), .A2(n11484), .ZN(n17593) );
  INV_X2 U12781 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15297) );
  AND2_X1 U12782 ( .A1(n11614), .A2(n11613), .ZN(n11316) );
  AND2_X1 U12783 ( .A1(n16052), .A2(n16049), .ZN(n11317) );
  NAND2_X1 U12784 ( .A1(n13229), .A2(n22168), .ZN(n11318) );
  AND2_X1 U12785 ( .A1(n11600), .A2(n15611), .ZN(n11319) );
  NAND2_X1 U12786 ( .A1(n11382), .A2(n12804), .ZN(n12795) );
  AND2_X1 U12787 ( .A1(n11548), .A2(n12649), .ZN(n11320) );
  INV_X1 U12788 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18071) );
  INV_X1 U12789 ( .A(n11488), .ZN(n11487) );
  NAND2_X1 U12790 ( .A1(n11494), .A2(n11489), .ZN(n11488) );
  INV_X2 U12791 ( .A(n22449), .ZN(n18186) );
  NAND2_X1 U12792 ( .A1(n14206), .A2(n14784), .ZN(n14215) );
  CLKBUF_X3 U12793 ( .A(n14215), .Z(n14293) );
  NOR2_X1 U12794 ( .A1(n17286), .A2(n17288), .ZN(n17279) );
  AND3_X1 U12795 ( .A1(n13360), .A2(n13361), .A3(n11283), .ZN(n11321) );
  NOR2_X1 U12796 ( .A1(n11757), .A2(n11520), .ZN(n11748) );
  NOR2_X1 U12797 ( .A1(n15634), .A2(n11672), .ZN(n15866) );
  NOR2_X1 U12798 ( .A1(n17860), .A2(n11597), .ZN(n15805) );
  NOR2_X1 U12799 ( .A1(n15937), .A2(n11701), .ZN(n16634) );
  NOR2_X1 U12800 ( .A1(n15634), .A2(n15849), .ZN(n15797) );
  NOR2_X1 U12801 ( .A1(n11751), .A2(n18081), .ZN(n11752) );
  NOR2_X1 U12802 ( .A1(n15903), .A2(n15902), .ZN(n15901) );
  OR2_X1 U12803 ( .A1(n11286), .A2(n15732), .ZN(n11322) );
  AND2_X1 U12804 ( .A1(n14236), .A2(n11566), .ZN(n11323) );
  AND2_X1 U12805 ( .A1(n11678), .A2(n15386), .ZN(n11324) );
  AND2_X1 U12806 ( .A1(n12416), .A2(n11602), .ZN(n11325) );
  NOR2_X1 U12807 ( .A1(n11749), .A2(n17626), .ZN(n11750) );
  XNOR2_X1 U12808 ( .A(n12555), .B(n15624), .ZN(n15546) );
  NAND2_X1 U12809 ( .A1(n11376), .A2(n12556), .ZN(n15618) );
  INV_X1 U12810 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13236) );
  AND2_X1 U12811 ( .A1(n11744), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11743) );
  AND2_X1 U12812 ( .A1(n11743), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11739) );
  AND3_X1 U12813 ( .A1(n13360), .A2(n13361), .A3(n11706), .ZN(n11326) );
  AND2_X1 U12814 ( .A1(n15981), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11327) );
  NOR2_X1 U12815 ( .A1(n11714), .A2(n11663), .ZN(n17274) );
  AND2_X1 U12816 ( .A1(n11624), .A2(n11623), .ZN(n11328) );
  AND2_X1 U12817 ( .A1(n11602), .A2(n15889), .ZN(n11329) );
  AND2_X1 U12818 ( .A1(n15984), .A2(n17707), .ZN(n11330) );
  AND2_X1 U12819 ( .A1(n15977), .A2(n17731), .ZN(n11331) );
  OR2_X1 U12820 ( .A1(n13235), .A2(n13139), .ZN(n11332) );
  OR2_X1 U12821 ( .A1(n16735), .A2(n11561), .ZN(n11333) );
  INV_X1 U12822 ( .A(n15937), .ZN(n11700) );
  INV_X1 U12823 ( .A(n11567), .ZN(n16557) );
  NOR2_X1 U12824 ( .A1(n16561), .A2(n16558), .ZN(n11567) );
  NOR2_X1 U12825 ( .A1(n18705), .A2(n11465), .ZN(n11334) );
  AND2_X1 U12826 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11335) );
  INV_X1 U12827 ( .A(n16624), .ZN(n13536) );
  INV_X1 U12828 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17542) );
  AND2_X1 U12829 ( .A1(n15387), .A2(n11618), .ZN(n15800) );
  NAND2_X1 U12830 ( .A1(n11903), .A2(n11549), .ZN(n11336) );
  NAND2_X1 U12831 ( .A1(n11704), .A2(n11703), .ZN(n11337) );
  AND2_X1 U12832 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11338) );
  OR2_X1 U12833 ( .A1(n13139), .A2(n13138), .ZN(n11339) );
  AND2_X1 U12834 ( .A1(n13235), .A2(n13233), .ZN(n11340) );
  AND2_X1 U12835 ( .A1(n17117), .A2(n17116), .ZN(n11341) );
  AND2_X1 U12836 ( .A1(n11324), .A2(n11677), .ZN(n11342) );
  AND2_X1 U12837 ( .A1(n11275), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11343) );
  INV_X1 U12838 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17487) );
  AND2_X1 U12839 ( .A1(n18816), .A2(n11284), .ZN(n11344) );
  NAND2_X1 U12840 ( .A1(n12860), .A2(n15324), .ZN(n19546) );
  INV_X1 U12841 ( .A(n19546), .ZN(n19530) );
  AND2_X1 U12842 ( .A1(n14967), .A2(n11316), .ZN(n15255) );
  NAND2_X1 U12843 ( .A1(n15251), .A2(n15254), .ZN(n15253) );
  OR2_X1 U12844 ( .A1(n17922), .A2(n17921), .ZN(n17220) );
  OR2_X1 U12845 ( .A1(n14811), .A2(n14810), .ZN(n22214) );
  INV_X1 U12846 ( .A(n22214), .ZN(n22199) );
  NAND2_X1 U12847 ( .A1(n14151), .A2(n11616), .ZN(n11345) );
  OR2_X1 U12848 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19019), .ZN(
        n11346) );
  NAND2_X1 U12849 ( .A1(n15716), .A2(n12276), .ZN(n17938) );
  AND2_X1 U12850 ( .A1(n11605), .A2(n11604), .ZN(n11347) );
  INV_X1 U12851 ( .A(n12634), .ZN(n11550) );
  AND2_X1 U12852 ( .A1(n20322), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11348) );
  NAND2_X1 U12853 ( .A1(n15251), .A2(n11324), .ZN(n15682) );
  OR2_X1 U12854 ( .A1(n17276), .A2(n11664), .ZN(n11349) );
  AND2_X1 U12855 ( .A1(n14043), .A2(n14042), .ZN(n11350) );
  NOR2_X1 U12856 ( .A1(n20311), .A2(n20360), .ZN(n11351) );
  NAND2_X1 U12857 ( .A1(n19281), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11352) );
  INV_X1 U12858 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21027) );
  INV_X1 U12859 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n21344) );
  INV_X1 U12860 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17468) );
  NAND2_X1 U12861 ( .A1(n11252), .A2(n11511), .ZN(n11353) );
  AND2_X1 U12862 ( .A1(n11736), .A2(n11500), .ZN(n11354) );
  AND2_X1 U12863 ( .A1(n11743), .A2(n11275), .ZN(n11355) );
  AND2_X1 U12864 ( .A1(n12261), .A2(n11600), .ZN(n11356) );
  AND2_X1 U12865 ( .A1(n11347), .A2(n17371), .ZN(n11357) );
  AND2_X1 U12866 ( .A1(n11655), .A2(n11654), .ZN(n11358) );
  AND2_X1 U12867 ( .A1(n11290), .A2(n15992), .ZN(n11359) );
  INV_X1 U12868 ( .A(n11507), .ZN(n11506) );
  NAND2_X1 U12869 ( .A1(n11353), .A2(n11509), .ZN(n11507) );
  INV_X1 U12870 ( .A(n18065), .ZN(n18089) );
  AND2_X1 U12871 ( .A1(n11730), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11726) );
  NOR2_X1 U12872 ( .A1(n11732), .A2(n17468), .ZN(n11733) );
  XNOR2_X1 U12873 ( .A(n18690), .B(n21699), .ZN(n19122) );
  NOR3_X1 U12874 ( .A1(n11732), .A2(n11513), .A3(n11512), .ZN(n11730) );
  AND2_X1 U12875 ( .A1(n18894), .A2(n11523), .ZN(n11360) );
  AND2_X1 U12876 ( .A1(n21842), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11361) );
  AND2_X1 U12877 ( .A1(n20967), .A2(n14534), .ZN(n11362) );
  NAND3_X1 U12878 ( .A1(n12359), .A2(n12358), .A3(n12357), .ZN(n11363) );
  OR3_X1 U12879 ( .A1(n11732), .A2(n11513), .A3(n11514), .ZN(n11364) );
  NAND2_X1 U12880 ( .A1(n11590), .A2(n11589), .ZN(n12728) );
  INV_X1 U12881 ( .A(n12728), .ZN(n11394) );
  INV_X1 U12882 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11527) );
  INV_X1 U12883 ( .A(n14096), .ZN(n11984) );
  INV_X1 U12884 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11514) );
  INV_X1 U12885 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19636) );
  INV_X1 U12886 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11526) );
  INV_X1 U12887 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11537) );
  INV_X1 U12888 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11524) );
  INV_X1 U12889 ( .A(n16031), .ZN(n11593) );
  INV_X1 U12890 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11501) );
  AND2_X1 U12891 ( .A1(n22418), .A2(n21998), .ZN(n11365) );
  INV_X1 U12892 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11502) );
  INV_X1 U12893 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11452) );
  INV_X1 U12894 ( .A(n17004), .ZN(n11437) );
  AND2_X1 U12895 ( .A1(n17657), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11366) );
  INV_X1 U12896 ( .A(n21400), .ZN(n11533) );
  OR3_X1 U12897 ( .A1(n22393), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14985), 
        .ZN(n15187) );
  OAI21_X2 U12898 ( .B1(n15186), .B2(n20934), .A(n15056), .ZN(n22845) );
  OAI21_X2 U12899 ( .B1(n15186), .B2(n20936), .A(n14997), .ZN(n22655) );
  OAI21_X2 U12900 ( .B1(n15186), .B2(n20922), .A(n15024), .ZN(n22688) );
  OAI21_X2 U12901 ( .B1(n15186), .B2(n20940), .A(n15023), .ZN(n22689) );
  NOR2_X2 U12902 ( .A1(n20322), .A2(n20454), .ZN(n20355) );
  NAND2_X1 U12903 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20257), .ZN(n20454) );
  NAND2_X1 U12904 ( .A1(n11367), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U12905 ( .A1(n11369), .A2(n12077), .ZN(n11367) );
  NAND3_X1 U12906 ( .A1(n12026), .A2(n12025), .A3(n11590), .ZN(n12831) );
  NAND2_X1 U12907 ( .A1(n12076), .A2(n12721), .ZN(n11369) );
  NAND2_X1 U12908 ( .A1(n12037), .A2(n12036), .ZN(n12076) );
  NAND3_X1 U12909 ( .A1(n12061), .A2(n11395), .A3(n11396), .ZN(n11372) );
  AND2_X2 U12910 ( .A1(n11371), .A2(n12086), .ZN(n12456) );
  NAND2_X2 U12911 ( .A1(n11370), .A2(n11374), .ZN(n12086) );
  NAND2_X1 U12912 ( .A1(n11373), .A2(n11372), .ZN(n11371) );
  NAND2_X1 U12913 ( .A1(n11375), .A2(n11276), .ZN(n12641) );
  NAND2_X1 U12914 ( .A1(n11375), .A2(n12638), .ZN(n17635) );
  NAND2_X1 U12915 ( .A1(n18075), .A2(n18076), .ZN(n11375) );
  INV_X1 U12916 ( .A(n12556), .ZN(n11380) );
  NAND3_X1 U12917 ( .A1(n12804), .A2(n11382), .A3(n16007), .ZN(n11381) );
  NAND2_X2 U12918 ( .A1(n11388), .A2(n15991), .ZN(n17456) );
  INV_X1 U12919 ( .A(n17451), .ZN(n11388) );
  OAI21_X1 U12920 ( .B1(n17451), .B2(n11389), .A(n16004), .ZN(n17433) );
  NAND2_X1 U12921 ( .A1(n11393), .A2(n11392), .ZN(n11391) );
  NAND2_X1 U12922 ( .A1(n14125), .A2(n15778), .ZN(n11392) );
  NAND2_X1 U12923 ( .A1(n11394), .A2(n12056), .ZN(n11393) );
  NAND2_X1 U12924 ( .A1(n17656), .A2(n11398), .ZN(P2_U3016) );
  NAND2_X1 U12925 ( .A1(n17430), .A2(n11399), .ZN(P2_U2984) );
  NAND2_X1 U12926 ( .A1(n18073), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11400) );
  NAND2_X1 U12927 ( .A1(n11583), .A2(n11582), .ZN(n11401) );
  AND2_X1 U12928 ( .A1(n16057), .A2(n11366), .ZN(n17435) );
  XNOR2_X1 U12929 ( .A(n17444), .B(n17660), .ZN(n16071) );
  NOR2_X2 U12930 ( .A1(n16620), .A2(n11337), .ZN(n16598) );
  INV_X1 U12931 ( .A(n15935), .ZN(n13467) );
  NAND2_X1 U12932 ( .A1(n13055), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11409) );
  OAI22_X1 U12933 ( .A1(n20848), .A2(n22385), .B1(n20877), .B2(n22321), .ZN(
        n20849) );
  NAND2_X1 U12934 ( .A1(n11415), .A2(n11412), .ZN(n11411) );
  OR2_X1 U12935 ( .A1(n17141), .A2(n11413), .ZN(n11412) );
  INV_X1 U12936 ( .A(n17137), .ZN(n11414) );
  NAND2_X1 U12937 ( .A1(n17141), .A2(n11160), .ZN(n11415) );
  AND2_X2 U12938 ( .A1(n13236), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12885) );
  NOR2_X2 U12939 ( .A1(n11418), .A2(n12609), .ZN(n12633) );
  NAND2_X2 U12940 ( .A1(n12566), .A2(n12785), .ZN(n11418) );
  NOR2_X2 U12941 ( .A1(n17571), .A2(n12811), .ZN(n17567) );
  NOR2_X1 U12942 ( .A1(n12797), .A2(n11419), .ZN(n11581) );
  NAND2_X1 U12943 ( .A1(n11421), .A2(n17134), .ZN(n11638) );
  INV_X1 U12944 ( .A(n11421), .ZN(n11420) );
  NOR2_X1 U12945 ( .A1(n16905), .A2(n11421), .ZN(n16897) );
  OR2_X1 U12946 ( .A1(n11640), .A2(n11421), .ZN(n11639) );
  NAND2_X1 U12947 ( .A1(n11422), .A2(n13026), .ZN(n13001) );
  OAI211_X1 U12948 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n11627), .A(
        n11424), .B(n11427), .ZN(n15380) );
  NAND2_X1 U12949 ( .A1(n11428), .A2(n14216), .ZN(n11427) );
  NAND2_X1 U12950 ( .A1(n11628), .A2(n13214), .ZN(n15644) );
  INV_X1 U12951 ( .A(n15643), .ZN(n11430) );
  NAND2_X1 U12952 ( .A1(n11438), .A2(n11432), .ZN(n16991) );
  NAND2_X1 U12953 ( .A1(n11433), .A2(n11434), .ZN(n11432) );
  NAND3_X1 U12954 ( .A1(n16839), .A2(n16840), .A3(n11435), .ZN(n11433) );
  NAND3_X1 U12955 ( .A1(n16839), .A2(n16840), .A3(n11436), .ZN(n11438) );
  AND2_X1 U12956 ( .A1(n16871), .A2(n17014), .ZN(n11439) );
  XNOR2_X2 U12957 ( .A(n13145), .B(n13144), .ZN(n13311) );
  INV_X2 U12958 ( .A(n18433), .ZN(n18682) );
  NAND3_X1 U12959 ( .A1(n18685), .A2(n18683), .A3(n11315), .ZN(n11444) );
  INV_X2 U12960 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21624) );
  NOR2_X2 U12961 ( .A1(n11454), .A2(n14340), .ZN(n18616) );
  OAI21_X1 U12962 ( .B1(n11461), .B2(n11457), .A(n11456), .ZN(n11455) );
  NOR2_X1 U12963 ( .A1(n11461), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11458) );
  NAND2_X1 U12964 ( .A1(n11461), .A2(n11460), .ZN(n11459) );
  NOR2_X1 U12965 ( .A1(n19636), .A2(n19653), .ZN(n11460) );
  NAND2_X1 U12966 ( .A1(n22059), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11462) );
  NAND2_X1 U12967 ( .A1(n14525), .A2(n21618), .ZN(n11463) );
  NAND3_X1 U12968 ( .A1(n22094), .A2(n14535), .A3(n19687), .ZN(n11473) );
  NOR2_X2 U12969 ( .A1(n11476), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U12970 ( .A1(n17456), .A2(n16049), .ZN(n16051) );
  NAND2_X1 U12971 ( .A1(n17443), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16054) );
  OAI211_X1 U12972 ( .C1(n17456), .C2(n16052), .A(n11479), .B(n11477), .ZN(
        n17443) );
  NAND2_X1 U12973 ( .A1(n11478), .A2(n16050), .ZN(n11477) );
  NAND2_X1 U12974 ( .A1(n17456), .A2(n11317), .ZN(n11479) );
  NAND2_X1 U12975 ( .A1(n15973), .A2(n15972), .ZN(n17493) );
  INV_X1 U12976 ( .A(n17494), .ZN(n11498) );
  NAND2_X1 U12977 ( .A1(n19485), .A2(n11504), .ZN(n11503) );
  NAND2_X1 U12978 ( .A1(n19485), .A2(n19486), .ZN(n19483) );
  OAI211_X1 U12979 ( .C1(n19485), .C2(n11507), .A(n11503), .B(n11277), .ZN(
        P2_U2825) );
  AOI21_X1 U12980 ( .B1(n17411), .B2(n17995), .A(n11516), .ZN(n11737) );
  NAND2_X1 U12981 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11517), .ZN(
        n11751) );
  NAND3_X1 U12982 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11753) );
  INV_X2 U12983 ( .A(n21214), .ZN(n21399) );
  NAND3_X1 U12984 ( .A1(n11543), .A2(n11546), .A3(n11542), .ZN(n11541) );
  INV_X2 U12985 ( .A(n12404), .ZN(n13951) );
  NAND2_X1 U12986 ( .A1(n11320), .A2(n11903), .ZN(n12653) );
  NOR2_X2 U12987 ( .A1(n11924), .A2(n11550), .ZN(n11549) );
  NAND2_X1 U12988 ( .A1(n11929), .A2(n11359), .ZN(n15997) );
  NAND2_X1 U12989 ( .A1(n11929), .A2(n11551), .ZN(n15986) );
  NAND2_X1 U12990 ( .A1(n11929), .A2(n15982), .ZN(n15990) );
  INV_X1 U12991 ( .A(n16647), .ZN(n11563) );
  NOR2_X1 U12992 ( .A1(n16561), .A2(n11568), .ZN(n16530) );
  NAND2_X1 U12993 ( .A1(n15548), .A2(n15549), .ZN(n11573) );
  XNOR2_X2 U12994 ( .A(n12564), .B(n12563), .ZN(n15548) );
  AND2_X2 U12995 ( .A1(n12513), .A2(n12512), .ZN(n12564) );
  OAI21_X1 U12996 ( .B1(n11230), .B2(n11579), .A(n11267), .ZN(n17624) );
  NAND2_X2 U12997 ( .A1(n11575), .A2(n11574), .ZN(n17580) );
  NAND2_X1 U12998 ( .A1(n17633), .A2(n11267), .ZN(n11575) );
  AOI21_X1 U12999 ( .B1(n11581), .B2(n12795), .A(n11274), .ZN(n11580) );
  AOI21_X1 U13000 ( .B1(n11586), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12795), .ZN(n11582) );
  AOI21_X1 U13001 ( .B1(n11587), .B2(n12453), .A(n12108), .ZN(n14883) );
  XNOR2_X2 U13002 ( .A(n11587), .B(n12453), .ZN(n12489) );
  INV_X1 U13003 ( .A(n17860), .ZN(n11594) );
  NAND2_X1 U13004 ( .A1(n11594), .A2(n11595), .ZN(n17815) );
  OR2_X1 U13005 ( .A1(n17922), .A2(n11286), .ZN(n17221) );
  NAND2_X1 U13006 ( .A1(n12425), .A2(n11357), .ZN(n17364) );
  NOR2_X1 U13007 ( .A1(n11264), .A2(n17177), .ZN(n16063) );
  OR3_X1 U13008 ( .A1(n11264), .A2(n11607), .A3(n17177), .ZN(n16039) );
  INV_X1 U13009 ( .A(n16064), .ZN(n11612) );
  INV_X2 U13010 ( .A(n14024), .ZN(n11994) );
  AND2_X2 U13011 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11781) );
  AND2_X2 U13012 ( .A1(n12016), .A2(n12015), .ZN(n12024) );
  INV_X1 U13013 ( .A(n12202), .ZN(n12203) );
  NOR2_X2 U13014 ( .A1(n17262), .A2(n17182), .ZN(n11617) );
  AND2_X2 U13015 ( .A1(n17305), .A2(n11622), .ZN(n17273) );
  OR2_X1 U13016 ( .A1(n16905), .A2(n11643), .ZN(n11640) );
  INV_X1 U13017 ( .A(n13051), .ZN(n13053) );
  NOR2_X2 U13018 ( .A1(n14339), .A2(n11646), .ZN(n14377) );
  INV_X2 U13019 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21618) );
  NAND2_X1 U13020 ( .A1(n18748), .A2(n18747), .ZN(n18868) );
  NOR2_X1 U13021 ( .A1(n18942), .A2(n18944), .ZN(n18908) );
  NAND3_X1 U13022 ( .A1(n11649), .A2(n21952), .A3(n21946), .ZN(n18902) );
  INV_X1 U13023 ( .A(n11655), .ZN(n19086) );
  INV_X1 U13024 ( .A(n18699), .ZN(n11654) );
  NAND2_X1 U13025 ( .A1(n11306), .A2(n19122), .ZN(n11656) );
  NAND3_X1 U13026 ( .A1(n11658), .A2(n11272), .A3(n11306), .ZN(n11657) );
  INV_X1 U13027 ( .A(n11658), .ZN(n19132) );
  XNOR2_X1 U13028 ( .A(n14021), .B(n14019), .ZN(n17266) );
  OAI21_X2 U13029 ( .B1(n17286), .B2(n11665), .A(n11349), .ZN(n14021) );
  AND2_X2 U13030 ( .A1(n15251), .A2(n11342), .ZN(n15632) );
  AND3_X4 U13031 ( .A1(n12054), .A2(n12833), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n12192) );
  AND2_X2 U13032 ( .A1(n12058), .A2(n12063), .ZN(n12159) );
  OAI21_X1 U13033 ( .B1(n17551), .B2(n11686), .A(n11684), .ZN(n11683) );
  OAI21_X1 U13034 ( .B1(n14786), .B2(n15016), .A(n14772), .ZN(n12930) );
  NAND2_X2 U13035 ( .A1(n12909), .A2(n11297), .ZN(n14786) );
  NAND2_X1 U13036 ( .A1(n13301), .A2(n13300), .ZN(n11693) );
  NAND2_X1 U13037 ( .A1(n11693), .A2(n11695), .ZN(n14911) );
  INV_X1 U13038 ( .A(n14911), .ZN(n11694) );
  NAND2_X1 U13039 ( .A1(n11694), .A2(n13319), .ZN(n14913) );
  INV_X1 U13040 ( .A(n15937), .ZN(n11699) );
  AND3_X2 U13041 ( .A1(n13360), .A2(n13361), .A3(n11287), .ZN(n15909) );
  NAND2_X1 U13042 ( .A1(n13360), .A2(n13361), .ZN(n15584) );
  INV_X1 U13043 ( .A(n15756), .ZN(n11706) );
  NOR2_X1 U13044 ( .A1(n16537), .A2(n11707), .ZN(n16517) );
  INV_X1 U13045 ( .A(n16041), .ZN(n12445) );
  INV_X1 U13046 ( .A(n15800), .ZN(n15882) );
  NAND2_X1 U13047 ( .A1(n19551), .A2(n12488), .ZN(n12575) );
  AND2_X1 U13048 ( .A1(n20322), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12692) );
  AND2_X1 U13049 ( .A1(n20322), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12667) );
  AND2_X1 U13050 ( .A1(n20322), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12662) );
  AND2_X1 U13051 ( .A1(n20322), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12652) );
  NAND2_X1 U13052 ( .A1(n17257), .A2(n14047), .ZN(n14090) );
  NAND2_X1 U13053 ( .A1(n14116), .A2(n14115), .ZN(n14157) );
  INV_X1 U13054 ( .A(n16037), .ZN(n16046) );
  AND2_X1 U13055 ( .A1(n20322), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12688) );
  AND2_X1 U13056 ( .A1(n20322), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12670) );
  NOR2_X1 U13057 ( .A1(n11261), .A2(n12483), .ZN(n12574) );
  NOR2_X2 U13058 ( .A1(n17459), .A2(n16034), .ZN(n17425) );
  AOI21_X2 U13059 ( .B1(n17556), .B2(n12682), .A(n12681), .ZN(n17551) );
  INV_X1 U13060 ( .A(n15963), .ZN(n17556) );
  NOR2_X1 U13061 ( .A1(n14699), .A2(n14674), .ZN(n18031) );
  NOR2_X1 U13062 ( .A1(n17266), .A2(n17268), .ZN(n17267) );
  AND2_X1 U13063 ( .A1(n11260), .A2(n19515), .ZN(n12496) );
  AND2_X1 U13064 ( .A1(n11261), .A2(n12481), .ZN(n12501) );
  OR2_X1 U13065 ( .A1(n19583), .A2(n19264), .ZN(n18065) );
  INV_X1 U13066 ( .A(n12219), .ZN(n13913) );
  OR2_X1 U13067 ( .A1(n17008), .A2(n22375), .ZN(n11712) );
  OR2_X1 U13068 ( .A1(n16534), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n11713) );
  AND2_X1 U13069 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n22464), .ZN(n22421) );
  AND2_X1 U13070 ( .A1(n13994), .A2(n19264), .ZN(n11714) );
  AND2_X1 U13071 ( .A1(n12038), .A2(n12046), .ZN(n11715) );
  NOR2_X1 U13072 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18577), .ZN(n22057) );
  AND2_X1 U13073 ( .A1(n11793), .A2(n11792), .ZN(n11716) );
  INV_X1 U13074 ( .A(n13404), .ZN(n13477) );
  NAND2_X1 U13075 ( .A1(n22556), .A2(n22393), .ZN(n22609) );
  INV_X1 U13076 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19509) );
  AND2_X1 U13077 ( .A1(n18572), .A2(n21533), .ZN(n18569) );
  INV_X2 U13078 ( .A(n18569), .ZN(n18565) );
  INV_X1 U13079 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18945) );
  OR2_X1 U13080 ( .A1(n14550), .A2(n14607), .ZN(n14615) );
  OR2_X1 U13081 ( .A1(n21619), .A2(n19143), .ZN(n20955) );
  OR2_X1 U13082 ( .A1(n15956), .A2(n15970), .ZN(n11718) );
  AND2_X1 U13083 ( .A1(n15962), .A2(n15961), .ZN(n11719) );
  INV_X1 U13084 ( .A(n16052), .ZN(n16050) );
  NAND2_X1 U13085 ( .A1(n18850), .A2(n19144), .ZN(n18937) );
  INV_X1 U13086 ( .A(n18937), .ZN(n18917) );
  INV_X1 U13087 ( .A(n19477), .ZN(n12449) );
  OR2_X1 U13088 ( .A1(n13830), .A2(n19509), .ZN(n11720) );
  INV_X1 U13089 ( .A(n20828), .ZN(n20825) );
  INV_X1 U13090 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22567) );
  AND4_X1 U13091 ( .A1(n12935), .A2(n12934), .A3(n12933), .A4(n12932), .ZN(
        n11721) );
  AND3_X1 U13092 ( .A1(n12897), .A2(n12896), .A3(n12895), .ZN(n11722) );
  AND2_X2 U13093 ( .A1(n14660), .A2(n12885), .ZN(n13028) );
  AND4_X1 U13094 ( .A1(n12974), .A2(n12973), .A3(n12972), .A4(n12971), .ZN(
        n11723) );
  AND4_X1 U13095 ( .A1(n12939), .A2(n12938), .A3(n12937), .A4(n12936), .ZN(
        n11724) );
  AND2_X1 U13096 ( .A1(n14770), .A2(n14784), .ZN(n13243) );
  INV_X1 U13097 ( .A(n13243), .ZN(n13258) );
  AND3_X1 U13098 ( .A1(n12516), .A2(n12515), .A3(n12514), .ZN(n11725) );
  NAND2_X1 U13099 ( .A1(n12574), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12523) );
  AND2_X1 U13100 ( .A1(n13288), .A2(n14193), .ZN(n13277) );
  INV_X1 U13101 ( .A(n13091), .ZN(n13768) );
  INV_X1 U13102 ( .A(n13216), .ZN(n13046) );
  NAND2_X1 U13103 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11950) );
  OR2_X1 U13104 ( .A1(n13252), .A2(n13259), .ZN(n13254) );
  INV_X1 U13105 ( .A(n13175), .ZN(n13111) );
  AND2_X1 U13106 ( .A1(n13050), .A2(n13216), .ZN(n13135) );
  OR2_X1 U13107 ( .A1(n13110), .A2(n13109), .ZN(n13186) );
  NAND2_X1 U13108 ( .A1(n14046), .A2(n11350), .ZN(n14047) );
  INV_X1 U13109 ( .A(n12608), .ZN(n12609) );
  AND4_X1 U13110 ( .A1(n12528), .A2(n12527), .A3(n12526), .A4(n12525), .ZN(
        n12531) );
  AND2_X1 U13111 ( .A1(n11993), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12000) );
  AND2_X1 U13112 ( .A1(n13254), .A2(n13253), .ZN(n14195) );
  NOR2_X1 U13113 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13245), .ZN(
        n13251) );
  INV_X1 U13114 ( .A(n16733), .ZN(n13485) );
  OR2_X1 U13115 ( .A1(n13133), .A2(n13132), .ZN(n13208) );
  OR2_X1 U13116 ( .A1(n13122), .A2(n13121), .ZN(n13189) );
  AOI22_X1 U13117 ( .A1(n13069), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12966), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12923) );
  INV_X1 U13118 ( .A(n14022), .ZN(n14019) );
  AND2_X1 U13119 ( .A1(n12632), .A2(n12631), .ZN(n12798) );
  NAND2_X1 U13120 ( .A1(n12013), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13830) );
  NAND2_X1 U13121 ( .A1(n14771), .A2(n11243), .ZN(n13068) );
  INV_X1 U13122 ( .A(n14286), .ZN(n14292) );
  AND2_X1 U13123 ( .A1(n16843), .A2(n13782), .ZN(n13783) );
  NOR2_X1 U13124 ( .A1(n13647), .A2(n16890), .ZN(n13648) );
  INV_X1 U13125 ( .A(n13345), .ZN(n13306) );
  NOR2_X1 U13126 ( .A1(n13136), .A2(n13258), .ZN(n13137) );
  INV_X1 U13127 ( .A(n14780), .ZN(n12978) );
  OR2_X1 U13128 ( .A1(n14674), .A2(n12982), .ZN(n12965) );
  INV_X1 U13129 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U13130 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11834) );
  INV_X1 U13131 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U13132 ( .A1(n13830), .A2(n20162), .ZN(n13820) );
  AND2_X1 U13133 ( .A1(n18866), .A2(n21960), .ZN(n18867) );
  AND2_X1 U13134 ( .A1(n18770), .A2(n18740), .ZN(n18741) );
  OR2_X1 U13135 ( .A1(n13791), .A2(n16845), .ZN(n13793) );
  AND2_X1 U13136 ( .A1(n16551), .A2(n13782), .ZN(n13684) );
  INV_X1 U13137 ( .A(n13306), .ZN(n13781) );
  NOR2_X1 U13138 ( .A1(n13486), .A2(n22336), .ZN(n13504) );
  NAND2_X1 U13139 ( .A1(n13450), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13468) );
  OR2_X1 U13140 ( .A1(n13097), .A2(n13096), .ZN(n13170) );
  NAND2_X1 U13141 ( .A1(n12979), .A2(n12978), .ZN(n14806) );
  NAND2_X1 U13142 ( .A1(n13086), .A2(n13085), .ZN(n15059) );
  INV_X1 U13143 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15199) );
  INV_X1 U13144 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n22553) );
  INV_X1 U13145 ( .A(n17818), .ZN(n12415) );
  INV_X1 U13146 ( .A(n14069), .ZN(n14042) );
  NAND2_X1 U13147 ( .A1(n13829), .A2(n13828), .ZN(n14900) );
  INV_X1 U13148 ( .A(n14157), .ZN(n14117) );
  INV_X1 U13149 ( .A(n13961), .ZN(n13917) );
  NAND2_X1 U13150 ( .A1(n12098), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12084) );
  AND2_X1 U13151 ( .A1(n18096), .A2(n19574), .ZN(n15767) );
  INV_X1 U13152 ( .A(n13950), .ZN(n15294) );
  NOR2_X1 U13153 ( .A1(n21470), .A2(n18696), .ZN(n18700) );
  NAND2_X1 U13154 ( .A1(n18868), .A2(n18867), .ZN(n18871) );
  NAND2_X1 U13155 ( .A1(n18744), .A2(n18743), .ZN(n18745) );
  INV_X1 U13156 ( .A(n18791), .ZN(n19040) );
  NOR2_X1 U13157 ( .A1(n20959), .A2(n21979), .ZN(n21932) );
  AND2_X1 U13158 ( .A1(n16098), .A2(n16097), .ZN(n16106) );
  OR2_X1 U13159 ( .A1(n16590), .A2(n20777), .ZN(n16578) );
  INV_X1 U13160 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n22336) );
  INV_X1 U13161 ( .A(n22339), .ZN(n16675) );
  AND2_X1 U13162 ( .A1(n14314), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14315) );
  AND2_X1 U13163 ( .A1(n14268), .A2(n14267), .ZN(n16636) );
  NAND2_X1 U13164 ( .A1(n13689), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13726) );
  INV_X1 U13165 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16890) );
  NOR2_X1 U13166 ( .A1(n13445), .A2(n13421), .ZN(n13450) );
  AND2_X1 U13167 ( .A1(n15911), .A2(n15910), .ZN(n16661) );
  AOI21_X1 U13168 ( .B1(n13350), .B2(n13477), .A(n13349), .ZN(n15538) );
  AND2_X1 U13169 ( .A1(n14282), .A2(n14281), .ZN(n16595) );
  INV_X1 U13170 ( .A(n17102), .ZN(n22118) );
  NOR2_X1 U13171 ( .A1(n22147), .A2(n17125), .ZN(n17103) );
  OR2_X1 U13172 ( .A1(n17152), .A2(n22609), .ZN(n17157) );
  INV_X1 U13173 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14688) );
  OR2_X1 U13174 ( .A1(n11254), .A2(n15044), .ZN(n15198) );
  NOR2_X1 U13175 ( .A1(n22632), .A2(n15435), .ZN(n22622) );
  AND2_X1 U13176 ( .A1(n15060), .A2(n13058), .ZN(n15399) );
  NOR2_X1 U13177 ( .A1(n22613), .A2(n15435), .ZN(n22639) );
  INV_X1 U13178 ( .A(n22748), .ZN(n22743) );
  INV_X1 U13179 ( .A(n22572), .ZN(n15205) );
  INV_X1 U13180 ( .A(n22434), .ZN(n18044) );
  NAND2_X1 U13181 ( .A1(n11928), .A2(n15978), .ZN(n15983) );
  INV_X1 U13182 ( .A(n17399), .ZN(n12424) );
  NOR2_X1 U13183 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U13184 ( .A1(n14042), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13825) );
  NAND2_X1 U13185 ( .A1(n13801), .A2(n13802), .ZN(n14069) );
  AND2_X1 U13186 ( .A1(n11589), .A2(n12045), .ZN(n14548) );
  INV_X1 U13187 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n19313) );
  OR2_X1 U13188 ( .A1(n19496), .A2(n19542), .ZN(n16045) );
  AND2_X1 U13189 ( .A1(n12434), .A2(n12433), .ZN(n17351) );
  INV_X1 U13190 ( .A(n15967), .ZN(n12707) );
  OR2_X1 U13191 ( .A1(n19347), .A2(n12686), .ZN(n17536) );
  AND3_X1 U13192 ( .A1(n12414), .A2(n12413), .A3(n12412), .ZN(n17818) );
  AND3_X1 U13193 ( .A1(n12312), .A2(n12311), .A3(n12310), .ZN(n17223) );
  NAND2_X1 U13194 ( .A1(n12771), .A2(n19570), .ZN(n12823) );
  NOR2_X2 U13195 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20222) );
  AND2_X1 U13196 ( .A1(n20257), .A2(n20222), .ZN(n20184) );
  AND2_X1 U13197 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20219) );
  OR2_X1 U13198 ( .A1(n20183), .A2(n20254), .ZN(n20233) );
  OR2_X1 U13199 ( .A1(n20132), .A2(n18109), .ZN(n20150) );
  INV_X1 U13200 ( .A(n13824), .ZN(n15765) );
  NOR2_X1 U13201 ( .A1(n21428), .A2(n20959), .ZN(n14485) );
  NOR2_X1 U13202 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n21262), .ZN(n21276) );
  NOR2_X1 U13203 ( .A1(n21224), .A2(n21226), .ZN(n21261) );
  NOR2_X1 U13204 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n21183), .ZN(n21199) );
  NOR2_X1 U13205 ( .A1(n21781), .A2(n21141), .ZN(n21170) );
  NOR2_X1 U13206 ( .A1(n19951), .A2(n20954), .ZN(n14453) );
  NOR2_X1 U13207 ( .A1(n18574), .A2(n14500), .ZN(n14455) );
  AOI211_X1 U13208 ( .C1(n11164), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n14390), .B(n14389), .ZN(n14391) );
  NOR4_X1 U13209 ( .A1(n21599), .A2(n21493), .A3(n21597), .A4(n21585), .ZN(
        n21494) );
  AOI211_X1 U13210 ( .C1(n11163), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n18623), .B(n18622), .ZN(n18624) );
  OAI21_X1 U13211 ( .B1(n14485), .B2(n20967), .A(n18573), .ZN(n14449) );
  INV_X1 U13212 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18835) );
  INV_X1 U13213 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21078) );
  NAND2_X1 U13214 ( .A1(n18871), .A2(n18870), .ZN(n18872) );
  OR2_X1 U13215 ( .A1(n22015), .A2(n21659), .ZN(n21660) );
  XNOR2_X1 U13216 ( .A(n18703), .B(n18767), .ZN(n19067) );
  NOR2_X1 U13217 ( .A1(n14359), .A2(n14358), .ZN(n19951) );
  INV_X1 U13218 ( .A(n19687), .ZN(n19670) );
  NAND2_X1 U13219 ( .A1(n14200), .A2(n14199), .ZN(n22104) );
  OR2_X1 U13220 ( .A1(n16541), .A2(n20787), .ZN(n16534) );
  NAND2_X1 U13221 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n13407), .ZN(
        n13445) );
  AND2_X1 U13222 ( .A1(n22255), .A2(n14205), .ZN(n22362) );
  NOR2_X1 U13223 ( .A1(n14313), .A2(n14311), .ZN(n22248) );
  AND2_X1 U13224 ( .A1(n16834), .A2(n16741), .ZN(n16742) );
  INV_X1 U13225 ( .A(n14809), .ZN(n18045) );
  INV_X1 U13226 ( .A(n22480), .ZN(n22521) );
  NAND2_X1 U13227 ( .A1(n13570), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13601) );
  NOR2_X1 U13228 ( .A1(n13569), .A2(n16919), .ZN(n13570) );
  INV_X1 U13229 ( .A(n20853), .ZN(n20873) );
  INV_X1 U13230 ( .A(n20842), .ZN(n20870) );
  INV_X1 U13231 ( .A(n22129), .ZN(n22202) );
  OR2_X1 U13232 ( .A1(n22188), .A2(n22123), .ZN(n22147) );
  INV_X1 U13233 ( .A(n22218), .ZN(n22200) );
  OAI211_X1 U13234 ( .C1(n17151), .C2(n15207), .A(n15206), .B(n15205), .ZN(
        n22545) );
  NAND2_X1 U13235 ( .A1(n15196), .A2(n13301), .ZN(n22562) );
  OAI21_X1 U13236 ( .B1(n22576), .B2(n22575), .A(n22574), .ZN(n22791) );
  NOR2_X2 U13237 ( .A1(n22562), .A2(n15392), .ZN(n22790) );
  AND2_X1 U13238 ( .A1(n15120), .A2(n15147), .ZN(n22802) );
  INV_X1 U13239 ( .A(n22602), .ZN(n22605) );
  INV_X1 U13240 ( .A(n22814), .ZN(n15469) );
  INV_X1 U13241 ( .A(n22830), .ZN(n22766) );
  OAI21_X1 U13242 ( .B1(n15039), .B2(n15040), .A(n15205), .ZN(n22827) );
  NOR2_X1 U13243 ( .A1(n15187), .A2(n15016), .ZN(n22748) );
  NOR2_X1 U13244 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14985), .ZN(n15397) );
  NOR2_X1 U13245 ( .A1(n15187), .A2(n13044), .ZN(n22652) );
  INV_X1 U13246 ( .A(n22650), .ZN(n22656) );
  INV_X1 U13247 ( .A(n22704), .ZN(n22709) );
  AND2_X1 U13248 ( .A1(n15149), .A2(n15057), .ZN(n22846) );
  NAND2_X1 U13249 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n22424) );
  AND2_X1 U13250 ( .A1(n22422), .A2(n12977), .ZN(n14305) );
  INV_X1 U13251 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n22433) );
  INV_X1 U13252 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n22437) );
  OR2_X1 U13253 ( .A1(n12738), .A2(n12736), .ZN(n15764) );
  OAI21_X1 U13254 ( .B1(n19440), .B2(n19441), .A(n11253), .ZN(n19456) );
  NOR2_X1 U13255 ( .A1(n19379), .A2(n19380), .ZN(n19400) );
  INV_X1 U13256 ( .A(n19462), .ZN(n19495) );
  OR2_X1 U13257 ( .A1(n19480), .A2(n15680), .ZN(n14154) );
  NAND2_X1 U13258 ( .A1(n15800), .A2(n12153), .ZN(n15903) );
  OR2_X1 U13259 ( .A1(n19479), .A2(n20548), .ZN(n14144) );
  AND2_X1 U13260 ( .A1(n15614), .A2(n15777), .ZN(n20050) );
  INV_X1 U13261 ( .A(n20081), .ZN(n20313) );
  AND2_X1 U13262 ( .A1(n17292), .A2(n17291), .ZN(n19404) );
  INV_X1 U13263 ( .A(n12823), .ZN(n12860) );
  INV_X1 U13264 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19512) );
  OAI21_X2 U13265 ( .B1(n17961), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15766), 
        .ZN(n20257) );
  NAND2_X1 U13266 ( .A1(n15764), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17961) );
  INV_X1 U13267 ( .A(n20257), .ZN(n20558) );
  OAI21_X1 U13268 ( .B1(n20236), .B2(n20235), .A(n20237), .ZN(n20648) );
  INV_X1 U13269 ( .A(n20639), .ZN(n20641) );
  OAI21_X1 U13270 ( .B1(n20215), .B2(n20214), .A(n20213), .ZN(n20635) );
  OAI21_X1 U13271 ( .B1(n20200), .B2(n20199), .A(n20198), .ZN(n20628) );
  AND2_X1 U13272 ( .A1(n20192), .A2(n20232), .ZN(n20627) );
  AND2_X1 U13273 ( .A1(n20132), .A2(n18109), .ZN(n20192) );
  INV_X1 U13274 ( .A(n20519), .ZN(n20608) );
  INV_X1 U13275 ( .A(n20606), .ZN(n20595) );
  OAI21_X1 U13276 ( .B1(n20125), .B2(n20124), .A(n20123), .ZN(n20584) );
  INV_X1 U13277 ( .A(n20150), .ZN(n20149) );
  INV_X1 U13278 ( .A(n20535), .ZN(n20540) );
  AND2_X1 U13279 ( .A1(n20108), .A2(n20554), .ZN(n20232) );
  INV_X1 U13280 ( .A(n20440), .ZN(n20442) );
  INV_X1 U13281 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17995) );
  NAND2_X1 U13282 ( .A1(n22097), .A2(n14494), .ZN(n18574) );
  NOR2_X1 U13283 ( .A1(n21419), .A2(n21356), .ZN(n21395) );
  NOR2_X1 U13284 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n21238), .ZN(n21257) );
  NOR2_X1 U13285 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n21158), .ZN(n21178) );
  AND2_X1 U13286 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n21033), .ZN(n21064) );
  NAND2_X1 U13287 ( .A1(n14534), .A2(n14453), .ZN(n21327) );
  AND2_X1 U13288 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18520), .ZN(n18446) );
  NOR2_X1 U13289 ( .A1(n21240), .A2(n18533), .ZN(n18547) );
  INV_X1 U13290 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n21117) );
  INV_X1 U13291 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n21068) );
  INV_X1 U13292 ( .A(n21552), .ZN(n21548) );
  NAND2_X1 U13293 ( .A1(n21534), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n21539) );
  NOR2_X1 U13294 ( .A1(n21496), .A2(n21495), .ZN(n21522) );
  NAND2_X1 U13295 ( .A1(n21590), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21581) );
  INV_X1 U13296 ( .A(n19951), .ZN(n21428) );
  INV_X1 U13297 ( .A(n14449), .ZN(n17988) );
  NOR2_X1 U13298 ( .A1(n21008), .A2(n20976), .ZN(n20987) );
  INV_X1 U13299 ( .A(n21022), .ZN(n20976) );
  AOI22_X1 U13300 ( .A1(n21766), .A2(n19000), .B1(n19072), .B2(n21769), .ZN(
        n19031) );
  NOR2_X2 U13301 ( .A1(n21661), .A2(n19147), .ZN(n19054) );
  OAI21_X1 U13302 ( .B1(n18735), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n22101), 
        .ZN(n19144) );
  INV_X1 U13303 ( .A(n19863), .ZN(n19948) );
  NAND2_X1 U13304 ( .A1(n21935), .A2(n18702), .ZN(n19019) );
  INV_X1 U13305 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n22039) );
  NOR2_X1 U13306 ( .A1(n19013), .A2(n21797), .ZN(n21783) );
  INV_X1 U13307 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21797) );
  NOR2_X2 U13308 ( .A1(n21661), .A2(n21707), .ZN(n22079) );
  NAND2_X2 U13309 ( .A1(n11250), .A2(n21894), .ZN(n21979) );
  INV_X1 U13310 ( .A(n22049), .ZN(n21869) );
  NOR2_X1 U13311 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19631), .ZN(
        n19639) );
  NOR2_X1 U13312 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n22084), .ZN(
        n22087) );
  CLKBUF_X1 U13313 ( .A(n19918), .Z(n20002) );
  CLKBUF_X1 U13314 ( .A(n19617), .Z(n20031) );
  INV_X1 U13315 ( .A(n19937), .ZN(n19939) );
  INV_X1 U13316 ( .A(n19778), .ZN(n19769) );
  INV_X1 U13317 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22464) );
  INV_X1 U13318 ( .A(n15777), .ZN(n15776) );
  AND2_X1 U13319 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22422), .ZN(n18059) );
  INV_X1 U13320 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22405) );
  INV_X1 U13321 ( .A(n22362), .ZN(n22377) );
  INV_X1 U13322 ( .A(n22327), .ZN(n22375) );
  NAND2_X1 U13323 ( .A1(n20833), .A2(n16741), .ZN(n20828) );
  NAND2_X1 U13324 ( .A1(n16740), .A2(n16757), .ZN(n16823) );
  NAND2_X2 U13325 ( .A1(n22480), .A2(n14929), .ZN(n16834) );
  NAND2_X1 U13326 ( .A1(n20709), .A2(n11243), .ZN(n14958) );
  NAND2_X1 U13327 ( .A1(n14783), .A2(n18045), .ZN(n22525) );
  OR3_X1 U13328 ( .A1(n16096), .A2(n14986), .A3(n22436), .ZN(n22480) );
  INV_X1 U13329 ( .A(n20862), .ZN(n20877) );
  INV_X1 U13330 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n22291) );
  INV_X1 U13331 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n22270) );
  OR2_X1 U13332 ( .A1(n18054), .A2(n22609), .ZN(n20853) );
  INV_X1 U13333 ( .A(n22190), .ZN(n22129) );
  OR2_X1 U13334 ( .A1(n14811), .A2(n14798), .ZN(n22218) );
  INV_X1 U13335 ( .A(n17155), .ZN(n18057) );
  INV_X1 U13336 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18038) );
  AOI22_X1 U13337 ( .A1(n22533), .A2(n22538), .B1(n22532), .B2(n22613), .ZN(
        n22780) );
  INV_X1 U13338 ( .A(n22776), .ZN(n15245) );
  AOI22_X1 U13339 ( .A1(n22551), .A2(n22558), .B1(n22613), .B2(n22586), .ZN(
        n22787) );
  AOI22_X1 U13340 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22570), .B1(n22571), 
        .B2(n22575), .ZN(n22794) );
  INV_X1 U13341 ( .A(n22581), .ZN(n15431) );
  NAND2_X1 U13342 ( .A1(n15120), .A2(n15148), .ZN(n22800) );
  AOI22_X1 U13343 ( .A1(n22587), .A2(n22592), .B1(n22632), .B2(n22586), .ZN(
        n22807) );
  INV_X1 U13344 ( .A(n22803), .ZN(n15250) );
  INV_X1 U13345 ( .A(n22606), .ZN(n15472) );
  INV_X1 U13346 ( .A(n22819), .ZN(n15240) );
  AOI22_X1 U13347 ( .A1(n22615), .A2(n22623), .B1(n22614), .B2(n22613), .ZN(
        n22823) );
  AND2_X1 U13348 ( .A1(n15006), .A2(n15005), .ZN(n22704) );
  NAND2_X1 U13349 ( .A1(n15045), .A2(n15038), .ZN(n22830) );
  AOI22_X1 U13350 ( .A1(n22633), .A2(n22640), .B1(n22632), .B2(n22631), .ZN(
        n22839) );
  INV_X1 U13351 ( .A(n22657), .ZN(n15536) );
  NAND2_X1 U13352 ( .A1(n15149), .A2(n15038), .ZN(n22850) );
  NAND2_X1 U13353 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n22391) );
  NOR2_X1 U13354 ( .A1(n18059), .A2(n22855), .ZN(n22408) );
  INV_X1 U13355 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20738) );
  CLKBUF_X1 U13356 ( .A(n20794), .Z(n22430) );
  OR2_X1 U13357 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22437), .ZN(n22852) );
  INV_X1 U13358 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22410) );
  NAND2_X1 U13359 ( .A1(n12450), .A2(n12449), .ZN(n12451) );
  NAND2_X1 U13360 ( .A1(n19275), .A2(n15354), .ZN(n19477) );
  XNOR2_X1 U13361 ( .A(n14716), .B(n14715), .ZN(n20108) );
  OAI21_X1 U13362 ( .B1(n14899), .B2(n14900), .A(n14902), .ZN(n20132) );
  XNOR2_X1 U13363 ( .A(n14764), .B(n14765), .ZN(n20447) );
  NAND2_X1 U13364 ( .A1(n20546), .A2(n20087), .ZN(n20548) );
  AND2_X2 U13365 ( .A1(n14124), .A2(n19570), .ZN(n20546) );
  INV_X1 U13366 ( .A(n20551), .ZN(n20405) );
  INV_X1 U13367 ( .A(n20072), .ZN(n20557) );
  NAND2_X1 U13368 ( .A1(n18127), .A2(n14653), .ZN(n14878) );
  INV_X1 U13369 ( .A(n18127), .ZN(n18156) );
  OR2_X1 U13370 ( .A1(n15339), .A2(n14549), .ZN(n14650) );
  INV_X1 U13371 ( .A(n12880), .ZN(n12881) );
  INV_X1 U13372 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18094) );
  INV_X1 U13373 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18081) );
  AOI21_X1 U13374 ( .B1(n16071), .B2(n19537), .A(n16070), .ZN(n16072) );
  INV_X1 U13375 ( .A(n12865), .ZN(n12866) );
  INV_X1 U13376 ( .A(n19537), .ZN(n17944) );
  NOR2_X1 U13377 ( .A1(n19539), .A2(n17919), .ZN(n19521) );
  INV_X1 U13378 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17998) );
  INV_X1 U13379 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20494) );
  INV_X1 U13380 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20311) );
  NAND2_X1 U13381 ( .A1(n20249), .A2(n20232), .ZN(n20659) );
  INV_X1 U13382 ( .A(n20649), .ZN(n20646) );
  NAND2_X1 U13383 ( .A1(n20249), .A2(n20203), .ZN(n20639) );
  NAND2_X1 U13384 ( .A1(n20192), .A2(n20191), .ZN(n20632) );
  INV_X1 U13385 ( .A(n20627), .ZN(n20528) );
  NAND2_X1 U13386 ( .A1(n20192), .A2(n20218), .ZN(n20625) );
  NAND2_X1 U13387 ( .A1(n20203), .A2(n20192), .ZN(n20619) );
  NAND2_X1 U13388 ( .A1(n20149), .A2(n20191), .ZN(n20519) );
  NAND2_X1 U13389 ( .A1(n20149), .A2(n20218), .ZN(n20600) );
  NAND2_X1 U13390 ( .A1(n20203), .A2(n20149), .ZN(n20593) );
  INV_X1 U13391 ( .A(n20357), .ZN(n20354) );
  AOI22_X1 U13392 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20563), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20564), .ZN(n20440) );
  AOI22_X1 U13393 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n20564), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n20563), .ZN(n20535) );
  NAND2_X1 U13394 ( .A1(n20114), .A2(n20218), .ZN(n20568) );
  INV_X1 U13395 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20235) );
  INV_X1 U13396 ( .A(n22413), .ZN(n18125) );
  NOR2_X1 U13397 ( .A1(n18192), .A2(n12207), .ZN(n22453) );
  INV_X1 U13398 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22414) );
  INV_X1 U13399 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21312) );
  INV_X1 U13400 ( .A(n21424), .ZN(n21359) );
  INV_X1 U13401 ( .A(n18473), .ZN(n18465) );
  NOR2_X1 U13402 ( .A1(n21331), .A2(n18479), .ZN(n18483) );
  INV_X1 U13403 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18402) );
  INV_X1 U13404 ( .A(n21579), .ZN(n21573) );
  OR2_X1 U13405 ( .A1(n21493), .A2(n21456), .ZN(n21451) );
  NOR2_X1 U13406 ( .A1(n21491), .A2(n21474), .ZN(n21468) );
  NAND2_X1 U13407 ( .A1(n19199), .A2(n21428), .ZN(n19218) );
  NAND3_X1 U13408 ( .A1(n17989), .A2(n17988), .A3(n20966), .ZN(n19198) );
  NAND2_X1 U13409 ( .A1(n21661), .A2(n19137), .ZN(n19052) );
  INV_X1 U13410 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n22028) );
  INV_X1 U13411 ( .A(n18964), .ZN(n18921) );
  INV_X1 U13412 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n22055) );
  NAND2_X1 U13413 ( .A1(n19948), .A2(n19648), .ZN(n19862) );
  INV_X1 U13414 ( .A(n19137), .ZN(n19147) );
  INV_X1 U13415 ( .A(n22049), .ZN(n22073) );
  INV_X1 U13416 ( .A(n22079), .ZN(n22044) );
  INV_X1 U13417 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21811) );
  INV_X1 U13418 ( .A(n22048), .ZN(n21947) );
  INV_X1 U13419 ( .A(n21962), .ZN(n21970) );
  INV_X1 U13420 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17987) );
  INV_X1 U13421 ( .A(n19952), .ZN(n20036) );
  INV_X1 U13422 ( .A(n20042), .ZN(n19849) );
  INV_X1 U13423 ( .A(n20032), .ZN(n20022) );
  INV_X1 U13424 ( .A(n19996), .ZN(n19989) );
  INV_X1 U13425 ( .A(n19991), .ZN(n19983) );
  INV_X1 U13426 ( .A(n19985), .ZN(n19977) );
  INV_X1 U13427 ( .A(n19979), .ZN(n19971) );
  INV_X1 U13428 ( .A(n19893), .ZN(n19902) );
  INV_X1 U13429 ( .A(n19974), .ZN(n19965) );
  INV_X1 U13430 ( .A(n19967), .ZN(n19956) );
  INV_X1 U13431 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n22095) );
  INV_X1 U13432 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n22084) );
  AND2_X1 U13433 ( .A1(n22469), .A2(n19219), .ZN(n22417) );
  INV_X1 U13434 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n21687) );
  INV_X1 U13435 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21127) );
  INV_X1 U13436 ( .A(n19254), .ZN(n19253) );
  NOR2_X1 U13437 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14335), .ZN(n19738)
         );
  INV_X1 U13438 ( .A(n20700), .ZN(n20699) );
  NAND2_X1 U13439 ( .A1(n11752), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U13440 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n11750), .ZN(
        n11757) );
  INV_X1 U13441 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n19461) );
  XNOR2_X1 U13442 ( .A(n11726), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n19500) );
  INV_X1 U13443 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11729) );
  INV_X1 U13444 ( .A(n11730), .ZN(n11731) );
  INV_X1 U13445 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17437) );
  AOI21_X1 U13446 ( .B1(n11731), .B2(n17437), .A(n11726), .ZN(n17439) );
  INV_X1 U13447 ( .A(n17439), .ZN(n19486) );
  AOI21_X1 U13448 ( .B1(n17468), .B2(n11732), .A(n11733), .ZN(n19440) );
  OAI21_X1 U13449 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n11734), .A(
        n11732), .ZN(n19431) );
  AOI21_X1 U13450 ( .B1(n11735), .B2(n19375), .A(n11736), .ZN(n19379) );
  OAI21_X1 U13451 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11355), .A(
        n11735), .ZN(n17525) );
  INV_X1 U13452 ( .A(n17525), .ZN(n19361) );
  AOI21_X1 U13453 ( .B1(n17542), .B2(n11738), .A(n11355), .ZN(n17540) );
  INV_X1 U13454 ( .A(n11739), .ZN(n11742) );
  INV_X1 U13455 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11741) );
  INV_X1 U13456 ( .A(n11738), .ZN(n11740) );
  AOI21_X1 U13457 ( .B1(n11742), .B2(n11741), .A(n11740), .ZN(n19352) );
  INV_X1 U13458 ( .A(n11743), .ZN(n11747) );
  INV_X1 U13459 ( .A(n11744), .ZN(n11762) );
  INV_X1 U13460 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11745) );
  NAND2_X1 U13461 ( .A1(n11762), .A2(n11745), .ZN(n11746) );
  NAND2_X1 U13462 ( .A1(n11747), .A2(n11746), .ZN(n19332) );
  INV_X1 U13463 ( .A(n19332), .ZN(n11763) );
  AOI21_X1 U13464 ( .B1(n11266), .B2(n19313), .A(n11748), .ZN(n19319) );
  AOI21_X1 U13465 ( .B1(n18094), .B2(n11757), .A(n11759), .ZN(n18082) );
  AOI21_X1 U13466 ( .B1(n17626), .B2(n11749), .A(n11750), .ZN(n19293) );
  AOI21_X1 U13467 ( .B1(n18081), .B2(n11751), .A(n11752), .ZN(n18072) );
  AOI21_X1 U13468 ( .B1(n18071), .B2(n11753), .A(n11754), .ZN(n18061) );
  INV_X1 U13469 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15708) );
  AOI21_X1 U13470 ( .B1(n11756), .B2(n15708), .A(n11755), .ZN(n15705) );
  AOI22_X1 U13471 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n11756), .B2(n17995), .ZN(
        n17230) );
  AOI22_X1 U13472 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17995), .ZN(n17229) );
  NAND2_X1 U13473 ( .A1(n17230), .A2(n17229), .ZN(n15703) );
  NOR2_X1 U13474 ( .A1(n15705), .A2(n15703), .ZN(n16081) );
  OAI21_X1 U13475 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11755), .A(
        n11753), .ZN(n16082) );
  NAND2_X1 U13476 ( .A1(n16081), .A2(n16082), .ZN(n15745) );
  NOR2_X1 U13477 ( .A1(n18061), .A2(n15745), .ZN(n15659) );
  OAI21_X1 U13478 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11754), .A(
        n11751), .ZN(n15827) );
  NAND2_X1 U13479 ( .A1(n15659), .A2(n15827), .ZN(n15719) );
  NOR2_X1 U13480 ( .A1(n18072), .A2(n15719), .ZN(n19278) );
  OAI21_X1 U13481 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11752), .A(
        n11749), .ZN(n19280) );
  NAND2_X1 U13482 ( .A1(n19278), .A2(n19280), .ZN(n19291) );
  NOR2_X1 U13483 ( .A1(n19293), .A2(n19291), .ZN(n17214) );
  OR2_X1 U13484 ( .A1(n11750), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U13485 ( .A1(n11758), .A2(n11757), .ZN(n17614) );
  NAND2_X1 U13486 ( .A1(n17214), .A2(n17614), .ZN(n15733) );
  NOR2_X1 U13487 ( .A1(n18082), .A2(n15733), .ZN(n19305) );
  OAI21_X1 U13488 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11759), .A(
        n11266), .ZN(n19312) );
  NAND2_X1 U13489 ( .A1(n19305), .A2(n19312), .ZN(n19304) );
  NOR2_X1 U13490 ( .A1(n19319), .A2(n19304), .ZN(n15811) );
  INV_X1 U13491 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15807) );
  INV_X1 U13492 ( .A(n11748), .ZN(n11760) );
  NAND2_X1 U13493 ( .A1(n15807), .A2(n11760), .ZN(n11761) );
  NAND2_X1 U13494 ( .A1(n11762), .A2(n11761), .ZN(n17588) );
  NAND2_X1 U13495 ( .A1(n15811), .A2(n17588), .ZN(n19325) );
  NOR2_X1 U13496 ( .A1(n11763), .A2(n19325), .ZN(n19336) );
  NOR2_X1 U13497 ( .A1(n11743), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11764) );
  NOR2_X1 U13498 ( .A1(n11739), .A2(n11764), .ZN(n19338) );
  INV_X1 U13499 ( .A(n19338), .ZN(n17566) );
  NOR2_X1 U13500 ( .A1(n19352), .A2(n19353), .ZN(n19351) );
  NOR2_X1 U13501 ( .A1(n19396), .A2(n19351), .ZN(n17204) );
  NOR2_X1 U13502 ( .A1(n17540), .A2(n17204), .ZN(n17203) );
  NOR2_X1 U13503 ( .A1(n19396), .A2(n17203), .ZN(n19360) );
  NOR2_X1 U13504 ( .A1(n19396), .A2(n19359), .ZN(n19380) );
  OR2_X1 U13505 ( .A1(n11736), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11766) );
  NAND2_X1 U13506 ( .A1(n11765), .A2(n11766), .ZN(n19397) );
  AOI21_X1 U13507 ( .B1(n19400), .B2(n19397), .A(n19396), .ZN(n17193) );
  AOI21_X1 U13508 ( .B1(n12874), .B2(n11765), .A(n11354), .ZN(n17194) );
  NAND2_X1 U13509 ( .A1(n17196), .A2(n11252), .ZN(n19411) );
  OAI21_X1 U13510 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11354), .A(
        n11767), .ZN(n19412) );
  NAND2_X1 U13511 ( .A1(n19411), .A2(n19412), .ZN(n19410) );
  NAND2_X1 U13512 ( .A1(n19410), .A2(n11252), .ZN(n19421) );
  AOI21_X1 U13513 ( .B1(n17487), .B2(n11767), .A(n11734), .ZN(n17490) );
  INV_X1 U13514 ( .A(n17490), .ZN(n19422) );
  NAND2_X1 U13515 ( .A1(n19421), .A2(n19422), .ZN(n19420) );
  NAND2_X1 U13516 ( .A1(n19420), .A2(n11253), .ZN(n19430) );
  NAND2_X1 U13517 ( .A1(n19431), .A2(n19430), .ZN(n19441) );
  INV_X1 U13518 ( .A(n11768), .ZN(n11771) );
  INV_X1 U13519 ( .A(n11733), .ZN(n11769) );
  NAND2_X1 U13520 ( .A1(n11514), .A2(n11769), .ZN(n11770) );
  NAND2_X1 U13521 ( .A1(n11771), .A2(n11770), .ZN(n19455) );
  NAND2_X1 U13522 ( .A1(n19456), .A2(n19455), .ZN(n19454) );
  NAND2_X1 U13523 ( .A1(n19454), .A2(n11253), .ZN(n17180) );
  OAI21_X1 U13524 ( .B1(n11768), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n11364), .ZN(n17446) );
  NAND2_X1 U13525 ( .A1(n17180), .A2(n17446), .ZN(n17179) );
  NAND2_X1 U13526 ( .A1(n17179), .A2(n11253), .ZN(n19472) );
  AND2_X1 U13527 ( .A1(n11364), .A2(n19461), .ZN(n11772) );
  OR2_X1 U13528 ( .A1(n11772), .A2(n11730), .ZN(n19473) );
  NAND2_X1 U13529 ( .A1(n19472), .A2(n19473), .ZN(n19471) );
  NAND2_X1 U13530 ( .A1(n19471), .A2(n11252), .ZN(n19485) );
  NAND4_X1 U13531 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n17995), .A3(n20235), 
        .A4(n22410), .ZN(n19563) );
  INV_X2 U13532 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11773) );
  AND2_X4 U13533 ( .A1(n15264), .A2(n15306), .ZN(n11995) );
  AND2_X4 U13534 ( .A1(n11781), .A2(n11237), .ZN(n11996) );
  AOI22_X1 U13535 ( .A1(n13946), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11779) );
  CLKBUF_X3 U13536 ( .A(n11985), .Z(n14160) );
  AOI22_X1 U13537 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13949), .B1(
        n13951), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11778) );
  AND2_X4 U13538 ( .A1(n15264), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11992) );
  AOI22_X1 U13539 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11777) );
  INV_X2 U13540 ( .A(n14024), .ZN(n14177) );
  AND2_X4 U13541 ( .A1(n11775), .A2(n15306), .ZN(n14163) );
  AOI22_X1 U13542 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n13961), .B1(
        n12219), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11776) );
  NAND4_X1 U13543 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11790) );
  AND2_X2 U13544 ( .A1(n11780), .A2(n13925), .ZN(n13958) );
  AOI22_X1 U13545 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11788) );
  NOR2_X1 U13546 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U13547 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U13548 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n13962), .B1(
        n13947), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11786) );
  AND2_X4 U13549 ( .A1(n15300), .A2(n11232), .ZN(n13935) );
  BUF_X1 U13550 ( .A(n13935), .Z(n11784) );
  AOI22_X1 U13551 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12228), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11785) );
  NAND4_X1 U13552 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(
        n11789) );
  NOR2_X1 U13553 ( .A1(n11790), .A2(n11789), .ZN(n12776) );
  AOI22_X1 U13554 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11255), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U13555 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U13556 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U13557 ( .A1(n11795), .A2(n11794), .A3(n11791), .A4(n11716), .ZN(
        n11803) );
  AOI22_X1 U13558 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U13559 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11800) );
  INV_X2 U13560 ( .A(n14096), .ZN(n13999) );
  AOI22_X1 U13561 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U13562 ( .A1(n11796), .A2(n15297), .ZN(n11797) );
  NOR2_X1 U13563 ( .A1(n11717), .A2(n11797), .ZN(n11798) );
  NAND4_X1 U13564 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        n11802) );
  INV_X1 U13565 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14719) );
  INV_X1 U13566 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12545) );
  NAND3_X1 U13567 ( .A1(n20322), .A2(n14719), .A3(n12545), .ZN(n11804) );
  NAND2_X1 U13568 ( .A1(n12247), .A2(n11804), .ZN(n12551) );
  AOI22_X1 U13569 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U13570 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U13571 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U13572 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11805) );
  NAND4_X1 U13573 ( .A1(n11808), .A2(n11807), .A3(n11806), .A4(n11805), .ZN(
        n11816) );
  NAND2_X1 U13574 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11810) );
  AOI22_X1 U13575 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11809) );
  AND2_X1 U13576 ( .A1(n11810), .A2(n11809), .ZN(n11814) );
  AOI22_X1 U13577 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U13578 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11812) );
  NAND2_X1 U13579 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11811) );
  NAND4_X1 U13580 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11815) );
  NOR2_X1 U13581 ( .A1(n11816), .A2(n11815), .ZN(n12778) );
  INV_X1 U13582 ( .A(n12778), .ZN(n11817) );
  INV_X1 U13583 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12089) );
  MUX2_X1 U13584 ( .A(n11817), .B(n12089), .S(n20322), .Z(n12550) );
  AOI22_X1 U13585 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U13586 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11820) );
  AOI22_X1 U13587 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U13588 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11818) );
  NAND4_X1 U13589 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11823) );
  INV_X1 U13590 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14034) );
  INV_X1 U13591 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14032) );
  OAI22_X1 U13592 ( .A1(n13919), .A2(n14034), .B1(n13917), .B2(n14032), .ZN(
        n11822) );
  NOR2_X1 U13593 ( .A1(n11823), .A2(n11822), .ZN(n11829) );
  AOI22_X1 U13594 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U13595 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11827) );
  INV_X1 U13596 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12469) );
  OAI22_X1 U13597 ( .A1(n12401), .A2(n12469), .B1(n12399), .B2(n15784), .ZN(
        n11825) );
  INV_X1 U13598 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12464) );
  INV_X1 U13599 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12335) );
  OAI22_X1 U13600 ( .A1(n12404), .A2(n12464), .B1(n15294), .B2(n12335), .ZN(
        n11824) );
  NOR2_X1 U13601 ( .A1(n11825), .A2(n11824), .ZN(n11826) );
  NAND4_X1 U13602 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n12511) );
  XNOR2_X1 U13603 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U13604 ( .A1(n12008), .A2(n12009), .ZN(n12010) );
  NAND2_X1 U13605 ( .A1(n20245), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11830) );
  NAND2_X1 U13606 ( .A1(n12010), .A2(n11830), .ZN(n12007) );
  XNOR2_X1 U13607 ( .A(n17957), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12006) );
  NAND2_X1 U13608 ( .A1(n12007), .A2(n12006), .ZN(n11832) );
  NAND2_X1 U13609 ( .A1(n20161), .A2(n17957), .ZN(n11831) );
  XNOR2_X1 U13610 ( .A(n11856), .B(n11857), .ZN(n12732) );
  AOI22_X1 U13611 ( .A1(n11248), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U13612 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11833) );
  NAND4_X1 U13613 ( .A1(n11836), .A2(n11835), .A3(n11834), .A4(n11833), .ZN(
        n11842) );
  AOI22_X1 U13614 ( .A1(n11248), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U13615 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U13616 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11837) );
  NAND4_X1 U13617 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(
        n11841) );
  AOI22_X1 U13618 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11968), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U13619 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U13620 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U13621 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11843) );
  NAND4_X1 U13622 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11847) );
  AOI22_X1 U13623 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U13624 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U13625 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11849) );
  NAND4_X1 U13626 ( .A1(n11852), .A2(n11851), .A3(n11850), .A4(n11849), .ZN(
        n11853) );
  NAND2_X1 U13627 ( .A1(n11853), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11854) );
  MUX2_X1 U13628 ( .A(n12511), .B(n12732), .S(n11245), .Z(n12717) );
  MUX2_X1 U13629 ( .A(n12717), .B(n16086), .S(n20322), .Z(n12537) );
  NAND2_X1 U13630 ( .A1(n12538), .A2(n12537), .ZN(n12557) );
  INV_X1 U13631 ( .A(n12557), .ZN(n11875) );
  NAND3_X1 U13632 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12005), .A3(
        n19509), .ZN(n12743) );
  INV_X1 U13633 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11860) );
  OAI22_X1 U13634 ( .A1(n12401), .A2(n11860), .B1(n12399), .B2(n20400), .ZN(
        n11862) );
  INV_X1 U13635 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14058) );
  INV_X1 U13636 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11861) );
  NAND2_X1 U13637 ( .A1(n12228), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11866) );
  NAND2_X1 U13638 ( .A1(n13946), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11865) );
  NAND2_X1 U13639 ( .A1(n13947), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U13640 ( .A1(n12300), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11863) );
  AOI22_X1 U13641 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U13642 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11869) );
  AOI22_X1 U13643 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11868) );
  NAND2_X1 U13644 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11867) );
  AND4_X1 U13645 ( .A1(n11870), .A2(n11869), .A3(n11868), .A4(n11867), .ZN(
        n11872) );
  AOI22_X1 U13646 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11871) );
  NAND4_X1 U13647 ( .A1(n11874), .A2(n11873), .A3(n11872), .A4(n11871), .ZN(
        n12785) );
  MUX2_X1 U13648 ( .A(n12743), .B(n12785), .S(n12721), .Z(n12718) );
  INV_X1 U13649 ( .A(n12602), .ZN(n11889) );
  AOI22_X1 U13650 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U13651 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11878) );
  INV_X1 U13652 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20360) );
  AOI22_X1 U13653 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U13654 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11876) );
  NAND4_X1 U13655 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11887) );
  NAND2_X1 U13656 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11881) );
  AOI22_X1 U13657 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11880) );
  AND2_X1 U13658 ( .A1(n11881), .A2(n11880), .ZN(n11885) );
  AOI22_X1 U13659 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U13660 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U13661 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11882) );
  NAND4_X1 U13662 ( .A1(n11885), .A2(n11884), .A3(n11883), .A4(n11882), .ZN(
        n11886) );
  NOR2_X1 U13663 ( .A1(n11887), .A2(n11886), .ZN(n12597) );
  INV_X1 U13664 ( .A(n12597), .ZN(n11888) );
  INV_X1 U13665 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12115) );
  MUX2_X1 U13666 ( .A(n11888), .B(n12115), .S(n20322), .Z(n12600) );
  NAND2_X1 U13667 ( .A1(n11889), .A2(n12600), .ZN(n12635) );
  INV_X1 U13668 ( .A(n12635), .ZN(n11903) );
  AOI22_X1 U13669 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U13670 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U13671 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U13672 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11890) );
  NAND4_X1 U13673 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n11890), .ZN(
        n11901) );
  NAND2_X1 U13674 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11895) );
  AOI22_X1 U13675 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11894) );
  AND2_X1 U13676 ( .A1(n11895), .A2(n11894), .ZN(n11899) );
  AOI22_X1 U13677 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U13678 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11897) );
  NAND2_X1 U13679 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11896) );
  NAND4_X1 U13680 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11900) );
  NOR2_X1 U13681 ( .A1(n11901), .A2(n11900), .ZN(n12630) );
  INV_X1 U13682 ( .A(n12630), .ZN(n11902) );
  INV_X1 U13683 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n15723) );
  MUX2_X1 U13684 ( .A(n11902), .B(n15723), .S(n20322), .Z(n12634) );
  AOI22_X1 U13685 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U13686 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11906) );
  AOI22_X1 U13687 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U13688 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11904) );
  NAND4_X1 U13689 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11911) );
  NAND2_X1 U13690 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11909) );
  NAND2_X1 U13691 ( .A1(n13961), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11908) );
  NAND2_X1 U13692 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  NOR2_X1 U13693 ( .A1(n11911), .A2(n11910), .ZN(n11922) );
  NAND2_X1 U13694 ( .A1(n12228), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11915) );
  NAND2_X1 U13695 ( .A1(n13946), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11914) );
  NAND2_X1 U13696 ( .A1(n13947), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11913) );
  NAND2_X1 U13697 ( .A1(n12300), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11912) );
  NAND2_X1 U13698 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11919) );
  NAND2_X1 U13699 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11918) );
  NAND2_X1 U13700 ( .A1(n13948), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U13701 ( .A1(n13950), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11916) );
  INV_X4 U13702 ( .A(n16007), .ZN(n16014) );
  INV_X1 U13703 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11923) );
  MUX2_X1 U13704 ( .A(n16014), .B(n11923), .S(n20322), .Z(n12639) );
  INV_X1 U13705 ( .A(n12639), .ZN(n11924) );
  NAND2_X1 U13706 ( .A1(n20322), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12642) );
  NAND2_X1 U13707 ( .A1(n20322), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12649) );
  OR2_X2 U13708 ( .A1(n12653), .A2(n12652), .ZN(n12660) );
  INV_X1 U13709 ( .A(n12660), .ZN(n11925) );
  NAND2_X1 U13710 ( .A1(n20322), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12659) );
  NAND2_X1 U13711 ( .A1(n11925), .A2(n12659), .ZN(n12663) );
  INV_X1 U13712 ( .A(n12663), .ZN(n11927) );
  INV_X1 U13713 ( .A(n12662), .ZN(n11926) );
  NAND2_X1 U13714 ( .A1(n11927), .A2(n11926), .ZN(n12671) );
  OR2_X2 U13715 ( .A1(n12671), .A2(n12670), .ZN(n12673) );
  NAND2_X1 U13716 ( .A1(n20322), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12683) );
  NOR2_X2 U13717 ( .A1(n11291), .A2(n12692), .ZN(n12695) );
  NAND2_X1 U13718 ( .A1(n20322), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12696) );
  NAND2_X1 U13719 ( .A1(n20322), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12703) );
  AND2_X1 U13720 ( .A1(n20322), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12710) );
  OR2_X2 U13721 ( .A1(n12711), .A2(n12710), .ZN(n15975) );
  AND2_X1 U13722 ( .A1(n20322), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15974) );
  OR2_X2 U13723 ( .A1(n15975), .A2(n15974), .ZN(n15979) );
  INV_X1 U13724 ( .A(n15979), .ZN(n11928) );
  NAND2_X1 U13725 ( .A1(n20322), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15978) );
  INV_X1 U13726 ( .A(n15983), .ZN(n11929) );
  NAND2_X1 U13727 ( .A1(n20322), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15982) );
  AND2_X1 U13728 ( .A1(n20322), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U13729 ( .A1(n20322), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15985) );
  NAND2_X1 U13730 ( .A1(n20322), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15992) );
  INV_X1 U13731 ( .A(n15997), .ZN(n11930) );
  NAND2_X1 U13732 ( .A1(n20322), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15996) );
  NAND2_X1 U13733 ( .A1(n20322), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16005) );
  NAND2_X1 U13734 ( .A1(n16006), .A2(n16005), .ZN(n16011) );
  NAND2_X1 U13735 ( .A1(n20322), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11931) );
  XNOR2_X1 U13736 ( .A(n16011), .B(n11931), .ZN(n16009) );
  AOI22_X1 U13737 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U13738 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U13739 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11932) );
  NAND4_X1 U13740 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11941) );
  AOI22_X1 U13741 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U13742 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U13743 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11937) );
  NAND4_X1 U13744 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11940) );
  AOI22_X1 U13745 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U13746 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U13747 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U13748 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11942) );
  NAND4_X1 U13749 ( .A1(n11945), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11946) );
  NAND2_X1 U13750 ( .A1(n11946), .A2(n15297), .ZN(n11955) );
  AOI22_X1 U13751 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U13752 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11948) );
  NAND3_X1 U13753 ( .A1(n11949), .A2(n11948), .A3(n11947), .ZN(n11953) );
  AOI22_X1 U13754 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U13755 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U13756 ( .A1(n11248), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U13757 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U13758 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  NAND2_X1 U13759 ( .A1(n11960), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11967) );
  AOI22_X1 U13760 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U13761 ( .A1(n11248), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11961) );
  NAND4_X1 U13762 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n11965) );
  NAND2_X1 U13763 ( .A1(n11965), .A2(n15297), .ZN(n11966) );
  NAND2_X2 U13764 ( .A1(n11967), .A2(n11966), .ZN(n12017) );
  AOI22_X1 U13765 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11968), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U13766 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U13767 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U13768 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U13769 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11973) );
  NAND2_X1 U13770 ( .A1(n11973), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11981) );
  AOI22_X1 U13771 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11978) );
  AOI21_X1 U13772 ( .B1(n11992), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n11974), .ZN(n11977) );
  AOI22_X1 U13773 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11255), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U13774 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U13775 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  NAND2_X1 U13776 ( .A1(n11979), .A2(n15297), .ZN(n11980) );
  AND2_X2 U13777 ( .A1(n11983), .A2(n11982), .ZN(n12040) );
  AOI22_X1 U13778 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U13779 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U13780 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14163), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U13781 ( .A1(n13935), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11995), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U13782 ( .A1(n13999), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11997) );
  NAND4_X1 U13783 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12001) );
  NAND2_X2 U13784 ( .A1(n12002), .A2(n12001), .ZN(n13800) );
  NAND2_X1 U13785 ( .A1(n13800), .A2(n12018), .ZN(n12031) );
  NAND2_X1 U13786 ( .A1(n12058), .A2(n12045), .ZN(n12857) );
  INV_X1 U13787 ( .A(n12857), .ZN(n12012) );
  NOR2_X1 U13788 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17998), .ZN(
        n12004) );
  XNOR2_X1 U13789 ( .A(n12007), .B(n12006), .ZN(n12727) );
  INV_X1 U13790 ( .A(n12727), .ZN(n12719) );
  AND2_X1 U13791 ( .A1(n12732), .A2(n12719), .ZN(n12742) );
  INV_X1 U13792 ( .A(n12008), .ZN(n12722) );
  INV_X1 U13793 ( .A(n12009), .ZN(n12543) );
  NAND2_X1 U13794 ( .A1(n12722), .A2(n12543), .ZN(n12757) );
  AND2_X1 U13795 ( .A1(n12757), .A2(n12010), .ZN(n12724) );
  AND3_X1 U13796 ( .A1(n12743), .A2(n12742), .A3(n12724), .ZN(n12011) );
  INV_X1 U13797 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17948) );
  INV_X1 U13798 ( .A(n19570), .ZN(n19580) );
  NAND2_X1 U13799 ( .A1(n12012), .A2(n12021), .ZN(n14547) );
  INV_X1 U13800 ( .A(n13800), .ZN(n12013) );
  NAND2_X2 U13801 ( .A1(n11241), .A2(n12017), .ZN(n12033) );
  NAND2_X1 U13802 ( .A1(n12027), .A2(n12033), .ZN(n12016) );
  NAND2_X1 U13803 ( .A1(n12030), .A2(n15778), .ZN(n12015) );
  INV_X1 U13804 ( .A(n12026), .ZN(n15342) );
  INV_X1 U13805 ( .A(n12019), .ZN(n12020) );
  NAND2_X1 U13806 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n22445) );
  INV_X1 U13807 ( .A(n22445), .ZN(n19566) );
  NOR2_X1 U13808 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19566), .ZN(n12208) );
  INV_X1 U13809 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n17243) );
  NOR2_X1 U13810 ( .A1(n12208), .A2(n17243), .ZN(n12022) );
  AND2_X1 U13811 ( .A1(n12721), .A2(n12022), .ZN(n12023) );
  NAND2_X1 U13812 ( .A1(n19275), .A2(n12023), .ZN(n19393) );
  INV_X1 U13813 ( .A(n13800), .ZN(n12047) );
  NAND2_X1 U13814 ( .A1(n12047), .A2(n12218), .ZN(n12038) );
  NAND2_X1 U13815 ( .A1(n12024), .A2(n11715), .ZN(n12025) );
  NOR2_X1 U13816 ( .A1(n11242), .A2(n12218), .ZN(n12028) );
  NAND2_X1 U13817 ( .A1(n12038), .A2(n12031), .ZN(n12749) );
  NAND2_X1 U13818 ( .A1(n12749), .A2(n11242), .ZN(n12748) );
  NAND2_X1 U13819 ( .A1(n12748), .A2(n12033), .ZN(n12034) );
  NAND2_X1 U13820 ( .A1(n12034), .A2(n12825), .ZN(n12035) );
  NAND2_X1 U13821 ( .A1(n12035), .A2(n15778), .ZN(n12037) );
  INV_X1 U13822 ( .A(n12038), .ZN(n12039) );
  NAND3_X1 U13823 ( .A1(n12773), .A2(n12046), .A3(n11259), .ZN(n12043) );
  AND2_X2 U13824 ( .A1(n12043), .A2(n12042), .ZN(n12855) );
  NAND2_X1 U13826 ( .A1(n12062), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12052) );
  NAND4_X1 U13827 ( .A1(n12832), .A2(n20322), .A3(n11242), .A4(n12047), .ZN(
        n12048) );
  AND2_X2 U13828 ( .A1(n12049), .A2(n12048), .ZN(n12060) );
  NAND2_X1 U13829 ( .A1(n12060), .A2(n12857), .ZN(n12816) );
  INV_X1 U13830 ( .A(n12033), .ZN(n12055) );
  NAND2_X1 U13831 ( .A1(n12058), .A2(n14548), .ZN(n12059) );
  INV_X1 U13833 ( .A(n12063), .ZN(n12065) );
  NOR2_X1 U13834 ( .A1(n12065), .A2(n12064), .ZN(n12066) );
  INV_X1 U13835 ( .A(n15261), .ZN(n12069) );
  INV_X1 U13836 ( .A(n12212), .ZN(n19556) );
  NOR2_X1 U13837 ( .A1(n19556), .A2(n20247), .ZN(n12068) );
  AOI21_X1 U13838 ( .B1(n12069), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12068), 
        .ZN(n12070) );
  NAND2_X1 U13839 ( .A1(n12071), .A2(n12070), .ZN(n12455) );
  NAND2_X1 U13840 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12072) );
  NAND2_X1 U13841 ( .A1(n19556), .A2(n12072), .ZN(n12073) );
  AOI21_X1 U13842 ( .B1(n12159), .B2(P2_REIP_REG_0__SCAN_IN), .A(n12073), .ZN(
        n12074) );
  INV_X1 U13843 ( .A(n12074), .ZN(n12083) );
  INV_X1 U13844 ( .A(n12192), .ZN(n12081) );
  NAND2_X1 U13845 ( .A1(n12076), .A2(n12075), .ZN(n12838) );
  NAND2_X1 U13846 ( .A1(n12077), .A2(n12838), .ZN(n12078) );
  NAND2_X1 U13847 ( .A1(n12078), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12080) );
  OAI211_X1 U13848 ( .C1(n12081), .C2(n12545), .A(n12080), .B(n12079), .ZN(
        n12082) );
  NOR2_X1 U13849 ( .A1(n12083), .A2(n12082), .ZN(n12085) );
  NAND2_X1 U13850 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12088) );
  NAND2_X1 U13851 ( .A1(n12159), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12087) );
  NAND2_X1 U13852 ( .A1(n12102), .A2(n17957), .ZN(n12093) );
  AOI21_X1 U13853 ( .B1(n17995), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12092) );
  INV_X1 U13854 ( .A(n12094), .ZN(n12096) );
  NAND2_X1 U13855 ( .A1(n12159), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12100) );
  NAND2_X1 U13856 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12099) );
  OAI211_X1 U13857 ( .C1(n16023), .C2(n16086), .A(n12100), .B(n12099), .ZN(
        n12101) );
  NAND2_X1 U13858 ( .A1(n12102), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12104) );
  NAND2_X1 U13859 ( .A1(n12212), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12103) );
  XNOR2_X2 U13860 ( .A(n12106), .B(n12105), .ZN(n12453) );
  INV_X1 U13861 ( .A(n12105), .ZN(n12107) );
  AND2_X1 U13862 ( .A1(n12107), .A2(n12106), .ZN(n12108) );
  NAND2_X1 U13863 ( .A1(n16025), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12112) );
  AOI22_X1 U13864 ( .A1(n12196), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12110) );
  NAND2_X1 U13865 ( .A1(n12192), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12109) );
  AND2_X1 U13866 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  NAND2_X1 U13867 ( .A1(n12112), .A2(n12111), .ZN(n14882) );
  NAND2_X1 U13868 ( .A1(n16025), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12114) );
  AOI22_X1 U13869 ( .A1(n12196), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12113) );
  OAI211_X1 U13870 ( .C1(n16023), .C2(n12115), .A(n12114), .B(n12113), .ZN(
        n14904) );
  NAND2_X1 U13871 ( .A1(n14905), .A2(n14904), .ZN(n14906) );
  AOI22_X1 U13872 ( .A1(n12196), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12117) );
  NAND2_X1 U13873 ( .A1(n12192), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12116) );
  NAND2_X1 U13874 ( .A1(n12117), .A2(n12116), .ZN(n12118) );
  AOI21_X1 U13875 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n12118), .ZN(n14966) );
  NAND2_X1 U13876 ( .A1(n16025), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12122) );
  AOI22_X1 U13877 ( .A1(n12196), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12120) );
  NAND2_X1 U13878 ( .A1(n12192), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n12119) );
  AND2_X1 U13879 ( .A1(n12120), .A2(n12119), .ZN(n12121) );
  NAND2_X1 U13880 ( .A1(n12122), .A2(n12121), .ZN(n14960) );
  INV_X1 U13881 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12125) );
  NAND2_X1 U13882 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U13883 ( .A1(n12196), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12123) );
  OAI211_X1 U13884 ( .C1(n16023), .C2(n12125), .A(n12124), .B(n12123), .ZN(
        n12126) );
  AOI21_X1 U13885 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12126), .ZN(n15370) );
  INV_X1 U13886 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U13887 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U13888 ( .A1(n12196), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12127) );
  OAI211_X1 U13889 ( .C1(n16023), .C2(n12129), .A(n12128), .B(n12127), .ZN(
        n12130) );
  AOI21_X1 U13890 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12130), .ZN(n15256) );
  INV_X1 U13891 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17894) );
  AOI22_X1 U13892 ( .A1(n12196), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12132) );
  NAND2_X1 U13893 ( .A1(n12192), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12131) );
  OAI211_X1 U13894 ( .C1(n12195), .C2(n17894), .A(n12132), .B(n12131), .ZN(
        n15589) );
  INV_X1 U13895 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12135) );
  NAND2_X1 U13896 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12134) );
  NAND2_X1 U13897 ( .A1(n12196), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12133) );
  OAI211_X1 U13898 ( .C1(n16023), .C2(n12135), .A(n12134), .B(n12133), .ZN(
        n12136) );
  AOI21_X1 U13899 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12136), .ZN(n15388) );
  NOR2_X4 U13900 ( .A1(n15588), .A2(n15388), .ZN(n15387) );
  AOI22_X1 U13901 ( .A1(n12196), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12138) );
  NAND2_X1 U13902 ( .A1(n12192), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12137) );
  NAND2_X1 U13903 ( .A1(n12138), .A2(n12137), .ZN(n12139) );
  AOI21_X1 U13904 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12139), .ZN(n15679) );
  INV_X1 U13905 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17847) );
  AOI22_X1 U13906 ( .A1(n12196), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12142) );
  NAND2_X1 U13907 ( .A1(n12192), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12141) );
  OAI211_X1 U13908 ( .C1(n12195), .C2(n17847), .A(n12142), .B(n12141), .ZN(
        n15638) );
  INV_X1 U13909 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U13910 ( .A1(n12196), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12144) );
  NAND2_X1 U13911 ( .A1(n12192), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12143) );
  OAI211_X1 U13912 ( .C1(n12195), .C2(n12811), .A(n12144), .B(n12143), .ZN(
        n15845) );
  INV_X1 U13913 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12147) );
  NAND2_X1 U13914 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U13915 ( .A1(n12196), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12145) );
  OAI211_X1 U13916 ( .C1(n16023), .C2(n12147), .A(n12146), .B(n12145), .ZN(
        n12148) );
  AOI21_X1 U13917 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12148), .ZN(n15801) );
  INV_X1 U13918 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U13919 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12150) );
  NAND2_X1 U13920 ( .A1(n12196), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12149) );
  OAI211_X1 U13921 ( .C1(n16023), .C2(n12151), .A(n12150), .B(n12149), .ZN(
        n12152) );
  AOI21_X1 U13922 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12152), .ZN(n15881) );
  INV_X1 U13923 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n17207) );
  NAND2_X1 U13924 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12155) );
  NAND2_X1 U13925 ( .A1(n12196), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12154) );
  OAI211_X1 U13926 ( .C1(n16023), .C2(n17207), .A(n12155), .B(n12154), .ZN(
        n12156) );
  AOI21_X1 U13927 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12156), .ZN(n15902) );
  INV_X1 U13928 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U13929 ( .A1(n12196), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12158) );
  NAND2_X1 U13930 ( .A1(n12192), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12157) );
  OAI211_X1 U13931 ( .C1(n12195), .C2(n12700), .A(n12158), .B(n12157), .ZN(
        n15930) );
  NAND2_X1 U13932 ( .A1(n15901), .A2(n15930), .ZN(n17312) );
  INV_X1 U13933 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12162) );
  NAND2_X1 U13934 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12161) );
  NAND2_X1 U13935 ( .A1(n12196), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12160) );
  OAI211_X1 U13936 ( .C1(n16023), .C2(n12162), .A(n12161), .B(n12160), .ZN(
        n12163) );
  AOI21_X1 U13937 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12163), .ZN(n17311) );
  INV_X1 U13938 ( .A(n12164), .ZN(n17304) );
  AOI22_X1 U13939 ( .A1(n12196), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12166) );
  NAND2_X1 U13940 ( .A1(n12192), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12165) );
  NAND2_X1 U13941 ( .A1(n12166), .A2(n12165), .ZN(n12167) );
  AOI21_X1 U13942 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12167), .ZN(n17306) );
  NOR2_X4 U13943 ( .A1(n17304), .A2(n17306), .ZN(n17305) );
  INV_X1 U13944 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U13945 ( .A1(n12196), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n12169) );
  NAND2_X1 U13946 ( .A1(n12192), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12168) );
  OAI211_X1 U13947 ( .C1(n12195), .C2(n12851), .A(n12169), .B(n12168), .ZN(
        n12814) );
  INV_X1 U13948 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12172) );
  NAND2_X1 U13949 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12171) );
  NAND2_X1 U13950 ( .A1(n12196), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12170) );
  OAI211_X1 U13951 ( .C1(n16023), .C2(n12172), .A(n12171), .B(n12170), .ZN(
        n12173) );
  AOI21_X1 U13952 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12173), .ZN(n17289) );
  INV_X1 U13953 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12176) );
  NAND2_X1 U13954 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12175) );
  NAND2_X1 U13955 ( .A1(n12196), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12174) );
  OAI211_X1 U13956 ( .C1(n16023), .C2(n12176), .A(n12175), .B(n12174), .ZN(
        n12177) );
  AOI21_X1 U13957 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12177), .ZN(n17281) );
  INV_X1 U13958 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17707) );
  AOI22_X1 U13959 ( .A1(n12196), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12179) );
  NAND2_X1 U13960 ( .A1(n12192), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12178) );
  OAI211_X1 U13961 ( .C1(n12195), .C2(n17707), .A(n12179), .B(n12178), .ZN(
        n17271) );
  INV_X1 U13962 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17700) );
  AOI22_X1 U13963 ( .A1(n12196), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12181) );
  NAND2_X1 U13964 ( .A1(n12192), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12180) );
  OAI211_X1 U13965 ( .C1(n12195), .C2(n17700), .A(n12181), .B(n12180), .ZN(
        n17265) );
  NAND2_X1 U13966 ( .A1(n17273), .A2(n17265), .ZN(n17259) );
  INV_X1 U13967 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12184) );
  NAND2_X1 U13968 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U13969 ( .A1(n12196), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12182) );
  OAI211_X1 U13970 ( .C1(n16023), .C2(n12184), .A(n12183), .B(n12182), .ZN(
        n12185) );
  AOI21_X1 U13971 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12185), .ZN(n17260) );
  OR2_X2 U13972 ( .A1(n17259), .A2(n17260), .ZN(n17262) );
  AOI22_X1 U13973 ( .A1(n12196), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12187) );
  NAND2_X1 U13974 ( .A1(n12192), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12186) );
  NAND2_X1 U13975 ( .A1(n12187), .A2(n12186), .ZN(n12188) );
  AOI21_X1 U13976 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12188), .ZN(n17182) );
  INV_X1 U13977 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n19463) );
  NAND2_X1 U13978 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12190) );
  NAND2_X1 U13979 ( .A1(n12196), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12189) );
  OAI211_X1 U13980 ( .C1(n16023), .C2(n19463), .A(n12190), .B(n12189), .ZN(
        n12191) );
  AOI21_X1 U13981 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12191), .ZN(n16058) );
  INV_X1 U13982 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17659) );
  AOI22_X1 U13983 ( .A1(n12196), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12194) );
  NAND2_X1 U13984 ( .A1(n12192), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12193) );
  OAI211_X1 U13985 ( .C1(n12195), .C2(n17659), .A(n12194), .B(n12193), .ZN(
        n14151) );
  INV_X1 U13986 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U13987 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12198) );
  NAND2_X1 U13988 ( .A1(n12196), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12197) );
  OAI211_X1 U13989 ( .C1(n16023), .C2(n12199), .A(n12198), .B(n12197), .ZN(
        n12200) );
  AOI21_X1 U13990 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12200), .ZN(n12204) );
  INV_X1 U13991 ( .A(n12204), .ZN(n12201) );
  NAND2_X1 U13992 ( .A1(n12203), .A2(n12204), .ZN(n12205) );
  AND2_X1 U13993 ( .A1(n12721), .A2(n12208), .ZN(n12206) );
  NOR2_X1 U13994 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n17993) );
  NAND2_X1 U13995 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17993), .ZN(n18158) );
  INV_X1 U13996 ( .A(n18158), .ZN(n12207) );
  NOR2_X1 U13997 ( .A1(n19566), .A2(n22453), .ZN(n15334) );
  INV_X1 U13998 ( .A(n15334), .ZN(n15275) );
  NOR2_X1 U13999 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15275), .ZN(n12448) );
  INV_X1 U14000 ( .A(n12208), .ZN(n12209) );
  NAND2_X1 U14001 ( .A1(n17243), .A2(n12209), .ZN(n12210) );
  AND2_X1 U14002 ( .A1(n11259), .A2(n12210), .ZN(n12211) );
  NOR2_X1 U14003 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n17995), .ZN(n19565) );
  NAND3_X1 U14004 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19565), .A3(n17948), 
        .ZN(n19577) );
  INV_X1 U14005 ( .A(n19577), .ZN(n12214) );
  NAND2_X1 U14006 ( .A1(n19301), .A2(n19563), .ZN(n12213) );
  AOI22_X1 U14007 ( .A1(n19491), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19495), .ZN(n12216) );
  NAND2_X1 U14008 ( .A1(n19494), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12215) );
  OAI211_X1 U14009 ( .C1(n17651), .C2(n19467), .A(n12216), .B(n12215), .ZN(
        n12217) );
  AOI21_X1 U14010 ( .B1(n16009), .B2(n19492), .A(n12217), .ZN(n12452) );
  NAND2_X1 U14011 ( .A1(n12239), .A2(n12218), .ZN(n12390) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12223) );
  NAND2_X1 U14013 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12222) );
  AOI22_X1 U14014 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U14015 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12220) );
  AND4_X1 U14016 ( .A1(n12223), .A2(n12222), .A3(n12221), .A4(n12220), .ZN(
        n12236) );
  NAND2_X1 U14017 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12227) );
  NAND2_X1 U14018 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12226) );
  INV_X1 U14019 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20671) );
  NAND2_X1 U14020 ( .A1(n13948), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12225) );
  NAND2_X1 U14021 ( .A1(n13950), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12224) );
  AND4_X1 U14022 ( .A1(n12227), .A2(n12226), .A3(n12225), .A4(n12224), .ZN(
        n12235) );
  NAND2_X1 U14023 ( .A1(n12228), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12232) );
  NAND2_X1 U14024 ( .A1(n13946), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12231) );
  NAND2_X1 U14025 ( .A1(n13947), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12230) );
  NAND2_X1 U14026 ( .A1(n12300), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12229) );
  AND4_X1 U14027 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12234) );
  AOI22_X1 U14028 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12233) );
  INV_X1 U14029 ( .A(n14542), .ZN(n12544) );
  NOR2_X1 U14030 ( .A1(n11242), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12255) );
  AND2_X1 U14031 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12237) );
  NOR2_X1 U14032 ( .A1(n12255), .A2(n12237), .ZN(n12238) );
  AND2_X2 U14033 ( .A1(n11259), .A2(n20162), .ZN(n12262) );
  NAND2_X1 U14034 ( .A1(n14125), .A2(n12262), .ZN(n12253) );
  NAND2_X1 U14035 ( .A1(n16041), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12243) );
  NAND2_X1 U14036 ( .A1(n11259), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12240) );
  OAI211_X1 U14037 ( .C1(n11242), .C2(n18129), .A(n12240), .B(n20162), .ZN(
        n12241) );
  INV_X1 U14038 ( .A(n12241), .ZN(n12242) );
  NAND2_X1 U14039 ( .A1(n12243), .A2(n12242), .ZN(n15602) );
  NAND2_X1 U14040 ( .A1(n15601), .A2(n15602), .ZN(n12250) );
  NAND2_X1 U14041 ( .A1(n16041), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U14042 ( .A1(n12255), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12262), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12244) );
  AND2_X1 U14043 ( .A1(n12245), .A2(n12244), .ZN(n12251) );
  INV_X1 U14044 ( .A(n12251), .ZN(n12246) );
  XNOR2_X1 U14045 ( .A(n12250), .B(n12246), .ZN(n14839) );
  INV_X1 U14046 ( .A(n11242), .ZN(n20087) );
  OAI22_X1 U14047 ( .A1(n12247), .A2(n11259), .B1(n20087), .B2(n14125), .ZN(
        n12248) );
  INV_X1 U14048 ( .A(n12248), .ZN(n12249) );
  NAND2_X1 U14049 ( .A1(n12251), .A2(n12250), .ZN(n12252) );
  NAND2_X1 U14050 ( .A1(n14838), .A2(n12252), .ZN(n12259) );
  OR2_X1 U14051 ( .A1(n12390), .A2(n12778), .ZN(n12254) );
  OAI211_X1 U14052 ( .C1(n20162), .C2(n20161), .A(n12254), .B(n12253), .ZN(
        n12258) );
  XNOR2_X1 U14053 ( .A(n12259), .B(n12258), .ZN(n15600) );
  NAND2_X1 U14054 ( .A1(n16041), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U14055 ( .A1(n16040), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12262), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12256) );
  AND2_X1 U14056 ( .A1(n12257), .A2(n12256), .ZN(n15599) );
  INV_X1 U14057 ( .A(n12258), .ZN(n12260) );
  NAND2_X1 U14058 ( .A1(n12260), .A2(n12259), .ZN(n12261) );
  NAND2_X1 U14059 ( .A1(n16041), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U14060 ( .A1(n12262), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12264) );
  NAND2_X1 U14061 ( .A1(n16040), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12263) );
  AND2_X1 U14062 ( .A1(n12264), .A2(n12263), .ZN(n12267) );
  INV_X1 U14063 ( .A(n12511), .ZN(n12265) );
  OR2_X1 U14064 ( .A1(n12390), .A2(n12265), .ZN(n12266) );
  INV_X1 U14065 ( .A(n12390), .ZN(n12411) );
  AOI22_X1 U14066 ( .A1(n12411), .A2(n12785), .B1(n16041), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U14067 ( .A1(n16040), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12262), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12269) );
  NAND2_X1 U14068 ( .A1(n12270), .A2(n12269), .ZN(n15611) );
  NAND2_X1 U14069 ( .A1(n16041), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U14070 ( .A1(n16040), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12262), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12271) );
  OAI211_X1 U14071 ( .C1(n12597), .C2(n12390), .A(n12272), .B(n12271), .ZN(
        n15657) );
  NAND2_X1 U14072 ( .A1(n15658), .A2(n15657), .ZN(n15656) );
  OR2_X1 U14073 ( .A1(n12390), .A2(n12630), .ZN(n12273) );
  NAND2_X1 U14074 ( .A1(n16041), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U14075 ( .A1(n16040), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12262), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12274) );
  NAND2_X1 U14076 ( .A1(n12275), .A2(n12274), .ZN(n15717) );
  NAND2_X1 U14077 ( .A1(n15718), .A2(n15717), .ZN(n15716) );
  OR2_X1 U14078 ( .A1(n12390), .A2(n16007), .ZN(n12276) );
  INV_X1 U14079 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n17640) );
  AOI22_X1 U14080 ( .A1(n16040), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12262), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12277) );
  OAI21_X1 U14081 ( .B1(n12445), .B2(n17640), .A(n12277), .ZN(n17939) );
  NAND2_X1 U14082 ( .A1(n17938), .A2(n17939), .ZN(n17922) );
  NAND2_X1 U14083 ( .A1(n16041), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U14084 ( .A1(n16040), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12262), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U14085 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n13946), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U14086 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n13949), .B1(
        n13951), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U14087 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13947), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U14088 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12278) );
  NAND4_X1 U14089 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12289) );
  NAND2_X1 U14090 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12283) );
  AOI22_X1 U14091 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12282) );
  AND2_X1 U14092 ( .A1(n12283), .A2(n12282), .ZN(n12287) );
  AOI22_X1 U14093 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13961), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U14094 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U14095 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12284) );
  NAND4_X1 U14096 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12288) );
  NOR2_X1 U14097 ( .A1(n12289), .A2(n12288), .ZN(n15375) );
  OR2_X1 U14098 ( .A1(n12390), .A2(n15375), .ZN(n12290) );
  NAND2_X1 U14099 ( .A1(n16041), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U14100 ( .A1(n16040), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12262), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U14101 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12296) );
  NAND2_X1 U14102 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12295) );
  AOI22_X1 U14103 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12294) );
  NAND2_X1 U14104 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12293) );
  NAND4_X1 U14105 ( .A1(n12296), .A2(n12295), .A3(n12294), .A4(n12293), .ZN(
        n12299) );
  INV_X1 U14106 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20545) );
  INV_X1 U14107 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12297) );
  OAI22_X1 U14108 ( .A1(n13919), .A2(n20545), .B1(n13917), .B2(n12297), .ZN(
        n12298) );
  NOR2_X1 U14109 ( .A1(n12299), .A2(n12298), .ZN(n12309) );
  AOI22_X1 U14110 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U14111 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12307) );
  INV_X1 U14112 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12302) );
  INV_X1 U14113 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12301) );
  OAI22_X1 U14114 ( .A1(n12401), .A2(n12302), .B1(n12399), .B2(n12301), .ZN(
        n12305) );
  INV_X1 U14115 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13983) );
  INV_X1 U14116 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12303) );
  OAI22_X1 U14117 ( .A1(n12404), .A2(n13983), .B1(n15294), .B2(n12303), .ZN(
        n12304) );
  NOR2_X1 U14118 ( .A1(n12305), .A2(n12304), .ZN(n12306) );
  NAND4_X1 U14119 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n15254) );
  NAND2_X1 U14120 ( .A1(n12411), .A2(n15254), .ZN(n12310) );
  NAND2_X1 U14121 ( .A1(n16041), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U14122 ( .A1(n16040), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U14123 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n12300), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U14124 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13946), .B1(
        n13947), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U14125 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n13948), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U14126 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12313) );
  NAND4_X1 U14127 ( .A1(n12316), .A2(n12315), .A3(n12314), .A4(n12313), .ZN(
        n12324) );
  AOI22_X1 U14128 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n13962), .B1(
        n13949), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U14129 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U14130 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12319) );
  AOI22_X1 U14131 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U14132 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12317) );
  AND4_X1 U14133 ( .A1(n12320), .A2(n12319), .A3(n12318), .A4(n12317), .ZN(
        n12321) );
  NAND2_X1 U14134 ( .A1(n12322), .A2(n12321), .ZN(n12323) );
  NOR2_X1 U14135 ( .A1(n12324), .A2(n12323), .ZN(n15590) );
  OR2_X1 U14136 ( .A1(n12390), .A2(n15590), .ZN(n12325) );
  INV_X1 U14137 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U14138 ( .A1(n16040), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U14139 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12331) );
  NAND2_X1 U14140 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12330) );
  AOI22_X1 U14141 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12329) );
  NAND2_X1 U14142 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12328) );
  NAND4_X1 U14143 ( .A1(n12331), .A2(n12330), .A3(n12329), .A4(n12328), .ZN(
        n12333) );
  INV_X1 U14144 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12502) );
  OAI22_X1 U14145 ( .A1(n13919), .A2(n15784), .B1(n13917), .B2(n12502), .ZN(
        n12332) );
  NOR2_X1 U14146 ( .A1(n12333), .A2(n12332), .ZN(n12341) );
  AOI22_X1 U14147 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U14148 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12339) );
  INV_X1 U14149 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12334) );
  OAI22_X1 U14150 ( .A1(n12401), .A2(n12335), .B1(n12399), .B2(n12334), .ZN(
        n12337) );
  INV_X1 U14151 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12465) );
  OAI22_X1 U14152 ( .A1(n12404), .A2(n14032), .B1(n15294), .B2(n12465), .ZN(
        n12336) );
  NOR2_X1 U14153 ( .A1(n12337), .A2(n12336), .ZN(n12338) );
  NAND4_X1 U14154 ( .A1(n12341), .A2(n12340), .A3(n12339), .A4(n12338), .ZN(
        n15386) );
  NAND2_X1 U14155 ( .A1(n12411), .A2(n15386), .ZN(n12342) );
  OAI211_X1 U14156 ( .C1(n12445), .C2(n12344), .A(n12343), .B(n12342), .ZN(
        n17873) );
  NAND2_X1 U14157 ( .A1(n17874), .A2(n17873), .ZN(n17860) );
  NAND2_X1 U14158 ( .A1(n16041), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U14159 ( .A1(n16040), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U14160 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12228), .B1(
        n13956), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U14161 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13949), .B1(
        n13951), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U14162 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13946), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U14163 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12345) );
  NAND4_X1 U14164 ( .A1(n12348), .A2(n12347), .A3(n12346), .A4(n12345), .ZN(
        n12356) );
  NAND2_X1 U14165 ( .A1(n13947), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12350) );
  AOI22_X1 U14166 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13964), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12349) );
  AND2_X1 U14167 ( .A1(n12350), .A2(n12349), .ZN(n12354) );
  AOI22_X1 U14168 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n13961), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U14169 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13958), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12352) );
  NAND2_X1 U14170 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12351) );
  NAND4_X1 U14171 ( .A1(n12354), .A2(n12353), .A3(n12352), .A4(n12351), .ZN(
        n12355) );
  NOR2_X1 U14172 ( .A1(n12356), .A2(n12355), .ZN(n15683) );
  OR2_X1 U14173 ( .A1(n12390), .A2(n15683), .ZN(n12357) );
  NAND2_X1 U14174 ( .A1(n16041), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U14175 ( .A1(n16040), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U14176 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12363) );
  NAND2_X1 U14177 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12362) );
  AOI22_X1 U14178 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12361) );
  NAND2_X1 U14179 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12360) );
  NAND4_X1 U14180 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n12365) );
  INV_X1 U14181 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12590) );
  OAI22_X1 U14182 ( .A1(n13919), .A2(n20360), .B1(n13917), .B2(n12590), .ZN(
        n12364) );
  NOR2_X1 U14183 ( .A1(n12365), .A2(n12364), .ZN(n12372) );
  AOI22_X1 U14184 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U14185 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12370) );
  INV_X1 U14186 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12366) );
  INV_X1 U14187 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13904) );
  OAI22_X1 U14188 ( .A1(n12401), .A2(n12366), .B1(n12399), .B2(n13904), .ZN(
        n12368) );
  INV_X1 U14189 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14079) );
  INV_X1 U14190 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12589) );
  OAI22_X1 U14191 ( .A1(n12404), .A2(n14079), .B1(n15294), .B2(n12589), .ZN(
        n12367) );
  NOR2_X1 U14192 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  NAND4_X1 U14193 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n15636) );
  NAND2_X1 U14194 ( .A1(n12411), .A2(n15636), .ZN(n12373) );
  AOI22_X1 U14195 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n13956), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U14196 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13947), .B1(
        n13946), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U14197 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n13948), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U14198 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12376) );
  NAND4_X1 U14199 ( .A1(n12379), .A2(n12378), .A3(n12377), .A4(n12376), .ZN(
        n12387) );
  AOI22_X1 U14200 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13962), .B1(
        n13949), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U14201 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13958), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12383) );
  NAND2_X1 U14202 ( .A1(n12300), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12382) );
  AOI22_X1 U14203 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13964), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12381) );
  NAND2_X1 U14204 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12380) );
  AND4_X1 U14205 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n12384) );
  NAND2_X1 U14206 ( .A1(n12385), .A2(n12384), .ZN(n12386) );
  NOR2_X1 U14207 ( .A1(n12387), .A2(n12386), .ZN(n15849) );
  NAND2_X1 U14208 ( .A1(n16041), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U14209 ( .A1(n16040), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12388) );
  OAI211_X1 U14210 ( .C1(n15849), .C2(n12390), .A(n12389), .B(n12388), .ZN(
        n17841) );
  NAND2_X1 U14211 ( .A1(n16041), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U14212 ( .A1(n16040), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U14213 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12394) );
  NAND2_X1 U14214 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12393) );
  AOI22_X1 U14215 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12392) );
  NAND2_X1 U14216 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12391) );
  NAND4_X1 U14217 ( .A1(n12394), .A2(n12393), .A3(n12392), .A4(n12391), .ZN(
        n12397) );
  INV_X1 U14218 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20268) );
  INV_X1 U14219 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12395) );
  OAI22_X1 U14220 ( .A1(n13919), .A2(n20268), .B1(n13917), .B2(n12395), .ZN(
        n12396) );
  NOR2_X1 U14221 ( .A1(n12397), .A2(n12396), .ZN(n12410) );
  AOI22_X1 U14222 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U14223 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12408) );
  INV_X1 U14224 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12400) );
  INV_X1 U14225 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12398) );
  OAI22_X1 U14226 ( .A1(n12401), .A2(n12400), .B1(n12399), .B2(n12398), .ZN(
        n12406) );
  INV_X1 U14227 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12403) );
  INV_X1 U14228 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12402) );
  OAI22_X1 U14229 ( .A1(n12404), .A2(n12403), .B1(n15294), .B2(n12402), .ZN(
        n12405) );
  NOR2_X1 U14230 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  NAND4_X1 U14231 ( .A1(n12410), .A2(n12409), .A3(n12408), .A4(n12407), .ZN(
        n15798) );
  NAND2_X1 U14232 ( .A1(n12411), .A2(n15798), .ZN(n12412) );
  NAND2_X1 U14233 ( .A1(n16041), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U14234 ( .A1(n16040), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12417) );
  INV_X1 U14235 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U14236 ( .A1(n16040), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12419) );
  OAI21_X1 U14237 ( .B1(n12445), .B2(n12420), .A(n12419), .ZN(n15889) );
  INV_X1 U14238 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19365) );
  AOI22_X1 U14239 ( .A1(n16040), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12421) );
  OAI21_X1 U14240 ( .B1(n12445), .B2(n19365), .A(n12421), .ZN(n15920) );
  NAND2_X1 U14241 ( .A1(n16041), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U14242 ( .A1(n16040), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12422) );
  AND2_X1 U14243 ( .A1(n12423), .A2(n12422), .ZN(n17399) );
  NAND2_X1 U14244 ( .A1(n16041), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U14245 ( .A1(n16040), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12426) );
  AND2_X1 U14246 ( .A1(n12427), .A2(n12426), .ZN(n17389) );
  NAND2_X1 U14247 ( .A1(n16041), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U14248 ( .A1(n16040), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12428) );
  INV_X1 U14249 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U14250 ( .A1(n16040), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12430) );
  OAI21_X1 U14251 ( .B1(n12445), .B2(n17496), .A(n12430), .ZN(n17371) );
  NAND2_X1 U14252 ( .A1(n16041), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U14253 ( .A1(n16040), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12431) );
  AND2_X1 U14254 ( .A1(n12432), .A2(n12431), .ZN(n17365) );
  NAND2_X1 U14255 ( .A1(n16041), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U14256 ( .A1(n16040), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12433) );
  INV_X1 U14257 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U14258 ( .A1(n16040), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12435) );
  OAI21_X1 U14259 ( .B1(n12445), .B2(n12436), .A(n12435), .ZN(n17340) );
  NAND2_X1 U14260 ( .A1(n17341), .A2(n17340), .ZN(n17330) );
  NAND2_X1 U14261 ( .A1(n16041), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U14262 ( .A1(n16040), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12437) );
  AND2_X1 U14263 ( .A1(n12438), .A2(n12437), .ZN(n17331) );
  NAND2_X1 U14264 ( .A1(n16041), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U14265 ( .A1(n16040), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12439) );
  INV_X1 U14266 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U14267 ( .A1(n16040), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12441) );
  OAI21_X1 U14268 ( .B1(n12445), .B2(n12442), .A(n12441), .ZN(n16064) );
  INV_X1 U14269 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U14270 ( .A1(n16040), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12443) );
  OAI21_X1 U14271 ( .B1(n12445), .B2(n12444), .A(n12443), .ZN(n14126) );
  NAND2_X1 U14272 ( .A1(n16041), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U14273 ( .A1(n16040), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12262), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12446) );
  AND2_X1 U14274 ( .A1(n12447), .A2(n12446), .ZN(n16038) );
  INV_X1 U14275 ( .A(n17652), .ZN(n12450) );
  AND2_X1 U14276 ( .A1(n14548), .A2(n12448), .ZN(n15354) );
  NAND2_X2 U14277 ( .A1(n12472), .A2(n12461), .ZN(n19515) );
  NAND2_X1 U14278 ( .A1(n11261), .A2(n12478), .ZN(n12500) );
  INV_X1 U14280 ( .A(n12461), .ZN(n12462) );
  NOR2_X1 U14281 ( .A1(n12476), .A2(n12462), .ZN(n12481) );
  OAI22_X1 U14282 ( .A1(n12465), .A2(n12622), .B1(n20128), .B2(n12464), .ZN(
        n12466) );
  INV_X1 U14283 ( .A(n12466), .ZN(n12487) );
  INV_X1 U14284 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12470) );
  NAND2_X1 U14285 ( .A1(n19551), .A2(n12478), .ZN(n12467) );
  OR2_X1 U14286 ( .A1(n11260), .A2(n12467), .ZN(n12576) );
  NAND2_X1 U14287 ( .A1(n19551), .A2(n12481), .ZN(n12468) );
  OAI22_X1 U14288 ( .A1(n12470), .A2(n12576), .B1(n12577), .B2(n12469), .ZN(
        n12471) );
  INV_X1 U14289 ( .A(n12471), .ZN(n12486) );
  INV_X1 U14290 ( .A(n12472), .ZN(n12474) );
  INV_X1 U14291 ( .A(n12456), .ZN(n12473) );
  NAND2_X1 U14292 ( .A1(n12474), .A2(n12473), .ZN(n12475) );
  INV_X1 U14293 ( .A(n17238), .ZN(n14646) );
  NAND2_X1 U14294 ( .A1(n12488), .A2(n12463), .ZN(n12529) );
  INV_X1 U14295 ( .A(n12529), .ZN(n12477) );
  NAND2_X1 U14296 ( .A1(n12477), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12485) );
  INV_X1 U14297 ( .A(n12478), .ZN(n12479) );
  OR2_X1 U14298 ( .A1(n19551), .A2(n12479), .ZN(n12480) );
  INV_X1 U14299 ( .A(n12481), .ZN(n12482) );
  AOI22_X1 U14300 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12573), .B1(
        n12574), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12484) );
  AND2_X1 U14301 ( .A1(n19551), .A2(n17238), .ZN(n12493) );
  AND2_X2 U14302 ( .A1(n12496), .A2(n12493), .ZN(n20100) );
  NAND2_X1 U14303 ( .A1(n20100), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12491) );
  INV_X1 U14304 ( .A(n19515), .ZN(n15700) );
  OR2_X1 U14305 ( .A1(n19551), .A2(n14646), .ZN(n12495) );
  NAND2_X1 U14306 ( .A1(n12519), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12490) );
  OAI211_X1 U14307 ( .C1(n12575), .C2(n14032), .A(n12491), .B(n12490), .ZN(
        n12492) );
  INV_X1 U14308 ( .A(n12492), .ZN(n12509) );
  INV_X1 U14309 ( .A(n12505), .ZN(n12494) );
  INV_X1 U14310 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12499) );
  INV_X1 U14311 ( .A(n12495), .ZN(n12497) );
  INV_X1 U14312 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12498) );
  OAI22_X1 U14313 ( .A1(n12568), .A2(n12499), .B1(n20138), .B2(n12498), .ZN(
        n12504) );
  OAI22_X1 U14314 ( .A1(n12502), .A2(n20111), .B1(n12621), .B2(n14034), .ZN(
        n12503) );
  NOR2_X1 U14315 ( .A1(n12504), .A2(n12503), .ZN(n12508) );
  AND2_X2 U14316 ( .A1(n12506), .A2(n12463), .ZN(n12585) );
  AOI22_X1 U14317 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12585), .B1(
        n12567), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12507) );
  NAND4_X1 U14318 ( .A1(n12510), .A2(n12509), .A3(n12508), .A4(n12507), .ZN(
        n12513) );
  OR2_X1 U14319 ( .A1(n11259), .A2(n12511), .ZN(n12512) );
  AOI22_X1 U14320 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12585), .B1(
        n12567), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U14321 ( .A1(n12573), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12515) );
  NAND2_X1 U14322 ( .A1(n20100), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12514) );
  AND2_X1 U14323 ( .A1(n12517), .A2(n11725), .ZN(n12533) );
  INV_X1 U14324 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13845) );
  INV_X1 U14325 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12518) );
  OAI22_X1 U14326 ( .A1(n12568), .A2(n13845), .B1(n20138), .B2(n12518), .ZN(
        n12522) );
  INV_X1 U14327 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12520) );
  INV_X1 U14328 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13985) );
  OAI22_X1 U14329 ( .A1(n12586), .A2(n12520), .B1(n20128), .B2(n13985), .ZN(
        n12521) );
  NOR2_X1 U14330 ( .A1(n12522), .A2(n12521), .ZN(n12532) );
  INV_X1 U14331 ( .A(n12576), .ZN(n20197) );
  AND2_X1 U14332 ( .A1(n12524), .A2(n12523), .ZN(n12528) );
  INV_X1 U14333 ( .A(n20111), .ZN(n20106) );
  NAND2_X1 U14334 ( .A1(n20106), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12527) );
  NAND2_X1 U14335 ( .A1(n20154), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12526) );
  NAND2_X1 U14336 ( .A1(n20088), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12525) );
  AOI22_X1 U14337 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20166), .B1(
        n20121), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12530) );
  NAND4_X1 U14338 ( .A1(n12533), .A2(n12532), .A3(n12531), .A4(n12530), .ZN(
        n12536) );
  NOR2_X1 U14339 ( .A1(n12544), .A2(n12776), .ZN(n12534) );
  NAND2_X1 U14340 ( .A1(n19264), .A2(n12534), .ZN(n12779) );
  NAND2_X1 U14341 ( .A1(n12779), .A2(n12778), .ZN(n12535) );
  NAND2_X1 U14342 ( .A1(n15548), .A2(n16007), .ZN(n12541) );
  INV_X1 U14343 ( .A(n12537), .ZN(n12539) );
  INV_X1 U14344 ( .A(n12538), .ZN(n12549) );
  NAND2_X1 U14345 ( .A1(n12539), .A2(n12549), .ZN(n12540) );
  NAND2_X1 U14346 ( .A1(n12557), .A2(n12540), .ZN(n16090) );
  INV_X1 U14347 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15624) );
  NAND2_X1 U14348 ( .A1(n15306), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12542) );
  NAND2_X1 U14349 ( .A1(n12543), .A2(n12542), .ZN(n12723) );
  MUX2_X1 U14350 ( .A(n12723), .B(n12544), .S(n12721), .Z(n12546) );
  MUX2_X1 U14351 ( .A(n12546), .B(n12545), .S(n20322), .Z(n15697) );
  NOR2_X1 U14352 ( .A1(n15697), .A2(n19512), .ZN(n12548) );
  AND3_X1 U14353 ( .A1(n20322), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12547) );
  NOR2_X1 U14354 ( .A1(n12551), .A2(n12547), .ZN(n17228) );
  NOR2_X1 U14355 ( .A1(n12548), .A2(n17228), .ZN(n14641) );
  AND2_X1 U14356 ( .A1(n12548), .A2(n17228), .ZN(n14640) );
  NOR2_X1 U14357 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14640), .ZN(
        n14639) );
  NOR2_X1 U14358 ( .A1(n14641), .A2(n14639), .ZN(n14634) );
  OAI21_X1 U14359 ( .B1(n12551), .B2(n12550), .A(n12549), .ZN(n12552) );
  XNOR2_X1 U14360 ( .A(n12552), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14633) );
  NAND2_X1 U14361 ( .A1(n14634), .A2(n14633), .ZN(n12554) );
  INV_X1 U14362 ( .A(n12552), .ZN(n15711) );
  NAND2_X1 U14363 ( .A1(n15711), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12553) );
  NAND2_X1 U14364 ( .A1(n12554), .A2(n12553), .ZN(n15547) );
  NAND2_X1 U14365 ( .A1(n12555), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12556) );
  NAND2_X1 U14366 ( .A1(n12558), .A2(n12557), .ZN(n12559) );
  NAND2_X1 U14367 ( .A1(n12602), .A2(n12559), .ZN(n12560) );
  XNOR2_X1 U14368 ( .A(n12560), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15619) );
  INV_X1 U14369 ( .A(n12560), .ZN(n15750) );
  NAND2_X1 U14370 ( .A1(n15750), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12561) );
  NAND2_X1 U14371 ( .A1(n12562), .A2(n12561), .ZN(n15825) );
  INV_X1 U14372 ( .A(n12563), .ZN(n12565) );
  NAND2_X1 U14373 ( .A1(n12565), .A2(n12564), .ZN(n12787) );
  INV_X1 U14374 ( .A(n12787), .ZN(n12566) );
  INV_X1 U14375 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12569) );
  INV_X1 U14376 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13903) );
  OAI22_X1 U14377 ( .A1(n12568), .A2(n12569), .B1(n20096), .B2(n13903), .ZN(
        n12570) );
  AOI21_X1 U14378 ( .B1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B2(n11228), .A(
        n12570), .ZN(n12596) );
  INV_X1 U14379 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14081) );
  INV_X1 U14380 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12571) );
  OAI22_X1 U14381 ( .A1(n14081), .A2(n20128), .B1(n12621), .B2(n12571), .ZN(
        n12572) );
  INV_X1 U14382 ( .A(n12572), .ZN(n12584) );
  AOI22_X1 U14383 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n12573), .B1(
        n20226), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12583) );
  OR2_X1 U14384 ( .A1(n12575), .A2(n14079), .ZN(n12582) );
  INV_X1 U14385 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12579) );
  INV_X1 U14386 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12578) );
  OAI22_X1 U14387 ( .A1(n12579), .A2(n12576), .B1(n12577), .B2(n12578), .ZN(
        n12580) );
  INV_X1 U14388 ( .A(n12580), .ZN(n12581) );
  AOI22_X1 U14389 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12585), .B1(
        n20166), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12594) );
  INV_X1 U14390 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12588) );
  INV_X1 U14391 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12587) );
  OAI22_X1 U14392 ( .A1(n12586), .A2(n12588), .B1(n20138), .B2(n12587), .ZN(
        n12592) );
  OAI22_X1 U14393 ( .A1(n12590), .A2(n20111), .B1(n12622), .B2(n12589), .ZN(
        n12591) );
  NOR2_X1 U14394 ( .A1(n12592), .A2(n12591), .ZN(n12593) );
  NAND4_X1 U14395 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12599) );
  NAND2_X1 U14396 ( .A1(n12597), .A2(n19264), .ZN(n12598) );
  NAND2_X1 U14397 ( .A1(n12792), .A2(n16007), .ZN(n12604) );
  INV_X1 U14398 ( .A(n12600), .ZN(n12601) );
  NAND2_X1 U14399 ( .A1(n12602), .A2(n12601), .ZN(n12603) );
  NAND2_X1 U14400 ( .A1(n12635), .A2(n12603), .ZN(n15665) );
  INV_X1 U14401 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15837) );
  XNOR2_X1 U14402 ( .A(n12605), .B(n15837), .ZN(n15826) );
  NAND2_X1 U14403 ( .A1(n15825), .A2(n15826), .ZN(n12607) );
  NAND2_X1 U14404 ( .A1(n12605), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12606) );
  NAND2_X1 U14405 ( .A1(n12607), .A2(n12606), .ZN(n18075) );
  INV_X1 U14406 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12610) );
  INV_X1 U14407 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13916) );
  OAI22_X1 U14408 ( .A1(n12568), .A2(n12610), .B1(n20096), .B2(n13916), .ZN(
        n12611) );
  AOI21_X1 U14409 ( .B1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n20166), .A(
        n12611), .ZN(n12629) );
  INV_X1 U14410 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12612) );
  INV_X1 U14411 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14106) );
  OAI22_X1 U14412 ( .A1(n12612), .A2(n20111), .B1(n20128), .B2(n14106), .ZN(
        n12613) );
  INV_X1 U14413 ( .A(n12613), .ZN(n12619) );
  INV_X1 U14414 ( .A(n11228), .ZN(n20210) );
  INV_X1 U14415 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14095) );
  OR2_X1 U14416 ( .A1(n20210), .A2(n14095), .ZN(n12618) );
  AOI22_X1 U14417 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12573), .B1(
        n20226), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12617) );
  INV_X1 U14418 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12614) );
  INV_X1 U14419 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14097) );
  OAI22_X1 U14420 ( .A1(n12614), .A2(n12576), .B1(n12577), .B2(n14097), .ZN(
        n12615) );
  INV_X1 U14421 ( .A(n12615), .ZN(n12616) );
  AOI22_X1 U14422 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12585), .B1(
        n20121), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12627) );
  INV_X1 U14423 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14098) );
  INV_X1 U14424 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14107) );
  OAI22_X1 U14425 ( .A1(n12586), .A2(n14098), .B1(n20138), .B2(n14107), .ZN(
        n12625) );
  INV_X1 U14426 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12623) );
  INV_X1 U14427 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12620) );
  OAI22_X1 U14428 ( .A1(n12623), .A2(n12622), .B1(n12621), .B2(n12620), .ZN(
        n12624) );
  NOR2_X1 U14429 ( .A1(n12625), .A2(n12624), .ZN(n12626) );
  NAND4_X1 U14430 ( .A1(n12629), .A2(n12628), .A3(n12627), .A4(n12626), .ZN(
        n12632) );
  NAND2_X1 U14431 ( .A1(n12630), .A2(n19264), .ZN(n12631) );
  NAND2_X1 U14432 ( .A1(n12635), .A2(n11550), .ZN(n12636) );
  NAND2_X1 U14433 ( .A1(n16013), .A2(n12636), .ZN(n15722) );
  INV_X1 U14434 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18074) );
  XNOR2_X1 U14435 ( .A(n12637), .B(n18074), .ZN(n18076) );
  NAND2_X1 U14436 ( .A1(n12637), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12638) );
  XNOR2_X1 U14437 ( .A(n16013), .B(n12639), .ZN(n19281) );
  INV_X1 U14438 ( .A(n19281), .ZN(n12640) );
  INV_X1 U14439 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17935) );
  NAND2_X1 U14440 ( .A1(n12640), .A2(n17935), .ZN(n17636) );
  INV_X1 U14441 ( .A(n12642), .ZN(n12643) );
  NAND2_X1 U14442 ( .A1(n11336), .A2(n12643), .ZN(n12644) );
  NAND2_X1 U14443 ( .A1(n12650), .A2(n12644), .ZN(n19289) );
  NOR2_X1 U14444 ( .A1(n19289), .A2(n16007), .ZN(n12645) );
  NAND2_X1 U14445 ( .A1(n12645), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17620) );
  INV_X1 U14446 ( .A(n12645), .ZN(n12647) );
  INV_X1 U14447 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U14448 ( .A1(n12647), .A2(n12646), .ZN(n17619) );
  XNOR2_X1 U14449 ( .A(n12650), .B(n12649), .ZN(n17217) );
  AOI21_X1 U14450 ( .B1(n17217), .B2(n16014), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17609) );
  INV_X1 U14451 ( .A(n17609), .ZN(n12651) );
  NAND2_X1 U14452 ( .A1(n12653), .A2(n12652), .ZN(n12654) );
  NAND2_X1 U14453 ( .A1(n12660), .A2(n12654), .ZN(n15739) );
  NOR2_X1 U14454 ( .A1(n15739), .A2(n16007), .ZN(n12656) );
  INV_X1 U14455 ( .A(n12656), .ZN(n12655) );
  NAND2_X1 U14456 ( .A1(n12656), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17888) );
  INV_X1 U14457 ( .A(n17217), .ZN(n12657) );
  INV_X1 U14458 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17904) );
  OR3_X1 U14459 ( .A1(n12657), .A2(n16007), .A3(n17904), .ZN(n17886) );
  AND2_X1 U14460 ( .A1(n17888), .A2(n17886), .ZN(n12658) );
  XNOR2_X1 U14461 ( .A(n12660), .B(n12659), .ZN(n19300) );
  NAND2_X1 U14462 ( .A1(n19300), .A2(n16014), .ZN(n17602) );
  INV_X1 U14463 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12661) );
  XNOR2_X1 U14464 ( .A(n12663), .B(n12662), .ZN(n19314) );
  INV_X1 U14465 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17865) );
  OR3_X1 U14466 ( .A1(n19314), .A2(n16007), .A3(n17865), .ZN(n17594) );
  NAND2_X1 U14467 ( .A1(n11298), .A2(n11348), .ZN(n12664) );
  NAND2_X1 U14468 ( .A1(n11268), .A2(n12664), .ZN(n19340) );
  INV_X1 U14469 ( .A(n19340), .ZN(n12666) );
  INV_X1 U14470 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17824) );
  NOR2_X1 U14471 ( .A1(n16007), .A2(n17824), .ZN(n12665) );
  NAND2_X1 U14472 ( .A1(n12666), .A2(n12665), .ZN(n17561) );
  NAND2_X1 U14473 ( .A1(n12673), .A2(n12667), .ZN(n12668) );
  NAND2_X1 U14474 ( .A1(n11298), .A2(n12668), .ZN(n19328) );
  OR2_X1 U14475 ( .A1(n16007), .A2(n12811), .ZN(n12669) );
  OR2_X1 U14476 ( .A1(n19328), .A2(n12669), .ZN(n17559) );
  NAND2_X1 U14477 ( .A1(n12671), .A2(n12670), .ZN(n12672) );
  NAND2_X1 U14478 ( .A1(n12673), .A2(n12672), .ZN(n12679) );
  INV_X1 U14479 ( .A(n12679), .ZN(n15809) );
  NOR2_X1 U14480 ( .A1(n16007), .A2(n17847), .ZN(n12674) );
  NAND2_X1 U14481 ( .A1(n15809), .A2(n12674), .ZN(n17583) );
  AND2_X1 U14482 ( .A1(n17559), .A2(n17583), .ZN(n12675) );
  NAND2_X1 U14483 ( .A1(n17561), .A2(n12675), .ZN(n15964) );
  INV_X1 U14484 ( .A(n15964), .ZN(n12682) );
  OR2_X1 U14485 ( .A1(n19328), .A2(n16007), .ZN(n12676) );
  NAND2_X1 U14486 ( .A1(n12676), .A2(n12811), .ZN(n17560) );
  INV_X1 U14487 ( .A(n19314), .ZN(n12677) );
  NAND2_X1 U14488 ( .A1(n12677), .A2(n16014), .ZN(n12678) );
  NAND2_X1 U14489 ( .A1(n12678), .A2(n17865), .ZN(n17595) );
  OAI21_X1 U14490 ( .B1(n12679), .B2(n16007), .A(n17847), .ZN(n17584) );
  AND3_X1 U14491 ( .A1(n17560), .A2(n17595), .A3(n17584), .ZN(n12680) );
  OAI21_X1 U14492 ( .B1(n19340), .B2(n16007), .A(n17824), .ZN(n17562) );
  AND2_X1 U14493 ( .A1(n12680), .A2(n17562), .ZN(n15957) );
  INV_X1 U14494 ( .A(n15957), .ZN(n12681) );
  INV_X1 U14495 ( .A(n12683), .ZN(n12684) );
  NAND2_X1 U14496 ( .A1(n11268), .A2(n12684), .ZN(n12685) );
  NAND2_X1 U14497 ( .A1(n11304), .A2(n12685), .ZN(n19347) );
  INV_X1 U14498 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17797) );
  OAI21_X1 U14499 ( .B1(n19347), .B2(n16007), .A(n17797), .ZN(n12687) );
  OR2_X1 U14500 ( .A1(n16007), .A2(n17797), .ZN(n12686) );
  NAND2_X1 U14501 ( .A1(n11304), .A2(n12688), .ZN(n12689) );
  AND2_X1 U14502 ( .A1(n11291), .A2(n12689), .ZN(n17211) );
  INV_X1 U14503 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17544) );
  NOR2_X1 U14504 ( .A1(n16007), .A2(n17544), .ZN(n12690) );
  NAND2_X1 U14505 ( .A1(n17211), .A2(n12690), .ZN(n17533) );
  NAND2_X1 U14506 ( .A1(n17533), .A2(n17536), .ZN(n15965) );
  NAND2_X1 U14507 ( .A1(n17211), .A2(n16014), .ZN(n12691) );
  NAND2_X1 U14508 ( .A1(n12691), .A2(n17544), .ZN(n17534) );
  INV_X1 U14509 ( .A(n12692), .ZN(n12693) );
  XNOR2_X1 U14510 ( .A(n11291), .B(n12693), .ZN(n19362) );
  NOR2_X1 U14511 ( .A1(n16007), .A2(n12700), .ZN(n12694) );
  NAND2_X1 U14512 ( .A1(n19362), .A2(n12694), .ZN(n17527) );
  INV_X1 U14513 ( .A(n12695), .ZN(n12697) );
  XNOR2_X1 U14514 ( .A(n12697), .B(n12696), .ZN(n19383) );
  NAND2_X1 U14515 ( .A1(n19383), .A2(n16014), .ZN(n12699) );
  INV_X1 U14516 ( .A(n12699), .ZN(n12698) );
  INV_X1 U14517 ( .A(n15968), .ZN(n17511) );
  INV_X1 U14518 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17762) );
  NAND2_X1 U14519 ( .A1(n12699), .A2(n17762), .ZN(n17510) );
  NAND2_X1 U14520 ( .A1(n19362), .A2(n16014), .ZN(n12701) );
  NAND2_X1 U14521 ( .A1(n12701), .A2(n12700), .ZN(n17529) );
  NAND2_X1 U14522 ( .A1(n17510), .A2(n17529), .ZN(n15959) );
  INV_X1 U14523 ( .A(n12702), .ZN(n12705) );
  INV_X1 U14524 ( .A(n12703), .ZN(n12704) );
  NAND2_X1 U14525 ( .A1(n12705), .A2(n12704), .ZN(n12706) );
  NAND2_X1 U14526 ( .A1(n12711), .A2(n12706), .ZN(n19394) );
  INV_X1 U14527 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17753) );
  NAND2_X1 U14528 ( .A1(n12708), .A2(n12707), .ZN(n12709) );
  OAI21_X1 U14529 ( .B1(n17503), .B2(n17753), .A(n12709), .ZN(n12715) );
  NAND2_X1 U14530 ( .A1(n12711), .A2(n12710), .ZN(n12712) );
  AND2_X1 U14531 ( .A1(n15975), .A2(n12712), .ZN(n17200) );
  AOI21_X1 U14532 ( .B1(n17200), .B2(n16014), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15956) );
  INV_X1 U14533 ( .A(n17200), .ZN(n12714) );
  OR2_X1 U14534 ( .A1(n16007), .A2(n12851), .ZN(n12713) );
  NOR2_X1 U14535 ( .A1(n12714), .A2(n12713), .ZN(n15970) );
  XNOR2_X1 U14536 ( .A(n12715), .B(n11718), .ZN(n12870) );
  NOR2_X1 U14537 ( .A1(n12743), .A2(n11245), .ZN(n12716) );
  OR2_X1 U14538 ( .A1(n12762), .A2(n12716), .ZN(n12734) );
  NAND2_X1 U14539 ( .A1(n12718), .A2(n12717), .ZN(n12761) );
  AND2_X1 U14540 ( .A1(n12772), .A2(n12719), .ZN(n12759) );
  INV_X1 U14541 ( .A(n14653), .ZN(n12720) );
  AOI21_X1 U14542 ( .B1(n12720), .B2(n11259), .A(n12719), .ZN(n12730) );
  OAI21_X1 U14543 ( .B1(n12722), .B2(n12723), .A(n12721), .ZN(n12726) );
  INV_X1 U14544 ( .A(n12723), .ZN(n12756) );
  OAI211_X1 U14545 ( .C1(n11259), .C2(n12756), .A(n11590), .B(n12724), .ZN(
        n12725) );
  OAI211_X1 U14546 ( .C1(n12728), .C2(n12727), .A(n12726), .B(n12725), .ZN(
        n12729) );
  OAI21_X1 U14547 ( .B1(n12759), .B2(n12730), .A(n12729), .ZN(n12731) );
  AOI22_X1 U14548 ( .A1(n12761), .A2(n11245), .B1(n12732), .B2(n12731), .ZN(
        n12733) );
  NOR2_X1 U14549 ( .A1(n12734), .A2(n12733), .ZN(n12735) );
  MUX2_X1 U14550 ( .A(n19509), .B(n12735), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12738) );
  AND2_X1 U14551 ( .A1(n12762), .A2(n14653), .ZN(n12736) );
  NAND2_X1 U14552 ( .A1(n15764), .A2(n11259), .ZN(n15274) );
  NAND2_X1 U14553 ( .A1(n12737), .A2(n15334), .ZN(n12770) );
  OAI21_X1 U14554 ( .B1(n12738), .B2(n12045), .A(n12017), .ZN(n12739) );
  INV_X1 U14555 ( .A(n12739), .ZN(n12740) );
  NAND2_X1 U14556 ( .A1(n12740), .A2(n15274), .ZN(n12769) );
  NOR2_X1 U14557 ( .A1(n12773), .A2(n19264), .ZN(n12767) );
  NAND2_X1 U14558 ( .A1(n17957), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13926) );
  OAI21_X1 U14559 ( .B1(n13926), .B2(n11476), .A(n19509), .ZN(n15340) );
  INV_X1 U14560 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12741) );
  OAI21_X1 U14561 ( .B1(n13956), .B2(n15340), .A(n12741), .ZN(n18095) );
  AND3_X1 U14562 ( .A1(n12743), .A2(n12756), .A3(n12742), .ZN(n12744) );
  NOR2_X1 U14563 ( .A1(n15339), .A2(n12744), .ZN(n12745) );
  MUX2_X1 U14564 ( .A(n18095), .B(n12745), .S(n17948), .Z(n19568) );
  MUX2_X1 U14565 ( .A(n12058), .B(n12737), .S(n19264), .Z(n12746) );
  NAND2_X1 U14566 ( .A1(n12746), .A2(n22445), .ZN(n12765) );
  NAND2_X1 U14567 ( .A1(n12058), .A2(n15334), .ZN(n12747) );
  OR2_X1 U14568 ( .A1(n15339), .A2(n12747), .ZN(n12755) );
  NAND2_X1 U14569 ( .A1(n12825), .A2(n12046), .ZN(n12753) );
  NAND2_X1 U14570 ( .A1(n12748), .A2(n14548), .ZN(n12828) );
  OR2_X1 U14571 ( .A1(n12749), .A2(n12017), .ZN(n12826) );
  NAND2_X1 U14572 ( .A1(n12045), .A2(n11242), .ZN(n12750) );
  OAI211_X1 U14573 ( .C1(n12033), .C2(n11259), .A(n12046), .B(n12750), .ZN(
        n12751) );
  NAND4_X1 U14574 ( .A1(n12828), .A2(n12064), .A3(n12826), .A4(n12751), .ZN(
        n12752) );
  AOI21_X1 U14575 ( .B1(n12019), .B2(n12753), .A(n12752), .ZN(n12754) );
  AND2_X1 U14576 ( .A1(n12757), .A2(n12756), .ZN(n12758) );
  NOR2_X1 U14577 ( .A1(n12759), .A2(n12758), .ZN(n12760) );
  NOR2_X1 U14578 ( .A1(n12761), .A2(n12760), .ZN(n12763) );
  OR2_X1 U14579 ( .A1(n12763), .A2(n12762), .ZN(n15325) );
  INV_X1 U14580 ( .A(n15325), .ZN(n12764) );
  INV_X1 U14581 ( .A(n14548), .ZN(n19265) );
  NOR2_X1 U14582 ( .A1(n12773), .A2(n19265), .ZN(n15326) );
  NAND2_X1 U14583 ( .A1(n12764), .A2(n15326), .ZN(n12868) );
  OAI211_X1 U14584 ( .C1(n15339), .C2(n12765), .A(n15280), .B(n12868), .ZN(
        n12766) );
  AOI21_X1 U14585 ( .B1(n12767), .B2(n19568), .A(n12766), .ZN(n12768) );
  OAI211_X1 U14586 ( .C1(n15274), .C2(n12770), .A(n12769), .B(n12768), .ZN(
        n12771) );
  NOR2_X1 U14587 ( .A1(n12773), .A2(n12772), .ZN(n15324) );
  NAND2_X1 U14588 ( .A1(n12870), .A2(n19530), .ZN(n12867) );
  NOR2_X1 U14589 ( .A1(n19512), .A2(n14542), .ZN(n14541) );
  INV_X1 U14590 ( .A(n12776), .ZN(n12774) );
  NAND2_X1 U14591 ( .A1(n14541), .A2(n12774), .ZN(n12777) );
  NOR2_X1 U14592 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14542), .ZN(
        n12775) );
  XOR2_X1 U14593 ( .A(n12776), .B(n12775), .Z(n14643) );
  NAND2_X1 U14594 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14643), .ZN(
        n14642) );
  NAND2_X1 U14595 ( .A1(n12777), .A2(n14642), .ZN(n12780) );
  XOR2_X1 U14596 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12780), .Z(
        n14630) );
  XNOR2_X1 U14597 ( .A(n12779), .B(n12778), .ZN(n14628) );
  NAND2_X1 U14598 ( .A1(n14630), .A2(n14628), .ZN(n12782) );
  NAND2_X1 U14599 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12780), .ZN(
        n12781) );
  NAND2_X1 U14600 ( .A1(n12782), .A2(n12781), .ZN(n12783) );
  XNOR2_X1 U14601 ( .A(n12783), .B(n15624), .ZN(n15549) );
  NAND2_X1 U14602 ( .A1(n12783), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12784) );
  INV_X1 U14603 ( .A(n12785), .ZN(n12786) );
  XNOR2_X1 U14604 ( .A(n12787), .B(n12786), .ZN(n12789) );
  XNOR2_X1 U14605 ( .A(n12788), .B(n12789), .ZN(n15627) );
  INV_X1 U14606 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15834) );
  INV_X1 U14607 ( .A(n11240), .ZN(n12790) );
  NAND2_X1 U14608 ( .A1(n12790), .A2(n12789), .ZN(n12791) );
  NAND2_X2 U14609 ( .A1(n15629), .A2(n12791), .ZN(n12797) );
  INV_X1 U14610 ( .A(n12797), .ZN(n12793) );
  NAND2_X1 U14611 ( .A1(n12793), .A2(n12800), .ZN(n12794) );
  INV_X1 U14612 ( .A(n12795), .ZN(n12801) );
  INV_X1 U14613 ( .A(n12798), .ZN(n12799) );
  NAND2_X1 U14614 ( .A1(n12802), .A2(n12801), .ZN(n12803) );
  NAND2_X1 U14615 ( .A1(n12804), .A2(n16007), .ZN(n12805) );
  NAND2_X1 U14616 ( .A1(n12807), .A2(n12805), .ZN(n12806) );
  NAND2_X1 U14617 ( .A1(n12806), .A2(n17935), .ZN(n17631) );
  XNOR2_X1 U14618 ( .A(n12807), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17622) );
  INV_X1 U14619 ( .A(n12807), .ZN(n12808) );
  AND3_X1 U14620 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17836) );
  AND2_X1 U14621 ( .A1(n17836), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17848) );
  INV_X1 U14622 ( .A(n17848), .ZN(n12809) );
  NOR2_X1 U14623 ( .A1(n12809), .A2(n17847), .ZN(n12810) );
  NAND2_X1 U14624 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17749) );
  NOR3_X1 U14625 ( .A1(n17797), .A2(n17824), .A3(n17544), .ZN(n17747) );
  NAND2_X1 U14626 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17747), .ZN(
        n12812) );
  NOR2_X1 U14627 ( .A1(n17749), .A2(n12812), .ZN(n12849) );
  INV_X1 U14628 ( .A(n12849), .ZN(n12813) );
  NOR2_X1 U14629 ( .A1(n17795), .A2(n12813), .ZN(n17507) );
  AND2_X1 U14630 ( .A1(n12849), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12843) );
  INV_X1 U14631 ( .A(n12843), .ZN(n16030) );
  OAI21_X1 U14632 ( .B1(n17507), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n17500), .ZN(n12879) );
  OR2_X1 U14633 ( .A1(n17305), .A2(n12814), .ZN(n12815) );
  NAND2_X1 U14634 ( .A1(n17290), .A2(n12815), .ZN(n17297) );
  INV_X1 U14635 ( .A(n17297), .ZN(n12863) );
  NAND2_X1 U14636 ( .A1(n12817), .A2(n19264), .ZN(n12818) );
  NAND2_X1 U14637 ( .A1(n12818), .A2(n15261), .ZN(n12819) );
  NOR3_X1 U14638 ( .A1(n20322), .A2(n12737), .A3(n11259), .ZN(n12821) );
  AND2_X1 U14639 ( .A1(n11236), .A2(n12821), .ZN(n14122) );
  INV_X1 U14640 ( .A(n14122), .ZN(n15333) );
  INV_X1 U14641 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14844) );
  NOR2_X1 U14642 ( .A1(n19512), .A2(n14844), .ZN(n15564) );
  NOR2_X1 U14643 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15564), .ZN(
        n15565) );
  NOR3_X1 U14644 ( .A1(n15624), .A2(n15834), .A3(n15837), .ZN(n19524) );
  NAND2_X1 U14645 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19524), .ZN(
        n17916) );
  NAND2_X1 U14646 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17925) );
  NOR3_X1 U14647 ( .A1(n15565), .A2(n17916), .A3(n17925), .ZN(n12846) );
  INV_X1 U14648 ( .A(n12846), .ZN(n12822) );
  NAND2_X1 U14649 ( .A1(n19539), .A2(n12822), .ZN(n12824) );
  NAND2_X1 U14650 ( .A1(n12823), .A2(n19301), .ZN(n19513) );
  NAND2_X1 U14651 ( .A1(n12824), .A2(n19513), .ZN(n17744) );
  NAND3_X1 U14652 ( .A1(n12826), .A2(n11242), .A3(n12825), .ZN(n12827) );
  NAND2_X1 U14653 ( .A1(n12827), .A2(n11259), .ZN(n15298) );
  AOI21_X1 U14654 ( .B1(n15298), .B2(n12828), .A(n11588), .ZN(n12836) );
  INV_X1 U14655 ( .A(n12829), .ZN(n14540) );
  NAND2_X1 U14656 ( .A1(n12064), .A2(n12014), .ZN(n12830) );
  AOI22_X1 U14657 ( .A1(n14540), .A2(n12830), .B1(n12045), .B2(n12737), .ZN(
        n12834) );
  NAND2_X1 U14658 ( .A1(n12833), .A2(n12832), .ZN(n14123) );
  NAND3_X1 U14659 ( .A1(n12834), .A2(n12831), .A3(n14123), .ZN(n12835) );
  NOR2_X1 U14660 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  OAI21_X1 U14661 ( .B1(n12838), .B2(n12064), .A(n12837), .ZN(n15304) );
  OR2_X1 U14662 ( .A1(n15304), .A2(n14148), .ZN(n12839) );
  INV_X1 U14663 ( .A(n17919), .ZN(n12840) );
  NAND2_X1 U14664 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15564), .ZN(
        n15561) );
  OR2_X1 U14665 ( .A1(n17916), .A2(n15561), .ZN(n17918) );
  NOR2_X1 U14666 ( .A1(n17925), .A2(n17918), .ZN(n17785) );
  NOR2_X1 U14667 ( .A1(n12840), .A2(n17785), .ZN(n12841) );
  OR2_X1 U14668 ( .A1(n17744), .A2(n12841), .ZN(n17875) );
  INV_X1 U14669 ( .A(n19521), .ZN(n17834) );
  OR2_X1 U14670 ( .A1(n17875), .A2(n17834), .ZN(n17685) );
  AND2_X1 U14671 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12842) );
  AND2_X1 U14672 ( .A1(n17848), .A2(n12842), .ZN(n17784) );
  NAND2_X1 U14673 ( .A1(n12843), .A2(n17784), .ZN(n12844) );
  OR2_X1 U14674 ( .A1(n17875), .A2(n12844), .ZN(n12845) );
  NAND2_X1 U14675 ( .A1(n17685), .A2(n12845), .ZN(n17732) );
  INV_X2 U14676 ( .A(n19301), .ZN(n19526) );
  NAND2_X1 U14677 ( .A1(n19526), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12873) );
  NAND2_X1 U14678 ( .A1(n19539), .A2(n12846), .ZN(n12848) );
  NAND2_X1 U14679 ( .A1(n17919), .A2(n17785), .ZN(n12847) );
  NAND2_X1 U14680 ( .A1(n12848), .A2(n12847), .ZN(n17877) );
  NAND2_X1 U14681 ( .A1(n17877), .A2(n17784), .ZN(n17794) );
  INV_X1 U14682 ( .A(n17794), .ZN(n17822) );
  NAND3_X1 U14683 ( .A1(n17822), .A2(n12849), .A3(n12851), .ZN(n12850) );
  OAI211_X1 U14684 ( .C1(n17732), .C2(n12851), .A(n12873), .B(n12850), .ZN(
        n12862) );
  INV_X1 U14685 ( .A(n17372), .ZN(n12854) );
  NAND2_X1 U14686 ( .A1(n17391), .A2(n12852), .ZN(n12853) );
  NAND2_X1 U14687 ( .A1(n12854), .A2(n12853), .ZN(n17385) );
  INV_X1 U14688 ( .A(n12855), .ZN(n12856) );
  AND2_X1 U14689 ( .A1(n11236), .A2(n12856), .ZN(n15330) );
  INV_X1 U14690 ( .A(n15330), .ZN(n15263) );
  NAND2_X1 U14691 ( .A1(n12857), .A2(n12019), .ZN(n15337) );
  NAND2_X1 U14692 ( .A1(n15337), .A2(n11259), .ZN(n12858) );
  NAND2_X1 U14693 ( .A1(n15263), .A2(n12858), .ZN(n12859) );
  NOR2_X1 U14694 ( .A1(n17385), .A2(n19542), .ZN(n12861) );
  AOI211_X1 U14695 ( .C1(n12863), .C2(n19550), .A(n12862), .B(n12861), .ZN(
        n12864) );
  NAND2_X1 U14696 ( .A1(n12867), .A2(n12866), .ZN(P2_U3025) );
  NAND2_X1 U14697 ( .A1(n19568), .A2(n15324), .ZN(n12869) );
  NAND2_X1 U14698 ( .A1(n12869), .A2(n12868), .ZN(n15345) );
  NAND2_X1 U14699 ( .A1(n12870), .A2(n18089), .ZN(n12882) );
  NAND2_X1 U14700 ( .A1(n20162), .A2(n18096), .ZN(n19273) );
  OR2_X1 U14701 ( .A1(n19273), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12871) );
  NAND2_X1 U14702 ( .A1(n22410), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12872) );
  NAND2_X1 U14703 ( .A1(n15765), .A2(n12872), .ZN(n14544) );
  OAI21_X1 U14704 ( .B1(n18093), .B2(n12874), .A(n12873), .ZN(n12877) );
  AND2_X1 U14705 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12875) );
  NOR2_X1 U14706 ( .A1(n17297), .A2(n17641), .ZN(n12876) );
  AOI211_X1 U14707 ( .C1(n18083), .C2(n17194), .A(n12877), .B(n12876), .ZN(
        n12878) );
  NAND2_X1 U14708 ( .A1(n12882), .A2(n12881), .ZN(P2_U2993) );
  AND2_X2 U14709 ( .A1(n12887), .A2(n14823), .ZN(n13434) );
  AND2_X2 U14710 ( .A1(n12885), .A2(n14818), .ZN(n13127) );
  AOI22_X1 U14711 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13759), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12884) );
  AND2_X2 U14712 ( .A1(n17162), .A2(n14823), .ZN(n13523) );
  AOI22_X1 U14713 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13034), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12883) );
  AND2_X2 U14714 ( .A1(n14823), .A2(n12885), .ZN(n12951) );
  AOI22_X1 U14715 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U14717 ( .A1(n13069), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12966), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U14718 ( .A1(n13027), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U14719 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U14720 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13034), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U14721 ( .A1(n13376), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U14722 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U14723 ( .A1(n13069), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12966), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U14724 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U14725 ( .A1(n13027), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U14726 ( .A1(n12900), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U14727 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12904) );
  AOI22_X1 U14728 ( .A1(n12900), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U14729 ( .A1(n13069), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12966), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U14730 ( .A1(n13027), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U14731 ( .A1(n13376), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U14732 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U14733 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U14734 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13034), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U14735 ( .A1(n13069), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13027), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U14736 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12912) );
  AOI22_X1 U14737 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U14738 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13034), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12910) );
  NAND4_X1 U14739 ( .A1(n12913), .A2(n12912), .A3(n12911), .A4(n12910), .ZN(
        n12919) );
  AOI22_X1 U14740 ( .A1(n13376), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U14741 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U14742 ( .A1(n12900), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12966), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U14743 ( .A1(n13028), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12914) );
  NAND4_X1 U14744 ( .A1(n12917), .A2(n12916), .A3(n12915), .A4(n12914), .ZN(
        n12918) );
  AOI21_X1 U14745 ( .B1(n14674), .B2(n14786), .A(n16741), .ZN(n12941) );
  AOI22_X1 U14746 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U14747 ( .A1(n12951), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U14748 ( .A1(n13027), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U14749 ( .A1(n13376), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U14750 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12900), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U14751 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U14752 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13034), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12924) );
  NAND2_X1 U14753 ( .A1(n12930), .A2(n12929), .ZN(n12940) );
  AOI22_X1 U14754 ( .A1(n12900), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13027), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U14755 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U14756 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13034), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U14757 ( .A1(n13069), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U14758 ( .A1(n13376), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U14759 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U14760 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12966), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U14761 ( .A1(n13028), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12936) );
  NAND2_X2 U14762 ( .A1(n11721), .A2(n11724), .ZN(n14206) );
  NAND2_X1 U14763 ( .A1(n13293), .A2(n14206), .ZN(n12993) );
  NAND2_X1 U14764 ( .A1(n13069), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12946) );
  NAND2_X1 U14765 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12945) );
  BUF_X8 U14766 ( .A(n12942), .Z(n13758) );
  NAND2_X1 U14767 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12944) );
  NAND2_X1 U14768 ( .A1(n12900), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12943) );
  NAND2_X1 U14769 ( .A1(n13376), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12950) );
  NAND2_X1 U14770 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12949) );
  NAND2_X1 U14771 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12948) );
  NAND2_X1 U14772 ( .A1(n13754), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12947) );
  NAND2_X1 U14773 ( .A1(n13027), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12955) );
  BUF_X4 U14774 ( .A(n12951), .Z(n13769) );
  NAND2_X1 U14775 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12954) );
  NAND2_X1 U14776 ( .A1(n13028), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12953) );
  NAND2_X1 U14777 ( .A1(n13033), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12952) );
  NAND2_X1 U14778 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12960) );
  NAND2_X1 U14779 ( .A1(n13759), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12959) );
  NAND2_X1 U14780 ( .A1(n12966), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12958) );
  NAND2_X1 U14781 ( .A1(n13034), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12957) );
  NOR2_X2 U14782 ( .A1(n12998), .A2(n12965), .ZN(n14198) );
  AOI22_X1 U14783 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U14784 ( .A1(n12900), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13028), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U14785 ( .A1(n13069), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12966), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U14786 ( .A1(n13027), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U14787 ( .A1(n13376), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U14788 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U14789 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U14790 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13034), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12971) );
  AND2_X2 U14791 ( .A1(n15025), .A2(n14206), .ZN(n14686) );
  NOR2_X1 U14792 ( .A1(n14772), .A2(n14771), .ZN(n12975) );
  NAND2_X1 U14793 ( .A1(n14696), .A2(n16494), .ZN(n12976) );
  NAND2_X1 U14794 ( .A1(n22433), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22422) );
  NAND2_X1 U14795 ( .A1(n22437), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n12977) );
  NOR2_X2 U14796 ( .A1(n14784), .A2(n12982), .ZN(n14706) );
  NOR2_X2 U14797 ( .A1(n14206), .A2(n14786), .ZN(n14819) );
  NAND3_X1 U14798 ( .A1(n14706), .A2(n15016), .A3(n14819), .ZN(n14682) );
  NAND2_X1 U14799 ( .A1(n14777), .A2(n14772), .ZN(n14780) );
  AND2_X1 U14800 ( .A1(n12980), .A2(n14777), .ZN(n13295) );
  NAND2_X1 U14801 ( .A1(n13295), .A2(n12981), .ZN(n12985) );
  AND2_X2 U14802 ( .A1(n14986), .A2(n11244), .ZN(n14721) );
  NAND2_X1 U14803 ( .A1(n12985), .A2(n14721), .ZN(n12984) );
  NAND2_X1 U14804 ( .A1(n13044), .A2(n14784), .ZN(n16690) );
  INV_X1 U14805 ( .A(n12985), .ZN(n12986) );
  INV_X1 U14806 ( .A(n13293), .ZN(n14671) );
  NAND2_X1 U14807 ( .A1(n12986), .A2(n13293), .ZN(n14673) );
  NAND2_X1 U14808 ( .A1(n14771), .A2(n14777), .ZN(n12987) );
  NAND2_X1 U14809 ( .A1(n14673), .A2(n14758), .ZN(n13000) );
  INV_X1 U14810 ( .A(n14819), .ZN(n14677) );
  INV_X1 U14811 ( .A(n14686), .ZN(n12988) );
  NAND2_X1 U14812 ( .A1(n17977), .A2(n22392), .ZN(n13789) );
  INV_X1 U14813 ( .A(n13789), .ZN(n13084) );
  XNOR2_X1 U14814 ( .A(n22567), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15491) );
  NAND2_X1 U14815 ( .A1(n13084), .A2(n15491), .ZN(n12989) );
  INV_X1 U14816 ( .A(n13292), .ZN(n18046) );
  NAND2_X1 U14817 ( .A1(n18046), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13061) );
  AND2_X1 U14818 ( .A1(n12989), .A2(n13061), .ZN(n12990) );
  MUX2_X1 U14819 ( .A(n13789), .B(n13292), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n12992) );
  INV_X1 U14820 ( .A(n12993), .ZN(n12996) );
  INV_X1 U14821 ( .A(n14706), .ZN(n16688) );
  NAND2_X1 U14822 ( .A1(n16688), .A2(n14293), .ZN(n14610) );
  NAND2_X1 U14823 ( .A1(n17977), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12994) );
  AOI21_X1 U14824 ( .B1(n14786), .B2(n11243), .A(n12994), .ZN(n12995) );
  NAND2_X1 U14825 ( .A1(n14819), .A2(n15033), .ZN(n14800) );
  OAI211_X1 U14826 ( .C1(n12996), .C2(n14610), .A(n12995), .B(n14800), .ZN(
        n12997) );
  NOR2_X1 U14827 ( .A1(n11166), .A2(n12997), .ZN(n12999) );
  NAND2_X1 U14828 ( .A1(n12998), .A2(n14706), .ZN(n14680) );
  AOI22_X1 U14829 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U14830 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13756), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U14831 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13003) );
  INV_X1 U14832 ( .A(n13033), .ZN(n13091) );
  AOI22_X1 U14833 ( .A1(n13757), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13002) );
  NAND4_X1 U14834 ( .A1(n13005), .A2(n13004), .A3(n13003), .A4(n13002), .ZN(
        n13011) );
  AOI22_X1 U14835 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13009) );
  AOI22_X1 U14836 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U14837 ( .A1(n13759), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U14838 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13006) );
  NAND4_X1 U14839 ( .A1(n13009), .A2(n13008), .A3(n13007), .A4(n13006), .ZN(
        n13010) );
  NAND2_X1 U14840 ( .A1(n13050), .A2(n13158), .ZN(n13012) );
  AOI22_X1 U14841 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13016) );
  AOI22_X1 U14842 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13015) );
  AOI22_X1 U14843 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U14844 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13013) );
  NAND4_X1 U14845 ( .A1(n13016), .A2(n13015), .A3(n13014), .A4(n13013), .ZN(
        n13022) );
  AOI22_X1 U14846 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U14847 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13019) );
  AOI22_X1 U14848 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U14849 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13017) );
  NAND4_X1 U14850 ( .A1(n13020), .A2(n13019), .A3(n13018), .A4(n13017), .ZN(
        n13021) );
  NOR2_X1 U14851 ( .A1(n11243), .A2(n22392), .ZN(n13023) );
  AOI22_X1 U14852 ( .A1(n13050), .A2(n13046), .B1(n13023), .B2(n13158), .ZN(
        n13025) );
  NAND2_X1 U14853 ( .A1(n13283), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13024) );
  AOI22_X1 U14854 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U14855 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U14856 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U14857 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13029) );
  NAND4_X1 U14858 ( .A1(n13032), .A2(n13031), .A3(n13030), .A4(n13029), .ZN(
        n13040) );
  AOI22_X1 U14859 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U14860 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U14861 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U14862 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13035) );
  NAND4_X1 U14863 ( .A1(n13038), .A2(n13037), .A3(n13036), .A4(n13035), .ZN(
        n13039) );
  XNOR2_X1 U14864 ( .A(n13046), .B(n13157), .ZN(n13041) );
  NAND2_X1 U14865 ( .A1(n13041), .A2(n13050), .ZN(n13042) );
  NAND2_X1 U14866 ( .A1(n13283), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13049) );
  NAND2_X1 U14867 ( .A1(n13044), .A2(n13157), .ZN(n13045) );
  OAI211_X1 U14868 ( .C1(n13046), .C2(n14771), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n13045), .ZN(n13047) );
  INV_X1 U14869 ( .A(n13047), .ZN(n13048) );
  NAND2_X1 U14870 ( .A1(n13055), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13060) );
  AND2_X1 U14871 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13056) );
  NAND2_X1 U14872 ( .A1(n13056), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15060) );
  INV_X1 U14873 ( .A(n13056), .ZN(n13057) );
  NAND2_X1 U14874 ( .A1(n13057), .A2(n22552), .ZN(n13058) );
  AOI22_X1 U14875 ( .A1(n15399), .A2(n13084), .B1(n18046), .B2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13059) );
  INV_X1 U14876 ( .A(n13061), .ZN(n13063) );
  OAI21_X1 U14877 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13063), .A(
        n13062), .ZN(n13064) );
  OAI21_X2 U14878 ( .B1(n13067), .B2(n13066), .A(n17974), .ZN(n17159) );
  AOI22_X1 U14879 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U14880 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13434), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U14881 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U14882 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13070) );
  NAND4_X1 U14883 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13079) );
  AOI22_X1 U14884 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U14885 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U14886 ( .A1(n12942), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U14887 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13074) );
  NAND4_X1 U14888 ( .A1(n13077), .A2(n13076), .A3(n13075), .A4(n13074), .ZN(
        n13078) );
  AOI22_X1 U14889 ( .A1(n13283), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13288), .B2(n13159), .ZN(n13080) );
  NAND2_X1 U14890 ( .A1(n13055), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13086) );
  INV_X1 U14891 ( .A(n15060), .ZN(n13081) );
  NAND2_X1 U14892 ( .A1(n13081), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22840) );
  NAND2_X1 U14893 ( .A1(n15060), .A2(n22553), .ZN(n13082) );
  NOR2_X1 U14894 ( .A1(n13292), .A2(n22553), .ZN(n13083) );
  AOI21_X1 U14895 ( .B1(n15437), .B2(n13084), .A(n13083), .ZN(n13085) );
  AOI22_X1 U14896 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U14897 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U14898 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U14899 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13087) );
  NAND4_X1 U14900 ( .A1(n13090), .A2(n13089), .A3(n13088), .A4(n13087), .ZN(
        n13097) );
  AOI22_X1 U14901 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U14902 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U14903 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U14904 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13092) );
  NAND4_X1 U14905 ( .A1(n13095), .A2(n13094), .A3(n13093), .A4(n13092), .ZN(
        n13096) );
  AOI22_X1 U14906 ( .A1(n13283), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13288), .B2(n13170), .ZN(n13098) );
  AOI22_X1 U14907 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U14908 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13734), .B1(
        n13755), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U14909 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n13767), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U14910 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13766), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13101) );
  NAND4_X1 U14911 ( .A1(n13104), .A2(n13103), .A3(n13102), .A4(n13101), .ZN(
        n13110) );
  AOI22_X1 U14912 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13756), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13108) );
  AOI22_X1 U14913 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U14914 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U14915 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13105) );
  NAND4_X1 U14916 ( .A1(n13108), .A2(n13107), .A3(n13106), .A4(n13105), .ZN(
        n13109) );
  AOI22_X1 U14917 ( .A1(n13283), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13288), .B2(n13186), .ZN(n13175) );
  AOI22_X1 U14918 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U14919 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13127), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U14920 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U14921 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13113) );
  NAND4_X1 U14922 ( .A1(n13116), .A2(n13115), .A3(n13114), .A4(n13113), .ZN(
        n13122) );
  AOI22_X1 U14923 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U14924 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U14925 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U14926 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13117) );
  NAND4_X1 U14927 ( .A1(n13120), .A2(n13119), .A3(n13118), .A4(n13117), .ZN(
        n13121) );
  AOI22_X1 U14928 ( .A1(n13283), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13288), .B2(n13189), .ZN(n13183) );
  AOI22_X1 U14929 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13126) );
  AOI22_X1 U14930 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13125) );
  AOI22_X1 U14931 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U14932 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13123) );
  NAND4_X1 U14933 ( .A1(n13126), .A2(n13125), .A3(n13124), .A4(n13123), .ZN(
        n13133) );
  AOI22_X1 U14934 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U14935 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U14936 ( .A1(n13759), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U14937 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13128) );
  NAND4_X1 U14938 ( .A1(n13131), .A2(n13130), .A3(n13129), .A4(n13128), .ZN(
        n13132) );
  AOI22_X1 U14939 ( .A1(n13283), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13288), .B2(n13208), .ZN(n13194) );
  INV_X1 U14940 ( .A(n13194), .ZN(n13134) );
  INV_X1 U14941 ( .A(n13135), .ZN(n13136) );
  OAI21_X1 U14942 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n17134), .ZN(n13234) );
  INV_X1 U14943 ( .A(n13234), .ZN(n13139) );
  INV_X1 U14944 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16995) );
  NAND2_X1 U14945 ( .A1(n11160), .A2(n16995), .ZN(n13233) );
  INV_X1 U14946 ( .A(n13233), .ZN(n13138) );
  INV_X1 U14947 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16987) );
  NAND2_X1 U14948 ( .A1(n13053), .A2(n13243), .ZN(n13143) );
  XNOR2_X1 U14949 ( .A(n13158), .B(n13157), .ZN(n13140) );
  INV_X1 U14950 ( .A(n14721), .ZN(n22109) );
  OAI211_X1 U14951 ( .C1(n13140), .C2(n22109), .A(n14686), .B(n14770), .ZN(
        n13141) );
  INV_X1 U14952 ( .A(n13141), .ZN(n13142) );
  NAND2_X1 U14953 ( .A1(n13143), .A2(n13142), .ZN(n13148) );
  NAND2_X1 U14954 ( .A1(n13044), .A2(n14206), .ZN(n13161) );
  OAI21_X1 U14955 ( .B1(n22109), .B2(n13157), .A(n13161), .ZN(n13146) );
  INV_X1 U14956 ( .A(n13146), .ZN(n13147) );
  OR2_X1 U14957 ( .A1(n14857), .A2(n11161), .ZN(n13149) );
  INV_X1 U14958 ( .A(n13151), .ZN(n13152) );
  NAND2_X1 U14959 ( .A1(n13153), .A2(n13152), .ZN(n13154) );
  INV_X1 U14960 ( .A(n13159), .ZN(n13156) );
  NAND2_X1 U14961 ( .A1(n13158), .A2(n13157), .ZN(n13155) );
  NAND2_X1 U14962 ( .A1(n13156), .A2(n13155), .ZN(n13169) );
  NAND3_X1 U14963 ( .A1(n13159), .A2(n13158), .A3(n13157), .ZN(n13160) );
  NAND2_X1 U14964 ( .A1(n13169), .A2(n13160), .ZN(n13163) );
  INV_X1 U14965 ( .A(n13161), .ZN(n13162) );
  AOI21_X1 U14966 ( .B1(n13163), .B2(n14721), .A(n13162), .ZN(n13164) );
  NAND2_X1 U14967 ( .A1(n13165), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13166) );
  INV_X1 U14968 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14216) );
  NAND2_X1 U14969 ( .A1(n13167), .A2(n13100), .ZN(n13168) );
  OR2_X1 U14970 ( .A1(n15196), .A2(n13258), .ZN(n13172) );
  NAND2_X1 U14971 ( .A1(n13169), .A2(n13170), .ZN(n13188) );
  OAI211_X1 U14972 ( .C1(n13170), .C2(n13169), .A(n13188), .B(n14721), .ZN(
        n13171) );
  NAND2_X1 U14973 ( .A1(n13172), .A2(n13171), .ZN(n15379) );
  NAND2_X1 U14974 ( .A1(n13173), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13174) );
  XNOR2_X1 U14975 ( .A(n13188), .B(n13186), .ZN(n13177) );
  NAND2_X1 U14976 ( .A1(n13177), .A2(n14721), .ZN(n13178) );
  INV_X1 U14977 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13179) );
  NAND2_X1 U14978 ( .A1(n15360), .A2(n15359), .ZN(n13182) );
  NAND2_X1 U14979 ( .A1(n13180), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13181) );
  NAND2_X1 U14980 ( .A1(n13184), .A2(n13183), .ZN(n13185) );
  NAND2_X1 U14981 ( .A1(n13195), .A2(n13185), .ZN(n13344) );
  INV_X1 U14982 ( .A(n13186), .ZN(n13187) );
  NOR2_X1 U14983 ( .A1(n13188), .A2(n13187), .ZN(n13190) );
  NAND2_X1 U14984 ( .A1(n13190), .A2(n13189), .ZN(n13207) );
  OAI211_X1 U14985 ( .C1(n13190), .C2(n13189), .A(n13207), .B(n14721), .ZN(
        n13191) );
  INV_X1 U14986 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15477) );
  XNOR2_X1 U14987 ( .A(n13192), .B(n15477), .ZN(n15473) );
  NAND2_X1 U14988 ( .A1(n13192), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13193) );
  NAND2_X1 U14989 ( .A1(n13195), .A2(n13194), .ZN(n13350) );
  NAND3_X1 U14990 ( .A1(n13196), .A2(n13243), .A3(n13350), .ZN(n13199) );
  XNOR2_X1 U14991 ( .A(n13207), .B(n13208), .ZN(n13197) );
  NAND2_X1 U14992 ( .A1(n13197), .A2(n14721), .ZN(n13198) );
  NAND2_X1 U14993 ( .A1(n13199), .A2(n13198), .ZN(n13200) );
  INV_X1 U14994 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15786) );
  INV_X1 U14995 ( .A(n13283), .ZN(n13204) );
  INV_X1 U14996 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13203) );
  NAND2_X1 U14997 ( .A1(n13288), .A2(n13216), .ZN(n13202) );
  OAI21_X1 U14998 ( .B1(n13204), .B2(n13203), .A(n13202), .ZN(n13205) );
  INV_X1 U14999 ( .A(n13359), .ZN(n13206) );
  OR2_X1 U15000 ( .A1(n13206), .A2(n13258), .ZN(n13212) );
  INV_X1 U15001 ( .A(n13207), .ZN(n13209) );
  NAND2_X1 U15002 ( .A1(n13209), .A2(n13208), .ZN(n13215) );
  XNOR2_X1 U15003 ( .A(n13215), .B(n13216), .ZN(n13210) );
  NAND2_X1 U15004 ( .A1(n13210), .A2(n14721), .ZN(n13211) );
  NAND2_X1 U15005 ( .A1(n13212), .A2(n13211), .ZN(n13213) );
  INV_X1 U15006 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15647) );
  XNOR2_X1 U15007 ( .A(n13213), .B(n15647), .ZN(n15671) );
  NAND2_X1 U15008 ( .A1(n13213), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13214) );
  INV_X1 U15009 ( .A(n13215), .ZN(n13217) );
  NAND3_X1 U15010 ( .A1(n13217), .A2(n14721), .A3(n13216), .ZN(n13218) );
  NAND2_X1 U15011 ( .A1(n13229), .A2(n13218), .ZN(n13219) );
  INV_X1 U15012 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15648) );
  XNOR2_X1 U15013 ( .A(n13219), .B(n15648), .ZN(n15643) );
  XNOR2_X1 U15014 ( .A(n11160), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15785) );
  INV_X1 U15015 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17144) );
  OR2_X1 U15016 ( .A1(n13229), .A2(n17144), .ZN(n13220) );
  INV_X1 U15017 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n22138) );
  NAND2_X1 U15018 ( .A1(n13229), .A2(n22138), .ZN(n13221) );
  INV_X1 U15019 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16970) );
  NAND3_X1 U15020 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13222) );
  AND2_X1 U15021 ( .A1(n13229), .A2(n13222), .ZN(n13223) );
  NOR2_X1 U15022 ( .A1(n16944), .A2(n13223), .ZN(n17089) );
  NAND2_X1 U15023 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n22178) );
  INV_X1 U15024 ( .A(n22178), .ZN(n13224) );
  NAND2_X1 U15025 ( .A1(n13224), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n22168) );
  INV_X1 U15026 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n22134) );
  OR2_X1 U15027 ( .A1(n13229), .A2(n22134), .ZN(n13225) );
  NAND2_X1 U15028 ( .A1(n16945), .A2(n13225), .ZN(n17093) );
  NOR2_X1 U15029 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16955) );
  AND2_X1 U15030 ( .A1(n16955), .A2(n16970), .ZN(n13226) );
  INV_X1 U15031 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17098) );
  INV_X1 U15032 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14256) );
  INV_X1 U15033 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17108) );
  AND3_X1 U15034 ( .A1(n17098), .A2(n14256), .A3(n17108), .ZN(n13227) );
  NOR2_X1 U15035 ( .A1(n11160), .A2(n13227), .ZN(n13228) );
  NAND3_X1 U15036 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16975) );
  INV_X1 U15037 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16915) );
  INV_X2 U15038 ( .A(n13229), .ZN(n17134) );
  INV_X1 U15039 ( .A(n16914), .ZN(n13232) );
  NOR4_X1 U15040 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13231) );
  NOR3_X1 U15041 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16858) );
  AND2_X1 U15042 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16984) );
  AOI21_X1 U15043 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16984), .A(
        n17134), .ZN(n16856) );
  NAND2_X1 U15044 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17004) );
  NOR2_X1 U15045 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17014) );
  XNOR2_X1 U15046 ( .A(n11160), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13235) );
  NAND2_X1 U15047 ( .A1(n15199), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13238) );
  NAND2_X1 U15048 ( .A1(n13236), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13237) );
  NAND2_X1 U15049 ( .A1(n13238), .A2(n13237), .ZN(n13252) );
  NAND2_X1 U15050 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n22567), .ZN(
        n13259) );
  NAND2_X1 U15051 ( .A1(n13254), .A2(n13238), .ZN(n13274) );
  NAND2_X1 U15052 ( .A1(n22552), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13241) );
  NAND2_X1 U15053 ( .A1(n14688), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13239) );
  NAND2_X1 U15054 ( .A1(n13241), .A2(n13239), .ZN(n13273) );
  INV_X1 U15055 ( .A(n13273), .ZN(n13240) );
  NAND2_X1 U15056 ( .A1(n13274), .A2(n13240), .ZN(n13242) );
  NAND2_X1 U15057 ( .A1(n13242), .A2(n13241), .ZN(n13247) );
  XNOR2_X1 U15058 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13246) );
  OAI222_X1 U15059 ( .A1(n18038), .A2(n13244), .B1(n18038), .B2(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n13244), .C2(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n13289) );
  INV_X1 U15060 ( .A(n13289), .ZN(n14197) );
  NAND2_X1 U15061 ( .A1(n13283), .A2(n13243), .ZN(n13287) );
  NAND2_X1 U15062 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13244), .ZN(
        n13245) );
  NOR2_X1 U15063 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  OR2_X1 U15064 ( .A1(n13249), .A2(n13248), .ZN(n13250) );
  INV_X1 U15065 ( .A(n13287), .ZN(n13264) );
  OAI21_X1 U15066 ( .B1(n13251), .B2(n13250), .A(n13264), .ZN(n13285) );
  NOR2_X1 U15067 ( .A1(n13251), .A2(n13250), .ZN(n14192) );
  INV_X1 U15068 ( .A(n13288), .ZN(n13256) );
  NAND2_X1 U15069 ( .A1(n13252), .A2(n13259), .ZN(n13253) );
  NOR2_X1 U15070 ( .A1(n14770), .A2(n22392), .ZN(n13266) );
  INV_X1 U15071 ( .A(n13266), .ZN(n13255) );
  OAI211_X1 U15072 ( .C1(n13256), .C2(n14986), .A(n14195), .B(n13255), .ZN(
        n13272) );
  INV_X1 U15073 ( .A(n14195), .ZN(n13257) );
  OAI21_X1 U15074 ( .B1(n13288), .B2(n13258), .A(n13257), .ZN(n13271) );
  INV_X1 U15075 ( .A(n14674), .ZN(n13263) );
  INV_X1 U15076 ( .A(n13259), .ZN(n13260) );
  AOI21_X1 U15077 ( .B1(n14761), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n13260), .ZN(n13265) );
  INV_X1 U15078 ( .A(n13265), .ZN(n13262) );
  NAND2_X1 U15079 ( .A1(n14986), .A2(n14770), .ZN(n13261) );
  NAND2_X1 U15080 ( .A1(n16688), .A2(n13261), .ZN(n13276) );
  AOI211_X1 U15081 ( .C1(n13263), .C2(n11244), .A(n13262), .B(n13276), .ZN(
        n13269) );
  AOI21_X1 U15082 ( .B1(n13288), .B2(n13265), .A(n13264), .ZN(n13268) );
  NOR3_X1 U15083 ( .A1(n13266), .A2(n14195), .A3(n14784), .ZN(n13267) );
  NOR3_X1 U15084 ( .A1(n13269), .A2(n13268), .A3(n13267), .ZN(n13270) );
  AOI21_X1 U15085 ( .B1(n13272), .B2(n13271), .A(n13270), .ZN(n13281) );
  XNOR2_X1 U15086 ( .A(n13274), .B(n13273), .ZN(n14193) );
  INV_X1 U15087 ( .A(n14193), .ZN(n13275) );
  AOI211_X1 U15088 ( .C1(n13283), .C2(n13275), .A(n13277), .B(n13276), .ZN(
        n13280) );
  INV_X1 U15089 ( .A(n13276), .ZN(n13279) );
  INV_X1 U15090 ( .A(n13277), .ZN(n13278) );
  OAI22_X1 U15091 ( .A1(n13281), .A2(n13280), .B1(n13279), .B2(n13278), .ZN(
        n13282) );
  OAI21_X1 U15092 ( .B1(n13283), .B2(n14192), .A(n13282), .ZN(n13284) );
  OAI211_X1 U15093 ( .C1(P1_STATE2_REG_0__SCAN_IN), .C2(n18038), .A(n13285), 
        .B(n13284), .ZN(n13286) );
  NAND2_X1 U15094 ( .A1(n13289), .A2(n13288), .ZN(n13290) );
  OR2_X1 U15095 ( .A1(n13293), .A2(n14771), .ZN(n13294) );
  AND2_X1 U15096 ( .A1(n13295), .A2(n13294), .ZN(n14669) );
  NAND2_X1 U15097 ( .A1(n14758), .A2(n13044), .ZN(n13296) );
  NAND3_X1 U15098 ( .A1(n14669), .A2(n14686), .A3(n13296), .ZN(n14699) );
  NAND2_X1 U15099 ( .A1(n12978), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13332) );
  XNOR2_X1 U15100 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n22231) );
  AOI21_X1 U15101 ( .B1(n13782), .B2(n22231), .A(n13786), .ZN(n13298) );
  NAND2_X1 U15102 ( .A1(n13781), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13297) );
  OAI211_X1 U15103 ( .C1(n13332), .C2(n14688), .A(n13298), .B(n13297), .ZN(
        n13299) );
  INV_X1 U15104 ( .A(n13299), .ZN(n13300) );
  NAND2_X1 U15105 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13320) );
  INV_X1 U15106 ( .A(n13302), .ZN(n13305) );
  INV_X1 U15107 ( .A(n13303), .ZN(n13304) );
  XNOR2_X1 U15108 ( .A(n13305), .B(n13304), .ZN(n14936) );
  NAND2_X1 U15109 ( .A1(n14936), .A2(n13477), .ZN(n13310) );
  AOI22_X1 U15110 ( .A1(n13781), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n22556), .ZN(n13308) );
  INV_X1 U15111 ( .A(n13332), .ZN(n13321) );
  NAND2_X1 U15112 ( .A1(n13321), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13307) );
  AND2_X1 U15113 ( .A1(n13308), .A2(n13307), .ZN(n13309) );
  NAND2_X1 U15114 ( .A1(n13311), .A2(n15033), .ZN(n13312) );
  NAND2_X1 U15115 ( .A1(n13312), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14851) );
  NAND2_X1 U15116 ( .A1(n22556), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13315) );
  NAND2_X1 U15117 ( .A1(n13345), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13314) );
  OAI211_X1 U15118 ( .C1(n13332), .C2(n14761), .A(n13315), .B(n13314), .ZN(
        n13316) );
  AOI21_X1 U15119 ( .B1(n13313), .B2(n13477), .A(n13316), .ZN(n14850) );
  OR2_X1 U15120 ( .A1(n14851), .A2(n14850), .ZN(n14853) );
  INV_X1 U15121 ( .A(n14850), .ZN(n13317) );
  OR2_X1 U15122 ( .A1(n13317), .A2(n13751), .ZN(n13318) );
  NAND2_X1 U15123 ( .A1(n14853), .A2(n13318), .ZN(n14767) );
  NAND2_X1 U15124 ( .A1(n13321), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13325) );
  NAND2_X1 U15125 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13322) );
  AOI21_X1 U15126 ( .B1(n15381), .B2(n13322), .A(n13329), .ZN(n22245) );
  INV_X1 U15127 ( .A(n13786), .ZN(n13341) );
  OAI22_X1 U15128 ( .A1(n22245), .A2(n13751), .B1(n13341), .B2(n15381), .ZN(
        n13323) );
  AOI21_X1 U15129 ( .B1(n13781), .B2(P1_EAX_REG_3__SCAN_IN), .A(n13323), .ZN(
        n13324) );
  AND2_X1 U15130 ( .A1(n13325), .A2(n13324), .ZN(n13326) );
  INV_X1 U15131 ( .A(n13328), .ZN(n13336) );
  OAI21_X1 U15132 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13329), .A(
        n13337), .ZN(n22258) );
  OAI21_X1 U15133 ( .B1(n22405), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22556), .ZN(n13331) );
  NAND2_X1 U15134 ( .A1(n13781), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13330) );
  OAI211_X1 U15135 ( .C1(n13332), .C2(n18038), .A(n13331), .B(n13330), .ZN(
        n13333) );
  OAI21_X1 U15136 ( .B1(n13751), .B2(n22258), .A(n13333), .ZN(n13334) );
  INV_X1 U15137 ( .A(n13337), .ZN(n13339) );
  INV_X1 U15138 ( .A(n13346), .ZN(n13338) );
  OAI21_X1 U15139 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13339), .A(
        n13338), .ZN(n22279) );
  NAND2_X1 U15140 ( .A1(n22279), .A2(n13782), .ZN(n13340) );
  OAI21_X1 U15141 ( .B1(n22270), .B2(n13341), .A(n13340), .ZN(n13342) );
  AOI21_X1 U15142 ( .B1(n13781), .B2(P1_EAX_REG_5__SCAN_IN), .A(n13342), .ZN(
        n13343) );
  NAND2_X1 U15143 ( .A1(n15112), .A2(n15367), .ZN(n15366) );
  INV_X1 U15144 ( .A(n15366), .ZN(n13352) );
  INV_X1 U15145 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13348) );
  OAI21_X1 U15146 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13346), .A(
        n13353), .ZN(n22290) );
  AOI22_X1 U15147 ( .A1(n13782), .A2(n22290), .B1(n13786), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13347) );
  OAI21_X1 U15148 ( .B1(n13306), .B2(n13348), .A(n13347), .ZN(n13349) );
  NAND2_X1 U15149 ( .A1(n13352), .A2(n13351), .ZN(n15537) );
  INV_X1 U15150 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13357) );
  INV_X1 U15151 ( .A(n13353), .ZN(n13355) );
  INV_X1 U15152 ( .A(n13375), .ZN(n13354) );
  OAI21_X1 U15153 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13355), .A(
        n13354), .ZN(n22301) );
  AOI22_X1 U15154 ( .A1(n13782), .A2(n22301), .B1(n13786), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13356) );
  OAI21_X1 U15155 ( .B1(n13306), .B2(n13357), .A(n13356), .ZN(n13358) );
  AOI21_X1 U15156 ( .B1(n13359), .B2(n13477), .A(n13358), .ZN(n15585) );
  INV_X1 U15157 ( .A(n15585), .ZN(n13360) );
  AOI22_X1 U15158 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U15159 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U15160 ( .A1(n13759), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13363) );
  AOI22_X1 U15161 ( .A1(n13757), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13362) );
  NAND4_X1 U15162 ( .A1(n13365), .A2(n13364), .A3(n13363), .A4(n13362), .ZN(
        n13371) );
  AOI22_X1 U15163 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13369) );
  AOI22_X1 U15164 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13368) );
  AOI22_X1 U15165 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U15166 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13366) );
  NAND4_X1 U15167 ( .A1(n13369), .A2(n13368), .A3(n13367), .A4(n13366), .ZN(
        n13370) );
  OAI21_X1 U15168 ( .B1(n13371), .B2(n13370), .A(n13477), .ZN(n13374) );
  XNOR2_X1 U15169 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13375), .ZN(
        n22303) );
  AOI22_X1 U15170 ( .A1(n13782), .A2(n22303), .B1(n13786), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13373) );
  NAND2_X1 U15171 ( .A1(n13781), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13372) );
  XOR2_X1 U15172 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13400), .Z(n16680) );
  AOI22_X1 U15173 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13380) );
  AOI22_X1 U15174 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U15175 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U15176 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13377) );
  NAND4_X1 U15177 ( .A1(n13380), .A2(n13379), .A3(n13378), .A4(n13377), .ZN(
        n13386) );
  AOI22_X1 U15178 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13384) );
  AOI22_X1 U15179 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13383) );
  AOI22_X1 U15180 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13382) );
  AOI22_X1 U15181 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13381) );
  NAND4_X1 U15182 ( .A1(n13384), .A2(n13383), .A3(n13382), .A4(n13381), .ZN(
        n13385) );
  OR2_X1 U15183 ( .A1(n13386), .A2(n13385), .ZN(n13387) );
  AOI22_X1 U15184 ( .A1(n13477), .A2(n13387), .B1(n13786), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13389) );
  NAND2_X1 U15185 ( .A1(n13781), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13388) );
  OAI211_X1 U15186 ( .C1(n16680), .C2(n13751), .A(n13389), .B(n13388), .ZN(
        n15687) );
  AOI22_X1 U15187 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13434), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U15188 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13392) );
  AOI22_X1 U15189 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13391) );
  AOI22_X1 U15190 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13390) );
  NAND4_X1 U15191 ( .A1(n13393), .A2(n13392), .A3(n13391), .A4(n13390), .ZN(
        n13399) );
  AOI22_X1 U15192 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13397) );
  AOI22_X1 U15193 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U15194 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13395) );
  AOI22_X1 U15195 ( .A1(n13757), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13394) );
  NAND4_X1 U15196 ( .A1(n13397), .A2(n13396), .A3(n13395), .A4(n13394), .ZN(
        n13398) );
  NOR2_X1 U15197 ( .A1(n13399), .A2(n13398), .ZN(n13405) );
  INV_X1 U15198 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13401) );
  XNOR2_X1 U15199 ( .A(n13406), .B(n13401), .ZN(n15858) );
  NAND2_X1 U15200 ( .A1(n15858), .A2(n13782), .ZN(n13403) );
  AOI22_X1 U15201 ( .A1(n13345), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13786), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13402) );
  OAI211_X1 U15202 ( .C1(n13405), .C2(n13404), .A(n13403), .B(n13402), .ZN(
        n15853) );
  NAND2_X1 U15203 ( .A1(n13781), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n13409) );
  OAI21_X1 U15204 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13407), .A(
        n13445), .ZN(n22321) );
  AOI22_X1 U15205 ( .A1(n13626), .A2(n22321), .B1(n13786), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13408) );
  NAND2_X1 U15206 ( .A1(n13409), .A2(n13408), .ZN(n15908) );
  AOI22_X1 U15207 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13755), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15208 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U15209 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U15210 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13410) );
  NAND4_X1 U15211 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13419) );
  AOI22_X1 U15212 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15213 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U15214 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U15215 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U15216 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13418) );
  OR2_X1 U15217 ( .A1(n13419), .A2(n13418), .ZN(n13420) );
  XOR2_X1 U15218 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n13450), .Z(
        n16965) );
  AOI22_X1 U15219 ( .A1(n13345), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n13786), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13433) );
  AOI22_X1 U15220 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13434), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U15221 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U15222 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U15223 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13422) );
  NAND4_X1 U15224 ( .A1(n13425), .A2(n13424), .A3(n13423), .A4(n13422), .ZN(
        n13431) );
  AOI22_X1 U15225 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13429) );
  AOI22_X1 U15226 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U15227 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U15228 ( .A1(n13757), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13426) );
  NAND4_X1 U15229 ( .A1(n13429), .A2(n13428), .A3(n13427), .A4(n13426), .ZN(
        n13430) );
  OAI21_X1 U15230 ( .B1(n13431), .B2(n13430), .A(n13477), .ZN(n13432) );
  OAI211_X1 U15231 ( .C1(n16965), .C2(n13751), .A(n13433), .B(n13432), .ZN(
        n16663) );
  INV_X1 U15232 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n16835) );
  AOI22_X1 U15233 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13767), .B1(
        n13755), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U15234 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U15235 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13436) );
  BUF_X1 U15236 ( .A(n13434), .Z(n13734) );
  AOI22_X1 U15237 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13435) );
  NAND4_X1 U15238 ( .A1(n13438), .A2(n13437), .A3(n13436), .A4(n13435), .ZN(
        n13444) );
  AOI22_X1 U15239 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13604), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U15240 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13758), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13441) );
  AOI22_X1 U15241 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U15242 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n13757), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13439) );
  NAND4_X1 U15243 ( .A1(n13442), .A2(n13441), .A3(n13440), .A4(n13439), .ZN(
        n13443) );
  OAI21_X1 U15244 ( .B1(n13444), .B2(n13443), .A(n13477), .ZN(n13448) );
  XNOR2_X1 U15245 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n13445), .ZN(
        n22329) );
  INV_X1 U15246 ( .A(n22329), .ZN(n13446) );
  AOI22_X1 U15247 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13626), .B2(n13446), .ZN(n13447) );
  OAI211_X1 U15248 ( .C1(n13306), .C2(n16835), .A(n13448), .B(n13447), .ZN(
        n16662) );
  AND2_X1 U15249 ( .A1(n16663), .A2(n16662), .ZN(n13449) );
  INV_X1 U15250 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13451) );
  XNOR2_X1 U15251 ( .A(n13468), .B(n13451), .ZN(n16951) );
  AOI22_X1 U15252 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U15253 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U15254 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U15255 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13452) );
  NAND4_X1 U15256 ( .A1(n13455), .A2(n13454), .A3(n13453), .A4(n13452), .ZN(
        n13461) );
  AOI22_X1 U15257 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13459) );
  AOI22_X1 U15258 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U15259 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U15260 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13456) );
  NAND4_X1 U15261 ( .A1(n13459), .A2(n13458), .A3(n13457), .A4(n13456), .ZN(
        n13460) );
  OAI21_X1 U15262 ( .B1(n13461), .B2(n13460), .A(n13477), .ZN(n13464) );
  NAND2_X1 U15263 ( .A1(n13781), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U15264 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13462) );
  NAND3_X1 U15265 ( .A1(n13464), .A2(n13463), .A3(n13462), .ZN(n13465) );
  AOI21_X1 U15266 ( .B1(n16951), .B2(n13626), .A(n13465), .ZN(n15938) );
  NAND2_X1 U15267 ( .A1(n13467), .A2(n13466), .ZN(n15937) );
  XNOR2_X1 U15268 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n13486), .ZN(
        n22344) );
  INV_X1 U15269 ( .A(n22344), .ZN(n13484) );
  AOI22_X1 U15270 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13472) );
  AOI22_X1 U15271 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U15272 ( .A1(n13757), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U15273 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13469) );
  NAND4_X1 U15274 ( .A1(n13472), .A2(n13471), .A3(n13470), .A4(n13469), .ZN(
        n13479) );
  AOI22_X1 U15275 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13476) );
  AOI22_X1 U15276 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13755), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13475) );
  AOI22_X1 U15277 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13474) );
  AOI22_X1 U15278 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13473) );
  NAND4_X1 U15279 ( .A1(n13476), .A2(n13475), .A3(n13474), .A4(n13473), .ZN(
        n13478) );
  OAI21_X1 U15280 ( .B1(n13479), .B2(n13478), .A(n13477), .ZN(n13482) );
  NAND2_X1 U15281 ( .A1(n13781), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U15282 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13480) );
  NAND3_X1 U15283 ( .A1(n13482), .A2(n13481), .A3(n13480), .ZN(n13483) );
  AOI21_X1 U15284 ( .B1(n13484), .B2(n13782), .A(n13483), .ZN(n16733) );
  INV_X1 U15285 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13487) );
  XNOR2_X1 U15286 ( .A(n13504), .B(n13487), .ZN(n16650) );
  NAND2_X1 U15287 ( .A1(n16650), .A2(n13626), .ZN(n13503) );
  AOI22_X1 U15288 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13755), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13491) );
  AOI22_X1 U15289 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13490) );
  AOI22_X1 U15290 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13489) );
  AOI22_X1 U15291 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13488) );
  NAND4_X1 U15292 ( .A1(n13491), .A2(n13490), .A3(n13489), .A4(n13488), .ZN(
        n13499) );
  AOI22_X1 U15293 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13497) );
  NAND2_X1 U15294 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13493) );
  NAND2_X1 U15295 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13492) );
  AND3_X1 U15296 ( .A1(n13493), .A2(n13492), .A3(n13751), .ZN(n13496) );
  AOI22_X1 U15297 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13495) );
  AOI22_X1 U15298 ( .A1(n13757), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13494) );
  NAND4_X1 U15299 ( .A1(n13497), .A2(n13496), .A3(n13495), .A4(n13494), .ZN(
        n13498) );
  NAND2_X1 U15300 ( .A1(n13748), .A2(n13751), .ZN(n13596) );
  OAI21_X1 U15301 ( .B1(n13499), .B2(n13498), .A(n13596), .ZN(n13501) );
  AOI22_X1 U15302 ( .A1(n13345), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n22556), .ZN(n13500) );
  NAND2_X1 U15303 ( .A1(n13501), .A2(n13500), .ZN(n13502) );
  NAND2_X1 U15304 ( .A1(n13503), .A2(n13502), .ZN(n16646) );
  XNOR2_X1 U15305 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n13517), .ZN(
        n20861) );
  AOI22_X1 U15306 ( .A1(n13345), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13786), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U15307 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13508) );
  AOI22_X1 U15308 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13507) );
  AOI22_X1 U15309 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U15310 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13505) );
  NAND4_X1 U15311 ( .A1(n13508), .A2(n13507), .A3(n13506), .A4(n13505), .ZN(
        n13514) );
  AOI22_X1 U15312 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13512) );
  AOI22_X1 U15313 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13511) );
  AOI22_X1 U15314 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13510) );
  AOI22_X1 U15315 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13509) );
  NAND4_X1 U15316 ( .A1(n13512), .A2(n13511), .A3(n13510), .A4(n13509), .ZN(
        n13513) );
  OAI21_X1 U15317 ( .B1(n13514), .B2(n13513), .A(n13778), .ZN(n13515) );
  OAI211_X1 U15318 ( .C1(n20861), .C2(n13751), .A(n13516), .B(n13515), .ZN(
        n16635) );
  INV_X1 U15319 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13518) );
  XNOR2_X1 U15320 ( .A(n13552), .B(n13518), .ZN(n16628) );
  NAND2_X1 U15321 ( .A1(n16628), .A2(n13626), .ZN(n13535) );
  AOI22_X1 U15322 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U15323 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U15324 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13520) );
  AOI22_X1 U15325 ( .A1(n13768), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13519) );
  NAND4_X1 U15326 ( .A1(n13522), .A2(n13521), .A3(n13520), .A4(n13519), .ZN(
        n13531) );
  NAND2_X1 U15327 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13525) );
  NAND2_X1 U15328 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13524) );
  AND3_X1 U15329 ( .A1(n13525), .A2(n13524), .A3(n13751), .ZN(n13529) );
  AOI22_X1 U15330 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13528) );
  AOI22_X1 U15331 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13759), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U15332 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13526) );
  NAND4_X1 U15333 ( .A1(n13529), .A2(n13528), .A3(n13527), .A4(n13526), .ZN(
        n13530) );
  OAI21_X1 U15334 ( .B1(n13531), .B2(n13530), .A(n13596), .ZN(n13533) );
  AOI22_X1 U15335 ( .A1(n13345), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n22556), .ZN(n13532) );
  NAND2_X1 U15336 ( .A1(n13533), .A2(n13532), .ZN(n13534) );
  NAND2_X1 U15337 ( .A1(n13535), .A2(n13534), .ZN(n16624) );
  AOI22_X1 U15338 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U15339 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U15340 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13759), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13539) );
  AOI22_X1 U15341 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13538) );
  NAND4_X1 U15342 ( .A1(n13541), .A2(n13540), .A3(n13539), .A4(n13538), .ZN(
        n13547) );
  AOI22_X1 U15343 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13545) );
  AOI22_X1 U15344 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13544) );
  AOI22_X1 U15345 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13543) );
  AOI22_X1 U15346 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13542) );
  NAND4_X1 U15347 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        n13546) );
  NOR2_X1 U15348 ( .A1(n13547), .A2(n13546), .ZN(n13551) );
  NAND2_X1 U15349 ( .A1(n22556), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13548) );
  NAND2_X1 U15350 ( .A1(n13751), .A2(n13548), .ZN(n13549) );
  AOI21_X1 U15351 ( .B1(n13781), .B2(P1_EAX_REG_19__SCAN_IN), .A(n13549), .ZN(
        n13550) );
  OAI21_X1 U15352 ( .B1(n13748), .B2(n13551), .A(n13550), .ZN(n13555) );
  OAI21_X1 U15353 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n13553), .A(
        n13569), .ZN(n22351) );
  OR2_X1 U15354 ( .A1(n13751), .A2(n22351), .ZN(n13554) );
  NAND2_X1 U15355 ( .A1(n13555), .A2(n13554), .ZN(n16726) );
  AOI22_X1 U15356 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13559) );
  AOI22_X1 U15357 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13558) );
  AOI22_X1 U15358 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13759), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13557) );
  AOI22_X1 U15359 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13556) );
  NAND4_X1 U15360 ( .A1(n13559), .A2(n13558), .A3(n13557), .A4(n13556), .ZN(
        n13565) );
  AOI22_X1 U15361 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13758), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U15362 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13755), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13562) );
  AOI22_X1 U15363 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U15364 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13560) );
  NAND4_X1 U15365 ( .A1(n13563), .A2(n13562), .A3(n13561), .A4(n13560), .ZN(
        n13564) );
  OAI21_X1 U15366 ( .B1(n13565), .B2(n13564), .A(n13778), .ZN(n13568) );
  INV_X1 U15367 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16919) );
  AOI21_X1 U15368 ( .B1(n16919), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13566) );
  AOI21_X1 U15369 ( .B1(n13781), .B2(P1_EAX_REG_20__SCAN_IN), .A(n13566), .ZN(
        n13567) );
  XNOR2_X1 U15370 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n13569), .ZN(
        n16921) );
  AOI22_X1 U15371 ( .A1(n13568), .A2(n13567), .B1(n13626), .B2(n16921), .ZN(
        n16612) );
  OAI21_X1 U15372 ( .B1(n13570), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n13601), .ZN(n22384) );
  INV_X1 U15373 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n16790) );
  AOI22_X1 U15374 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13574) );
  AOI22_X1 U15375 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13573) );
  AOI22_X1 U15376 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13572) );
  AOI22_X1 U15377 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13571) );
  NAND4_X1 U15378 ( .A1(n13574), .A2(n13573), .A3(n13572), .A4(n13571), .ZN(
        n13580) );
  AOI22_X1 U15379 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13578) );
  AOI22_X1 U15380 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13577) );
  AOI22_X1 U15381 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13759), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13576) );
  AOI22_X1 U15382 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13575) );
  NAND4_X1 U15383 ( .A1(n13578), .A2(n13577), .A3(n13576), .A4(n13575), .ZN(
        n13579) );
  OAI21_X1 U15384 ( .B1(n13580), .B2(n13579), .A(n13778), .ZN(n13582) );
  OAI21_X1 U15385 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n22405), .A(
        n22556), .ZN(n13581) );
  OAI211_X1 U15386 ( .C1(n13306), .C2(n16790), .A(n13582), .B(n13581), .ZN(
        n13583) );
  OAI21_X1 U15387 ( .B1(n22384), .B2(n13751), .A(n13583), .ZN(n16721) );
  AOI22_X1 U15388 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U15389 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13604), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13587) );
  AOI22_X1 U15390 ( .A1(n13434), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13584), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13586) );
  AOI22_X1 U15391 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13585) );
  NAND4_X1 U15392 ( .A1(n13588), .A2(n13587), .A3(n13586), .A4(n13585), .ZN(
        n13598) );
  INV_X1 U15393 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13591) );
  AOI22_X1 U15394 ( .A1(n13757), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13590) );
  AOI21_X1 U15395 ( .B1(n13765), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n13626), .ZN(n13589) );
  OAI211_X1 U15396 ( .C1(n13091), .C2(n13591), .A(n13590), .B(n13589), .ZN(
        n13592) );
  INV_X1 U15397 ( .A(n13592), .ZN(n13595) );
  AOI22_X1 U15398 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U15399 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13593) );
  NAND3_X1 U15400 ( .A1(n13595), .A2(n13594), .A3(n13593), .ZN(n13597) );
  OAI21_X1 U15401 ( .B1(n13598), .B2(n13597), .A(n13596), .ZN(n13600) );
  AOI22_X1 U15402 ( .A1(n13345), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n22556), .ZN(n13599) );
  XNOR2_X1 U15403 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n13601), .ZN(
        n16908) );
  AOI22_X1 U15404 ( .A1(n13600), .A2(n13599), .B1(n13626), .B2(n16908), .ZN(
        n16600) );
  OAI21_X1 U15405 ( .B1(n13603), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n13647), .ZN(n16900) );
  AOI22_X1 U15406 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U15407 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13604), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13607) );
  AOI22_X1 U15408 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13606) );
  AOI22_X1 U15409 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13605) );
  NAND4_X1 U15410 ( .A1(n13608), .A2(n13607), .A3(n13606), .A4(n13605), .ZN(
        n13614) );
  AOI22_X1 U15411 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13612) );
  AOI22_X1 U15412 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U15413 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U15414 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13609) );
  NAND4_X1 U15415 ( .A1(n13612), .A2(n13611), .A3(n13610), .A4(n13609), .ZN(
        n13613) );
  NOR2_X1 U15416 ( .A1(n13614), .A2(n13613), .ZN(n13641) );
  AOI22_X1 U15417 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U15418 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13617) );
  AOI22_X1 U15419 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13616) );
  AOI22_X1 U15420 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13615) );
  NAND4_X1 U15421 ( .A1(n13618), .A2(n13617), .A3(n13616), .A4(n13615), .ZN(
        n13625) );
  AOI22_X1 U15422 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13623) );
  AOI22_X1 U15423 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13622) );
  AOI22_X1 U15424 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13621) );
  AOI22_X1 U15425 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13620) );
  NAND4_X1 U15426 ( .A1(n13623), .A2(n13622), .A3(n13621), .A4(n13620), .ZN(
        n13624) );
  NOR2_X1 U15427 ( .A1(n13625), .A2(n13624), .ZN(n13642) );
  XNOR2_X1 U15428 ( .A(n13641), .B(n13642), .ZN(n13629) );
  AOI21_X1 U15429 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n22556), .A(
        n13626), .ZN(n13628) );
  NAND2_X1 U15430 ( .A1(n13345), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n13627) );
  OAI211_X1 U15431 ( .C1(n13748), .C2(n13629), .A(n13628), .B(n13627), .ZN(
        n13630) );
  OAI21_X1 U15432 ( .B1(n13751), .B2(n16900), .A(n13630), .ZN(n16586) );
  XNOR2_X1 U15433 ( .A(n13647), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16894) );
  AOI22_X1 U15434 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U15435 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13633) );
  AOI22_X1 U15436 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13632) );
  AOI22_X1 U15437 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13631) );
  NAND4_X1 U15438 ( .A1(n13634), .A2(n13633), .A3(n13632), .A4(n13631), .ZN(
        n13640) );
  AOI22_X1 U15439 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13769), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13638) );
  AOI22_X1 U15440 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13637) );
  AOI22_X1 U15441 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U15442 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13635) );
  NAND4_X1 U15443 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13635), .ZN(
        n13639) );
  OR2_X1 U15444 ( .A1(n13640), .A2(n13639), .ZN(n13663) );
  NOR2_X1 U15445 ( .A1(n13642), .A2(n13641), .ZN(n13664) );
  XOR2_X1 U15446 ( .A(n13663), .B(n13664), .Z(n13645) );
  INV_X1 U15447 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n22482) );
  OAI21_X1 U15448 ( .B1(n22405), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n22556), .ZN(n13643) );
  OAI21_X1 U15449 ( .B1(n13306), .B2(n22482), .A(n13643), .ZN(n13644) );
  AOI21_X1 U15450 ( .B1(n13645), .B2(n13778), .A(n13644), .ZN(n13646) );
  AOI21_X1 U15451 ( .B1(n13782), .B2(n16894), .A(n13646), .ZN(n16574) );
  NAND2_X1 U15452 ( .A1(n16573), .A2(n16574), .ZN(n16563) );
  INV_X1 U15453 ( .A(n13648), .ZN(n13649) );
  INV_X1 U15454 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16566) );
  NAND2_X1 U15455 ( .A1(n13649), .A2(n16566), .ZN(n13650) );
  NAND2_X1 U15456 ( .A1(n13687), .A2(n13650), .ZN(n16883) );
  AOI22_X1 U15457 ( .A1(n13651), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13655) );
  AOI22_X1 U15458 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U15459 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U15460 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13652) );
  NAND4_X1 U15461 ( .A1(n13655), .A2(n13654), .A3(n13653), .A4(n13652), .ZN(
        n13662) );
  AOI22_X1 U15462 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U15463 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U15464 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13656), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U15465 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13657) );
  NAND4_X1 U15466 ( .A1(n13660), .A2(n13659), .A3(n13658), .A4(n13657), .ZN(
        n13661) );
  NOR2_X1 U15467 ( .A1(n13662), .A2(n13661), .ZN(n13670) );
  NAND2_X1 U15468 ( .A1(n13664), .A2(n13663), .ZN(n13669) );
  XNOR2_X1 U15469 ( .A(n13670), .B(n13669), .ZN(n13667) );
  OAI21_X1 U15470 ( .B1(n22405), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n22556), .ZN(n13666) );
  NAND2_X1 U15471 ( .A1(n13345), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n13665) );
  OAI211_X1 U15472 ( .C1(n13667), .C2(n13748), .A(n13666), .B(n13665), .ZN(
        n13668) );
  OAI21_X1 U15473 ( .B1(n13751), .B2(n16883), .A(n13668), .ZN(n16565) );
  NOR2_X1 U15474 ( .A1(n13670), .A2(n13669), .ZN(n13693) );
  AOI22_X1 U15475 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U15476 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U15477 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13672) );
  AOI22_X1 U15478 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13671) );
  NAND4_X1 U15479 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13680) );
  AOI22_X1 U15480 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U15481 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U15482 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13676) );
  AOI22_X1 U15483 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13675) );
  NAND4_X1 U15484 ( .A1(n13678), .A2(n13677), .A3(n13676), .A4(n13675), .ZN(
        n13679) );
  OR2_X1 U15485 ( .A1(n13680), .A2(n13679), .ZN(n13692) );
  INV_X1 U15486 ( .A(n13692), .ZN(n13681) );
  XNOR2_X1 U15487 ( .A(n13693), .B(n13681), .ZN(n13682) );
  NAND2_X1 U15488 ( .A1(n13682), .A2(n13778), .ZN(n13686) );
  INV_X1 U15489 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16552) );
  AOI21_X1 U15490 ( .B1(n16552), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13683) );
  AOI21_X1 U15491 ( .B1(n13781), .B2(P1_EAX_REG_26__SCAN_IN), .A(n13683), .ZN(
        n13685) );
  XNOR2_X1 U15492 ( .A(n13687), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16551) );
  AOI21_X1 U15493 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(n16550) );
  INV_X1 U15494 ( .A(n13687), .ZN(n13688) );
  INV_X1 U15495 ( .A(n13689), .ZN(n13690) );
  INV_X1 U15496 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16542) );
  NAND2_X1 U15497 ( .A1(n13690), .A2(n16542), .ZN(n13691) );
  NAND2_X1 U15498 ( .A1(n13726), .A2(n13691), .ZN(n16867) );
  NAND2_X1 U15499 ( .A1(n13693), .A2(n13692), .ZN(n13720) );
  AOI22_X1 U15500 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13758), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U15501 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13709), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U15502 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13766), .B1(
        n13694), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U15503 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13695) );
  NAND4_X1 U15504 ( .A1(n13698), .A2(n13697), .A3(n13696), .A4(n13695), .ZN(
        n13704) );
  AOI22_X1 U15505 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13756), .B1(
        n13755), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U15506 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U15507 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U15508 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13033), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13699) );
  NAND4_X1 U15509 ( .A1(n13702), .A2(n13701), .A3(n13700), .A4(n13699), .ZN(
        n13703) );
  NOR2_X1 U15510 ( .A1(n13704), .A2(n13703), .ZN(n13721) );
  XNOR2_X1 U15511 ( .A(n13720), .B(n13721), .ZN(n13707) );
  AOI21_X1 U15512 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n22556), .A(
        n13782), .ZN(n13706) );
  NAND2_X1 U15513 ( .A1(n13345), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n13705) );
  OAI211_X1 U15514 ( .C1(n13707), .C2(n13748), .A(n13706), .B(n13705), .ZN(
        n13708) );
  OAI21_X1 U15515 ( .B1(n13751), .B2(n16867), .A(n13708), .ZN(n16538) );
  XNOR2_X1 U15516 ( .A(n13726), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16863) );
  AOI22_X1 U15517 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U15518 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U15519 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13759), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U15520 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13710) );
  NAND4_X1 U15521 ( .A1(n13713), .A2(n13712), .A3(n13711), .A4(n13710), .ZN(
        n13719) );
  AOI22_X1 U15522 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U15523 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13716) );
  AOI22_X1 U15524 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U15525 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13714) );
  NAND4_X1 U15526 ( .A1(n13717), .A2(n13716), .A3(n13715), .A4(n13714), .ZN(
        n13718) );
  OR2_X1 U15527 ( .A1(n13719), .A2(n13718), .ZN(n13732) );
  NOR2_X1 U15528 ( .A1(n13721), .A2(n13720), .ZN(n13733) );
  XOR2_X1 U15529 ( .A(n13732), .B(n13733), .Z(n13724) );
  INV_X1 U15530 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n22509) );
  OAI21_X1 U15531 ( .B1(n22405), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n22556), .ZN(n13722) );
  OAI21_X1 U15532 ( .B1(n13306), .B2(n22509), .A(n13722), .ZN(n13723) );
  AOI21_X1 U15533 ( .B1(n13724), .B2(n13778), .A(n13723), .ZN(n13725) );
  INV_X1 U15534 ( .A(n13726), .ZN(n13727) );
  INV_X1 U15535 ( .A(n13728), .ZN(n13730) );
  INV_X1 U15536 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13729) );
  NAND2_X1 U15537 ( .A1(n13730), .A2(n13729), .ZN(n13731) );
  NAND2_X1 U15538 ( .A1(n13791), .A2(n13731), .ZN(n16852) );
  NAND2_X1 U15539 ( .A1(n13733), .A2(n13732), .ZN(n13752) );
  AOI22_X1 U15540 ( .A1(n13755), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13767), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13738) );
  AOI22_X1 U15541 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U15542 ( .A1(n13765), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13759), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13736) );
  AOI22_X1 U15543 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13735) );
  NAND4_X1 U15544 ( .A1(n13738), .A2(n13737), .A3(n13736), .A4(n13735), .ZN(
        n13745) );
  AOI22_X1 U15545 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13743) );
  AOI22_X1 U15546 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U15547 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13741) );
  AOI22_X1 U15548 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13740) );
  NAND4_X1 U15549 ( .A1(n13743), .A2(n13742), .A3(n13741), .A4(n13740), .ZN(
        n13744) );
  NOR2_X1 U15550 ( .A1(n13745), .A2(n13744), .ZN(n13753) );
  XNOR2_X1 U15551 ( .A(n13752), .B(n13753), .ZN(n13749) );
  AOI21_X1 U15552 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n22556), .A(
        n13782), .ZN(n13747) );
  NAND2_X1 U15553 ( .A1(n13781), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13746) );
  OAI211_X1 U15554 ( .C1(n13749), .C2(n13748), .A(n13747), .B(n13746), .ZN(
        n13750) );
  OAI21_X1 U15555 ( .B1(n13751), .B2(n16852), .A(n13750), .ZN(n14190) );
  NOR2_X1 U15556 ( .A1(n13753), .A2(n13752), .ZN(n13777) );
  AOI22_X1 U15557 ( .A1(n13734), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13754), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U15558 ( .A1(n13756), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13755), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13762) );
  AOI22_X1 U15559 ( .A1(n13758), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13757), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U15560 ( .A1(n13759), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13739), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13760) );
  NAND4_X1 U15561 ( .A1(n13763), .A2(n13762), .A3(n13761), .A4(n13760), .ZN(
        n13775) );
  AOI22_X1 U15562 ( .A1(n13764), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13651), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U15563 ( .A1(n13766), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13765), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13772) );
  AOI22_X1 U15564 ( .A1(n13767), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13619), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U15565 ( .A1(n13769), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13768), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13770) );
  NAND4_X1 U15566 ( .A1(n13773), .A2(n13772), .A3(n13771), .A4(n13770), .ZN(
        n13774) );
  NOR2_X1 U15567 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  XNOR2_X1 U15568 ( .A(n13777), .B(n13776), .ZN(n13779) );
  NAND2_X1 U15569 ( .A1(n13779), .A2(n13778), .ZN(n13785) );
  INV_X1 U15570 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16845) );
  AOI21_X1 U15571 ( .B1(n16845), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13780) );
  AOI21_X1 U15572 ( .B1(n13781), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13780), .ZN(
        n13784) );
  XNOR2_X1 U15573 ( .A(n13791), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16843) );
  AOI21_X1 U15574 ( .B1(n13785), .B2(n13784), .A(n13783), .ZN(n16515) );
  AOI22_X1 U15575 ( .A1(n13781), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13786), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13787) );
  NAND3_X1 U15576 ( .A1(n22392), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n18054) );
  NAND2_X1 U15577 ( .A1(n16743), .A2(n20873), .ZN(n13797) );
  NAND2_X1 U15578 ( .A1(n13789), .A2(n22609), .ZN(n22105) );
  NAND2_X1 U15579 ( .A1(n22105), .A2(n22392), .ZN(n13790) );
  NAND2_X1 U15580 ( .A1(n22392), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n18047) );
  NAND2_X1 U15581 ( .A1(n22405), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14201) );
  NAND2_X1 U15582 ( .A1(n18047), .A2(n14201), .ZN(n14858) );
  INV_X1 U15583 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13792) );
  OR2_X1 U15584 ( .A1(n22609), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20881) );
  INV_X1 U15585 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20791) );
  NOR2_X1 U15586 ( .A1(n22129), .A2(n20791), .ZN(n16989) );
  AOI21_X1 U15587 ( .B1(n20870), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16989), .ZN(n13794) );
  OAI21_X1 U15588 ( .B1(n20877), .B2(n14314), .A(n13794), .ZN(n13795) );
  INV_X1 U15589 ( .A(n13795), .ZN(n13796) );
  OAI211_X1 U15590 ( .C1(n16991), .C2(n22385), .A(n13797), .B(n13796), .ZN(
        P1_U2968) );
  NAND2_X1 U15591 ( .A1(n20219), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15315) );
  AOI21_X1 U15592 ( .B1(n15315), .B2(n20140), .A(n20254), .ZN(n13799) );
  INV_X1 U15593 ( .A(n15315), .ZN(n13798) );
  NAND2_X1 U15594 ( .A1(n13798), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15763) );
  AOI22_X1 U15595 ( .A1(n13820), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13799), .B2(n15763), .ZN(n13805) );
  INV_X1 U15596 ( .A(n13805), .ZN(n13803) );
  NOR2_X1 U15597 ( .A1(n14069), .A2(n15784), .ZN(n13804) );
  NAND2_X1 U15598 ( .A1(n13803), .A2(n13804), .ZN(n13831) );
  NAND2_X1 U15599 ( .A1(n11261), .A2(n13824), .ZN(n13808) );
  INV_X1 U15600 ( .A(n13804), .ZN(n13806) );
  AND2_X1 U15601 ( .A1(n13806), .A2(n13805), .ZN(n13807) );
  NAND2_X1 U15602 ( .A1(n13808), .A2(n13807), .ZN(n13809) );
  NAND2_X1 U15603 ( .A1(n13810), .A2(n13824), .ZN(n13813) );
  INV_X1 U15604 ( .A(n20219), .ZN(n15314) );
  NAND2_X1 U15605 ( .A1(n15314), .A2(n20161), .ZN(n13811) );
  AND2_X1 U15606 ( .A1(n15315), .A2(n13811), .ZN(n20117) );
  AOI22_X1 U15607 ( .A1(n13820), .A2(n17957), .B1(n20222), .B2(n20117), .ZN(
        n13812) );
  NAND2_X1 U15608 ( .A1(n13813), .A2(n13812), .ZN(n13815) );
  NOR2_X1 U15609 ( .A1(n14069), .A2(n20494), .ZN(n13814) );
  OR2_X1 U15610 ( .A1(n13815), .A2(n13814), .ZN(n13816) );
  NAND2_X1 U15611 ( .A1(n13815), .A2(n13814), .ZN(n13828) );
  NOR2_X1 U15613 ( .A1(n20254), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13817) );
  AOI21_X1 U15614 ( .B1(n13820), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13817), .ZN(n13818) );
  NAND2_X1 U15617 ( .A1(n13820), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13822) );
  NOR2_X1 U15618 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20205) );
  INV_X1 U15619 ( .A(n20205), .ZN(n13821) );
  NAND2_X1 U15620 ( .A1(n15314), .A2(n13821), .ZN(n20183) );
  NAND2_X1 U15621 ( .A1(n13822), .A2(n20233), .ZN(n13823) );
  INV_X1 U15622 ( .A(n13825), .ZN(n13826) );
  NOR2_X1 U15623 ( .A1(n14658), .A2(n13826), .ZN(n13827) );
  AOI21_X2 U15624 ( .B1(n14715), .B2(n14714), .A(n13827), .ZN(n14765) );
  NAND2_X1 U15625 ( .A1(n14764), .A2(n14765), .ZN(n13829) );
  NAND2_X1 U15626 ( .A1(n14899), .A2(n14900), .ZN(n14901) );
  NOR2_X1 U15627 ( .A1(n14069), .A2(n20400), .ZN(n14881) );
  NAND2_X1 U15628 ( .A1(n15632), .A2(n15636), .ZN(n15634) );
  INV_X1 U15629 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13924) );
  INV_X1 U15630 ( .A(n13964), .ZN(n13895) );
  INV_X1 U15631 ( .A(n13963), .ZN(n13894) );
  INV_X1 U15632 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13929) );
  OAI22_X1 U15633 ( .A1(n13924), .A2(n13895), .B1(n13894), .B2(n13929), .ZN(
        n13833) );
  AOI21_X1 U15634 ( .B1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n12219), .A(
        n13833), .ZN(n13835) );
  AOI22_X1 U15635 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13834) );
  OAI211_X1 U15636 ( .C1(n20671), .C2(n13915), .A(n13835), .B(n13834), .ZN(
        n13844) );
  AOI22_X1 U15637 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13839) );
  AOI22_X1 U15638 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13838) );
  AOI22_X1 U15639 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13837) );
  AOI22_X1 U15640 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13836) );
  NAND4_X1 U15641 ( .A1(n13839), .A2(n13838), .A3(n13837), .A4(n13836), .ZN(
        n13843) );
  INV_X1 U15642 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13841) );
  INV_X1 U15643 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13840) );
  OAI22_X1 U15644 ( .A1(n13919), .A2(n13841), .B1(n13917), .B2(n13840), .ZN(
        n13842) );
  NOR3_X1 U15645 ( .A1(n13844), .A2(n13843), .A3(n13842), .ZN(n15867) );
  INV_X1 U15646 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13848) );
  INV_X1 U15647 ( .A(n13958), .ZN(n13847) );
  INV_X1 U15648 ( .A(n13957), .ZN(n13846) );
  OAI22_X1 U15649 ( .A1(n13848), .A2(n13847), .B1(n13846), .B2(n13845), .ZN(
        n13851) );
  AOI22_X1 U15650 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13849) );
  OAI21_X1 U15651 ( .B1(n13985), .B2(n13913), .A(n13849), .ZN(n13850) );
  AOI211_X1 U15652 ( .C1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .C2(n13956), .A(
        n13851), .B(n13850), .ZN(n13858) );
  AOI22_X1 U15653 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13857) );
  AOI22_X1 U15654 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U15655 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U15656 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U15657 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13852) );
  AND4_X1 U15658 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13856) );
  NAND3_X1 U15659 ( .A1(n13858), .A2(n13857), .A3(n13856), .ZN(n15888) );
  AOI22_X1 U15660 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13862) );
  AOI22_X1 U15661 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13861) );
  AOI22_X1 U15662 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13860) );
  AOI22_X1 U15663 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13859) );
  NAND4_X1 U15664 ( .A1(n13862), .A2(n13861), .A3(n13860), .A4(n13859), .ZN(
        n13870) );
  INV_X1 U15665 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14010) );
  AOI22_X1 U15666 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13863) );
  OAI21_X1 U15667 ( .B1(n14010), .B2(n13913), .A(n13863), .ZN(n13869) );
  AOI22_X1 U15668 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13864) );
  OAI21_X1 U15669 ( .B1(n20494), .B2(n13915), .A(n13864), .ZN(n13868) );
  INV_X1 U15670 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13866) );
  INV_X1 U15671 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13865) );
  OAI22_X1 U15672 ( .A1(n13919), .A2(n13866), .B1(n13917), .B2(n13865), .ZN(
        n13867) );
  NOR4_X1 U15673 ( .A1(n13870), .A2(n13869), .A3(n13868), .A4(n13867), .ZN(
        n15919) );
  INV_X1 U15674 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14025) );
  INV_X1 U15675 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13871) );
  OAI22_X1 U15676 ( .A1(n14025), .A2(n13895), .B1(n13894), .B2(n13871), .ZN(
        n13874) );
  AOI22_X1 U15677 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13872) );
  OAI21_X1 U15678 ( .B1(n15784), .B2(n13915), .A(n13872), .ZN(n13873) );
  AOI211_X1 U15679 ( .C1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .C2(n12219), .A(
        n13874), .B(n13873), .ZN(n13881) );
  AOI22_X1 U15680 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U15681 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U15682 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U15683 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U15684 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13875) );
  AND4_X1 U15685 ( .A1(n13878), .A2(n13877), .A3(n13876), .A4(n13875), .ZN(
        n13879) );
  NAND3_X1 U15686 ( .A1(n13881), .A2(n13880), .A3(n13879), .ZN(n17310) );
  NAND2_X1 U15687 ( .A1(n15918), .A2(n17310), .ZN(n17300) );
  INV_X1 U15688 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14048) );
  INV_X1 U15689 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14050) );
  OAI22_X1 U15690 ( .A1(n14048), .A2(n13895), .B1(n13894), .B2(n14050), .ZN(
        n13882) );
  AOI21_X1 U15691 ( .B1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n12219), .A(
        n13882), .ZN(n13884) );
  AOI22_X1 U15692 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13883) );
  OAI211_X1 U15693 ( .C1(n20400), .C2(n13915), .A(n13884), .B(n13883), .ZN(
        n13893) );
  AOI22_X1 U15694 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U15695 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13887) );
  AOI22_X1 U15696 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U15697 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13885) );
  NAND4_X1 U15698 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n13892) );
  INV_X1 U15699 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13890) );
  INV_X1 U15700 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13889) );
  OAI22_X1 U15701 ( .A1(n13919), .A2(n13890), .B1(n13917), .B2(n13889), .ZN(
        n13891) );
  NOR3_X1 U15702 ( .A1(n13893), .A2(n13892), .A3(n13891), .ZN(n17302) );
  INV_X1 U15703 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14071) );
  INV_X1 U15704 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14073) );
  OAI22_X1 U15705 ( .A1(n14071), .A2(n13895), .B1(n13894), .B2(n14073), .ZN(
        n13896) );
  AOI21_X1 U15706 ( .B1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B2(n12219), .A(
        n13896), .ZN(n13898) );
  AOI22_X1 U15707 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13897) );
  OAI211_X1 U15708 ( .C1(n20360), .C2(n13915), .A(n13898), .B(n13897), .ZN(
        n13907) );
  AOI22_X1 U15709 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U15710 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U15711 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U15712 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13899) );
  NAND4_X1 U15713 ( .A1(n13902), .A2(n13901), .A3(n13900), .A4(n13899), .ZN(
        n13906) );
  OAI22_X1 U15714 ( .A1(n13919), .A2(n13904), .B1(n13917), .B2(n13903), .ZN(
        n13905) );
  AOI22_X1 U15715 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U15716 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13910) );
  AOI22_X1 U15717 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U15718 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13908) );
  NAND4_X1 U15719 ( .A1(n13911), .A2(n13910), .A3(n13909), .A4(n13908), .ZN(
        n13923) );
  AOI22_X1 U15720 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13912) );
  OAI21_X1 U15721 ( .B1(n14106), .B2(n13913), .A(n13912), .ZN(n13922) );
  AOI22_X1 U15722 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13914) );
  OAI21_X1 U15723 ( .B1(n20311), .B2(n13915), .A(n13914), .ZN(n13921) );
  INV_X1 U15724 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13918) );
  OAI22_X1 U15725 ( .A1(n13919), .A2(n13918), .B1(n13917), .B2(n13916), .ZN(
        n13920) );
  NOR4_X1 U15726 ( .A1(n13923), .A2(n13922), .A3(n13921), .A4(n13920), .ZN(
        n17288) );
  AOI22_X1 U15727 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13934) );
  AOI22_X1 U15728 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U15729 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13932) );
  INV_X1 U15730 ( .A(n11996), .ZN(n15285) );
  INV_X1 U15731 ( .A(n14163), .ZN(n14169) );
  OR2_X1 U15732 ( .A1(n14169), .A2(n13924), .ZN(n13928) );
  INV_X1 U15733 ( .A(n13925), .ZN(n13927) );
  NAND2_X1 U15734 ( .A1(n13927), .A2(n13926), .ZN(n14167) );
  OAI211_X1 U15735 ( .C1(n15285), .C2(n13929), .A(n13928), .B(n14167), .ZN(
        n13930) );
  INV_X1 U15736 ( .A(n13930), .ZN(n13931) );
  NAND4_X1 U15737 ( .A1(n13934), .A2(n13933), .A3(n13932), .A4(n13931), .ZN(
        n13945) );
  AOI22_X1 U15738 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13943) );
  AOI22_X1 U15739 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13942) );
  AOI22_X1 U15740 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13941) );
  INV_X1 U15741 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13938) );
  INV_X1 U15742 ( .A(n14167), .ZN(n14104) );
  INV_X1 U15743 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13936) );
  OR2_X1 U15744 ( .A1(n14169), .A2(n13936), .ZN(n13937) );
  OAI211_X1 U15745 ( .C1(n15285), .C2(n13938), .A(n14104), .B(n13937), .ZN(
        n13939) );
  INV_X1 U15746 ( .A(n13939), .ZN(n13940) );
  NAND4_X1 U15747 ( .A1(n13943), .A2(n13942), .A3(n13941), .A4(n13940), .ZN(
        n13944) );
  NAND2_X1 U15748 ( .A1(n13945), .A2(n13944), .ZN(n13972) );
  AOI22_X1 U15749 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13946), .B1(
        n12228), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U15750 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n13947), .B1(
        n12300), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U15751 ( .A1(n13949), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13948), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U15752 ( .A1(n13951), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13950), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13952) );
  NAND4_X1 U15753 ( .A1(n13955), .A2(n13954), .A3(n13953), .A4(n13952), .ZN(
        n13970) );
  NAND2_X1 U15754 ( .A1(n13956), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13960) );
  AOI22_X1 U15755 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13958), .B1(
        n13957), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13959) );
  AND2_X1 U15756 ( .A1(n13960), .A2(n13959), .ZN(n13968) );
  AOI22_X1 U15757 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13961), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U15758 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13964), .B1(
        n13963), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U15759 ( .A1(n12219), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13965) );
  NAND4_X1 U15760 ( .A1(n13968), .A2(n13967), .A3(n13966), .A4(n13965), .ZN(
        n13969) );
  NOR2_X1 U15761 ( .A1(n13970), .A2(n13969), .ZN(n13971) );
  XOR2_X1 U15762 ( .A(n13972), .B(n13971), .Z(n17280) );
  INV_X1 U15763 ( .A(n13971), .ZN(n13974) );
  INV_X1 U15764 ( .A(n13972), .ZN(n13973) );
  AND2_X1 U15765 ( .A1(n13974), .A2(n13973), .ZN(n13994) );
  AOI22_X1 U15766 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13982) );
  AOI22_X1 U15767 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13981) );
  AOI22_X1 U15768 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13980) );
  INV_X1 U15769 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13977) );
  INV_X1 U15770 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13975) );
  OR2_X1 U15771 ( .A1(n14169), .A2(n13975), .ZN(n13976) );
  OAI211_X1 U15772 ( .C1(n15285), .C2(n13977), .A(n13976), .B(n14167), .ZN(
        n13978) );
  INV_X1 U15773 ( .A(n13978), .ZN(n13979) );
  NAND4_X1 U15774 ( .A1(n13982), .A2(n13981), .A3(n13980), .A4(n13979), .ZN(
        n13992) );
  AOI22_X1 U15775 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14175), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U15776 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13989) );
  AOI22_X1 U15777 ( .A1(n14176), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11255), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13988) );
  OR2_X1 U15778 ( .A1(n14169), .A2(n13983), .ZN(n13984) );
  OAI211_X1 U15779 ( .C1(n15285), .C2(n13985), .A(n14104), .B(n13984), .ZN(
        n13986) );
  INV_X1 U15780 ( .A(n13986), .ZN(n13987) );
  NAND4_X1 U15781 ( .A1(n13990), .A2(n13989), .A3(n13988), .A4(n13987), .ZN(
        n13991) );
  NAND2_X1 U15782 ( .A1(n13992), .A2(n13991), .ZN(n13995) );
  INV_X1 U15783 ( .A(n13995), .ZN(n13993) );
  NAND2_X1 U15784 ( .A1(n13994), .A2(n13993), .ZN(n13998) );
  INV_X1 U15785 ( .A(n13994), .ZN(n13996) );
  OAI21_X1 U15786 ( .B1(n14069), .B2(n13996), .A(n13995), .ZN(n13997) );
  OAI21_X1 U15787 ( .B1(n13998), .B2(n19264), .A(n13997), .ZN(n17276) );
  INV_X1 U15788 ( .A(n13998), .ZN(n14018) );
  AOI22_X1 U15789 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14007) );
  AOI22_X1 U15790 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U15791 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11255), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14005) );
  INV_X1 U15792 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14002) );
  INV_X1 U15793 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14000) );
  OR2_X1 U15794 ( .A1(n14169), .A2(n14000), .ZN(n14001) );
  OAI211_X1 U15795 ( .C1(n15285), .C2(n14002), .A(n14001), .B(n14167), .ZN(
        n14003) );
  INV_X1 U15796 ( .A(n14003), .ZN(n14004) );
  NAND4_X1 U15797 ( .A1(n14007), .A2(n14006), .A3(n14005), .A4(n14004), .ZN(
        n14017) );
  AOI22_X1 U15798 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14015) );
  AOI22_X1 U15799 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14014) );
  AOI22_X1 U15800 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14013) );
  INV_X1 U15801 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14008) );
  OR2_X1 U15802 ( .A1(n14169), .A2(n14008), .ZN(n14009) );
  OAI211_X1 U15803 ( .C1(n15285), .C2(n14010), .A(n14104), .B(n14009), .ZN(
        n14011) );
  INV_X1 U15804 ( .A(n14011), .ZN(n14012) );
  NAND4_X1 U15805 ( .A1(n14015), .A2(n14014), .A3(n14013), .A4(n14012), .ZN(
        n14016) );
  AND2_X1 U15806 ( .A1(n14017), .A2(n14016), .ZN(n14020) );
  NAND2_X1 U15807 ( .A1(n14018), .A2(n14020), .ZN(n14066) );
  OAI211_X1 U15808 ( .C1(n14018), .C2(n14020), .A(n14042), .B(n14066), .ZN(
        n14022) );
  NAND2_X1 U15809 ( .A1(n19264), .A2(n14020), .ZN(n17268) );
  AOI22_X1 U15810 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14031) );
  AOI22_X1 U15811 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U15812 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14029) );
  OR2_X1 U15813 ( .A1(n14169), .A2(n14025), .ZN(n14026) );
  OAI211_X1 U15814 ( .C1(n11256), .C2(n12469), .A(n14026), .B(n14167), .ZN(
        n14027) );
  INV_X1 U15815 ( .A(n14027), .ZN(n14028) );
  NAND4_X1 U15816 ( .A1(n14031), .A2(n14030), .A3(n14029), .A4(n14028), .ZN(
        n14041) );
  AOI22_X1 U15817 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U15818 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14038) );
  AOI22_X1 U15819 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14037) );
  OR2_X1 U15820 ( .A1(n14169), .A2(n14032), .ZN(n14033) );
  OAI211_X1 U15821 ( .C1(n11257), .C2(n14034), .A(n14104), .B(n14033), .ZN(
        n14035) );
  INV_X1 U15822 ( .A(n14035), .ZN(n14036) );
  NAND4_X1 U15823 ( .A1(n14039), .A2(n14038), .A3(n14037), .A4(n14036), .ZN(
        n14040) );
  AND2_X1 U15824 ( .A1(n14041), .A2(n14040), .ZN(n14067) );
  XNOR2_X1 U15825 ( .A(n14066), .B(n14067), .ZN(n14043) );
  XNOR2_X1 U15826 ( .A(n14045), .B(n11350), .ZN(n17256) );
  INV_X1 U15827 ( .A(n14067), .ZN(n14044) );
  NOR2_X1 U15828 ( .A1(n11259), .A2(n14044), .ZN(n17258) );
  NAND2_X1 U15829 ( .A1(n17256), .A2(n17258), .ZN(n17257) );
  INV_X1 U15830 ( .A(n14045), .ZN(n14046) );
  AOI22_X1 U15831 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U15832 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U15833 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14053) );
  OR2_X1 U15834 ( .A1(n14169), .A2(n14048), .ZN(n14049) );
  OAI211_X1 U15835 ( .C1(n15285), .C2(n14050), .A(n14049), .B(n14167), .ZN(
        n14051) );
  INV_X1 U15836 ( .A(n14051), .ZN(n14052) );
  NAND4_X1 U15837 ( .A1(n14055), .A2(n14054), .A3(n14053), .A4(n14052), .ZN(
        n14065) );
  AOI22_X1 U15838 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U15839 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U15840 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11994), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14061) );
  INV_X1 U15841 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14056) );
  OR2_X1 U15842 ( .A1(n14169), .A2(n14056), .ZN(n14057) );
  OAI211_X1 U15843 ( .C1(n15285), .C2(n14058), .A(n14104), .B(n14057), .ZN(
        n14059) );
  INV_X1 U15844 ( .A(n14059), .ZN(n14060) );
  NAND4_X1 U15845 ( .A1(n14063), .A2(n14062), .A3(n14061), .A4(n14060), .ZN(
        n14064) );
  NAND2_X1 U15846 ( .A1(n14065), .A2(n14064), .ZN(n14091) );
  INV_X1 U15847 ( .A(n14066), .ZN(n14068) );
  NAND2_X1 U15848 ( .A1(n14068), .A2(n14067), .ZN(n14070) );
  NOR2_X1 U15849 ( .A1(n14070), .A2(n14091), .ZN(n17245) );
  NOR2_X1 U15850 ( .A1(n14090), .A2(n14089), .ZN(n17250) );
  AOI22_X1 U15851 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U15852 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U15853 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14076) );
  OR2_X1 U15854 ( .A1(n14169), .A2(n14071), .ZN(n14072) );
  OAI211_X1 U15855 ( .C1(n15285), .C2(n14073), .A(n14072), .B(n14167), .ZN(
        n14074) );
  INV_X1 U15856 ( .A(n14074), .ZN(n14075) );
  NAND4_X1 U15857 ( .A1(n14078), .A2(n14077), .A3(n14076), .A4(n14075), .ZN(
        n14088) );
  AOI22_X1 U15858 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U15859 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14085) );
  AOI22_X1 U15860 ( .A1(n14175), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14084) );
  OR2_X1 U15861 ( .A1(n14169), .A2(n14079), .ZN(n14080) );
  OAI211_X1 U15862 ( .C1(n15285), .C2(n14081), .A(n14104), .B(n14080), .ZN(
        n14082) );
  INV_X1 U15863 ( .A(n14082), .ZN(n14083) );
  NAND4_X1 U15864 ( .A1(n14086), .A2(n14085), .A3(n14084), .A4(n14083), .ZN(
        n14087) );
  NAND2_X1 U15865 ( .A1(n14088), .A2(n14087), .ZN(n14118) );
  NOR2_X1 U15866 ( .A1(n17250), .A2(n14118), .ZN(n14094) );
  NAND2_X1 U15867 ( .A1(n14090), .A2(n14089), .ZN(n17244) );
  INV_X1 U15868 ( .A(n14091), .ZN(n14092) );
  NAND2_X1 U15869 ( .A1(n19264), .A2(n14092), .ZN(n17252) );
  OAI21_X1 U15870 ( .B1(n14169), .B2(n14095), .A(n14167), .ZN(n14100) );
  OAI22_X1 U15871 ( .A1(n14096), .A2(n14098), .B1(n11258), .B2(n14097), .ZN(
        n14099) );
  AOI211_X1 U15872 ( .C1(n11996), .C2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n14100), .B(n14099), .ZN(n14103) );
  AOI22_X1 U15873 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U15874 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14101) );
  NAND3_X1 U15875 ( .A1(n14103), .A2(n14102), .A3(n14101), .ZN(n14114) );
  INV_X1 U15876 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14105) );
  OAI21_X1 U15877 ( .B1(n14169), .B2(n14105), .A(n14104), .ZN(n14109) );
  OAI22_X1 U15878 ( .A1(n14096), .A2(n14107), .B1(n15285), .B2(n14106), .ZN(
        n14108) );
  AOI211_X1 U15879 ( .C1(n14160), .C2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n14109), .B(n14108), .ZN(n14112) );
  AOI22_X1 U15880 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U15881 ( .A1(n14176), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11255), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14110) );
  NAND3_X1 U15882 ( .A1(n14112), .A2(n14111), .A3(n14110), .ZN(n14113) );
  NOR2_X1 U15883 ( .A1(n14116), .A2(n14115), .ZN(n14159) );
  NOR2_X1 U15884 ( .A1(n14117), .A2(n14159), .ZN(n14119) );
  INV_X1 U15885 ( .A(n14118), .ZN(n17246) );
  NAND3_X1 U15886 ( .A1(n17245), .A2(n17246), .A3(n11259), .ZN(n14158) );
  XNOR2_X1 U15887 ( .A(n14119), .B(n14158), .ZN(n14150) );
  AND2_X1 U15888 ( .A1(n12829), .A2(n22445), .ZN(n15335) );
  NAND2_X1 U15889 ( .A1(n15337), .A2(n15335), .ZN(n14120) );
  NOR2_X1 U15890 ( .A1(n15339), .A2(n14120), .ZN(n14121) );
  AOI21_X1 U15891 ( .B1(n15764), .B2(n14122), .A(n14121), .ZN(n15279) );
  NAND2_X1 U15892 ( .A1(n15279), .A2(n14123), .ZN(n14124) );
  NAND2_X1 U15893 ( .A1(n14150), .A2(n20551), .ZN(n14146) );
  OAI21_X1 U15894 ( .B1(n14127), .B2(n14126), .A(n16039), .ZN(n19479) );
  NOR2_X1 U15895 ( .A1(n20087), .A2(n13801), .ZN(n14128) );
  NOR4_X1 U15896 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14132) );
  NOR4_X1 U15897 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14131) );
  NOR4_X1 U15898 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14130) );
  NOR4_X1 U15899 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14129) );
  NAND4_X1 U15900 ( .A1(n14132), .A2(n14131), .A3(n14130), .A4(n14129), .ZN(
        n14137) );
  NOR4_X1 U15901 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n14135) );
  NOR4_X1 U15902 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14134) );
  NOR4_X1 U15903 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14133) );
  NAND4_X1 U15904 ( .A1(n14135), .A2(n14134), .A3(n14133), .A4(n20675), .ZN(
        n14136) );
  NAND2_X1 U15905 ( .A1(n20546), .A2(n14139), .ZN(n17404) );
  AOI22_X1 U15906 ( .A1(n15777), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n15776), .ZN(n20061) );
  INV_X1 U15907 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14869) );
  OAI22_X1 U15908 ( .A1(n17404), .A2(n20061), .B1(n20546), .B2(n14869), .ZN(
        n14142) );
  INV_X1 U15909 ( .A(n20048), .ZN(n17355) );
  INV_X1 U15910 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n14140) );
  NOR2_X1 U15911 ( .A1(n17355), .A2(n14140), .ZN(n14141) );
  AOI211_X1 U15912 ( .C1(BUF1_REG_29__SCAN_IN), .C2(n20050), .A(n14142), .B(
        n14141), .ZN(n14143) );
  NAND2_X1 U15913 ( .A1(n14146), .A2(n14145), .ZN(P2_U2890) );
  INV_X1 U15914 ( .A(n15764), .ZN(n14147) );
  NAND2_X1 U15915 ( .A1(n14147), .A2(n15330), .ZN(n15278) );
  INV_X1 U15916 ( .A(n14148), .ZN(n15260) );
  NAND2_X1 U15917 ( .A1(n15278), .A2(n15260), .ZN(n14149) );
  NAND2_X1 U15918 ( .A1(n14150), .A2(n17303), .ZN(n14156) );
  OAI21_X1 U15919 ( .B1(n14152), .B2(n14151), .A(n12203), .ZN(n19480) );
  NAND2_X1 U15920 ( .A1(n15680), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14153) );
  NAND2_X1 U15921 ( .A1(n14156), .A2(n14155), .ZN(P2_U2858) );
  OAI21_X1 U15922 ( .B1(n14159), .B2(n14158), .A(n14157), .ZN(n14185) );
  AOI22_X1 U15923 ( .A1(n11992), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U15924 ( .A1(n14160), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14161) );
  NAND2_X1 U15925 ( .A1(n14162), .A2(n14161), .ZN(n14183) );
  INV_X1 U15926 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14166) );
  AOI22_X1 U15927 ( .A1(n11255), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14165) );
  AOI21_X1 U15928 ( .B1(n14163), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n14167), .ZN(n14164) );
  OAI211_X1 U15929 ( .C1(n14096), .C2(n14166), .A(n14165), .B(n14164), .ZN(
        n14182) );
  INV_X1 U15930 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14168) );
  OAI21_X1 U15931 ( .B1(n14169), .B2(n14168), .A(n14167), .ZN(n14174) );
  INV_X1 U15932 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14172) );
  INV_X1 U15933 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14171) );
  OAI22_X1 U15934 ( .A1(n11247), .A2(n14172), .B1(n15285), .B2(n14171), .ZN(
        n14173) );
  AOI211_X1 U15935 ( .C1(n14175), .C2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n14174), .B(n14173), .ZN(n14180) );
  AOI22_X1 U15936 ( .A1(n11784), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14176), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14179) );
  AOI22_X1 U15937 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14177), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14178) );
  NAND3_X1 U15938 ( .A1(n14180), .A2(n14179), .A3(n14178), .ZN(n14181) );
  OAI21_X1 U15939 ( .B1(n14183), .B2(n14182), .A(n14181), .ZN(n14184) );
  XNOR2_X1 U15940 ( .A(n14185), .B(n14184), .ZN(n16079) );
  NAND2_X1 U15941 ( .A1(n16079), .A2(n17303), .ZN(n14189) );
  NAND2_X1 U15942 ( .A1(n15680), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14186) );
  NAND2_X1 U15943 ( .A1(n14189), .A2(n14188), .ZN(P2_U2857) );
  INV_X1 U15944 ( .A(n14722), .ZN(n14191) );
  NAND2_X1 U15945 ( .A1(n14783), .A2(n14191), .ZN(n14200) );
  AND2_X1 U15946 ( .A1(n14193), .A2(n14192), .ZN(n14194) );
  NAND2_X1 U15947 ( .A1(n14195), .A2(n14194), .ZN(n14196) );
  AND2_X1 U15948 ( .A1(n14197), .A2(n14196), .ZN(n16098) );
  NAND2_X1 U15949 ( .A1(n14927), .A2(n16106), .ZN(n14199) );
  NAND2_X1 U15950 ( .A1(n22388), .A2(n22556), .ZN(n18051) );
  OAI22_X1 U15951 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .B1(n18051), .B2(n22393), .ZN(n14203) );
  INV_X1 U15952 ( .A(n17977), .ZN(n17175) );
  NAND3_X1 U15953 ( .A1(n17175), .A2(n22392), .A3(n14201), .ZN(n14202) );
  AND2_X1 U15954 ( .A1(n14203), .A2(n14202), .ZN(n14204) );
  INV_X1 U15955 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14895) );
  INV_X1 U15956 ( .A(n14206), .ZN(n15007) );
  NAND2_X1 U15957 ( .A1(n14895), .A2(n16495), .ZN(n14208) );
  MUX2_X1 U15958 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n14207) );
  NAND2_X1 U15959 ( .A1(n14208), .A2(n14207), .ZN(n14210) );
  MUX2_X1 U15960 ( .A(n14293), .B(n14295), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n14849) );
  INV_X1 U15961 ( .A(n14849), .ZN(n14209) );
  XNOR2_X1 U15962 ( .A(n14210), .B(n14209), .ZN(n14778) );
  AOI21_X1 U15963 ( .B1(n14778), .B2(n11155), .A(n14210), .ZN(n14893) );
  INV_X1 U15964 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n22228) );
  NAND2_X1 U15965 ( .A1(n14292), .A2(n22228), .ZN(n14214) );
  NAND2_X1 U15966 ( .A1(n11155), .A2(n22228), .ZN(n14212) );
  NAND2_X1 U15967 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14211) );
  NAND3_X1 U15968 ( .A1(n14212), .A2(n14295), .A3(n14211), .ZN(n14213) );
  AND2_X1 U15969 ( .A1(n14214), .A2(n14213), .ZN(n14892) );
  INV_X1 U15970 ( .A(n14215), .ZN(n16496) );
  OR2_X1 U15971 ( .A1(n14301), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n14221) );
  NAND2_X1 U15972 ( .A1(n14295), .A2(n14216), .ZN(n14219) );
  INV_X1 U15973 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14217) );
  NAND2_X1 U15974 ( .A1(n11155), .A2(n14217), .ZN(n14218) );
  NAND3_X1 U15975 ( .A1(n14219), .A2(n14293), .A3(n14218), .ZN(n14220) );
  NAND2_X1 U15976 ( .A1(n14221), .A2(n14220), .ZN(n14975) );
  NAND2_X1 U15977 ( .A1(n14976), .A2(n14975), .ZN(n15115) );
  MUX2_X1 U15978 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n14222) );
  OAI21_X1 U15979 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16499), .A(
        n14222), .ZN(n15114) );
  MUX2_X1 U15980 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n14224) );
  OR2_X1 U15981 ( .A1(n16499), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14223) );
  NAND2_X1 U15982 ( .A1(n14224), .A2(n14223), .ZN(n15540) );
  INV_X1 U15983 ( .A(n15540), .ZN(n14229) );
  MUX2_X1 U15984 ( .A(n14301), .B(n14295), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n14228) );
  INV_X1 U15985 ( .A(n14295), .ZN(n14225) );
  NAND2_X1 U15986 ( .A1(n14225), .A2(n16498), .ZN(n14273) );
  NAND2_X1 U15987 ( .A1(n16498), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14226) );
  AND2_X1 U15988 ( .A1(n14273), .A2(n14226), .ZN(n14227) );
  NAND2_X1 U15989 ( .A1(n14228), .A2(n14227), .ZN(n15483) );
  NAND2_X1 U15990 ( .A1(n14229), .A2(n15483), .ZN(n14230) );
  NOR2_X1 U15991 ( .A1(n15542), .A2(n14230), .ZN(n15595) );
  MUX2_X1 U15992 ( .A(n14301), .B(n14295), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n14233) );
  NAND2_X1 U15993 ( .A1(n16498), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14231) );
  AND2_X1 U15994 ( .A1(n14273), .A2(n14231), .ZN(n14232) );
  NAND2_X1 U15995 ( .A1(n14233), .A2(n14232), .ZN(n15594) );
  MUX2_X1 U15996 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n14235) );
  OR2_X1 U15997 ( .A1(n16499), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14234) );
  NAND2_X1 U15998 ( .A1(n14235), .A2(n14234), .ZN(n15653) );
  INV_X1 U15999 ( .A(n15653), .ZN(n14236) );
  OR2_X1 U16000 ( .A1(n14301), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n14240) );
  NAND2_X1 U16001 ( .A1(n14295), .A2(n17144), .ZN(n14238) );
  INV_X1 U16002 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n16682) );
  NAND2_X1 U16003 ( .A1(n11155), .A2(n16682), .ZN(n14237) );
  NAND3_X1 U16004 ( .A1(n14238), .A2(n14293), .A3(n14237), .ZN(n14239) );
  INV_X1 U16005 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n20819) );
  NAND2_X1 U16006 ( .A1(n11155), .A2(n20819), .ZN(n14242) );
  NAND2_X1 U16007 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14241) );
  NAND3_X1 U16008 ( .A1(n14242), .A2(n14295), .A3(n14241), .ZN(n14243) );
  OAI21_X1 U16009 ( .B1(n14286), .B2(P1_EBX_REG_10__SCAN_IN), .A(n14243), .ZN(
        n15855) );
  MUX2_X1 U16010 ( .A(n14301), .B(n14295), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n14246) );
  NAND2_X1 U16011 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16498), .ZN(
        n14244) );
  AND2_X1 U16012 ( .A1(n14273), .A2(n14244), .ZN(n14245) );
  NAND2_X1 U16013 ( .A1(n14246), .A2(n14245), .ZN(n17117) );
  INV_X1 U16014 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n20815) );
  NAND2_X1 U16015 ( .A1(n14292), .A2(n20815), .ZN(n14250) );
  NAND2_X1 U16016 ( .A1(n11155), .A2(n20815), .ZN(n14248) );
  NAND2_X1 U16017 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14247) );
  NAND3_X1 U16018 ( .A1(n14248), .A2(n14295), .A3(n14247), .ZN(n14249) );
  AND2_X1 U16019 ( .A1(n14250), .A2(n14249), .ZN(n17116) );
  OR2_X1 U16020 ( .A1(n14301), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n14254) );
  NAND2_X1 U16021 ( .A1(n14295), .A2(n22138), .ZN(n14252) );
  INV_X1 U16022 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n16739) );
  NAND2_X1 U16023 ( .A1(n11155), .A2(n16739), .ZN(n14251) );
  NAND3_X1 U16024 ( .A1(n14252), .A2(n14293), .A3(n14251), .ZN(n14253) );
  NAND2_X1 U16025 ( .A1(n14254), .A2(n14253), .ZN(n16664) );
  NAND2_X1 U16026 ( .A1(n17119), .A2(n16664), .ZN(n16666) );
  MUX2_X1 U16027 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n14255) );
  OAI21_X1 U16028 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16499), .A(
        n14255), .ZN(n15944) );
  OR2_X1 U16029 ( .A1(n14301), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U16030 ( .A1(n14295), .A2(n14256), .ZN(n14258) );
  INV_X1 U16031 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n16738) );
  NAND2_X1 U16032 ( .A1(n11155), .A2(n16738), .ZN(n14257) );
  NAND3_X1 U16033 ( .A1(n14258), .A2(n14293), .A3(n14257), .ZN(n14259) );
  INV_X1 U16034 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16731) );
  NAND2_X1 U16035 ( .A1(n14292), .A2(n16731), .ZN(n14264) );
  NAND2_X1 U16036 ( .A1(n11155), .A2(n16731), .ZN(n14262) );
  NAND2_X1 U16037 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14261) );
  NAND3_X1 U16038 ( .A1(n14262), .A2(n14295), .A3(n14261), .ZN(n14263) );
  OR2_X1 U16039 ( .A1(n14301), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14268) );
  NAND2_X1 U16040 ( .A1(n14295), .A2(n17108), .ZN(n14266) );
  INV_X1 U16041 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n20824) );
  NAND2_X1 U16042 ( .A1(n11155), .A2(n20824), .ZN(n14265) );
  NAND3_X1 U16043 ( .A1(n14266), .A2(n14293), .A3(n14265), .ZN(n14267) );
  MUX2_X1 U16044 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n14270) );
  OR2_X1 U16045 ( .A1(n16499), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14269) );
  NAND2_X1 U16046 ( .A1(n14270), .A2(n14269), .ZN(n16626) );
  NOR2_X1 U16047 ( .A1(n16636), .A2(n16626), .ZN(n14271) );
  MUX2_X1 U16048 ( .A(n14301), .B(n14295), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14274) );
  NAND2_X1 U16049 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16498), .ZN(
        n14272) );
  MUX2_X1 U16050 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14275) );
  OAI21_X1 U16051 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n16499), .A(
        n14275), .ZN(n16614) );
  MUX2_X1 U16052 ( .A(n14301), .B(n14295), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14277) );
  NAND2_X1 U16053 ( .A1(n16498), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14276) );
  NAND2_X1 U16054 ( .A1(n14277), .A2(n14276), .ZN(n16719) );
  NAND2_X1 U16055 ( .A1(n16720), .A2(n16719), .ZN(n16718) );
  MUX2_X1 U16056 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14278) );
  OAI21_X1 U16057 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16499), .A(
        n14278), .ZN(n16601) );
  OR2_X1 U16058 ( .A1(n14301), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n14282) );
  INV_X1 U16059 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17052) );
  NAND2_X1 U16060 ( .A1(n14295), .A2(n17052), .ZN(n14280) );
  INV_X1 U16061 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n16435) );
  NAND2_X1 U16062 ( .A1(n11155), .A2(n16435), .ZN(n14279) );
  NAND3_X1 U16063 ( .A1(n14280), .A2(n14293), .A3(n14279), .ZN(n14281) );
  MUX2_X1 U16064 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14283) );
  OAI21_X1 U16065 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16499), .A(
        n14283), .ZN(n16581) );
  MUX2_X1 U16066 ( .A(n14301), .B(n14295), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14285) );
  NAND2_X1 U16067 ( .A1(n16498), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14284) );
  NAND2_X1 U16068 ( .A1(n14285), .A2(n14284), .ZN(n16562) );
  NAND2_X1 U16069 ( .A1(n16580), .A2(n16562), .ZN(n16561) );
  MUX2_X1 U16070 ( .A(n14286), .B(n14293), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14287) );
  OAI21_X1 U16071 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n16499), .A(
        n14287), .ZN(n16558) );
  OR2_X1 U16072 ( .A1(n14301), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14291) );
  INV_X1 U16073 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17024) );
  NAND2_X1 U16074 ( .A1(n14295), .A2(n17024), .ZN(n14289) );
  INV_X1 U16075 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n16427) );
  NAND2_X1 U16076 ( .A1(n11155), .A2(n16427), .ZN(n14288) );
  NAND3_X1 U16077 ( .A1(n14289), .A2(n14293), .A3(n14288), .ZN(n14290) );
  INV_X1 U16078 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n16709) );
  NAND2_X1 U16079 ( .A1(n14292), .A2(n16709), .ZN(n14298) );
  NAND2_X1 U16080 ( .A1(n11155), .A2(n16709), .ZN(n14296) );
  NAND2_X1 U16081 ( .A1(n14293), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14294) );
  NAND3_X1 U16082 ( .A1(n14296), .A2(n14295), .A3(n14294), .ZN(n14297) );
  AND2_X1 U16083 ( .A1(n14298), .A2(n14297), .ZN(n16528) );
  OR2_X1 U16084 ( .A1(n16499), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14300) );
  INV_X1 U16085 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16708) );
  NAND2_X1 U16086 ( .A1(n11155), .A2(n16708), .ZN(n14299) );
  NAND2_X1 U16087 ( .A1(n14300), .A2(n14299), .ZN(n16511) );
  OAI22_X1 U16088 ( .A1(n16511), .A2(n16496), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14301), .ZN(n14302) );
  OR2_X1 U16089 ( .A1(n16530), .A2(n14302), .ZN(n14303) );
  NAND2_X1 U16090 ( .A1(n16497), .A2(n14303), .ZN(n17008) );
  OR2_X1 U16091 ( .A1(n16691), .A2(n13044), .ZN(n14313) );
  NAND2_X1 U16092 ( .A1(n22424), .A2(n22405), .ZN(n14306) );
  NAND3_X1 U16093 ( .A1(n14784), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n14306), 
        .ZN(n14304) );
  OR2_X1 U16094 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n14305), .ZN(n22434) );
  NAND2_X1 U16095 ( .A1(n14986), .A2(n22434), .ZN(n14694) );
  INV_X1 U16096 ( .A(n14306), .ZN(n18043) );
  NAND2_X1 U16097 ( .A1(n14694), .A2(n18043), .ZN(n14311) );
  INV_X1 U16098 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20771) );
  INV_X1 U16099 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20757) );
  INV_X1 U16100 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20753) );
  INV_X1 U16101 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20749) );
  INV_X1 U16102 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n22284) );
  INV_X1 U16103 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22296) );
  INV_X1 U16104 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20743) );
  NAND3_X1 U16105 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n22253) );
  NOR2_X1 U16106 ( .A1(n20743), .A2(n22253), .ZN(n22272) );
  NAND2_X1 U16107 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22272), .ZN(n22285) );
  NOR4_X1 U16108 ( .A1(n20749), .A2(n22284), .A3(n22296), .A4(n22285), .ZN(
        n16678) );
  NAND2_X1 U16109 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n16678), .ZN(n15854) );
  NOR2_X1 U16110 ( .A1(n20753), .A2(n15854), .ZN(n22312) );
  NAND2_X1 U16111 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22312), .ZN(n22322) );
  NOR2_X1 U16112 ( .A1(n20757), .A2(n22322), .ZN(n16669) );
  NAND2_X1 U16113 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16669), .ZN(n16668) );
  INV_X1 U16114 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20765) );
  INV_X1 U16115 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20764) );
  INV_X1 U16116 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20762) );
  INV_X1 U16117 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20760) );
  NOR4_X1 U16118 ( .A1(n20765), .A2(n20764), .A3(n20762), .A4(n20760), .ZN(
        n14307) );
  NAND3_X1 U16119 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(n14307), .ZN(n16606) );
  NOR3_X1 U16120 ( .A1(n20771), .A2(n16668), .A3(n16606), .ZN(n22370) );
  AND3_X1 U16121 ( .A1(n22370), .A2(P1_REIP_REG_21__SCAN_IN), .A3(
        P1_REIP_REG_22__SCAN_IN), .ZN(n14308) );
  NAND2_X1 U16122 ( .A1(n22248), .A2(n14308), .ZN(n16590) );
  INV_X1 U16123 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20777) );
  NAND2_X1 U16124 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14309) );
  INV_X1 U16125 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20784) );
  NOR2_X1 U16126 ( .A1(n16569), .A2(n20784), .ZN(n16553) );
  NAND2_X1 U16127 ( .A1(n16553), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16541) );
  INV_X1 U16128 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20787) );
  NAND2_X1 U16129 ( .A1(n14784), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U16130 ( .A1(n14311), .A2(n14310), .ZN(n14312) );
  NOR2_X2 U16131 ( .A1(n14313), .A2(n14312), .ZN(n22358) );
  INV_X1 U16132 ( .A(n22255), .ZN(n22238) );
  NAND3_X1 U16133 ( .A1(n16534), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n22339), 
        .ZN(n14318) );
  AND2_X2 U16134 ( .A1(n22255), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22371) );
  INV_X1 U16135 ( .A(n16852), .ZN(n14316) );
  AOI22_X1 U16136 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n22371), .B1(
        n22353), .B2(n14316), .ZN(n14317) );
  OAI211_X1 U16137 ( .C1(n16708), .C2(n22374), .A(n14318), .B(n14317), .ZN(
        n14319) );
  INV_X1 U16138 ( .A(n14319), .ZN(n14320) );
  NAND4_X1 U16139 ( .A1(n11303), .A2(n11712), .A3(n11713), .A4(n14320), .ZN(
        P1_U2811) );
  NOR2_X1 U16140 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14322) );
  NOR4_X1 U16141 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14321) );
  NAND4_X1 U16142 ( .A1(n14322), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14321), .ZN(n14335) );
  NOR4_X1 U16143 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n14326) );
  NOR4_X1 U16144 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n14325) );
  NOR4_X1 U16145 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n14324) );
  NOR4_X1 U16146 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14323) );
  NAND4_X1 U16147 ( .A1(n14326), .A2(n14325), .A3(n14324), .A4(n14323), .ZN(
        n14331) );
  NOR4_X1 U16148 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n14329) );
  NOR4_X1 U16149 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n14328) );
  NOR4_X1 U16150 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n14327) );
  NAND4_X1 U16151 ( .A1(n14329), .A2(n14328), .A3(n14327), .A4(n20738), .ZN(
        n14330) );
  INV_X1 U16152 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22853) );
  INV_X1 U16153 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20953) );
  NOR4_X1 U16154 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n22853), .A4(n20953), .ZN(n14334) );
  NOR4_X1 U16155 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14333) );
  NAND3_X1 U16156 ( .A1(n15793), .A2(n14334), .A3(n14333), .ZN(U214) );
  NOR2_X1 U16157 ( .A1(n15776), .A2(n14335), .ZN(n20884) );
  NAND2_X1 U16158 ( .A1(n20884), .A2(U214), .ZN(U212) );
  INV_X1 U16159 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19223) );
  NOR2_X1 U16160 ( .A1(n19223), .A2(n21687), .ZN(n21033) );
  INV_X1 U16161 ( .A(n18677), .ZN(n14336) );
  INV_X1 U16162 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18629) );
  AOI22_X1 U16163 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14338) );
  OAI21_X1 U16164 ( .B1(n14336), .B2(n18629), .A(n14338), .ZN(n14346) );
  AOI22_X1 U16165 ( .A1(n18658), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14344) );
  BUF_X4 U16166 ( .A(n14377), .Z(n18678) );
  AOI22_X1 U16167 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14343) );
  AOI22_X1 U16168 ( .A1(n18647), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14342) );
  INV_X2 U16169 ( .A(n11293), .ZN(n21043) );
  AOI22_X1 U16170 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14341) );
  NAND4_X1 U16171 ( .A1(n14344), .A2(n14343), .A3(n14342), .A4(n14341), .ZN(
        n14345) );
  INV_X1 U16172 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22463) );
  INV_X1 U16173 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n17980) );
  NOR2_X2 U16174 ( .A1(n22463), .A2(n22469), .ZN(n19254) );
  INV_X1 U16175 ( .A(n17989), .ZN(n20958) );
  NAND2_X1 U16176 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n22470) );
  AOI22_X1 U16177 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14353) );
  AOI22_X1 U16178 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18664), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14352) );
  AOI22_X1 U16179 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14351) );
  BUF_X4 U16180 ( .A(n18612), .Z(n18660) );
  AOI22_X1 U16181 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14350) );
  NAND4_X1 U16182 ( .A1(n14353), .A2(n14352), .A3(n14351), .A4(n14350), .ZN(
        n14359) );
  AOI22_X1 U16183 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U16184 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U16185 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14355) );
  CLKBUF_X3 U16186 ( .A(n18630), .Z(n18665) );
  AOI22_X1 U16187 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14354) );
  NAND4_X1 U16188 ( .A1(n14357), .A2(n14356), .A3(n14355), .A4(n14354), .ZN(
        n14358) );
  XNOR2_X1 U16189 ( .A(n14475), .B(n14476), .ZN(n14371) );
  AOI22_X1 U16190 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n19609), .B2(n14501), .ZN(
        n14365) );
  OAI21_X1 U16191 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14501), .A(
        n14361), .ZN(n14362) );
  OAI22_X1 U16192 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17987), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14362), .ZN(n14368) );
  NOR2_X1 U16193 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17987), .ZN(
        n14363) );
  NAND2_X1 U16194 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14362), .ZN(
        n14369) );
  AOI22_X1 U16195 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14368), .B1(
        n14363), .B2(n14369), .ZN(n14477) );
  OAI21_X1 U16196 ( .B1(n14366), .B2(n14365), .A(n14477), .ZN(n14364) );
  AOI21_X1 U16197 ( .B1(n14366), .B2(n14365), .A(n14364), .ZN(n14367) );
  AOI21_X1 U16198 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14369), .A(
        n14368), .ZN(n14370) );
  AOI22_X1 U16199 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U16200 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18630), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U16201 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14374) );
  AOI22_X1 U16202 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14373) );
  NAND4_X1 U16203 ( .A1(n14376), .A2(n14375), .A3(n14374), .A4(n14373), .ZN(
        n14383) );
  AOI22_X1 U16204 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14381) );
  AOI22_X1 U16205 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14380) );
  AOI22_X1 U16206 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14379) );
  AOI22_X1 U16207 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14378) );
  NAND4_X1 U16208 ( .A1(n14381), .A2(n14380), .A3(n14379), .A4(n14378), .ZN(
        n14382) );
  AOI22_X1 U16209 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14393) );
  AOI22_X1 U16210 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14392) );
  AOI22_X1 U16211 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14384) );
  OAI21_X1 U16212 ( .B1(n14336), .B2(n18402), .A(n14384), .ZN(n14390) );
  AOI22_X1 U16213 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U16214 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U16215 ( .A1(n18665), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14386) );
  AOI22_X1 U16216 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14385) );
  NAND4_X1 U16217 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14385), .ZN(
        n14389) );
  AOI22_X1 U16218 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U16219 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14396) );
  AOI22_X1 U16220 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14395) );
  AOI22_X1 U16221 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14394) );
  NAND4_X1 U16222 ( .A1(n14397), .A2(n14396), .A3(n14395), .A4(n14394), .ZN(
        n14403) );
  AOI22_X1 U16223 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U16224 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18630), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14400) );
  INV_X4 U16225 ( .A(n18496), .ZN(n18647) );
  AOI22_X1 U16226 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14399) );
  INV_X2 U16227 ( .A(n14336), .ZN(n18666) );
  AOI22_X1 U16228 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14398) );
  NAND4_X1 U16229 ( .A1(n14401), .A2(n14400), .A3(n14399), .A4(n14398), .ZN(
        n14402) );
  AOI22_X1 U16230 ( .A1(n18658), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18630), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U16231 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U16232 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U16233 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14405) );
  NAND4_X1 U16234 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        n14414) );
  AOI22_X1 U16235 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14412) );
  AOI22_X1 U16236 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14411) );
  AOI22_X1 U16237 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14410) );
  AOI22_X1 U16238 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14409) );
  NAND4_X1 U16239 ( .A1(n14412), .A2(n14411), .A3(n14410), .A4(n14409), .ZN(
        n14413) );
  NOR2_X1 U16240 ( .A1(n19819), .A2(n21648), .ZN(n14438) );
  AOI22_X1 U16241 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U16242 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U16243 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14416) );
  AOI22_X1 U16244 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14415) );
  NAND4_X1 U16245 ( .A1(n14418), .A2(n14417), .A3(n14416), .A4(n14415), .ZN(
        n14425) );
  AOI22_X1 U16246 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14423) );
  AOI22_X1 U16247 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18664), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14422) );
  AOI22_X1 U16248 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U16249 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14420) );
  NAND4_X1 U16250 ( .A1(n14423), .A2(n14422), .A3(n14421), .A4(n14420), .ZN(
        n14424) );
  INV_X1 U16251 ( .A(n21656), .ZN(n14443) );
  NOR2_X1 U16252 ( .A1(n14440), .A2(n14443), .ZN(n14466) );
  AOI22_X1 U16253 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14435) );
  AOI22_X1 U16254 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14434) );
  AOI22_X1 U16255 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14426) );
  OAI21_X1 U16256 ( .B1(n14336), .B2(n18662), .A(n14426), .ZN(n14432) );
  AOI22_X1 U16257 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14430) );
  AOI22_X1 U16258 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14429) );
  AOI22_X1 U16259 ( .A1(n18658), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U16260 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14427) );
  NAND4_X1 U16261 ( .A1(n14430), .A2(n14429), .A3(n14428), .A4(n14427), .ZN(
        n14431) );
  AOI211_X1 U16262 ( .C1(n18664), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n14432), .B(n14431), .ZN(n14433) );
  NAND3_X1 U16263 ( .A1(n14435), .A2(n14434), .A3(n14433), .ZN(n19698) );
  NAND2_X1 U16264 ( .A1(n19739), .A2(n19698), .ZN(n14467) );
  NAND2_X1 U16265 ( .A1(n14466), .A2(n14467), .ZN(n14437) );
  AOI21_X1 U16266 ( .B1(n19951), .B2(n21652), .A(n21439), .ZN(n14474) );
  NOR2_X1 U16267 ( .A1(n21656), .A2(n19698), .ZN(n14505) );
  NOR2_X1 U16268 ( .A1(n14474), .A2(n14505), .ZN(n14436) );
  AOI22_X1 U16269 ( .A1(n14438), .A2(n14437), .B1(n14436), .B2(n14467), .ZN(
        n14447) );
  NAND3_X1 U16270 ( .A1(n19739), .A2(n14489), .A3(n14447), .ZN(n14439) );
  NAND2_X1 U16271 ( .A1(n19951), .A2(n21533), .ZN(n14441) );
  INV_X1 U16272 ( .A(n14441), .ZN(n14448) );
  INV_X1 U16273 ( .A(n19739), .ZN(n21497) );
  NAND2_X1 U16274 ( .A1(n21497), .A2(n19698), .ZN(n21643) );
  INV_X1 U16275 ( .A(n21643), .ZN(n14444) );
  NAND4_X1 U16276 ( .A1(n19819), .A2(n21656), .A3(n14448), .A4(n14444), .ZN(
        n14488) );
  INV_X1 U16277 ( .A(n14488), .ZN(n14450) );
  NAND2_X1 U16278 ( .A1(n14450), .A2(n14440), .ZN(n14468) );
  NAND2_X1 U16279 ( .A1(n14468), .A2(n14439), .ZN(n18573) );
  OR2_X1 U16280 ( .A1(n14440), .A2(n14485), .ZN(n14470) );
  AOI22_X1 U16281 ( .A1(n19819), .A2(n14441), .B1(n21643), .B2(n14470), .ZN(
        n14446) );
  NOR2_X1 U16282 ( .A1(n19951), .A2(n21641), .ZN(n14486) );
  INV_X1 U16283 ( .A(n21439), .ZN(n14442) );
  NAND2_X1 U16284 ( .A1(n21533), .A2(n14442), .ZN(n21433) );
  NAND2_X1 U16285 ( .A1(n14486), .A2(n21433), .ZN(n14472) );
  OAI21_X1 U16286 ( .B1(n21435), .B2(n14444), .A(n14443), .ZN(n14445) );
  NAND4_X1 U16287 ( .A1(n14447), .A2(n14446), .A3(n14472), .A4(n14445), .ZN(
        n14516) );
  NAND2_X1 U16288 ( .A1(n21652), .A2(n19819), .ZN(n14509) );
  NOR2_X1 U16289 ( .A1(n14467), .A2(n14509), .ZN(n18200) );
  NAND3_X1 U16290 ( .A1(n20959), .A2(n14448), .A3(n18200), .ZN(n14499) );
  NAND2_X1 U16291 ( .A1(n14450), .A2(n14506), .ZN(n14495) );
  AOI211_X1 U16292 ( .C1(n19223), .C2(n21687), .A(n21033), .B(n21327), .ZN(
        n14465) );
  INV_X1 U16293 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18571) );
  INV_X1 U16294 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18566) );
  NAND2_X1 U16295 ( .A1(n18571), .A2(n18566), .ZN(n14452) );
  NOR3_X1 U16296 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n21038) );
  NAND2_X1 U16297 ( .A1(n22470), .A2(n22414), .ZN(n14451) );
  NAND4_X1 U16298 ( .A1(n14453), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n21641), 
        .A4(n14451), .ZN(n21397) );
  AOI211_X1 U16299 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n14452), .A(n21038), .B(
        n21397), .ZN(n14464) );
  INV_X1 U16300 ( .A(n14453), .ZN(n14454) );
  AOI211_X4 U16301 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n21641), .A(n14534), .B(
        n14454), .ZN(n21424) );
  INV_X1 U16302 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n18203) );
  INV_X1 U16303 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19130) );
  NOR2_X1 U16304 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n22088) );
  NAND2_X1 U16305 ( .A1(n22088), .A2(n22084), .ZN(n18577) );
  INV_X2 U16306 ( .A(n22057), .ZN(n22049) );
  NOR4_X1 U16307 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n21619), .ZN(n21249) );
  INV_X1 U16308 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21998) );
  NAND2_X1 U16309 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21998), .ZN(n19687) );
  AND2_X1 U16310 ( .A1(n14535), .A2(n19670), .ZN(n22090) );
  OAI22_X1 U16311 ( .A1(n21359), .A2(n18203), .B1(n19130), .B2(n21357), .ZN(
        n14463) );
  NAND4_X1 U16312 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19025) );
  NOR2_X1 U16313 ( .A1(n19025), .A2(n21149), .ZN(n18993) );
  NAND2_X1 U16314 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19104) );
  NAND2_X1 U16315 ( .A1(n19088), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19079) );
  NAND2_X1 U16316 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18995) );
  NAND2_X1 U16317 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n21229) );
  INV_X1 U16318 ( .A(n18890), .ZN(n18909) );
  INV_X1 U16319 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21358) );
  INV_X1 U16320 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14456) );
  INV_X1 U16321 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18953) );
  XNOR2_X2 U16322 ( .A(n14457), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n21214) );
  NAND2_X1 U16323 ( .A1(n11533), .A2(n21214), .ZN(n21171) );
  NOR2_X1 U16324 ( .A1(n19130), .A2(n21027), .ZN(n19114) );
  AOI21_X1 U16325 ( .B1(n19130), .B2(n21027), .A(n19114), .ZN(n14458) );
  INV_X1 U16326 ( .A(n14458), .ZN(n19127) );
  NOR2_X1 U16327 ( .A1(n21428), .A2(n20954), .ZN(n21421) );
  NAND2_X1 U16328 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n14522), .ZN(
        n21629) );
  NAND2_X1 U16329 ( .A1(n14459), .A2(n21629), .ZN(n14521) );
  AOI22_X1 U16330 ( .A1(n11262), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n21421), 
        .B2(n14521), .ZN(n14461) );
  NOR2_X1 U16331 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21027), .ZN(
        n21195) );
  INV_X1 U16332 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21113) );
  AOI21_X1 U16333 ( .B1(n19114), .B2(n21113), .A(n21214), .ZN(n21035) );
  OAI211_X1 U16334 ( .C1(n21195), .C2(n19127), .A(n21249), .B(n21035), .ZN(
        n14460) );
  OAI211_X1 U16335 ( .C1(n21171), .C2(n19127), .A(n14461), .B(n14460), .ZN(
        n14462) );
  OR4_X1 U16336 ( .A1(n14465), .A2(n14464), .A3(n14463), .A4(n14462), .ZN(
        P3_U2669) );
  NOR2_X1 U16337 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21998), .ZN(n18850) );
  INV_X1 U16338 ( .A(n18850), .ZN(n19143) );
  NOR2_X1 U16339 ( .A1(n22470), .A2(n20955), .ZN(n22086) );
  NOR4_X1 U16340 ( .A1(n21619), .A2(n22095), .A3(n22470), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17984) );
  INV_X1 U16341 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17972) );
  AOI21_X1 U16342 ( .B1(n17989), .B2(n17988), .A(n21429), .ZN(n14484) );
  NAND2_X1 U16343 ( .A1(n14494), .A2(n22470), .ZN(n14483) );
  INV_X1 U16344 ( .A(n14466), .ZN(n14473) );
  OAI211_X1 U16345 ( .C1(n21439), .C2(n21656), .A(n14489), .B(n14467), .ZN(
        n14469) );
  OAI21_X1 U16346 ( .B1(n14470), .B2(n14469), .A(n14468), .ZN(n14471) );
  OAI211_X1 U16347 ( .C1(n14474), .C2(n14473), .A(n14472), .B(n14471), .ZN(
        n21649) );
  INV_X1 U16348 ( .A(n21649), .ZN(n14482) );
  OAI21_X1 U16349 ( .B1(n19653), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n14475), .ZN(n14490) );
  INV_X1 U16350 ( .A(n14476), .ZN(n14478) );
  NAND2_X1 U16351 ( .A1(n14478), .A2(n14477), .ZN(n14480) );
  INV_X1 U16352 ( .A(n21654), .ZN(n14481) );
  NAND2_X1 U16353 ( .A1(n14481), .A2(n14487), .ZN(n18202) );
  OR2_X1 U16354 ( .A1(n20959), .A2(n14489), .ZN(n14507) );
  NOR2_X4 U16355 ( .A1(n21641), .A2(n21979), .ZN(n21964) );
  OAI21_X1 U16356 ( .B1(n14491), .B2(n14490), .A(n14494), .ZN(n14496) );
  INV_X1 U16357 ( .A(n14496), .ZN(n21642) );
  AOI221_X1 U16358 ( .B1(n14494), .B2(n21657), .C1(n14500), .C2(n21657), .A(
        n21642), .ZN(n14492) );
  INV_X1 U16359 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n22102) );
  INV_X1 U16360 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n22099) );
  XOR2_X1 U16361 ( .A(n20959), .B(n21652), .Z(n14493) );
  OAI21_X1 U16362 ( .B1(n14493), .B2(n17989), .A(n22470), .ZN(n21646) );
  NAND3_X1 U16363 ( .A1(n14494), .A2(n21646), .A3(n18573), .ZN(n22096) );
  AOI21_X1 U16364 ( .B1(n22102), .B2(n22099), .A(n22096), .ZN(n14532) );
  AOI21_X1 U16365 ( .B1(n17963), .B2(n17972), .A(n14495), .ZN(n17970) );
  INV_X1 U16366 ( .A(n17969), .ZN(n14527) );
  NAND2_X1 U16367 ( .A1(n14500), .A2(n14499), .ZN(n22071) );
  AOI21_X1 U16368 ( .B1(n21892), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n22071), .ZN(n14524) );
  OR2_X1 U16369 ( .A1(n21624), .A2(n14524), .ZN(n14519) );
  AND2_X1 U16370 ( .A1(n14501), .A2(n14522), .ZN(n14502) );
  XNOR2_X1 U16371 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14502), .ZN(
        n14504) );
  NOR2_X1 U16372 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21638), .ZN(
        n14503) );
  AOI22_X1 U16373 ( .A1(n22016), .A2(n14504), .B1(n14503), .B2(n14516), .ZN(
        n14514) );
  AOI21_X1 U16374 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n21638), .ZN(n14512) );
  INV_X1 U16375 ( .A(n14505), .ZN(n14510) );
  INV_X1 U16376 ( .A(n14506), .ZN(n14508) );
  OAI22_X1 U16377 ( .A1(n14510), .A2(n14509), .B1(n14508), .B2(n14507), .ZN(
        n14517) );
  AOI21_X1 U16378 ( .B1(n21618), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14512), .ZN(n14511) );
  INV_X1 U16379 ( .A(n14511), .ZN(n21031) );
  AOI22_X1 U16380 ( .A1(n14512), .A2(n14518), .B1(n14517), .B2(n21031), .ZN(
        n14513) );
  OAI211_X1 U16381 ( .C1(n14515), .C2(n14519), .A(n14514), .B(n14513), .ZN(
        n21633) );
  AOI22_X1 U16382 ( .A1(n14527), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21633), .B2(n17969), .ZN(n14531) );
  AOI211_X1 U16383 ( .C1(n14518), .C2(n21624), .A(n14517), .B(n14516), .ZN(
        n14520) );
  OAI222_X1 U16384 ( .A1(n21894), .A2(n14521), .B1(n21629), .B2(n14520), .C1(
        n14519), .C2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21628) );
  MUX2_X1 U16385 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n21628), .S(
        n17969), .Z(n14529) );
  INV_X1 U16386 ( .A(n22071), .ZN(n22059) );
  NOR2_X1 U16387 ( .A1(n21439), .A2(n21892), .ZN(n14525) );
  NAND2_X1 U16388 ( .A1(n14523), .A2(n14522), .ZN(n21023) );
  OAI22_X1 U16389 ( .A1(n14525), .A2(n21023), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n14524), .ZN(n21622) );
  NAND2_X1 U16390 ( .A1(n19636), .A2(n19653), .ZN(n19671) );
  OAI21_X1 U16391 ( .B1(n14527), .B2(n14526), .A(n19671), .ZN(n14528) );
  INV_X1 U16392 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19631) );
  AOI21_X1 U16393 ( .B1(n17987), .B2(n19631), .A(n14529), .ZN(n14530) );
  OAI211_X1 U16394 ( .C1(n17972), .C2(n17969), .A(n22100), .B(n14533), .ZN(
        n22091) );
  OAI21_X1 U16395 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n20254), .A(n14547), 
        .ZN(n14538) );
  AOI21_X1 U16396 ( .B1(P2_MEMORYFETCH_REG_SCAN_IN), .B2(n17240), .A(n14538), 
        .ZN(n14536) );
  INV_X1 U16397 ( .A(n14536), .ZN(P2_U2814) );
  INV_X1 U16398 ( .A(n17240), .ZN(n14537) );
  NOR3_X1 U16399 ( .A1(n14538), .A2(n14537), .A3(P2_READREQUEST_REG_SCAN_IN), 
        .ZN(n14539) );
  AOI21_X1 U16400 ( .B1(n14540), .B2(n19275), .A(n14539), .ZN(P2_U3612) );
  XNOR2_X1 U16401 ( .A(n15697), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19511) );
  INV_X1 U16402 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18010) );
  NOR2_X1 U16403 ( .A1(n19301), .A2(n18010), .ZN(n19517) );
  AOI21_X1 U16404 ( .B1(n19512), .B2(n14542), .A(n14541), .ZN(n19518) );
  AND2_X1 U16405 ( .A1(n18086), .A2(n19518), .ZN(n14543) );
  AOI211_X1 U16406 ( .C1(n18089), .C2(n19511), .A(n19517), .B(n14543), .ZN(
        n14546) );
  OAI21_X1 U16407 ( .B1(n17612), .B2(n14544), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14545) );
  OAI211_X1 U16408 ( .C1(n17641), .C2(n19515), .A(n14546), .B(n14545), .ZN(
        P2_U3014) );
  NOR2_X1 U16409 ( .A1(n14547), .A2(n19566), .ZN(n14550) );
  NAND3_X1 U16410 ( .A1(n12058), .A2(n19570), .A3(n14548), .ZN(n14549) );
  INV_X2 U16411 ( .A(n14615), .ZN(n14625) );
  AOI22_X1 U16412 ( .A1(n14625), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n14607), .ZN(n14554) );
  INV_X1 U16413 ( .A(n14550), .ZN(n14551) );
  INV_X1 U16414 ( .A(n20061), .ZN(n14553) );
  NAND2_X1 U16415 ( .A1(n14552), .A2(n14553), .ZN(n14573) );
  NAND2_X1 U16416 ( .A1(n14554), .A2(n14573), .ZN(P2_U2965) );
  AOI22_X1 U16417 ( .A1(n14625), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n14607), .ZN(n14556) );
  AOI22_X1 U16418 ( .A1(n15777), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n15776), .ZN(n20056) );
  INV_X1 U16419 ( .A(n20056), .ZN(n14555) );
  NAND2_X1 U16420 ( .A1(n14552), .A2(n14555), .ZN(n14569) );
  NAND2_X1 U16421 ( .A1(n14556), .A2(n14569), .ZN(P2_U2966) );
  AOI22_X1 U16422 ( .A1(n14625), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n14607), .ZN(n14560) );
  INV_X1 U16423 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20906) );
  OR2_X1 U16424 ( .A1(n15776), .A2(n20906), .ZN(n14558) );
  NAND2_X1 U16425 ( .A1(n15776), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14557) );
  AND2_X1 U16426 ( .A1(n14558), .A2(n14557), .ZN(n20071) );
  INV_X1 U16427 ( .A(n20071), .ZN(n14559) );
  NAND2_X1 U16428 ( .A1(n14552), .A2(n14559), .ZN(n14575) );
  NAND2_X1 U16429 ( .A1(n14560), .A2(n14575), .ZN(P2_U2962) );
  AOI22_X1 U16430 ( .A1(n14625), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n14607), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n14562) );
  AOI22_X1 U16431 ( .A1(n15777), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15776), .ZN(n20077) );
  INV_X1 U16432 ( .A(n20077), .ZN(n14561) );
  NAND2_X1 U16433 ( .A1(n14552), .A2(n14561), .ZN(n14571) );
  NAND2_X1 U16434 ( .A1(n14562), .A2(n14571), .ZN(P2_U2960) );
  AOI22_X1 U16435 ( .A1(n14625), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n14607), .ZN(n14566) );
  INV_X1 U16436 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20910) );
  OR2_X1 U16437 ( .A1(n15776), .A2(n20910), .ZN(n14564) );
  NAND2_X1 U16438 ( .A1(n15776), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14563) );
  AND2_X1 U16439 ( .A1(n14564), .A2(n14563), .ZN(n20062) );
  INV_X1 U16440 ( .A(n20062), .ZN(n14565) );
  NAND2_X1 U16441 ( .A1(n14552), .A2(n14565), .ZN(n14567) );
  NAND2_X1 U16442 ( .A1(n14566), .A2(n14567), .ZN(P2_U2979) );
  AOI22_X1 U16443 ( .A1(n14625), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n14607), .ZN(n14568) );
  NAND2_X1 U16444 ( .A1(n14568), .A2(n14567), .ZN(P2_U2964) );
  AOI22_X1 U16445 ( .A1(n14625), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n14607), .ZN(n14570) );
  NAND2_X1 U16446 ( .A1(n14570), .A2(n14569), .ZN(P2_U2981) );
  AOI22_X1 U16447 ( .A1(n14625), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n14607), .ZN(n14572) );
  NAND2_X1 U16448 ( .A1(n14572), .A2(n14571), .ZN(P2_U2975) );
  AOI22_X1 U16449 ( .A1(n14625), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n14607), .ZN(n14574) );
  NAND2_X1 U16450 ( .A1(n14574), .A2(n14573), .ZN(P2_U2980) );
  AOI22_X1 U16451 ( .A1(n14625), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n14607), .ZN(n14576) );
  NAND2_X1 U16452 ( .A1(n14576), .A2(n14575), .ZN(P2_U2977) );
  AOI22_X1 U16453 ( .A1(n14625), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n14607), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n14578) );
  AOI22_X1 U16454 ( .A1(n15777), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15776), .ZN(n20271) );
  INV_X1 U16455 ( .A(n20271), .ZN(n14577) );
  NAND2_X1 U16456 ( .A1(n14552), .A2(n14577), .ZN(n14591) );
  NAND2_X1 U16457 ( .A1(n14578), .A2(n14591), .ZN(P2_U2958) );
  AOI22_X1 U16458 ( .A1(n14625), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n14607), .ZN(n14580) );
  AOI22_X1 U16459 ( .A1(n15777), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15776), .ZN(n20320) );
  INV_X1 U16460 ( .A(n20320), .ZN(n14579) );
  NAND2_X1 U16461 ( .A1(n14552), .A2(n14579), .ZN(n14589) );
  NAND2_X1 U16462 ( .A1(n14580), .A2(n14589), .ZN(P2_U2957) );
  AOI22_X1 U16463 ( .A1(n14625), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n14607), .ZN(n14582) );
  AOI22_X1 U16464 ( .A1(n15777), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15776), .ZN(n20409) );
  INV_X1 U16465 ( .A(n20409), .ZN(n14581) );
  NAND2_X1 U16466 ( .A1(n14552), .A2(n14581), .ZN(n14595) );
  NAND2_X1 U16467 ( .A1(n14582), .A2(n14595), .ZN(P2_U2955) );
  AOI22_X1 U16468 ( .A1(n14625), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n14607), .ZN(n14584) );
  AOI22_X1 U16469 ( .A1(n15777), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15776), .ZN(n20361) );
  INV_X1 U16470 ( .A(n20361), .ZN(n14583) );
  NAND2_X1 U16471 ( .A1(n14552), .A2(n14583), .ZN(n14597) );
  NAND2_X1 U16472 ( .A1(n14584), .A2(n14597), .ZN(P2_U2956) );
  AOI22_X1 U16473 ( .A1(n14625), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n14607), .ZN(n14586) );
  AOI22_X1 U16474 ( .A1(n15777), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15776), .ZN(n20085) );
  INV_X1 U16475 ( .A(n20085), .ZN(n14585) );
  NAND2_X1 U16476 ( .A1(n14552), .A2(n14585), .ZN(n14593) );
  NAND2_X1 U16477 ( .A1(n14586), .A2(n14593), .ZN(P2_U2959) );
  AOI22_X1 U16478 ( .A1(n14625), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n14607), .ZN(n14588) );
  AOI22_X1 U16479 ( .A1(n15777), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15776), .ZN(n20452) );
  INV_X1 U16480 ( .A(n20452), .ZN(n14587) );
  NAND2_X1 U16481 ( .A1(n14552), .A2(n14587), .ZN(n14599) );
  NAND2_X1 U16482 ( .A1(n14588), .A2(n14599), .ZN(P2_U2969) );
  AOI22_X1 U16483 ( .A1(n14625), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n14607), .ZN(n14590) );
  NAND2_X1 U16484 ( .A1(n14590), .A2(n14589), .ZN(P2_U2972) );
  AOI22_X1 U16485 ( .A1(n14625), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n14607), .ZN(n14592) );
  NAND2_X1 U16486 ( .A1(n14592), .A2(n14591), .ZN(P2_U2973) );
  AOI22_X1 U16487 ( .A1(n14625), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n14607), .ZN(n14594) );
  NAND2_X1 U16488 ( .A1(n14594), .A2(n14593), .ZN(P2_U2974) );
  AOI22_X1 U16489 ( .A1(n14625), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n14607), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U16490 ( .A1(n14596), .A2(n14595), .ZN(P2_U2970) );
  AOI22_X1 U16491 ( .A1(n14625), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n14607), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n14598) );
  NAND2_X1 U16492 ( .A1(n14598), .A2(n14597), .ZN(P2_U2971) );
  AOI22_X1 U16493 ( .A1(n14625), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n14607), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n14600) );
  NAND2_X1 U16494 ( .A1(n14600), .A2(n14599), .ZN(P2_U2954) );
  AOI22_X1 U16495 ( .A1(n14625), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n14607), .ZN(n14602) );
  AOI22_X1 U16496 ( .A1(n15777), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15776), .ZN(n20502) );
  INV_X1 U16497 ( .A(n20502), .ZN(n14601) );
  NAND2_X1 U16498 ( .A1(n14552), .A2(n14601), .ZN(n14608) );
  NAND2_X1 U16499 ( .A1(n14602), .A2(n14608), .ZN(P2_U2953) );
  AOI22_X1 U16500 ( .A1(n14625), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n14607), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n14604) );
  AOI22_X1 U16501 ( .A1(n15777), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15776), .ZN(n20559) );
  INV_X1 U16502 ( .A(n20559), .ZN(n14603) );
  NAND2_X1 U16503 ( .A1(n14552), .A2(n14603), .ZN(n14605) );
  NAND2_X1 U16504 ( .A1(n14604), .A2(n14605), .ZN(P2_U2952) );
  AOI22_X1 U16505 ( .A1(n14625), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n14607), .ZN(n14606) );
  NAND2_X1 U16506 ( .A1(n14606), .A2(n14605), .ZN(P2_U2967) );
  AOI22_X1 U16507 ( .A1(n14625), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n14607), .ZN(n14609) );
  NAND2_X1 U16508 ( .A1(n14609), .A2(n14608), .ZN(P2_U2968) );
  INV_X1 U16509 ( .A(n14610), .ZN(n14613) );
  INV_X1 U16510 ( .A(n22104), .ZN(n14612) );
  INV_X1 U16511 ( .A(n20881), .ZN(n15859) );
  OAI21_X1 U16512 ( .B1(n15859), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n14612), 
        .ZN(n14611) );
  OAI21_X1 U16513 ( .B1(n14613), .B2(n14612), .A(n14611), .ZN(P1_U3487) );
  INV_X1 U16514 ( .A(n14552), .ZN(n14616) );
  AOI22_X1 U16515 ( .A1(n15777), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15776), .ZN(n20055) );
  INV_X1 U16516 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14614) );
  INV_X1 U16517 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n18157) );
  OAI222_X1 U16518 ( .A1(n14616), .A2(n20055), .B1(n14615), .B2(n14614), .C1(
        n14650), .C2(n18157), .ZN(P2_U2982) );
  INV_X1 U16519 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14864) );
  NAND2_X1 U16520 ( .A1(n15776), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14618) );
  INV_X1 U16521 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20904) );
  OR2_X1 U16522 ( .A1(n15776), .A2(n20904), .ZN(n14617) );
  NAND2_X1 U16523 ( .A1(n14618), .A2(n14617), .ZN(n20073) );
  NAND2_X1 U16524 ( .A1(n14552), .A2(n20073), .ZN(n14621) );
  NAND2_X1 U16525 ( .A1(n14625), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14619) );
  OAI211_X1 U16526 ( .C1(n14864), .C2(n14650), .A(n14621), .B(n14619), .ZN(
        P2_U2961) );
  INV_X1 U16527 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20076) );
  NAND2_X1 U16528 ( .A1(n14625), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n14620) );
  OAI211_X1 U16529 ( .C1(n20076), .C2(n14650), .A(n14621), .B(n14620), .ZN(
        P2_U2976) );
  INV_X1 U16530 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14872) );
  NAND2_X1 U16531 ( .A1(n15776), .A2(BUF2_REG_11__SCAN_IN), .ZN(n14623) );
  INV_X1 U16532 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20908) );
  OR2_X1 U16533 ( .A1(n15776), .A2(n20908), .ZN(n14622) );
  NAND2_X1 U16534 ( .A1(n14623), .A2(n14622), .ZN(n20065) );
  NAND2_X1 U16535 ( .A1(n14552), .A2(n20065), .ZN(n14627) );
  NAND2_X1 U16536 ( .A1(n14625), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14624) );
  OAI211_X1 U16537 ( .C1(n14872), .C2(n14650), .A(n14627), .B(n14624), .ZN(
        P2_U2963) );
  INV_X1 U16538 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20068) );
  NAND2_X1 U16539 ( .A1(n14625), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n14626) );
  OAI211_X1 U16540 ( .C1(n20068), .C2(n14650), .A(n14627), .B(n14626), .ZN(
        P2_U2978) );
  INV_X1 U16541 ( .A(n14628), .ZN(n14629) );
  XNOR2_X1 U16542 ( .A(n14630), .B(n14629), .ZN(n19536) );
  INV_X1 U16543 ( .A(n19536), .ZN(n14632) );
  OR2_X1 U16544 ( .A1(n18093), .A2(n15708), .ZN(n14631) );
  INV_X1 U16545 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n15707) );
  OR2_X1 U16546 ( .A1(n19301), .A2(n15707), .ZN(n19540) );
  OAI211_X1 U16547 ( .C1(n18063), .C2(n14632), .A(n14631), .B(n19540), .ZN(
        n14636) );
  XNOR2_X1 U16548 ( .A(n14634), .B(n14633), .ZN(n19547) );
  NOR2_X1 U16549 ( .A1(n19547), .A2(n18065), .ZN(n14635) );
  AOI211_X1 U16550 ( .C1(n18083), .C2(n15705), .A(n14636), .B(n14635), .ZN(
        n14637) );
  OAI21_X1 U16551 ( .B1(n12463), .B2(n17641), .A(n14637), .ZN(P2_U3012) );
  INV_X1 U16552 ( .A(n14641), .ZN(n14638) );
  AOI222_X1 U16553 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14641), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14640), .C1(n14639), .C2(
        n14638), .ZN(n14835) );
  OAI21_X1 U16554 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14643), .A(
        n14642), .ZN(n14836) );
  INV_X1 U16555 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n14644) );
  NOR2_X1 U16556 ( .A1(n19301), .A2(n14644), .ZN(n14841) );
  INV_X1 U16557 ( .A(n14841), .ZN(n14645) );
  OAI21_X1 U16558 ( .B1(n18063), .B2(n14836), .A(n14645), .ZN(n14648) );
  OAI22_X1 U16559 ( .A1(n14646), .A2(n17641), .B1(n17638), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14647) );
  AOI211_X1 U16560 ( .C1(n17612), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14648), .B(n14647), .ZN(n14649) );
  OAI21_X1 U16561 ( .B1(n14835), .B2(n18065), .A(n14649), .ZN(P2_U3013) );
  INV_X1 U16562 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15891) );
  OR2_X1 U16563 ( .A1(n12019), .A2(n19580), .ZN(n14651) );
  OAI21_X1 U16564 ( .B1(n15274), .B2(n14651), .A(n14650), .ZN(n14652) );
  INV_X1 U16565 ( .A(n22453), .ZN(n19266) );
  NOR2_X1 U16566 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18096), .ZN(n18146) );
  NOR2_X4 U16567 ( .A1(n18127), .A2(n18154), .ZN(n18145) );
  AOI22_X1 U16568 ( .A1(n18146), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14654) );
  OAI21_X1 U16569 ( .B1(n15891), .B2(n14878), .A(n14654), .ZN(P2_U2934) );
  INV_X1 U16570 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15923) );
  AOI22_X1 U16571 ( .A1(n18146), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14655) );
  OAI21_X1 U16572 ( .B1(n15923), .B2(n14878), .A(n14655), .ZN(P2_U2933) );
  NAND2_X1 U16573 ( .A1(n11259), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14656) );
  AND4_X1 U16574 ( .A1(n13801), .A2(n14656), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20162), .ZN(n14657) );
  MUX2_X1 U16575 ( .A(n12545), .B(n19515), .S(n17309), .Z(n14659) );
  OAI21_X1 U16576 ( .B1(n17316), .B2(n18098), .A(n14659), .ZN(P2_U2887) );
  INV_X1 U16577 ( .A(n14660), .ZN(n14661) );
  OAI21_X1 U16578 ( .B1(n14661), .B2(n17162), .A(n18038), .ZN(n14662) );
  INV_X1 U16579 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22386) );
  NAND2_X1 U16580 ( .A1(n14662), .A2(n22386), .ZN(n14664) );
  OR2_X1 U16581 ( .A1(n22392), .A2(n22391), .ZN(n14711) );
  AOI21_X1 U16582 ( .B1(n14664), .B2(n22386), .A(n14711), .ZN(n14663) );
  OR2_X1 U16583 ( .A1(n15397), .A2(n14663), .ZN(n17155) );
  NAND2_X1 U16584 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22393), .ZN(n17153) );
  INV_X1 U16585 ( .A(n14664), .ZN(n14665) );
  NOR2_X1 U16586 ( .A1(n14665), .A2(n22391), .ZN(n22400) );
  AOI21_X1 U16587 ( .B1(n13313), .B2(n17153), .A(n22400), .ZN(n14666) );
  OAI21_X1 U16588 ( .B1(n13311), .B2(n22609), .A(n14666), .ZN(n14667) );
  NAND2_X1 U16589 ( .A1(n17155), .A2(n14667), .ZN(n14668) );
  OAI21_X1 U16590 ( .B1(n17155), .B2(n22567), .A(n14668), .ZN(P1_U3478) );
  OAI22_X1 U16591 ( .A1(n14669), .A2(n14293), .B1(n13044), .B2(n14686), .ZN(
        n14670) );
  INV_X1 U16592 ( .A(n14670), .ZN(n14681) );
  AOI21_X1 U16593 ( .B1(n14671), .B2(n14784), .A(n13044), .ZN(n14672) );
  NAND2_X1 U16594 ( .A1(n14673), .A2(n14672), .ZN(n14701) );
  AOI21_X1 U16595 ( .B1(n15033), .B2(n14786), .A(n16741), .ZN(n14676) );
  NAND2_X1 U16596 ( .A1(n14674), .A2(n13044), .ZN(n14675) );
  NAND3_X1 U16597 ( .A1(n14677), .A2(n14676), .A3(n14675), .ZN(n14678) );
  NAND2_X1 U16598 ( .A1(n14678), .A2(n14784), .ZN(n14679) );
  NAND4_X1 U16599 ( .A1(n14681), .A2(n14680), .A3(n14701), .A4(n14679), .ZN(
        n14803) );
  INV_X1 U16600 ( .A(n14696), .ZN(n14683) );
  NAND3_X1 U16601 ( .A1(n14683), .A2(n14682), .A3(n14801), .ZN(n14684) );
  NOR2_X1 U16602 ( .A1(n14803), .A2(n14684), .ZN(n14685) );
  INV_X1 U16603 ( .A(n17167), .ZN(n14820) );
  NAND2_X1 U16604 ( .A1(n16097), .A2(n14784), .ZN(n17165) );
  INV_X1 U16605 ( .A(n17165), .ZN(n18019) );
  XNOR2_X1 U16606 ( .A(n13236), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14690) );
  AND2_X1 U16607 ( .A1(n17163), .A2(n14686), .ZN(n14769) );
  INV_X1 U16608 ( .A(n16690), .ZN(n14687) );
  NOR2_X1 U16609 ( .A1(n14687), .A2(n14721), .ZN(n16109) );
  AND2_X1 U16610 ( .A1(n14769), .A2(n16109), .ZN(n14824) );
  XNOR2_X1 U16611 ( .A(n14822), .B(n14688), .ZN(n14693) );
  INV_X1 U16612 ( .A(n14693), .ZN(n14689) );
  AOI22_X1 U16613 ( .A1(n18019), .A2(n14690), .B1(n14824), .B2(n14689), .ZN(
        n14692) );
  NAND3_X1 U16614 ( .A1(n14820), .A2(n14819), .A3(n14693), .ZN(n14691) );
  OAI211_X1 U16615 ( .C1(n17159), .C2(n14820), .A(n14692), .B(n14691), .ZN(
        n18014) );
  INV_X1 U16616 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U16617 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14895), .B2(n16979), .ZN(
        n17168) );
  NOR2_X1 U16618 ( .A1(n22388), .A2(n11214), .ZN(n17170) );
  AOI222_X1 U16619 ( .A1(n18014), .A2(n17977), .B1(n17168), .B2(n17170), .C1(
        n22396), .C2(n14693), .ZN(n14713) );
  INV_X1 U16620 ( .A(n16108), .ZN(n14705) );
  AND2_X1 U16621 ( .A1(n14694), .A2(n22424), .ZN(n14695) );
  NAND2_X1 U16622 ( .A1(n14696), .A2(n14695), .ZN(n14781) );
  NAND2_X1 U16623 ( .A1(n18044), .A2(n22424), .ZN(n14697) );
  AOI22_X1 U16624 ( .A1(n17165), .A2(n14781), .B1(n14722), .B2(n14697), .ZN(
        n14704) );
  INV_X1 U16625 ( .A(n22424), .ZN(n22436) );
  NOR2_X1 U16626 ( .A1(n14784), .A2(n22436), .ZN(n14698) );
  NAND2_X1 U16627 ( .A1(n16106), .A2(n14698), .ZN(n14924) );
  INV_X1 U16628 ( .A(n14699), .ZN(n14700) );
  OR2_X1 U16629 ( .A1(n14700), .A2(n16097), .ZN(n14702) );
  OAI211_X1 U16630 ( .C1(n16690), .C2(n14786), .A(n14924), .B(n14788), .ZN(
        n14703) );
  AOI21_X1 U16631 ( .B1(n14705), .B2(n14704), .A(n14703), .ZN(n14710) );
  NAND2_X1 U16632 ( .A1(n14769), .A2(n14706), .ZN(n14793) );
  OR2_X1 U16633 ( .A1(n16108), .A2(n14793), .ZN(n14925) );
  NAND2_X1 U16634 ( .A1(n14769), .A2(n11155), .ZN(n16105) );
  INV_X1 U16635 ( .A(n16105), .ZN(n14707) );
  NAND2_X1 U16636 ( .A1(n16108), .A2(n14707), .ZN(n14708) );
  AND2_X1 U16637 ( .A1(n14925), .A2(n14708), .ZN(n14709) );
  NAND2_X1 U16638 ( .A1(n14710), .A2(n14709), .ZN(n18037) );
  OAI22_X1 U16639 ( .A1(n18017), .A2(n22402), .B1(n14711), .B2(n22386), .ZN(
        n17976) );
  AOI21_X1 U16640 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22392), .A(n17976), 
        .ZN(n14832) );
  NAND2_X1 U16641 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n14832), .ZN(
        n14712) );
  OAI21_X1 U16642 ( .B1(n14713), .B2(n14832), .A(n14712), .ZN(P1_U3472) );
  INV_X1 U16643 ( .A(n14714), .ZN(n14716) );
  INV_X1 U16644 ( .A(n20108), .ZN(n18106) );
  NAND2_X1 U16645 ( .A1(n18106), .A2(n17303), .ZN(n14718) );
  NAND2_X1 U16646 ( .A1(n17309), .A2(n17238), .ZN(n14717) );
  OAI211_X1 U16647 ( .C1(n14719), .C2(n17309), .A(n14718), .B(n14717), .ZN(
        P2_U2886) );
  NAND2_X1 U16648 ( .A1(n14783), .A2(n14191), .ZN(n16096) );
  INV_X1 U16649 ( .A(n16096), .ZN(n14720) );
  OR2_X1 U16650 ( .A1(n14722), .A2(n14784), .ZN(n14809) );
  AOI22_X1 U16651 ( .A1(n22523), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n22527), .ZN(n14723) );
  INV_X1 U16652 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20890) );
  INV_X1 U16653 ( .A(DATAI_2_), .ZN(n16344) );
  AOI22_X1 U16654 ( .A1(n15793), .A2(n20890), .B1(n16344), .B2(n16757), .ZN(
        n16808) );
  INV_X1 U16655 ( .A(n16808), .ZN(n14933) );
  OR2_X1 U16656 ( .A1(n22480), .A2(n14933), .ZN(n14728) );
  NAND2_X1 U16657 ( .A1(n14723), .A2(n14728), .ZN(P1_U2939) );
  AOI22_X1 U16658 ( .A1(n22523), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n22527), .ZN(n14724) );
  INV_X1 U16659 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20896) );
  INV_X1 U16660 ( .A(DATAI_5_), .ZN(n16339) );
  AOI22_X1 U16661 ( .A1(n15793), .A2(n20896), .B1(n16339), .B2(n16757), .ZN(
        n15017) );
  INV_X1 U16662 ( .A(n15017), .ZN(n16791) );
  OR2_X1 U16663 ( .A1(n22480), .A2(n16791), .ZN(n14733) );
  NAND2_X1 U16664 ( .A1(n14724), .A2(n14733), .ZN(P1_U2942) );
  AOI22_X1 U16665 ( .A1(n22523), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n22527), .ZN(n14725) );
  INV_X1 U16666 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20892) );
  INV_X1 U16667 ( .A(DATAI_3_), .ZN(n16343) );
  AOI22_X1 U16668 ( .A1(n15793), .A2(n20892), .B1(n16343), .B2(n16757), .ZN(
        n16802) );
  INV_X1 U16669 ( .A(n16802), .ZN(n15055) );
  OR2_X1 U16670 ( .A1(n22480), .A2(n15055), .ZN(n14730) );
  NAND2_X1 U16671 ( .A1(n14725), .A2(n14730), .ZN(P1_U2940) );
  AOI22_X1 U16672 ( .A1(n22523), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(
        P1_EAX_REG_7__SCAN_IN), .B2(n22527), .ZN(n14727) );
  INV_X1 U16673 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20900) );
  INV_X1 U16674 ( .A(DATAI_7_), .ZN(n14726) );
  AOI22_X1 U16675 ( .A1(n15793), .A2(n20900), .B1(n14726), .B2(n16757), .ZN(
        n16779) );
  INV_X1 U16676 ( .A(n16779), .ZN(n15587) );
  OR2_X1 U16677 ( .A1(n22480), .A2(n15587), .ZN(n14738) );
  NAND2_X1 U16678 ( .A1(n14727), .A2(n14738), .ZN(P1_U2959) );
  AOI22_X1 U16679 ( .A1(n22523), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(
        P1_EAX_REG_2__SCAN_IN), .B2(n22527), .ZN(n14729) );
  NAND2_X1 U16680 ( .A1(n14729), .A2(n14728), .ZN(P1_U2954) );
  AOI22_X1 U16681 ( .A1(n22523), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(
        P1_EAX_REG_3__SCAN_IN), .B2(n22527), .ZN(n14731) );
  NAND2_X1 U16682 ( .A1(n14731), .A2(n14730), .ZN(P1_U2955) );
  AOI22_X1 U16683 ( .A1(n22523), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(
        P1_EAX_REG_6__SCAN_IN), .B2(n22527), .ZN(n14732) );
  INV_X1 U16684 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20898) );
  INV_X1 U16685 ( .A(DATAI_6_), .ZN(n16335) );
  AOI22_X1 U16686 ( .A1(n15793), .A2(n20898), .B1(n16335), .B2(n16757), .ZN(
        n16785) );
  INV_X1 U16687 ( .A(n16785), .ZN(n15539) );
  OR2_X1 U16688 ( .A1(n22480), .A2(n15539), .ZN(n14740) );
  NAND2_X1 U16689 ( .A1(n14732), .A2(n14740), .ZN(P1_U2958) );
  AOI22_X1 U16690 ( .A1(n22523), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(
        P1_EAX_REG_5__SCAN_IN), .B2(n22527), .ZN(n14734) );
  NAND2_X1 U16691 ( .A1(n14734), .A2(n14733), .ZN(P1_U2957) );
  AOI22_X1 U16692 ( .A1(n22523), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n22527), .ZN(n14735) );
  INV_X1 U16693 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20888) );
  INV_X1 U16694 ( .A(DATAI_1_), .ZN(n16348) );
  AOI22_X1 U16695 ( .A1(n15793), .A2(n20888), .B1(n16348), .B2(n16757), .ZN(
        n16814) );
  INV_X1 U16696 ( .A(n16814), .ZN(n14934) );
  OR2_X1 U16697 ( .A1(n22480), .A2(n14934), .ZN(n14736) );
  NAND2_X1 U16698 ( .A1(n14735), .A2(n14736), .ZN(P1_U2938) );
  AOI22_X1 U16699 ( .A1(n22523), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(
        P1_EAX_REG_1__SCAN_IN), .B2(n22527), .ZN(n14737) );
  NAND2_X1 U16700 ( .A1(n14737), .A2(n14736), .ZN(P1_U2953) );
  AOI22_X1 U16701 ( .A1(n22523), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n22527), .ZN(n14739) );
  NAND2_X1 U16702 ( .A1(n14739), .A2(n14738), .ZN(P1_U2944) );
  AOI22_X1 U16703 ( .A1(n22523), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n22527), .ZN(n14741) );
  NAND2_X1 U16704 ( .A1(n14741), .A2(n14740), .ZN(P1_U2943) );
  AOI22_X1 U16705 ( .A1(n22523), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n22527), .ZN(n14742) );
  OAI22_X1 U16706 ( .A1(n16757), .A2(BUF1_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        n15793), .ZN(n14932) );
  INV_X1 U16707 ( .A(n14932), .ZN(n16820) );
  NAND2_X1 U16708 ( .A1(n22521), .A2(n16820), .ZN(n14746) );
  NAND2_X1 U16709 ( .A1(n14742), .A2(n14746), .ZN(P1_U2937) );
  AOI22_X1 U16710 ( .A1(n22523), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(
        P1_EAX_REG_4__SCAN_IN), .B2(n22527), .ZN(n14743) );
  OAI22_X1 U16711 ( .A1(n16757), .A2(BUF1_REG_4__SCAN_IN), .B1(DATAI_4_), .B2(
        n15793), .ZN(n15117) );
  INV_X1 U16712 ( .A(n15117), .ZN(n16797) );
  NAND2_X1 U16713 ( .A1(n22521), .A2(n16797), .ZN(n14744) );
  NAND2_X1 U16714 ( .A1(n14743), .A2(n14744), .ZN(P1_U2956) );
  AOI22_X1 U16715 ( .A1(n22523), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n22527), .ZN(n14745) );
  NAND2_X1 U16716 ( .A1(n14745), .A2(n14744), .ZN(P1_U2941) );
  AOI22_X1 U16717 ( .A1(n22523), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(
        P1_EAX_REG_0__SCAN_IN), .B2(n22527), .ZN(n14747) );
  NAND2_X1 U16718 ( .A1(n14747), .A2(n14746), .ZN(P1_U2952) );
  INV_X1 U16719 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U16720 ( .A1(n14783), .A2(n18019), .ZN(n14748) );
  NAND2_X1 U16721 ( .A1(n22525), .A2(n14748), .ZN(n14749) );
  NOR2_X1 U16722 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22391), .ZN(n20725) );
  AOI22_X1 U16723 ( .A1(n20725), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14750) );
  OAI21_X1 U16724 ( .B1(n14751), .B2(n14958), .A(n14750), .ZN(P1_U2913) );
  INV_X1 U16725 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n22489) );
  AOI22_X1 U16726 ( .A1(n22106), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14752) );
  OAI21_X1 U16727 ( .B1(n22489), .B2(n14958), .A(n14752), .ZN(P1_U2911) );
  INV_X1 U16728 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U16729 ( .A1(n22106), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14753) );
  OAI21_X1 U16730 ( .B1(n14754), .B2(n14958), .A(n14753), .ZN(P1_U2914) );
  AOI22_X1 U16731 ( .A1(n22106), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14755) );
  OAI21_X1 U16732 ( .B1(n16790), .B2(n14958), .A(n14755), .ZN(P1_U2915) );
  AOI22_X1 U16733 ( .A1(n22106), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14756) );
  OAI21_X1 U16734 ( .B1(n22482), .B2(n14958), .A(n14756), .ZN(P1_U2912) );
  AOI22_X1 U16735 ( .A1(n15793), .A2(BUF1_REG_15__SCAN_IN), .B1(DATAI_15_), 
        .B2(n16757), .ZN(n16828) );
  AOI22_X1 U16736 ( .A1(n22528), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(
        P1_EAX_REG_15__SCAN_IN), .B2(n22527), .ZN(n14757) );
  OAI21_X1 U16737 ( .B1(n16828), .B2(n22480), .A(n14757), .ZN(P1_U2967) );
  INV_X1 U16738 ( .A(n13313), .ZN(n16700) );
  OAI22_X1 U16739 ( .A1(n16700), .A2(n14820), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14758), .ZN(n18018) );
  INV_X1 U16740 ( .A(n22396), .ZN(n14759) );
  OAI22_X1 U16741 ( .A1(n22388), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14759), .ZN(n14760) );
  AOI21_X1 U16742 ( .B1(n18018), .B2(n17977), .A(n14760), .ZN(n14763) );
  AOI21_X1 U16743 ( .B1(n18019), .B2(n17977), .A(n14832), .ZN(n14762) );
  OAI22_X1 U16744 ( .A1(n14763), .A2(n14832), .B1(n14762), .B2(n14761), .ZN(
        P1_U3474) );
  MUX2_X1 U16745 ( .A(n12463), .B(n12089), .S(n15680), .Z(n14766) );
  OAI21_X1 U16746 ( .B1(n20447), .B2(n17316), .A(n14766), .ZN(P2_U2885) );
  OAI21_X1 U16747 ( .B1(n14768), .B2(n14767), .A(n14910), .ZN(n16698) );
  NAND2_X1 U16748 ( .A1(n16108), .A2(n14769), .ZN(n14774) );
  NOR2_X1 U16749 ( .A1(n14771), .A2(n14770), .ZN(n14773) );
  NAND4_X1 U16750 ( .A1(n14819), .A2(n16741), .A3(n14773), .A4(n14772), .ZN(
        n14926) );
  NAND2_X1 U16751 ( .A1(n14774), .A2(n14926), .ZN(n14776) );
  NAND2_X2 U16752 ( .A1(n14777), .A2(n20833), .ZN(n20812) );
  XNOR2_X1 U16753 ( .A(n14778), .B(n11155), .ZN(n16695) );
  AOI22_X1 U16754 ( .A1(n20825), .A2(n16695), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n16714), .ZN(n14779) );
  OAI21_X1 U16755 ( .B1(n16698), .B2(n20812), .A(n14779), .ZN(P1_U2871) );
  NAND3_X1 U16756 ( .A1(n14781), .A2(n11244), .A3(n14780), .ZN(n14782) );
  NAND3_X1 U16757 ( .A1(n14783), .A2(n15025), .A3(n14782), .ZN(n14792) );
  NAND3_X1 U16758 ( .A1(n16108), .A2(n17163), .A3(n14784), .ZN(n14789) );
  NAND2_X1 U16759 ( .A1(n14784), .A2(n22434), .ZN(n14785) );
  NAND4_X1 U16760 ( .A1(n16098), .A2(n14786), .A3(n22424), .A4(n14785), .ZN(
        n14787) );
  NAND3_X1 U16761 ( .A1(n14789), .A2(n14788), .A3(n14787), .ZN(n14790) );
  NAND2_X1 U16762 ( .A1(n14790), .A2(n14927), .ZN(n14791) );
  INV_X1 U16763 ( .A(n14793), .ZN(n14794) );
  NOR2_X1 U16764 ( .A1(n18031), .A2(n14794), .ZN(n16101) );
  INV_X1 U16765 ( .A(n14795), .ZN(n14796) );
  OAI211_X1 U16766 ( .C1(n12981), .C2(n14806), .A(n16101), .B(n14796), .ZN(
        n14797) );
  INV_X1 U16767 ( .A(n14797), .ZN(n14798) );
  XOR2_X1 U16768 ( .A(n14799), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n14921) );
  OAI21_X1 U16769 ( .B1(n14801), .B2(n11244), .A(n14800), .ZN(n14802) );
  NOR2_X1 U16770 ( .A1(n14803), .A2(n14802), .ZN(n14804) );
  OR2_X1 U16771 ( .A1(n17125), .A2(n22123), .ZN(n14805) );
  NAND2_X1 U16772 ( .A1(n14805), .A2(n11214), .ZN(n22217) );
  NAND2_X1 U16773 ( .A1(n22129), .A2(n14811), .ZN(n22222) );
  AOI21_X1 U16774 ( .B1(n22217), .B2(n22222), .A(n14895), .ZN(n14815) );
  OR2_X1 U16775 ( .A1(n14811), .A2(n17165), .ZN(n22223) );
  OAI21_X1 U16776 ( .B1(n22188), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14895), .ZN(n14813) );
  INV_X1 U16777 ( .A(n14806), .ZN(n14807) );
  NAND2_X1 U16778 ( .A1(n14807), .A2(n12981), .ZN(n14808) );
  AND2_X1 U16779 ( .A1(n14809), .A2(n14808), .ZN(n14810) );
  AND2_X1 U16780 ( .A1(n22202), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14920) );
  AOI21_X1 U16781 ( .B1(n22199), .B2(n16695), .A(n14920), .ZN(n14812) );
  OAI21_X1 U16782 ( .B1(n17103), .B2(n14813), .A(n14812), .ZN(n14814) );
  AOI211_X1 U16783 ( .C1(n22200), .C2(n14921), .A(n14815), .B(n14814), .ZN(
        n14816) );
  INV_X1 U16784 ( .A(n14816), .ZN(P1_U3030) );
  NAND2_X1 U16785 ( .A1(n22237), .A2(n17167), .ZN(n14830) );
  INV_X1 U16786 ( .A(n14822), .ZN(n17171) );
  AOI211_X1 U16787 ( .C1(n11416), .C2(n17171), .A(n14818), .B(n13739), .ZN(
        n14831) );
  NAND3_X1 U16788 ( .A1(n14820), .A2(n14819), .A3(n14831), .ZN(n14829) );
  MUX2_X1 U16789 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14826), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n14821) );
  OAI21_X1 U16790 ( .B1(n14823), .B2(n14821), .A(n18019), .ZN(n14828) );
  MUX2_X1 U16791 ( .A(n14823), .B(n11416), .S(n14822), .Z(n14825) );
  OAI21_X1 U16792 ( .B1(n14826), .B2(n14825), .A(n14824), .ZN(n14827) );
  NAND4_X1 U16793 ( .A1(n14830), .A2(n14829), .A3(n14828), .A4(n14827), .ZN(
        n18015) );
  AOI22_X1 U16794 ( .A1(n18015), .A2(n17977), .B1(n14831), .B2(n22396), .ZN(
        n14833) );
  INV_X1 U16795 ( .A(n14832), .ZN(n17979) );
  MUX2_X1 U16796 ( .A(n11416), .B(n14833), .S(n17979), .Z(n14834) );
  INV_X1 U16797 ( .A(n14834), .ZN(P1_U3469) );
  AOI211_X1 U16798 ( .C1(n19512), .C2(n14844), .A(n15564), .B(n19521), .ZN(
        n14847) );
  NOR2_X1 U16799 ( .A1(n14835), .A2(n19546), .ZN(n14846) );
  INV_X1 U16800 ( .A(n14836), .ZN(n14837) );
  AOI22_X1 U16801 ( .A1(n19550), .A2(n17238), .B1(n19537), .B2(n14837), .ZN(
        n14843) );
  OAI21_X1 U16802 ( .B1(n14840), .B2(n14839), .A(n14838), .ZN(n20496) );
  AOI21_X1 U16803 ( .B1(n19527), .B2(n20496), .A(n14841), .ZN(n14842) );
  OAI211_X1 U16804 ( .C1(n14844), .C2(n19513), .A(n14843), .B(n14842), .ZN(
        n14845) );
  OR3_X1 U16805 ( .A1(n14847), .A2(n14846), .A3(n14845), .ZN(P2_U3045) );
  NAND2_X1 U16806 ( .A1(n16495), .A2(n11214), .ZN(n14848) );
  NAND2_X1 U16807 ( .A1(n14849), .A2(n14848), .ZN(n22213) );
  INV_X1 U16808 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14854) );
  NAND2_X1 U16809 ( .A1(n14851), .A2(n14850), .ZN(n14852) );
  NAND2_X1 U16810 ( .A1(n14853), .A2(n14852), .ZN(n16705) );
  OAI222_X1 U16811 ( .A1(n22213), .A2(n20828), .B1(n14854), .B2(n20833), .C1(
        n16705), .C2(n20812), .ZN(P1_U2872) );
  OR2_X1 U16812 ( .A1(n14855), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14856) );
  NAND2_X1 U16813 ( .A1(n14857), .A2(n14856), .ZN(n22219) );
  NAND2_X1 U16814 ( .A1(n22202), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n22212) );
  OAI21_X1 U16815 ( .B1(n20870), .B2(n14858), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14859) );
  OAI211_X1 U16816 ( .C1(n22219), .C2(n22385), .A(n22212), .B(n14859), .ZN(
        n14860) );
  INV_X1 U16817 ( .A(n14860), .ZN(n14861) );
  OAI21_X1 U16818 ( .B1(n20853), .B2(n16705), .A(n14861), .ZN(P1_U2999) );
  INV_X1 U16819 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n15870) );
  AOI22_X1 U16820 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n18154), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n18145), .ZN(n14862) );
  OAI21_X1 U16821 ( .B1(n15870), .B2(n14878), .A(n14862), .ZN(P2_U2935) );
  AOI22_X1 U16822 ( .A1(n18154), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14863) );
  OAI21_X1 U16823 ( .B1(n14864), .B2(n14878), .A(n14863), .ZN(P2_U2926) );
  INV_X1 U16824 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U16825 ( .A1(n18154), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14865) );
  OAI21_X1 U16826 ( .B1(n17353), .B2(n14878), .A(n14865), .ZN(P2_U2927) );
  INV_X1 U16827 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U16828 ( .A1(n18154), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14866) );
  OAI21_X1 U16829 ( .B1(n17362), .B2(n14878), .A(n14866), .ZN(P2_U2928) );
  INV_X1 U16830 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U16831 ( .A1(n18154), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14867) );
  OAI21_X1 U16832 ( .B1(n17392), .B2(n14878), .A(n14867), .ZN(P2_U2931) );
  AOI22_X1 U16833 ( .A1(n18154), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14868) );
  OAI21_X1 U16834 ( .B1(n14869), .B2(n14878), .A(n14868), .ZN(P2_U2922) );
  INV_X1 U16835 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n17317) );
  AOI22_X1 U16836 ( .A1(n18154), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14870) );
  OAI21_X1 U16837 ( .B1(n17317), .B2(n14878), .A(n14870), .ZN(P2_U2923) );
  AOI22_X1 U16838 ( .A1(n18154), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14871) );
  OAI21_X1 U16839 ( .B1(n14872), .B2(n14878), .A(n14871), .ZN(P2_U2924) );
  INV_X1 U16840 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n17333) );
  AOI22_X1 U16841 ( .A1(n18154), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14873) );
  OAI21_X1 U16842 ( .B1(n17333), .B2(n14878), .A(n14873), .ZN(P2_U2925) );
  INV_X1 U16843 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U16844 ( .A1(n18154), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14874) );
  OAI21_X1 U16845 ( .B1(n17381), .B2(n14878), .A(n14874), .ZN(P2_U2930) );
  INV_X1 U16846 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U16847 ( .A1(n18154), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14875) );
  OAI21_X1 U16848 ( .B1(n17374), .B2(n14878), .A(n14875), .ZN(P2_U2929) );
  INV_X1 U16849 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n17403) );
  AOI22_X1 U16850 ( .A1(n18146), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14876) );
  OAI21_X1 U16851 ( .B1(n17403), .B2(n14878), .A(n14876), .ZN(P2_U2932) );
  INV_X1 U16852 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U16853 ( .A1(n18146), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14877) );
  OAI21_X1 U16854 ( .B1(n16074), .B2(n14878), .A(n14877), .ZN(P2_U2921) );
  OAI21_X1 U16855 ( .B1(n14879), .B2(n14881), .A(n14880), .ZN(n20315) );
  NOR2_X1 U16856 ( .A1(n14883), .A2(n14882), .ZN(n14884) );
  OR2_X1 U16857 ( .A1(n14905), .A2(n14884), .ZN(n18062) );
  INV_X1 U16858 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14885) );
  MUX2_X1 U16859 ( .A(n18062), .B(n14885), .S(n15680), .Z(n14886) );
  OAI21_X1 U16860 ( .B1(n20315), .B2(n17316), .A(n14886), .ZN(P2_U2883) );
  XOR2_X1 U16861 ( .A(n14888), .B(n14887), .Z(n14914) );
  INV_X1 U16862 ( .A(n14914), .ZN(n14898) );
  NAND2_X1 U16863 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n22123), .ZN(
        n22114) );
  NAND2_X1 U16864 ( .A1(n22223), .A2(n22114), .ZN(n17105) );
  AND2_X1 U16865 ( .A1(n17105), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15475) );
  INV_X1 U16866 ( .A(n15475), .ZN(n14891) );
  NOR3_X1 U16867 ( .A1(n11214), .A2(n14895), .A3(n22119), .ZN(n15476) );
  NAND2_X1 U16868 ( .A1(n22123), .A2(n11214), .ZN(n14889) );
  NAND2_X1 U16869 ( .A1(n22222), .A2(n14889), .ZN(n17102) );
  OAI21_X1 U16870 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17122), .A(
        n22118), .ZN(n22145) );
  NOR2_X1 U16871 ( .A1(n15476), .A2(n22145), .ZN(n14890) );
  MUX2_X1 U16872 ( .A(n14891), .B(n14890), .S(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n14897) );
  NOR2_X1 U16873 ( .A1(n14893), .A2(n14892), .ZN(n14894) );
  OR2_X1 U16874 ( .A1(n14976), .A2(n14894), .ZN(n20809) );
  INV_X1 U16875 ( .A(n20809), .ZN(n22230) );
  INV_X1 U16876 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n22246) );
  NOR2_X1 U16877 ( .A1(n22129), .A2(n22246), .ZN(n14916) );
  INV_X1 U16878 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n22148) );
  OAI21_X1 U16879 ( .B1(n11214), .B2(n14895), .A(n22148), .ZN(n15480) );
  NOR2_X1 U16880 ( .A1(n22119), .A2(n15480), .ZN(n22146) );
  AOI211_X1 U16881 ( .C1(n22199), .C2(n22230), .A(n14916), .B(n22146), .ZN(
        n14896) );
  OAI211_X1 U16882 ( .C1(n14898), .C2(n22218), .A(n14897), .B(n14896), .ZN(
        P1_U3029) );
  INV_X1 U16883 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n16086) );
  INV_X1 U16884 ( .A(n11260), .ZN(n15559) );
  MUX2_X1 U16885 ( .A(n16086), .B(n15559), .S(n17309), .Z(n14903) );
  OAI21_X1 U16886 ( .B1(n20132), .B2(n17316), .A(n14903), .ZN(P2_U2884) );
  XOR2_X1 U16887 ( .A(n14880), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14909)
         );
  OR2_X1 U16888 ( .A1(n14905), .A2(n14904), .ZN(n14907) );
  NAND2_X1 U16889 ( .A1(n14907), .A2(n14906), .ZN(n15839) );
  MUX2_X1 U16890 ( .A(n15839), .B(n12115), .S(n15680), .Z(n14908) );
  OAI21_X1 U16891 ( .B1(n14909), .B2(n17316), .A(n14908), .ZN(P2_U2882) );
  NAND2_X1 U16892 ( .A1(n14911), .A2(n14910), .ZN(n14912) );
  NAND2_X1 U16893 ( .A1(n14913), .A2(n14912), .ZN(n22232) );
  INV_X1 U16894 ( .A(n22385), .ZN(n20872) );
  NAND2_X1 U16895 ( .A1(n14914), .A2(n20872), .ZN(n14918) );
  NOR2_X1 U16896 ( .A1(n20877), .A2(n22231), .ZN(n14915) );
  AOI211_X1 U16897 ( .C1(n20870), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14916), .B(n14915), .ZN(n14917) );
  OAI211_X1 U16898 ( .C1(n20853), .C2(n22232), .A(n14918), .B(n14917), .ZN(
        P1_U2997) );
  NOR2_X1 U16899 ( .A1(n20877), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14919) );
  AOI211_X1 U16900 ( .C1(n20870), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14920), .B(n14919), .ZN(n14923) );
  NAND2_X1 U16901 ( .A1(n14921), .A2(n20872), .ZN(n14922) );
  OAI211_X1 U16902 ( .C1(n20853), .C2(n16698), .A(n14923), .B(n14922), .ZN(
        P1_U2998) );
  OAI211_X1 U16903 ( .C1(n16688), .C2(n14926), .A(n14925), .B(n14924), .ZN(
        n14928) );
  NAND2_X1 U16904 ( .A1(n14928), .A2(n14927), .ZN(n14929) );
  NOR2_X1 U16905 ( .A1(n14931), .A2(n12978), .ZN(n14930) );
  INV_X1 U16906 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20711) );
  OAI222_X1 U16907 ( .A1(n16705), .A2(n16837), .B1(n16836), .B2(n14932), .C1(
        n16834), .C2(n20711), .ZN(P1_U2904) );
  INV_X1 U16908 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20715) );
  OAI222_X1 U16909 ( .A1(n22232), .A2(n16837), .B1(n16836), .B2(n14933), .C1(
        n16834), .C2(n20715), .ZN(P1_U2902) );
  INV_X1 U16910 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20713) );
  OAI222_X1 U16911 ( .A1(n16698), .A2(n16837), .B1(n16836), .B2(n14934), .C1(
        n16834), .C2(n20713), .ZN(P1_U2903) );
  NAND2_X1 U16912 ( .A1(n11254), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n17152) );
  INV_X1 U16913 ( .A(n13301), .ZN(n14937) );
  INV_X1 U16914 ( .A(n15196), .ZN(n14938) );
  NAND2_X1 U16915 ( .A1(n14938), .A2(n17152), .ZN(n14939) );
  OAI211_X1 U16916 ( .C1(n15118), .C2(n17152), .A(n15050), .B(n14939), .ZN(
        n14940) );
  AOI22_X1 U16917 ( .A1(n14940), .A2(n17151), .B1(n17153), .B2(n22237), .ZN(
        n14942) );
  NAND2_X1 U16918 ( .A1(n18057), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14941) );
  OAI21_X1 U16919 ( .B1(n14942), .B2(n18057), .A(n14941), .ZN(P1_U3475) );
  INV_X1 U16920 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U16921 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20734), .B1(n20725), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14943) );
  OAI21_X1 U16922 ( .B1(n14944), .B2(n14958), .A(n14943), .ZN(P1_U2920) );
  INV_X1 U16923 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14946) );
  AOI22_X1 U16924 ( .A1(n20725), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14945) );
  OAI21_X1 U16925 ( .B1(n14946), .B2(n14958), .A(n14945), .ZN(P1_U2919) );
  INV_X1 U16926 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14948) );
  AOI22_X1 U16927 ( .A1(n22106), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14947) );
  OAI21_X1 U16928 ( .B1(n14948), .B2(n14958), .A(n14947), .ZN(P1_U2917) );
  INV_X1 U16929 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14950) );
  AOI22_X1 U16930 ( .A1(n22106), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14949) );
  OAI21_X1 U16931 ( .B1(n14950), .B2(n14958), .A(n14949), .ZN(P1_U2918) );
  INV_X1 U16932 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n22496) );
  AOI22_X1 U16933 ( .A1(n22106), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14951) );
  OAI21_X1 U16934 ( .B1(n22496), .B2(n14958), .A(n14951), .ZN(P1_U2910) );
  INV_X1 U16935 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n22516) );
  AOI22_X1 U16936 ( .A1(n22106), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14952) );
  OAI21_X1 U16937 ( .B1(n22516), .B2(n14958), .A(n14952), .ZN(P1_U2907) );
  INV_X1 U16938 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n22502) );
  AOI22_X1 U16939 ( .A1(n22106), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14953) );
  OAI21_X1 U16940 ( .B1(n22502), .B2(n14958), .A(n14953), .ZN(P1_U2909) );
  AOI22_X1 U16941 ( .A1(n22106), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14954) );
  OAI21_X1 U16942 ( .B1(n22509), .B2(n14958), .A(n14954), .ZN(P1_U2908) );
  INV_X1 U16943 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14956) );
  AOI22_X1 U16944 ( .A1(n22106), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14955) );
  OAI21_X1 U16945 ( .B1(n14956), .B2(n14958), .A(n14955), .ZN(P1_U2916) );
  INV_X1 U16946 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n22526) );
  AOI22_X1 U16947 ( .A1(n22106), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14957) );
  OAI21_X1 U16948 ( .B1(n22526), .B2(n14958), .A(n14957), .ZN(P1_U2906) );
  XNOR2_X1 U16949 ( .A(n14959), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14963) );
  OR2_X1 U16950 ( .A1(n14960), .A2(n14967), .ZN(n14961) );
  NAND2_X1 U16951 ( .A1(n15371), .A2(n14961), .ZN(n19283) );
  MUX2_X1 U16952 ( .A(n11923), .B(n19283), .S(n17309), .Z(n14962) );
  OAI21_X1 U16953 ( .B1(n14963), .B2(n17316), .A(n14962), .ZN(P2_U2880) );
  NOR2_X1 U16954 ( .A1(n14880), .A2(n20360), .ZN(n14965) );
  INV_X1 U16955 ( .A(n14959), .ZN(n14964) );
  OAI211_X1 U16956 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14965), .A(
        n14964), .B(n17303), .ZN(n14971) );
  NAND2_X1 U16957 ( .A1(n14966), .A2(n14906), .ZN(n14969) );
  INV_X1 U16958 ( .A(n14967), .ZN(n14968) );
  AND2_X1 U16959 ( .A1(n14969), .A2(n14968), .ZN(n19531) );
  NAND2_X1 U16960 ( .A1(n17309), .A2(n19531), .ZN(n14970) );
  OAI211_X1 U16961 ( .C1(n17309), .C2(n15723), .A(n14971), .B(n14970), .ZN(
        P2_U2881) );
  OAI21_X1 U16962 ( .B1(n14974), .B2(n14973), .A(n14972), .ZN(n22243) );
  OR2_X1 U16963 ( .A1(n14976), .A2(n14975), .ZN(n14977) );
  NAND2_X1 U16964 ( .A1(n15115), .A2(n14977), .ZN(n22252) );
  INV_X1 U16965 ( .A(n22252), .ZN(n14978) );
  AOI22_X1 U16966 ( .A1(n20825), .A2(n14978), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n16714), .ZN(n14979) );
  OAI21_X1 U16967 ( .B1(n22243), .B2(n20812), .A(n14979), .ZN(P1_U2869) );
  INV_X1 U16968 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20938) );
  INV_X1 U16969 ( .A(DATAI_25_), .ZN(n14980) );
  OR2_X1 U16970 ( .A1(n15184), .A2(n14980), .ZN(n14981) );
  OAI21_X1 U16971 ( .B1(n15186), .B2(n20938), .A(n14981), .ZN(n22673) );
  INV_X1 U16972 ( .A(n11149), .ZN(n15449) );
  INV_X1 U16973 ( .A(n22548), .ZN(n15038) );
  INV_X1 U16974 ( .A(n15149), .ZN(n15145) );
  NOR2_X1 U16975 ( .A1(n15145), .A2(n17157), .ZN(n14983) );
  NAND3_X1 U16976 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15490) );
  INV_X1 U16977 ( .A(n15490), .ZN(n14982) );
  OAI21_X1 U16978 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n22393), .A(
        n15397), .ZN(n22572) );
  NAND2_X1 U16979 ( .A1(n22847), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14995) );
  INV_X1 U16980 ( .A(n15392), .ZN(n15057) );
  INV_X1 U16981 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20920) );
  INV_X1 U16982 ( .A(DATAI_17_), .ZN(n16816) );
  OR2_X1 U16983 ( .A1(n15184), .A2(n16816), .ZN(n14984) );
  OAI21_X1 U16984 ( .B1(n15186), .B2(n20920), .A(n14984), .ZN(n22672) );
  INV_X1 U16985 ( .A(n22671), .ZN(n15223) );
  NAND2_X1 U16986 ( .A1(n15397), .A2(n16814), .ZN(n22676) );
  INV_X1 U16987 ( .A(n22676), .ZN(n15524) );
  INV_X1 U16988 ( .A(n15059), .ZN(n17973) );
  OR2_X1 U16989 ( .A1(n17159), .A2(n17973), .ZN(n22630) );
  NOR2_X1 U16990 ( .A1(n14987), .A2(n22609), .ZN(n14988) );
  AND2_X1 U16991 ( .A1(n14988), .A2(n13313), .ZN(n15061) );
  INV_X1 U16992 ( .A(n15061), .ZN(n14991) );
  OAI22_X1 U16993 ( .A1(n22840), .A2(n22609), .B1(n15490), .B2(n22556), .ZN(
        n14989) );
  INV_X1 U16994 ( .A(n14989), .ZN(n14990) );
  OAI21_X1 U16995 ( .B1(n22630), .B2(n14991), .A(n14990), .ZN(n22843) );
  NAND2_X1 U16996 ( .A1(n15524), .A2(n22843), .ZN(n14992) );
  OAI21_X1 U16997 ( .B1(n15223), .B2(n22840), .A(n14992), .ZN(n14993) );
  AOI21_X1 U16998 ( .B1(n22846), .B2(n22672), .A(n14993), .ZN(n14994) );
  OAI211_X1 U16999 ( .C1(n15449), .C2(n22850), .A(n14995), .B(n14994), .ZN(
        P1_U3154) );
  INV_X1 U17000 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20936) );
  INV_X1 U17001 ( .A(DATAI_24_), .ZN(n14996) );
  OR2_X1 U17002 ( .A1(n15184), .A2(n14996), .ZN(n14997) );
  INV_X1 U17003 ( .A(n22655), .ZN(n22554) );
  NAND2_X1 U17004 ( .A1(n22847), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n15002) );
  INV_X1 U17005 ( .A(DATAI_16_), .ZN(n14998) );
  INV_X1 U17006 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20918) );
  OAI22_X1 U17007 ( .A1(n14998), .A2(n15184), .B1(n20918), .B2(n15186), .ZN(
        n22635) );
  INV_X1 U17008 ( .A(n22652), .ZN(n22617) );
  NAND2_X1 U17009 ( .A1(n15397), .A2(n16820), .ZN(n22644) );
  INV_X1 U17010 ( .A(n22644), .ZN(n22654) );
  NAND2_X1 U17011 ( .A1(n22654), .A2(n22843), .ZN(n14999) );
  OAI21_X1 U17012 ( .B1(n22617), .B2(n22840), .A(n14999), .ZN(n15000) );
  AOI21_X1 U17013 ( .B1(n22846), .B2(n22635), .A(n15000), .ZN(n15001) );
  OAI211_X1 U17014 ( .C1(n22554), .C2(n22850), .A(n15002), .B(n15001), .ZN(
        P1_U3153) );
  INV_X1 U17015 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20942) );
  INV_X1 U17016 ( .A(DATAI_27_), .ZN(n16764) );
  OR2_X1 U17017 ( .A1(n15184), .A2(n16764), .ZN(n15003) );
  OAI21_X1 U17018 ( .B1(n15186), .B2(n20942), .A(n15003), .ZN(n22710) );
  INV_X1 U17019 ( .A(n22710), .ZN(n15463) );
  NAND2_X1 U17020 ( .A1(n22847), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n15011) );
  INV_X1 U17021 ( .A(n15186), .ZN(n15004) );
  NAND2_X1 U17022 ( .A1(n15004), .A2(BUF1_REG_19__SCAN_IN), .ZN(n15006) );
  INV_X1 U17023 ( .A(DATAI_19_), .ZN(n16804) );
  OR2_X1 U17024 ( .A1(n15184), .A2(n16804), .ZN(n15005) );
  INV_X1 U17025 ( .A(n22708), .ZN(n22703) );
  NAND2_X1 U17026 ( .A1(n15397), .A2(n16802), .ZN(n22713) );
  INV_X1 U17027 ( .A(n22713), .ZN(n15502) );
  NAND2_X1 U17028 ( .A1(n15502), .A2(n22843), .ZN(n15008) );
  OAI21_X1 U17029 ( .B1(n22703), .B2(n22840), .A(n15008), .ZN(n15009) );
  AOI21_X1 U17030 ( .B1(n22846), .B2(n22709), .A(n15009), .ZN(n15010) );
  OAI211_X1 U17031 ( .C1(n15463), .C2(n22850), .A(n15011), .B(n15010), .ZN(
        P1_U3156) );
  INV_X1 U17032 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20946) );
  INV_X1 U17033 ( .A(DATAI_29_), .ZN(n15012) );
  OR2_X1 U17034 ( .A1(n15184), .A2(n15012), .ZN(n15013) );
  OAI21_X1 U17035 ( .B1(n15186), .B2(n20946), .A(n15013), .ZN(n22750) );
  INV_X1 U17036 ( .A(n22750), .ZN(n22735) );
  NAND2_X1 U17037 ( .A1(n22847), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n15021) );
  INV_X1 U17038 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20928) );
  INV_X1 U17039 ( .A(DATAI_21_), .ZN(n15014) );
  OR2_X1 U17040 ( .A1(n15184), .A2(n15014), .ZN(n15015) );
  OAI21_X1 U17041 ( .B1(n15186), .B2(n20928), .A(n15015), .ZN(n22749) );
  NAND2_X1 U17042 ( .A1(n15397), .A2(n15017), .ZN(n22753) );
  INV_X1 U17043 ( .A(n22753), .ZN(n15497) );
  NAND2_X1 U17044 ( .A1(n15497), .A2(n22843), .ZN(n15018) );
  OAI21_X1 U17045 ( .B1(n22743), .B2(n22840), .A(n15018), .ZN(n15019) );
  AOI21_X1 U17046 ( .B1(n22846), .B2(n22749), .A(n15019), .ZN(n15020) );
  OAI211_X1 U17047 ( .C1(n22735), .C2(n22850), .A(n15021), .B(n15020), .ZN(
        P1_U3158) );
  INV_X1 U17048 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20940) );
  INV_X1 U17049 ( .A(DATAI_26_), .ZN(n15022) );
  OR2_X1 U17050 ( .A1(n15184), .A2(n15022), .ZN(n15023) );
  INV_X1 U17051 ( .A(n22689), .ZN(n15454) );
  NAND2_X1 U17052 ( .A1(n22847), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n15029) );
  INV_X1 U17053 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20922) );
  INV_X1 U17054 ( .A(DATAI_18_), .ZN(n16810) );
  OR2_X1 U17055 ( .A1(n15184), .A2(n16810), .ZN(n15024) );
  INV_X1 U17056 ( .A(n22687), .ZN(n15219) );
  NAND2_X1 U17057 ( .A1(n15397), .A2(n16808), .ZN(n22692) );
  INV_X1 U17058 ( .A(n22692), .ZN(n15530) );
  NAND2_X1 U17059 ( .A1(n15530), .A2(n22843), .ZN(n15026) );
  OAI21_X1 U17060 ( .B1(n15219), .B2(n22840), .A(n15026), .ZN(n15027) );
  AOI21_X1 U17061 ( .B1(n22846), .B2(n22688), .A(n15027), .ZN(n15028) );
  OAI211_X1 U17062 ( .C1(n15454), .C2(n22850), .A(n15029), .B(n15028), .ZN(
        P1_U3155) );
  INV_X1 U17063 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20949) );
  INV_X1 U17064 ( .A(DATAI_30_), .ZN(n15030) );
  OR2_X1 U17065 ( .A1(n15184), .A2(n15030), .ZN(n15031) );
  OAI21_X1 U17066 ( .B1(n15186), .B2(n20949), .A(n15031), .ZN(n22771) );
  INV_X1 U17067 ( .A(n22771), .ZN(n22757) );
  NAND2_X1 U17068 ( .A1(n22847), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n15037) );
  INV_X1 U17069 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20930) );
  INV_X1 U17070 ( .A(DATAI_22_), .ZN(n16787) );
  OR2_X1 U17071 ( .A1(n15184), .A2(n16787), .ZN(n15032) );
  OAI21_X1 U17072 ( .B1(n15186), .B2(n20930), .A(n15032), .ZN(n22770) );
  INV_X1 U17073 ( .A(n22769), .ZN(n22756) );
  NAND2_X1 U17074 ( .A1(n15397), .A2(n16785), .ZN(n22774) );
  INV_X1 U17075 ( .A(n22774), .ZN(n15518) );
  NAND2_X1 U17076 ( .A1(n15518), .A2(n22843), .ZN(n15034) );
  OAI21_X1 U17077 ( .B1(n22756), .B2(n22840), .A(n15034), .ZN(n15035) );
  AOI21_X1 U17078 ( .B1(n22846), .B2(n11150), .A(n15035), .ZN(n15036) );
  OAI211_X1 U17079 ( .C1(n22757), .C2(n22850), .A(n15037), .B(n15036), .ZN(
        P1_U3159) );
  NOR2_X1 U17080 ( .A1(n15050), .A2(n17157), .ZN(n15039) );
  NAND3_X1 U17081 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n22552), .ZN(n22616) );
  INV_X1 U17082 ( .A(n22616), .ZN(n15040) );
  NAND2_X1 U17083 ( .A1(n22827), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n15043) );
  NAND2_X1 U17084 ( .A1(n22237), .A2(n17159), .ZN(n22612) );
  INV_X1 U17085 ( .A(n22612), .ZN(n15433) );
  NOR2_X1 U17086 ( .A1(n22567), .A2(n22616), .ZN(n22825) );
  INV_X1 U17087 ( .A(n22825), .ZN(n15231) );
  OAI22_X1 U17088 ( .A1(n22824), .A2(n22644), .B1(n22617), .B2(n15231), .ZN(
        n15041) );
  AOI21_X1 U17089 ( .B1(n22834), .B2(n22635), .A(n15041), .ZN(n15042) );
  OAI211_X1 U17090 ( .C1(n22554), .C2(n22830), .A(n15043), .B(n15042), .ZN(
        P1_U3121) );
  OR2_X1 U17091 ( .A1(n11254), .A2(n13311), .ZN(n15197) );
  INV_X1 U17092 ( .A(n15046), .ZN(n15200) );
  NAND3_X1 U17093 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n22552), .A3(
        n15199), .ZN(n15432) );
  NOR2_X1 U17094 ( .A1(n22567), .A2(n15432), .ZN(n22809) );
  AOI21_X1 U17095 ( .B1(n15433), .B2(n15200), .A(n22809), .ZN(n15049) );
  INV_X1 U17096 ( .A(n15049), .ZN(n15047) );
  INV_X1 U17097 ( .A(n15432), .ZN(n15052) );
  AOI22_X1 U17098 ( .A1(n15047), .A2(n17151), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15052), .ZN(n22808) );
  INV_X1 U17099 ( .A(n22809), .ZN(n15236) );
  OAI22_X1 U17100 ( .A1(n22808), .A2(n22644), .B1(n22617), .B2(n15236), .ZN(
        n15048) );
  AOI21_X1 U17101 ( .B1(n22819), .B2(n22635), .A(n15048), .ZN(n15054) );
  OAI211_X1 U17102 ( .C1(n15050), .C2(n22405), .A(n17151), .B(n15049), .ZN(
        n15051) );
  NAND2_X1 U17103 ( .A1(n22811), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n15053) );
  OAI211_X1 U17104 ( .C1(n22554), .C2(n22814), .A(n15054), .B(n15053), .ZN(
        P1_U3105) );
  INV_X1 U17105 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20717) );
  OAI222_X1 U17106 ( .A1(n22243), .A2(n16837), .B1(n16836), .B2(n15055), .C1(
        n16834), .C2(n20717), .ZN(P1_U2901) );
  INV_X1 U17107 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20934) );
  INV_X1 U17108 ( .A(DATAI_23_), .ZN(n16781) );
  OR2_X1 U17109 ( .A1(n15184), .A2(n16781), .ZN(n15056) );
  INV_X1 U17110 ( .A(n22845), .ZN(n22817) );
  INV_X1 U17111 ( .A(DATAI_31_), .ZN(n15058) );
  INV_X1 U17112 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20951) );
  OAI22_X1 U17113 ( .A1(n15058), .A2(n15184), .B1(n20951), .B2(n15186), .ZN(
        n22833) );
  NAND3_X1 U17114 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n22553), .ZN(n22588) );
  INV_X1 U17115 ( .A(n22588), .ZN(n15062) );
  NOR2_X1 U17116 ( .A1(n17159), .A2(n15059), .ZN(n22585) );
  NOR2_X1 U17117 ( .A1(n15060), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22597) );
  NAND2_X1 U17118 ( .A1(n15397), .A2(n16779), .ZN(n22838) );
  NOR2_X2 U17119 ( .A1(n15187), .A2(n16741), .ZN(n22841) );
  INV_X1 U17120 ( .A(n22841), .ZN(n22815) );
  INV_X1 U17121 ( .A(n22597), .ZN(n15246) );
  OAI22_X1 U17122 ( .A1(n22596), .A2(n22838), .B1(n22815), .B2(n15246), .ZN(
        n15063) );
  AOI21_X1 U17123 ( .B1(n22803), .B2(n22833), .A(n15063), .ZN(n15066) );
  OAI21_X1 U17124 ( .B1(n15118), .B2(n17157), .A(n22588), .ZN(n15064) );
  NAND2_X1 U17125 ( .A1(n15064), .A2(n15205), .ZN(n22599) );
  NAND2_X1 U17126 ( .A1(n22599), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n15065) );
  OAI211_X1 U17127 ( .C1(n22817), .C2(n22602), .A(n15066), .B(n15065), .ZN(
        P1_U3096) );
  INV_X1 U17128 ( .A(n22749), .ZN(n22744) );
  OAI22_X1 U17129 ( .A1(n22808), .A2(n22753), .B1(n22743), .B2(n15236), .ZN(
        n15067) );
  AOI21_X1 U17130 ( .B1(n15469), .B2(n22750), .A(n15067), .ZN(n15069) );
  NAND2_X1 U17131 ( .A1(n22811), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n15068) );
  OAI211_X1 U17132 ( .C1(n22744), .C2(n15240), .A(n15069), .B(n15068), .ZN(
        P1_U3110) );
  INV_X1 U17133 ( .A(n11150), .ZN(n15520) );
  OAI22_X1 U17134 ( .A1(n22808), .A2(n22774), .B1(n22756), .B2(n15236), .ZN(
        n15070) );
  AOI21_X1 U17135 ( .B1(n15469), .B2(n22771), .A(n15070), .ZN(n15072) );
  NAND2_X1 U17136 ( .A1(n22811), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n15071) );
  OAI211_X1 U17137 ( .C1(n15520), .C2(n15240), .A(n15072), .B(n15071), .ZN(
        P1_U3111) );
  INV_X1 U17138 ( .A(n22688), .ZN(n15532) );
  OAI22_X1 U17139 ( .A1(n22808), .A2(n22692), .B1(n15219), .B2(n15236), .ZN(
        n15073) );
  AOI21_X1 U17140 ( .B1(n15469), .B2(n22689), .A(n15073), .ZN(n15075) );
  NAND2_X1 U17141 ( .A1(n22811), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n15074) );
  OAI211_X1 U17142 ( .C1(n15532), .C2(n15240), .A(n15075), .B(n15074), .ZN(
        P1_U3107) );
  INV_X1 U17143 ( .A(n22672), .ZN(n15526) );
  OAI22_X1 U17144 ( .A1(n22808), .A2(n22676), .B1(n15223), .B2(n15236), .ZN(
        n15076) );
  AOI21_X1 U17145 ( .B1(n15469), .B2(n11149), .A(n15076), .ZN(n15078) );
  NAND2_X1 U17146 ( .A1(n22811), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n15077) );
  OAI211_X1 U17147 ( .C1(n15526), .C2(n15240), .A(n15078), .B(n15077), .ZN(
        P1_U3106) );
  OAI22_X1 U17148 ( .A1(n22808), .A2(n22713), .B1(n22703), .B2(n15236), .ZN(
        n15079) );
  AOI21_X1 U17149 ( .B1(n15469), .B2(n22710), .A(n15079), .ZN(n15081) );
  NAND2_X1 U17150 ( .A1(n22811), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n15080) );
  OAI211_X1 U17151 ( .C1(n22704), .C2(n15240), .A(n15081), .B(n15080), .ZN(
        P1_U3108) );
  OAI22_X1 U17152 ( .A1(n22596), .A2(n22676), .B1(n15223), .B2(n15246), .ZN(
        n15082) );
  AOI21_X1 U17153 ( .B1(n22605), .B2(n22672), .A(n15082), .ZN(n15084) );
  NAND2_X1 U17154 ( .A1(n22599), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n15083) );
  OAI211_X1 U17155 ( .C1(n15250), .C2(n15449), .A(n15084), .B(n15083), .ZN(
        P1_U3090) );
  OAI22_X1 U17156 ( .A1(n22596), .A2(n22713), .B1(n22703), .B2(n15246), .ZN(
        n15085) );
  AOI21_X1 U17157 ( .B1(n22605), .B2(n22709), .A(n15085), .ZN(n15087) );
  NAND2_X1 U17158 ( .A1(n22599), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n15086) );
  OAI211_X1 U17159 ( .C1(n15250), .C2(n15463), .A(n15087), .B(n15086), .ZN(
        P1_U3092) );
  OAI22_X1 U17160 ( .A1(n22596), .A2(n22692), .B1(n15219), .B2(n15246), .ZN(
        n15088) );
  AOI21_X1 U17161 ( .B1(n22605), .B2(n22688), .A(n15088), .ZN(n15090) );
  NAND2_X1 U17162 ( .A1(n22599), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n15089) );
  OAI211_X1 U17163 ( .C1(n15250), .C2(n15454), .A(n15090), .B(n15089), .ZN(
        P1_U3091) );
  OAI22_X1 U17164 ( .A1(n22596), .A2(n22774), .B1(n22756), .B2(n15246), .ZN(
        n15091) );
  AOI21_X1 U17165 ( .B1(n22605), .B2(n11150), .A(n15091), .ZN(n15093) );
  NAND2_X1 U17166 ( .A1(n22599), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n15092) );
  OAI211_X1 U17167 ( .C1(n15250), .C2(n22757), .A(n15093), .B(n15092), .ZN(
        P1_U3095) );
  OAI22_X1 U17168 ( .A1(n22596), .A2(n22753), .B1(n22743), .B2(n15246), .ZN(
        n15094) );
  AOI21_X1 U17169 ( .B1(n22605), .B2(n22749), .A(n15094), .ZN(n15096) );
  NAND2_X1 U17170 ( .A1(n22599), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n15095) );
  OAI211_X1 U17171 ( .C1(n15250), .C2(n22735), .A(n15096), .B(n15095), .ZN(
        P1_U3094) );
  INV_X1 U17172 ( .A(n22834), .ZN(n15235) );
  OAI22_X1 U17173 ( .A1(n22824), .A2(n22692), .B1(n15219), .B2(n15231), .ZN(
        n15097) );
  AOI21_X1 U17174 ( .B1(n22766), .B2(n22689), .A(n15097), .ZN(n15099) );
  NAND2_X1 U17175 ( .A1(n22827), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n15098) );
  OAI211_X1 U17176 ( .C1(n15532), .C2(n15235), .A(n15099), .B(n15098), .ZN(
        P1_U3123) );
  OAI22_X1 U17177 ( .A1(n22824), .A2(n22753), .B1(n22743), .B2(n15231), .ZN(
        n15100) );
  AOI21_X1 U17178 ( .B1(n22766), .B2(n22750), .A(n15100), .ZN(n15102) );
  NAND2_X1 U17179 ( .A1(n22827), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n15101) );
  OAI211_X1 U17180 ( .C1(n22744), .C2(n15235), .A(n15102), .B(n15101), .ZN(
        P1_U3126) );
  OAI22_X1 U17181 ( .A1(n22824), .A2(n22676), .B1(n15223), .B2(n15231), .ZN(
        n15103) );
  AOI21_X1 U17182 ( .B1(n22766), .B2(n11149), .A(n15103), .ZN(n15105) );
  NAND2_X1 U17183 ( .A1(n22827), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n15104) );
  OAI211_X1 U17184 ( .C1(n15526), .C2(n15235), .A(n15105), .B(n15104), .ZN(
        P1_U3122) );
  OAI22_X1 U17185 ( .A1(n22824), .A2(n22713), .B1(n22703), .B2(n15231), .ZN(
        n15106) );
  AOI21_X1 U17186 ( .B1(n22766), .B2(n22710), .A(n15106), .ZN(n15108) );
  NAND2_X1 U17187 ( .A1(n22827), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n15107) );
  OAI211_X1 U17188 ( .C1(n22704), .C2(n15235), .A(n15108), .B(n15107), .ZN(
        P1_U3124) );
  OAI22_X1 U17189 ( .A1(n22824), .A2(n22774), .B1(n22756), .B2(n15231), .ZN(
        n15109) );
  AOI21_X1 U17190 ( .B1(n22766), .B2(n22771), .A(n15109), .ZN(n15111) );
  NAND2_X1 U17191 ( .A1(n22827), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n15110) );
  OAI211_X1 U17192 ( .C1(n15520), .C2(n15235), .A(n15111), .B(n15110), .ZN(
        P1_U3127) );
  AOI21_X1 U17193 ( .B1(n15113), .B2(n14972), .A(n15112), .ZN(n15363) );
  INV_X1 U17194 ( .A(n15363), .ZN(n22260) );
  INV_X1 U17195 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n22256) );
  NAND2_X1 U17196 ( .A1(n15115), .A2(n15114), .ZN(n15116) );
  NAND2_X1 U17197 ( .A1(n15542), .A2(n15116), .ZN(n22257) );
  OAI222_X1 U17198 ( .A1(n22260), .A2(n20812), .B1(n22256), .B2(n20833), .C1(
        n22257), .C2(n20828), .ZN(P1_U2868) );
  INV_X1 U17199 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20719) );
  OAI222_X1 U17200 ( .A1(n22260), .A2(n16837), .B1(n16836), .B2(n15117), .C1(
        n20719), .C2(n16834), .ZN(P1_U2900) );
  NAND3_X1 U17201 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n22553), .A3(
        n15199), .ZN(n15396) );
  INV_X1 U17202 ( .A(n15396), .ZN(n15122) );
  NOR2_X1 U17203 ( .A1(n22567), .A2(n15396), .ZN(n22795) );
  AOI21_X1 U17204 ( .B1(n22585), .B2(n15200), .A(n22795), .ZN(n15121) );
  OAI211_X1 U17205 ( .C1(n15118), .C2(n22405), .A(n17151), .B(n15121), .ZN(
        n15119) );
  OAI211_X1 U17206 ( .C1(n17151), .C2(n15122), .A(n15119), .B(n15205), .ZN(
        n22797) );
  NAND2_X1 U17207 ( .A1(n22802), .A2(n22709), .ZN(n15126) );
  OR2_X1 U17208 ( .A1(n15121), .A2(n22609), .ZN(n15124) );
  NAND2_X1 U17209 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15122), .ZN(n15123) );
  NAND2_X1 U17210 ( .A1(n15124), .A2(n15123), .ZN(n22796) );
  AOI22_X1 U17211 ( .A1(n15502), .A2(n22796), .B1(n22708), .B2(n22795), .ZN(
        n15125) );
  OAI211_X1 U17212 ( .C1(n15463), .C2(n22800), .A(n15126), .B(n15125), .ZN(
        n15127) );
  AOI21_X1 U17213 ( .B1(n22797), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n15127), .ZN(n15128) );
  INV_X1 U17214 ( .A(n15128), .ZN(P1_U3076) );
  NAND2_X1 U17215 ( .A1(n22802), .A2(n22749), .ZN(n15130) );
  AOI22_X1 U17216 ( .A1(n15497), .A2(n22796), .B1(n22748), .B2(n22795), .ZN(
        n15129) );
  OAI211_X1 U17217 ( .C1(n22735), .C2(n22800), .A(n15130), .B(n15129), .ZN(
        n15131) );
  AOI21_X1 U17218 ( .B1(n22797), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15131), .ZN(n15132) );
  INV_X1 U17219 ( .A(n15132), .ZN(P1_U3078) );
  NAND2_X1 U17220 ( .A1(n11150), .A2(n22802), .ZN(n15134) );
  AOI22_X1 U17221 ( .A1(n15518), .A2(n22796), .B1(n22769), .B2(n22795), .ZN(
        n15133) );
  OAI211_X1 U17222 ( .C1(n22757), .C2(n22800), .A(n15134), .B(n15133), .ZN(
        n15135) );
  AOI21_X1 U17223 ( .B1(n22797), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n15135), .ZN(n15136) );
  INV_X1 U17224 ( .A(n15136), .ZN(P1_U3079) );
  NAND2_X1 U17225 ( .A1(n22672), .A2(n22802), .ZN(n15138) );
  AOI22_X1 U17226 ( .A1(n15524), .A2(n22796), .B1(n22671), .B2(n22795), .ZN(
        n15137) );
  OAI211_X1 U17227 ( .C1(n15449), .C2(n22800), .A(n15138), .B(n15137), .ZN(
        n15139) );
  AOI21_X1 U17228 ( .B1(n22797), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n15139), .ZN(n15140) );
  INV_X1 U17229 ( .A(n15140), .ZN(P1_U3074) );
  NAND2_X1 U17230 ( .A1(n22802), .A2(n22688), .ZN(n15142) );
  AOI22_X1 U17231 ( .A1(n15530), .A2(n22796), .B1(n22687), .B2(n22795), .ZN(
        n15141) );
  OAI211_X1 U17232 ( .C1(n15454), .C2(n22800), .A(n15142), .B(n15141), .ZN(
        n15143) );
  AOI21_X1 U17233 ( .B1(n22797), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n15143), .ZN(n15144) );
  INV_X1 U17234 ( .A(n15144), .ZN(P1_U3075) );
  NAND3_X1 U17235 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n15199), .ZN(n22634) );
  INV_X1 U17236 ( .A(n22634), .ZN(n15151) );
  INV_X1 U17237 ( .A(n22630), .ZN(n15488) );
  NOR2_X1 U17238 ( .A1(n22567), .A2(n22634), .ZN(n22645) );
  AOI21_X1 U17239 ( .B1(n15488), .B2(n15200), .A(n22645), .ZN(n15150) );
  OAI211_X1 U17240 ( .C1(n15145), .C2(n22405), .A(n17151), .B(n15150), .ZN(
        n15146) );
  OAI211_X1 U17241 ( .C1(n17151), .C2(n15151), .A(n15146), .B(n15205), .ZN(
        n22647) );
  NAND2_X1 U17242 ( .A1(n22832), .A2(n22771), .ZN(n15155) );
  OR2_X1 U17243 ( .A1(n15150), .A2(n22609), .ZN(n15153) );
  NAND2_X1 U17244 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15151), .ZN(n15152) );
  NAND2_X1 U17245 ( .A1(n15153), .A2(n15152), .ZN(n22646) );
  AOI22_X1 U17246 ( .A1(n15518), .A2(n22646), .B1(n22769), .B2(n22645), .ZN(
        n15154) );
  OAI211_X1 U17247 ( .C1(n15520), .C2(n22650), .A(n15155), .B(n15154), .ZN(
        n15156) );
  AOI21_X1 U17248 ( .B1(n22647), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n15156), .ZN(n15157) );
  INV_X1 U17249 ( .A(n15157), .ZN(P1_U3143) );
  NAND2_X1 U17250 ( .A1(n22832), .A2(n22750), .ZN(n15159) );
  AOI22_X1 U17251 ( .A1(n15497), .A2(n22646), .B1(n22748), .B2(n22645), .ZN(
        n15158) );
  OAI211_X1 U17252 ( .C1(n22744), .C2(n22650), .A(n15159), .B(n15158), .ZN(
        n15160) );
  AOI21_X1 U17253 ( .B1(n22647), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15160), .ZN(n15161) );
  INV_X1 U17254 ( .A(n15161), .ZN(P1_U3142) );
  NAND2_X1 U17255 ( .A1(n22832), .A2(n22689), .ZN(n15163) );
  AOI22_X1 U17256 ( .A1(n15530), .A2(n22646), .B1(n22687), .B2(n22645), .ZN(
        n15162) );
  OAI211_X1 U17257 ( .C1(n15532), .C2(n22650), .A(n15163), .B(n15162), .ZN(
        n15164) );
  AOI21_X1 U17258 ( .B1(n22647), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n15164), .ZN(n15165) );
  INV_X1 U17259 ( .A(n15165), .ZN(P1_U3139) );
  NAND2_X1 U17260 ( .A1(n11149), .A2(n22832), .ZN(n15167) );
  AOI22_X1 U17261 ( .A1(n15524), .A2(n22646), .B1(n22671), .B2(n22645), .ZN(
        n15166) );
  OAI211_X1 U17262 ( .C1(n15526), .C2(n22650), .A(n15167), .B(n15166), .ZN(
        n15168) );
  AOI21_X1 U17263 ( .B1(n22647), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n15168), .ZN(n15169) );
  INV_X1 U17264 ( .A(n15169), .ZN(P1_U3138) );
  NAND2_X1 U17265 ( .A1(n22710), .A2(n22832), .ZN(n15171) );
  AOI22_X1 U17266 ( .A1(n15502), .A2(n22646), .B1(n22708), .B2(n22645), .ZN(
        n15170) );
  OAI211_X1 U17267 ( .C1(n22704), .C2(n22650), .A(n15171), .B(n15170), .ZN(
        n15172) );
  AOI21_X1 U17268 ( .B1(n22647), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n15172), .ZN(n15173) );
  INV_X1 U17269 ( .A(n15173), .ZN(P1_U3140) );
  NAND2_X1 U17270 ( .A1(n22802), .A2(n22635), .ZN(n15175) );
  AOI22_X1 U17271 ( .A1(n22654), .A2(n22796), .B1(n22652), .B2(n22795), .ZN(
        n15174) );
  OAI211_X1 U17272 ( .C1(n22554), .C2(n22800), .A(n15175), .B(n15174), .ZN(
        n15176) );
  AOI21_X1 U17273 ( .B1(n22797), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n15176), .ZN(n15177) );
  INV_X1 U17274 ( .A(n15177), .ZN(P1_U3073) );
  NAND2_X1 U17275 ( .A1(n22832), .A2(n22833), .ZN(n15179) );
  AOI22_X1 U17276 ( .A1(n22844), .A2(n22646), .B1(n22841), .B2(n22645), .ZN(
        n15178) );
  OAI211_X1 U17277 ( .C1(n22817), .C2(n22650), .A(n15179), .B(n15178), .ZN(
        n15180) );
  AOI21_X1 U17278 ( .B1(n22647), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n15180), .ZN(n15181) );
  INV_X1 U17279 ( .A(n15181), .ZN(P1_U3144) );
  INV_X1 U17280 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20926) );
  INV_X1 U17281 ( .A(DATAI_20_), .ZN(n16799) );
  OR2_X1 U17282 ( .A1(n15184), .A2(n16799), .ZN(n15182) );
  OAI21_X1 U17283 ( .B1(n15186), .B2(n20926), .A(n15182), .ZN(n22728) );
  INV_X1 U17284 ( .A(n22728), .ZN(n15509) );
  INV_X1 U17285 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20944) );
  INV_X1 U17286 ( .A(DATAI_28_), .ZN(n15183) );
  OR2_X1 U17287 ( .A1(n15184), .A2(n15183), .ZN(n15185) );
  OAI21_X1 U17288 ( .B1(n15186), .B2(n20944), .A(n15185), .ZN(n22729) );
  NAND2_X1 U17289 ( .A1(n22832), .A2(n22729), .ZN(n15189) );
  NAND2_X1 U17290 ( .A1(n15397), .A2(n16797), .ZN(n22732) );
  INV_X1 U17291 ( .A(n22732), .ZN(n15507) );
  NOR2_X1 U17292 ( .A1(n15187), .A2(n12981), .ZN(n22727) );
  AOI22_X1 U17293 ( .A1(n15507), .A2(n22646), .B1(n22727), .B2(n22645), .ZN(
        n15188) );
  OAI211_X1 U17294 ( .C1(n15509), .C2(n22650), .A(n15189), .B(n15188), .ZN(
        n15190) );
  AOI21_X1 U17295 ( .B1(n22647), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n15190), .ZN(n15191) );
  INV_X1 U17296 ( .A(n15191), .ZN(P1_U3141) );
  INV_X1 U17297 ( .A(n22729), .ZN(n22717) );
  NAND2_X1 U17298 ( .A1(n22728), .A2(n22802), .ZN(n15193) );
  AOI22_X1 U17299 ( .A1(n15507), .A2(n22796), .B1(n22727), .B2(n22795), .ZN(
        n15192) );
  OAI211_X1 U17300 ( .C1(n22717), .C2(n22800), .A(n15193), .B(n15192), .ZN(
        n15194) );
  AOI21_X1 U17301 ( .B1(n22797), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n15194), .ZN(n15195) );
  INV_X1 U17302 ( .A(n15195), .ZN(P1_U3077) );
  INV_X1 U17303 ( .A(n17159), .ZN(n22224) );
  INV_X1 U17304 ( .A(n22566), .ZN(n15201) );
  NAND3_X1 U17305 ( .A1(n22553), .A2(n22552), .A3(n15199), .ZN(n22534) );
  NOR2_X1 U17306 ( .A1(n22567), .A2(n22534), .ZN(n22543) );
  AOI21_X1 U17307 ( .B1(n15201), .B2(n15200), .A(n22543), .ZN(n15204) );
  INV_X1 U17308 ( .A(n15204), .ZN(n15202) );
  INV_X1 U17309 ( .A(n22534), .ZN(n15207) );
  AOI22_X1 U17310 ( .A1(n15202), .A2(n17151), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15207), .ZN(n22542) );
  INV_X1 U17311 ( .A(n22543), .ZN(n15241) );
  OAI22_X1 U17312 ( .A1(n22542), .A2(n22838), .B1(n22815), .B2(n15241), .ZN(
        n15203) );
  AOI21_X1 U17313 ( .B1(n22776), .B2(n22833), .A(n15203), .ZN(n15209) );
  OAI211_X1 U17314 ( .C1(n22562), .C2(n22405), .A(n17151), .B(n15204), .ZN(
        n15206) );
  NAND2_X1 U17315 ( .A1(n22545), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n15208) );
  OAI211_X1 U17316 ( .C1(n22817), .C2(n22782), .A(n15209), .B(n15208), .ZN(
        P1_U3048) );
  OAI22_X1 U17317 ( .A1(n22542), .A2(n22713), .B1(n22703), .B2(n15241), .ZN(
        n15210) );
  AOI21_X1 U17318 ( .B1(n22696), .B2(n22709), .A(n15210), .ZN(n15212) );
  NAND2_X1 U17319 ( .A1(n22545), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15211) );
  OAI211_X1 U17320 ( .C1(n15245), .C2(n15463), .A(n15212), .B(n15211), .ZN(
        P1_U3044) );
  OAI22_X1 U17321 ( .A1(n22542), .A2(n22753), .B1(n22743), .B2(n15241), .ZN(
        n15213) );
  AOI21_X1 U17322 ( .B1(n22696), .B2(n22749), .A(n15213), .ZN(n15215) );
  NAND2_X1 U17323 ( .A1(n22545), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15214) );
  OAI211_X1 U17324 ( .C1(n15245), .C2(n22735), .A(n15215), .B(n15214), .ZN(
        P1_U3046) );
  OAI22_X1 U17325 ( .A1(n22542), .A2(n22774), .B1(n22756), .B2(n15241), .ZN(
        n15216) );
  AOI21_X1 U17326 ( .B1(n22696), .B2(n11150), .A(n15216), .ZN(n15218) );
  NAND2_X1 U17327 ( .A1(n22545), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n15217) );
  OAI211_X1 U17328 ( .C1(n15245), .C2(n22757), .A(n15218), .B(n15217), .ZN(
        P1_U3047) );
  OAI22_X1 U17329 ( .A1(n22542), .A2(n22692), .B1(n15219), .B2(n15241), .ZN(
        n15220) );
  AOI21_X1 U17330 ( .B1(n22696), .B2(n22688), .A(n15220), .ZN(n15222) );
  NAND2_X1 U17331 ( .A1(n22545), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n15221) );
  OAI211_X1 U17332 ( .C1(n15245), .C2(n15454), .A(n15222), .B(n15221), .ZN(
        P1_U3043) );
  OAI22_X1 U17333 ( .A1(n22542), .A2(n22676), .B1(n15223), .B2(n15241), .ZN(
        n15224) );
  AOI21_X1 U17334 ( .B1(n22696), .B2(n22672), .A(n15224), .ZN(n15226) );
  NAND2_X1 U17335 ( .A1(n22545), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n15225) );
  OAI211_X1 U17336 ( .C1(n15245), .C2(n15449), .A(n15226), .B(n15225), .ZN(
        P1_U3042) );
  NAND2_X1 U17337 ( .A1(n22847), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n15230) );
  INV_X1 U17338 ( .A(n22727), .ZN(n22716) );
  NAND2_X1 U17339 ( .A1(n15507), .A2(n22843), .ZN(n15227) );
  OAI21_X1 U17340 ( .B1(n22716), .B2(n22840), .A(n15227), .ZN(n15228) );
  AOI21_X1 U17341 ( .B1(n22846), .B2(n22728), .A(n15228), .ZN(n15229) );
  OAI211_X1 U17342 ( .C1(n22717), .C2(n22850), .A(n15230), .B(n15229), .ZN(
        P1_U3157) );
  OAI22_X1 U17343 ( .A1(n22824), .A2(n22732), .B1(n22716), .B2(n15231), .ZN(
        n15232) );
  AOI21_X1 U17344 ( .B1(n22766), .B2(n22729), .A(n15232), .ZN(n15234) );
  NAND2_X1 U17345 ( .A1(n22827), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n15233) );
  OAI211_X1 U17346 ( .C1(n15509), .C2(n15235), .A(n15234), .B(n15233), .ZN(
        P1_U3125) );
  OAI22_X1 U17347 ( .A1(n22808), .A2(n22732), .B1(n22716), .B2(n15236), .ZN(
        n15237) );
  AOI21_X1 U17348 ( .B1(n15469), .B2(n22729), .A(n15237), .ZN(n15239) );
  NAND2_X1 U17349 ( .A1(n22811), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n15238) );
  OAI211_X1 U17350 ( .C1(n15509), .C2(n15240), .A(n15239), .B(n15238), .ZN(
        P1_U3109) );
  OAI22_X1 U17351 ( .A1(n22542), .A2(n22732), .B1(n22716), .B2(n15241), .ZN(
        n15242) );
  AOI21_X1 U17352 ( .B1(n22696), .B2(n22728), .A(n15242), .ZN(n15244) );
  NAND2_X1 U17353 ( .A1(n22545), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n15243) );
  OAI211_X1 U17354 ( .C1(n15245), .C2(n22717), .A(n15244), .B(n15243), .ZN(
        P1_U3045) );
  OAI22_X1 U17355 ( .A1(n22596), .A2(n22732), .B1(n22716), .B2(n15246), .ZN(
        n15247) );
  AOI21_X1 U17356 ( .B1(n22605), .B2(n22728), .A(n15247), .ZN(n15249) );
  NAND2_X1 U17357 ( .A1(n22599), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n15248) );
  OAI211_X1 U17358 ( .C1(n15250), .C2(n22717), .A(n15249), .B(n15248), .ZN(
        P1_U3093) );
  OAI211_X1 U17359 ( .C1(n15252), .C2(n15254), .A(n15253), .B(n17303), .ZN(
        n15259) );
  AND2_X1 U17360 ( .A1(n15373), .A2(n15256), .ZN(n15257) );
  NOR2_X1 U17361 ( .A1(n15255), .A2(n15257), .ZN(n17906) );
  NAND2_X1 U17362 ( .A1(n17906), .A2(n17309), .ZN(n15258) );
  OAI211_X1 U17363 ( .C1(n17309), .C2(n12129), .A(n15259), .B(n15258), .ZN(
        P2_U2878) );
  NAND2_X1 U17364 ( .A1(n19551), .A2(n15304), .ZN(n15273) );
  NAND2_X1 U17365 ( .A1(n15261), .A2(n15260), .ZN(n15286) );
  INV_X1 U17366 ( .A(n15286), .ZN(n15270) );
  INV_X1 U17367 ( .A(n11781), .ZN(n15262) );
  NAND2_X1 U17368 ( .A1(n15262), .A2(n11232), .ZN(n15290) );
  NAND2_X1 U17369 ( .A1(n15285), .A2(n15290), .ZN(n15269) );
  NAND2_X1 U17370 ( .A1(n15263), .A2(n15333), .ZN(n15291) );
  NAND2_X1 U17371 ( .A1(n15291), .A2(n15269), .ZN(n15268) );
  INV_X1 U17372 ( .A(n15264), .ZN(n15265) );
  OAI21_X1 U17373 ( .B1(n17957), .B2(n11476), .A(n15265), .ZN(n15266) );
  NAND2_X1 U17374 ( .A1(n12817), .A2(n15266), .ZN(n15267) );
  OAI211_X1 U17375 ( .C1(n15270), .C2(n15269), .A(n15268), .B(n15267), .ZN(
        n15271) );
  INV_X1 U17376 ( .A(n15271), .ZN(n15272) );
  NAND2_X1 U17377 ( .A1(n15273), .A2(n15272), .ZN(n17956) );
  INV_X1 U17378 ( .A(n15274), .ZN(n15277) );
  NOR2_X1 U17379 ( .A1(n12019), .A2(n15275), .ZN(n15276) );
  NAND2_X1 U17380 ( .A1(n15277), .A2(n15276), .ZN(n15281) );
  NAND4_X1 U17381 ( .A1(n15281), .A2(n15280), .A3(n15279), .A4(n15278), .ZN(
        n15819) );
  INV_X1 U17382 ( .A(n15819), .ZN(n15313) );
  OR2_X1 U17383 ( .A1(n17956), .A2(n15313), .ZN(n15283) );
  NAND2_X1 U17384 ( .A1(n15313), .A2(n11232), .ZN(n15282) );
  NAND2_X1 U17385 ( .A1(n15283), .A2(n15282), .ZN(n15352) );
  AND2_X1 U17386 ( .A1(n17957), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15289) );
  INV_X1 U17387 ( .A(n15289), .ZN(n15284) );
  NAND2_X1 U17388 ( .A1(n12817), .A2(n15284), .ZN(n15288) );
  NAND2_X1 U17389 ( .A1(n15286), .A2(n15285), .ZN(n15287) );
  AND3_X1 U17390 ( .A1(n15288), .A2(n15287), .A3(n15290), .ZN(n15293) );
  AOI22_X1 U17391 ( .A1(n15291), .A2(n15290), .B1(n15289), .B2(n12817), .ZN(
        n15292) );
  MUX2_X1 U17392 ( .A(n15293), .B(n15292), .S(n15297), .Z(n15295) );
  NAND2_X1 U17393 ( .A1(n15295), .A2(n15294), .ZN(n15296) );
  AOI21_X1 U17394 ( .B1(n11261), .B2(n15304), .A(n15296), .ZN(n17960) );
  MUX2_X1 U17395 ( .A(n15297), .B(n17960), .S(n15819), .Z(n15351) );
  INV_X1 U17396 ( .A(n15298), .ZN(n15299) );
  NOR2_X1 U17397 ( .A1(n15299), .A2(n11236), .ZN(n15307) );
  NOR2_X1 U17398 ( .A1(n11780), .A2(n15300), .ZN(n15302) );
  NAND2_X1 U17399 ( .A1(n12817), .A2(n11476), .ZN(n15301) );
  OAI21_X1 U17400 ( .B1(n15307), .B2(n15302), .A(n15301), .ZN(n15303) );
  AOI21_X1 U17401 ( .B1(n17238), .B2(n15304), .A(n15303), .ZN(n17950) );
  INV_X1 U17402 ( .A(n15304), .ZN(n15305) );
  OR2_X1 U17403 ( .A1(n19515), .A2(n15305), .ZN(n15310) );
  INV_X1 U17404 ( .A(n12817), .ZN(n15308) );
  MUX2_X1 U17405 ( .A(n15308), .B(n15307), .S(n15306), .Z(n15309) );
  NAND2_X1 U17406 ( .A1(n15310), .A2(n15309), .ZN(n15818) );
  AOI21_X1 U17407 ( .B1(n15818), .B2(n20245), .A(n20205), .ZN(n15311) );
  AND2_X1 U17408 ( .A1(n17950), .A2(n15311), .ZN(n15312) );
  OAI22_X1 U17409 ( .A1(n15352), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n15313), .B2(n15312), .ZN(n15319) );
  OAI21_X1 U17410 ( .B1(n15818), .B2(n15314), .A(n20161), .ZN(n15317) );
  NOR2_X1 U17411 ( .A1(n15818), .A2(n15315), .ZN(n15316) );
  AOI21_X1 U17412 ( .B1(n15352), .B2(n15317), .A(n15316), .ZN(n15318) );
  NAND2_X1 U17413 ( .A1(n15319), .A2(n15318), .ZN(n15320) );
  NAND2_X1 U17414 ( .A1(n15320), .A2(n15351), .ZN(n15323) );
  OR2_X1 U17415 ( .A1(n15320), .A2(n15351), .ZN(n15321) );
  AOI21_X1 U17416 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15321), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15322) );
  NAND2_X1 U17417 ( .A1(n15323), .A2(n15322), .ZN(n15350) );
  INV_X1 U17418 ( .A(n15324), .ZN(n15328) );
  AOI22_X1 U17419 ( .A1(n15326), .A2(n15325), .B1(n15339), .B2(n15337), .ZN(
        n15327) );
  OAI21_X1 U17420 ( .B1(n19568), .B2(n15328), .A(n15327), .ZN(n15329) );
  INV_X1 U17421 ( .A(n15329), .ZN(n15332) );
  NAND2_X1 U17422 ( .A1(n15764), .A2(n15330), .ZN(n15331) );
  OAI211_X1 U17423 ( .C1(n15333), .C2(n15764), .A(n15332), .B(n15331), .ZN(
        n19582) );
  INV_X1 U17424 ( .A(n19582), .ZN(n15347) );
  NOR2_X1 U17425 ( .A1(n15335), .A2(n15334), .ZN(n15336) );
  NAND2_X1 U17426 ( .A1(n15337), .A2(n15336), .ZN(n15338) );
  NOR2_X1 U17427 ( .A1(n15339), .A2(n15338), .ZN(n19581) );
  OAI21_X1 U17428 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19581), .ZN(n15343) );
  AND2_X1 U17429 ( .A1(n11394), .A2(n15340), .ZN(n15341) );
  NAND2_X1 U17430 ( .A1(n15342), .A2(n15341), .ZN(n19506) );
  NAND2_X1 U17431 ( .A1(n15343), .A2(n19506), .ZN(n15344) );
  NOR2_X1 U17432 ( .A1(n15345), .A2(n15344), .ZN(n15346) );
  OAI211_X1 U17433 ( .C1(n15819), .C2(n19509), .A(n15347), .B(n15346), .ZN(
        n15348) );
  INV_X1 U17434 ( .A(n15348), .ZN(n15349) );
  OAI211_X1 U17435 ( .C1(n15352), .C2(n15351), .A(n15350), .B(n15349), .ZN(
        n19569) );
  NAND2_X1 U17436 ( .A1(n17948), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15353) );
  OAI21_X1 U17437 ( .B1(n19569), .B2(n15353), .A(n15765), .ZN(n15356) );
  NAND2_X1 U17438 ( .A1(n12058), .A2(n15354), .ZN(n15355) );
  OAI21_X1 U17439 ( .B1(n19571), .B2(n17995), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n15358) );
  NOR2_X1 U17440 ( .A1(n17995), .A2(n18096), .ZN(n19567) );
  INV_X1 U17441 ( .A(n19567), .ZN(n15357) );
  NAND2_X1 U17442 ( .A1(n15358), .A2(n15357), .ZN(P2_U3593) );
  XOR2_X1 U17443 ( .A(n15360), .B(n15359), .Z(n22153) );
  INV_X1 U17444 ( .A(n22153), .ZN(n15365) );
  NAND2_X1 U17445 ( .A1(n22202), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n22150) );
  NAND2_X1 U17446 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15361) );
  OAI211_X1 U17447 ( .C1(n20877), .C2(n22258), .A(n22150), .B(n15361), .ZN(
        n15362) );
  AOI21_X1 U17448 ( .B1(n15363), .B2(n20873), .A(n15362), .ZN(n15364) );
  OAI21_X1 U17449 ( .B1(n15365), .B2(n22385), .A(n15364), .ZN(P1_U2995) );
  OR2_X1 U17450 ( .A1(n15112), .A2(n15367), .ZN(n15368) );
  AND2_X1 U17451 ( .A1(n15366), .A2(n15368), .ZN(n22276) );
  INV_X1 U17452 ( .A(n22276), .ZN(n15369) );
  INV_X1 U17453 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20721) );
  OAI222_X1 U17454 ( .A1(n15369), .A2(n16837), .B1(n16836), .B2(n16791), .C1(
        n16834), .C2(n20721), .ZN(P1_U2899) );
  NAND2_X1 U17455 ( .A1(n15371), .A2(n15370), .ZN(n15372) );
  NAND2_X1 U17456 ( .A1(n15373), .A2(n15372), .ZN(n19294) );
  NOR2_X1 U17457 ( .A1(n15680), .A2(n19294), .ZN(n15377) );
  AOI211_X1 U17458 ( .C1(n15375), .C2(n15374), .A(n17316), .B(n15252), .ZN(
        n15376) );
  AOI211_X1 U17459 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n15680), .A(n15377), .B(
        n15376), .ZN(n15378) );
  INV_X1 U17460 ( .A(n15378), .ZN(P2_U2879) );
  XNOR2_X1 U17461 ( .A(n15380), .B(n15379), .ZN(n22156) );
  NAND2_X1 U17462 ( .A1(n22202), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n22157) );
  OAI21_X1 U17463 ( .B1(n20842), .B2(n15381), .A(n22157), .ZN(n15383) );
  NOR2_X1 U17464 ( .A1(n22243), .A2(n20853), .ZN(n15382) );
  AOI211_X1 U17465 ( .C1(n20862), .C2(n22245), .A(n15383), .B(n15382), .ZN(
        n15384) );
  OAI21_X1 U17466 ( .B1(n22385), .B2(n22156), .A(n15384), .ZN(P1_U2996) );
  XNOR2_X1 U17467 ( .A(n15385), .B(n15386), .ZN(n15391) );
  INV_X1 U17468 ( .A(n15387), .ZN(n15678) );
  NAND2_X1 U17469 ( .A1(n15588), .A2(n15388), .ZN(n15389) );
  NAND2_X1 U17470 ( .A1(n15678), .A2(n15389), .ZN(n19306) );
  MUX2_X1 U17471 ( .A(n19306), .B(n12135), .S(n15680), .Z(n15390) );
  OAI21_X1 U17472 ( .B1(n15391), .B2(n17316), .A(n15390), .ZN(P2_U2876) );
  INV_X1 U17473 ( .A(n22800), .ZN(n15393) );
  OAI21_X1 U17474 ( .B1(n22790), .B2(n15393), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15395) );
  NAND2_X1 U17475 ( .A1(n22585), .A2(n22611), .ZN(n15402) );
  AOI21_X1 U17476 ( .B1(n15395), .B2(n15402), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15398) );
  NOR2_X1 U17477 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15396), .ZN(
        n22579) );
  NOR2_X1 U17478 ( .A1(n15399), .A2(n22556), .ZN(n22613) );
  INV_X1 U17479 ( .A(n15397), .ZN(n15435) );
  OAI21_X1 U17480 ( .B1(n15398), .B2(n22579), .A(n22639), .ZN(n22581) );
  INV_X1 U17481 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15406) );
  AND2_X1 U17482 ( .A1(n15399), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22632) );
  INV_X1 U17483 ( .A(n22632), .ZN(n15401) );
  INV_X1 U17484 ( .A(n15437), .ZN(n15400) );
  INV_X1 U17485 ( .A(n15491), .ZN(n22550) );
  NAND2_X1 U17486 ( .A1(n15400), .A2(n22550), .ZN(n22536) );
  OAI22_X1 U17487 ( .A1(n15402), .A2(n22609), .B1(n15401), .B2(n22536), .ZN(
        n22580) );
  AOI22_X1 U17488 ( .A1(n15502), .A2(n22580), .B1(n22708), .B2(n22579), .ZN(
        n15403) );
  OAI21_X1 U17489 ( .B1(n22800), .B2(n22704), .A(n15403), .ZN(n15404) );
  AOI21_X1 U17490 ( .B1(n22790), .B2(n22710), .A(n15404), .ZN(n15405) );
  OAI21_X1 U17491 ( .B1(n15431), .B2(n15406), .A(n15405), .ZN(P1_U3068) );
  INV_X1 U17492 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U17493 ( .A1(n22844), .A2(n22580), .B1(n22841), .B2(n22579), .ZN(
        n15407) );
  OAI21_X1 U17494 ( .B1(n22800), .B2(n22817), .A(n15407), .ZN(n15408) );
  AOI21_X1 U17495 ( .B1(n22790), .B2(n22833), .A(n15408), .ZN(n15409) );
  OAI21_X1 U17496 ( .B1(n15431), .B2(n15410), .A(n15409), .ZN(P1_U3072) );
  INV_X1 U17497 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U17498 ( .A1(n15530), .A2(n22580), .B1(n22687), .B2(n22579), .ZN(
        n15411) );
  OAI21_X1 U17499 ( .B1(n22800), .B2(n15532), .A(n15411), .ZN(n15412) );
  AOI21_X1 U17500 ( .B1(n22790), .B2(n22689), .A(n15412), .ZN(n15413) );
  OAI21_X1 U17501 ( .B1(n15431), .B2(n15414), .A(n15413), .ZN(P1_U3067) );
  INV_X1 U17502 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U17503 ( .A1(n15507), .A2(n22580), .B1(n22727), .B2(n22579), .ZN(
        n15415) );
  OAI21_X1 U17504 ( .B1(n22800), .B2(n15509), .A(n15415), .ZN(n15416) );
  AOI21_X1 U17505 ( .B1(n22790), .B2(n22729), .A(n15416), .ZN(n15417) );
  OAI21_X1 U17506 ( .B1(n15431), .B2(n15418), .A(n15417), .ZN(P1_U3069) );
  INV_X1 U17507 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U17508 ( .A1(n15497), .A2(n22580), .B1(n22748), .B2(n22579), .ZN(
        n15419) );
  OAI21_X1 U17509 ( .B1(n22800), .B2(n22744), .A(n15419), .ZN(n15420) );
  AOI21_X1 U17510 ( .B1(n22790), .B2(n22750), .A(n15420), .ZN(n15421) );
  OAI21_X1 U17511 ( .B1(n15431), .B2(n15422), .A(n15421), .ZN(P1_U3070) );
  INV_X1 U17512 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15426) );
  AOI22_X1 U17513 ( .A1(n15518), .A2(n22580), .B1(n22769), .B2(n22579), .ZN(
        n15423) );
  OAI21_X1 U17514 ( .B1(n22800), .B2(n15520), .A(n15423), .ZN(n15424) );
  AOI21_X1 U17515 ( .B1(n22790), .B2(n22771), .A(n15424), .ZN(n15425) );
  OAI21_X1 U17516 ( .B1(n15431), .B2(n15426), .A(n15425), .ZN(P1_U3071) );
  INV_X1 U17517 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U17518 ( .A1(n15524), .A2(n22580), .B1(n22671), .B2(n22579), .ZN(
        n15427) );
  OAI21_X1 U17519 ( .B1(n22800), .B2(n15526), .A(n15427), .ZN(n15428) );
  AOI21_X1 U17520 ( .B1(n22790), .B2(n11149), .A(n15428), .ZN(n15429) );
  OAI21_X1 U17521 ( .B1(n15431), .B2(n15430), .A(n15429), .ZN(P1_U3066) );
  NOR2_X1 U17522 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15432), .ZN(
        n22603) );
  OAI21_X1 U17523 ( .B1(n15469), .B2(n22605), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15434) );
  AOI21_X1 U17524 ( .B1(n15433), .B2(n22611), .A(n22603), .ZN(n15439) );
  NAND2_X1 U17525 ( .A1(n15434), .A2(n15439), .ZN(n15436) );
  OAI211_X1 U17526 ( .C1(n22603), .C2(n22393), .A(n15436), .B(n22622), .ZN(
        n22606) );
  INV_X1 U17527 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15443) );
  NAND2_X1 U17528 ( .A1(n15437), .A2(n22550), .ZN(n22637) );
  INV_X1 U17529 ( .A(n22613), .ZN(n15438) );
  OAI22_X1 U17530 ( .A1(n15439), .A2(n22609), .B1(n22637), .B2(n15438), .ZN(
        n22604) );
  AOI22_X1 U17531 ( .A1(n22604), .A2(n15518), .B1(n22769), .B2(n22603), .ZN(
        n15440) );
  OAI21_X1 U17532 ( .B1(n22602), .B2(n22757), .A(n15440), .ZN(n15441) );
  AOI21_X1 U17533 ( .B1(n15469), .B2(n11150), .A(n15441), .ZN(n15442) );
  OAI21_X1 U17534 ( .B1(n15472), .B2(n15443), .A(n15442), .ZN(P1_U3103) );
  INV_X1 U17535 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15447) );
  INV_X1 U17536 ( .A(n22833), .ZN(n22851) );
  AOI22_X1 U17537 ( .A1(n22604), .A2(n22844), .B1(n22841), .B2(n22603), .ZN(
        n15444) );
  OAI21_X1 U17538 ( .B1(n22602), .B2(n22851), .A(n15444), .ZN(n15445) );
  AOI21_X1 U17539 ( .B1(n15469), .B2(n22845), .A(n15445), .ZN(n15446) );
  OAI21_X1 U17540 ( .B1(n15472), .B2(n15447), .A(n15446), .ZN(P1_U3104) );
  INV_X1 U17541 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U17542 ( .A1(n22604), .A2(n15524), .B1(n22671), .B2(n22603), .ZN(
        n15448) );
  OAI21_X1 U17543 ( .B1(n22602), .B2(n15449), .A(n15448), .ZN(n15450) );
  AOI21_X1 U17544 ( .B1(n15469), .B2(n22672), .A(n15450), .ZN(n15451) );
  OAI21_X1 U17545 ( .B1(n15472), .B2(n15452), .A(n15451), .ZN(P1_U3098) );
  INV_X1 U17546 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U17547 ( .A1(n22604), .A2(n15530), .B1(n22687), .B2(n22603), .ZN(
        n15453) );
  OAI21_X1 U17548 ( .B1(n22602), .B2(n15454), .A(n15453), .ZN(n15455) );
  AOI21_X1 U17549 ( .B1(n15469), .B2(n22688), .A(n15455), .ZN(n15456) );
  OAI21_X1 U17550 ( .B1(n15472), .B2(n15457), .A(n15456), .ZN(P1_U3099) );
  INV_X1 U17551 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15461) );
  AOI22_X1 U17552 ( .A1(n22604), .A2(n15507), .B1(n22727), .B2(n22603), .ZN(
        n15458) );
  OAI21_X1 U17553 ( .B1(n22602), .B2(n22717), .A(n15458), .ZN(n15459) );
  AOI21_X1 U17554 ( .B1(n15469), .B2(n22728), .A(n15459), .ZN(n15460) );
  OAI21_X1 U17555 ( .B1(n15472), .B2(n15461), .A(n15460), .ZN(P1_U3101) );
  INV_X1 U17556 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U17557 ( .A1(n22604), .A2(n15502), .B1(n22708), .B2(n22603), .ZN(
        n15462) );
  OAI21_X1 U17558 ( .B1(n22602), .B2(n15463), .A(n15462), .ZN(n15464) );
  AOI21_X1 U17559 ( .B1(n15469), .B2(n22709), .A(n15464), .ZN(n15465) );
  OAI21_X1 U17560 ( .B1(n15472), .B2(n15466), .A(n15465), .ZN(P1_U3100) );
  INV_X1 U17561 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U17562 ( .A1(n22604), .A2(n15497), .B1(n22748), .B2(n22603), .ZN(
        n15467) );
  OAI21_X1 U17563 ( .B1(n22602), .B2(n22735), .A(n15467), .ZN(n15468) );
  AOI21_X1 U17564 ( .B1(n15469), .B2(n22749), .A(n15468), .ZN(n15470) );
  OAI21_X1 U17565 ( .B1(n15472), .B2(n15471), .A(n15470), .ZN(P1_U3102) );
  XOR2_X1 U17566 ( .A(n15474), .B(n15473), .Z(n20835) );
  INV_X1 U17567 ( .A(n20835), .ZN(n15487) );
  NAND2_X1 U17568 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n22144) );
  OAI22_X1 U17569 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15476), .B1(
        n17125), .B2(n15475), .ZN(n22162) );
  OAI21_X1 U17570 ( .B1(n22144), .B2(n22162), .A(n15477), .ZN(n15485) );
  NOR2_X1 U17571 ( .A1(n15477), .A2(n22144), .ZN(n15573) );
  NAND3_X1 U17572 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n15573), .ZN(n16973) );
  INV_X1 U17573 ( .A(n16973), .ZN(n15478) );
  OAI21_X1 U17574 ( .B1(n17122), .B2(n15478), .A(n22118), .ZN(n15479) );
  INV_X1 U17575 ( .A(n15479), .ZN(n15482) );
  NAND2_X1 U17576 ( .A1(n15573), .A2(n15480), .ZN(n16969) );
  NAND2_X1 U17577 ( .A1(n17125), .A2(n16969), .ZN(n15481) );
  NAND2_X1 U17578 ( .A1(n15482), .A2(n15481), .ZN(n15645) );
  INV_X1 U17579 ( .A(n15483), .ZN(n15541) );
  XNOR2_X1 U17580 ( .A(n15542), .B(n15541), .ZN(n22267) );
  NAND2_X1 U17581 ( .A1(n22202), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n20836) );
  OAI21_X1 U17582 ( .B1(n22214), .B2(n22267), .A(n20836), .ZN(n15484) );
  AOI21_X1 U17583 ( .B1(n15485), .B2(n15645), .A(n15484), .ZN(n15486) );
  OAI21_X1 U17584 ( .B1(n15487), .B2(n22218), .A(n15486), .ZN(P1_U3026) );
  INV_X1 U17585 ( .A(n22850), .ZN(n15515) );
  OAI21_X1 U17586 ( .B1(n22656), .B2(n15515), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15489) );
  INV_X1 U17587 ( .A(n22611), .ZN(n22629) );
  NAND2_X1 U17588 ( .A1(n15488), .A2(n22629), .ZN(n15493) );
  AOI21_X1 U17589 ( .B1(n15489), .B2(n15493), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15492) );
  NOR2_X1 U17590 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15490), .ZN(
        n22651) );
  NAND2_X1 U17591 ( .A1(n15491), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15494) );
  NAND2_X1 U17592 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15494), .ZN(n22619) );
  OAI211_X1 U17593 ( .C1(n15492), .C2(n22651), .A(n22619), .B(n22639), .ZN(
        n22657) );
  INV_X1 U17594 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15501) );
  OR2_X1 U17595 ( .A1(n15493), .A2(n22609), .ZN(n15496) );
  INV_X1 U17596 ( .A(n15494), .ZN(n22614) );
  NAND2_X1 U17597 ( .A1(n22632), .A2(n22614), .ZN(n15495) );
  NAND2_X1 U17598 ( .A1(n15496), .A2(n15495), .ZN(n22653) );
  AOI22_X1 U17599 ( .A1(n15497), .A2(n22653), .B1(n22748), .B2(n22651), .ZN(
        n15498) );
  OAI21_X1 U17600 ( .B1(n22850), .B2(n22744), .A(n15498), .ZN(n15499) );
  AOI21_X1 U17601 ( .B1(n22656), .B2(n22750), .A(n15499), .ZN(n15500) );
  OAI21_X1 U17602 ( .B1(n15536), .B2(n15501), .A(n15500), .ZN(P1_U3150) );
  INV_X1 U17603 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U17604 ( .A1(n15502), .A2(n22653), .B1(n22708), .B2(n22651), .ZN(
        n15503) );
  OAI21_X1 U17605 ( .B1(n22850), .B2(n22704), .A(n15503), .ZN(n15504) );
  AOI21_X1 U17606 ( .B1(n22656), .B2(n22710), .A(n15504), .ZN(n15505) );
  OAI21_X1 U17607 ( .B1(n15536), .B2(n15506), .A(n15505), .ZN(P1_U3148) );
  INV_X1 U17608 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15512) );
  AOI22_X1 U17609 ( .A1(n15507), .A2(n22653), .B1(n22727), .B2(n22651), .ZN(
        n15508) );
  OAI21_X1 U17610 ( .B1(n22850), .B2(n15509), .A(n15508), .ZN(n15510) );
  AOI21_X1 U17611 ( .B1(n22656), .B2(n22729), .A(n15510), .ZN(n15511) );
  OAI21_X1 U17612 ( .B1(n15536), .B2(n15512), .A(n15511), .ZN(P1_U3149) );
  INV_X1 U17613 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15517) );
  AOI22_X1 U17614 ( .A1(n22844), .A2(n22653), .B1(n22841), .B2(n22651), .ZN(
        n15513) );
  OAI21_X1 U17615 ( .B1(n22650), .B2(n22851), .A(n15513), .ZN(n15514) );
  AOI21_X1 U17616 ( .B1(n15515), .B2(n22845), .A(n15514), .ZN(n15516) );
  OAI21_X1 U17617 ( .B1(n15536), .B2(n15517), .A(n15516), .ZN(P1_U3152) );
  INV_X1 U17618 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15523) );
  AOI22_X1 U17619 ( .A1(n15518), .A2(n22653), .B1(n22769), .B2(n22651), .ZN(
        n15519) );
  OAI21_X1 U17620 ( .B1(n22850), .B2(n15520), .A(n15519), .ZN(n15521) );
  AOI21_X1 U17621 ( .B1(n22656), .B2(n22771), .A(n15521), .ZN(n15522) );
  OAI21_X1 U17622 ( .B1(n15536), .B2(n15523), .A(n15522), .ZN(P1_U3151) );
  INV_X1 U17623 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15529) );
  AOI22_X1 U17624 ( .A1(n15524), .A2(n22653), .B1(n22671), .B2(n22651), .ZN(
        n15525) );
  OAI21_X1 U17625 ( .B1(n22850), .B2(n15526), .A(n15525), .ZN(n15527) );
  AOI21_X1 U17626 ( .B1(n22656), .B2(n11149), .A(n15527), .ZN(n15528) );
  OAI21_X1 U17627 ( .B1(n15536), .B2(n15529), .A(n15528), .ZN(P1_U3146) );
  INV_X1 U17628 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15535) );
  AOI22_X1 U17629 ( .A1(n15530), .A2(n22653), .B1(n22687), .B2(n22651), .ZN(
        n15531) );
  OAI21_X1 U17630 ( .B1(n22850), .B2(n15532), .A(n15531), .ZN(n15533) );
  AOI21_X1 U17631 ( .B1(n22656), .B2(n22689), .A(n15533), .ZN(n15534) );
  OAI21_X1 U17632 ( .B1(n15536), .B2(n15535), .A(n15534), .ZN(P1_U3147) );
  AOI21_X1 U17633 ( .B1(n15538), .B2(n15366), .A(n13361), .ZN(n22287) );
  INV_X1 U17634 ( .A(n22287), .ZN(n15545) );
  OAI222_X1 U17635 ( .A1(n15545), .A2(n16837), .B1(n16836), .B2(n15539), .C1(
        n16834), .C2(n13348), .ZN(P1_U2898) );
  INV_X1 U17636 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n22280) );
  OAI21_X1 U17637 ( .B1(n15542), .B2(n15541), .A(n15540), .ZN(n15543) );
  INV_X1 U17638 ( .A(n15543), .ZN(n15544) );
  OR2_X1 U17639 ( .A1(n15544), .A2(n15595), .ZN(n22281) );
  OAI222_X1 U17640 ( .A1(n15545), .A2(n20812), .B1(n22280), .B2(n20833), .C1(
        n22281), .C2(n20828), .ZN(P1_U2866) );
  XNOR2_X1 U17641 ( .A(n15546), .B(n15547), .ZN(n15570) );
  XOR2_X1 U17642 ( .A(n15548), .B(n15549), .Z(n15568) );
  NAND2_X1 U17643 ( .A1(n11261), .A2(n18088), .ZN(n15551) );
  INV_X1 U17644 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n16085) );
  NOR2_X1 U17645 ( .A1(n19301), .A2(n16085), .ZN(n15557) );
  AOI21_X1 U17646 ( .B1(n17612), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15557), .ZN(n15550) );
  OAI211_X1 U17647 ( .C1(n16082), .C2(n17638), .A(n15551), .B(n15550), .ZN(
        n15552) );
  AOI21_X1 U17648 ( .B1(n15568), .B2(n18086), .A(n15552), .ZN(n15553) );
  OAI21_X1 U17649 ( .B1(n15570), .B2(n18065), .A(n15553), .ZN(P2_U3011) );
  AOI21_X1 U17650 ( .B1(n15556), .B2(n15555), .A(n15554), .ZN(n20401) );
  AOI21_X1 U17651 ( .B1(n19527), .B2(n20401), .A(n15557), .ZN(n15558) );
  OAI21_X1 U17652 ( .B1(n15559), .B2(n19514), .A(n15558), .ZN(n15567) );
  INV_X1 U17653 ( .A(n15565), .ZN(n15560) );
  NAND2_X1 U17654 ( .A1(n19539), .A2(n15560), .ZN(n15563) );
  INV_X1 U17655 ( .A(n15561), .ZN(n19538) );
  NAND2_X1 U17656 ( .A1(n17919), .A2(n19538), .ZN(n15562) );
  NAND2_X1 U17657 ( .A1(n15563), .A2(n15562), .ZN(n17924) );
  INV_X1 U17658 ( .A(n15564), .ZN(n19545) );
  NAND2_X1 U17659 ( .A1(n19539), .A2(n15565), .ZN(n19553) );
  NAND2_X1 U17660 ( .A1(n19513), .A2(n19553), .ZN(n17917) );
  AOI21_X1 U17661 ( .B1(n17919), .B2(n19545), .A(n17917), .ZN(n19555) );
  INV_X1 U17662 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19554) );
  NAND2_X1 U17663 ( .A1(n17919), .A2(n19554), .ZN(n19544) );
  NAND2_X1 U17664 ( .A1(n19555), .A2(n19544), .ZN(n15623) );
  MUX2_X1 U17665 ( .A(n17924), .B(n15623), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n15566) );
  AOI211_X1 U17666 ( .C1(n19537), .C2(n15568), .A(n15567), .B(n15566), .ZN(
        n15569) );
  OAI21_X1 U17667 ( .B1(n15570), .B2(n19546), .A(n15569), .ZN(P2_U3043) );
  XOR2_X1 U17668 ( .A(n15572), .B(n15571), .Z(n15578) );
  INV_X1 U17669 ( .A(n15573), .ZN(n15574) );
  NOR2_X1 U17670 ( .A1(n15574), .A2(n22162), .ZN(n15646) );
  AOI22_X1 U17671 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15645), .B1(
        n15646), .B2(n15786), .ZN(n15575) );
  NAND2_X1 U17672 ( .A1(n22202), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n15580) );
  OAI211_X1 U17673 ( .C1(n22214), .C2(n22281), .A(n15575), .B(n15580), .ZN(
        n15576) );
  AOI21_X1 U17674 ( .B1(n15578), .B2(n22200), .A(n15576), .ZN(n15577) );
  INV_X1 U17675 ( .A(n15577), .ZN(P1_U3025) );
  INV_X1 U17676 ( .A(n15578), .ZN(n15583) );
  NAND2_X1 U17677 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15579) );
  OAI211_X1 U17678 ( .C1(n20877), .C2(n22290), .A(n15580), .B(n15579), .ZN(
        n15581) );
  AOI21_X1 U17679 ( .B1(n22287), .B2(n20873), .A(n15581), .ZN(n15582) );
  OAI21_X1 U17680 ( .B1(n15583), .B2(n22385), .A(n15582), .ZN(P1_U2993) );
  NAND2_X1 U17681 ( .A1(n15537), .A2(n15585), .ZN(n15586) );
  AND2_X1 U17682 ( .A1(n15584), .A2(n15586), .ZN(n22298) );
  INV_X1 U17683 ( .A(n22298), .ZN(n15597) );
  OAI222_X1 U17684 ( .A1(n15597), .A2(n16837), .B1(n16836), .B2(n15587), .C1(
        n16834), .C2(n13357), .ZN(P1_U2897) );
  OAI21_X1 U17685 ( .B1(n15255), .B2(n15589), .A(n15588), .ZN(n15736) );
  NOR2_X1 U17686 ( .A1(n15680), .A2(n15736), .ZN(n15592) );
  AOI211_X1 U17687 ( .C1(n15590), .C2(n15253), .A(n17316), .B(n15385), .ZN(
        n15591) );
  AOI211_X1 U17688 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n15680), .A(n15592), .B(
        n15591), .ZN(n15593) );
  INV_X1 U17689 ( .A(n15593), .ZN(P2_U2877) );
  NOR2_X1 U17690 ( .A1(n15595), .A2(n15594), .ZN(n15596) );
  OR2_X1 U17691 ( .A1(n15650), .A2(n15596), .ZN(n22293) );
  INV_X1 U17692 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n22292) );
  OAI222_X1 U17693 ( .A1(n22293), .A2(n20828), .B1(n22292), .B2(n20833), .C1(
        n15597), .C2(n20812), .ZN(P1_U2865) );
  OAI21_X1 U17694 ( .B1(n15600), .B2(n15599), .A(n15598), .ZN(n20446) );
  INV_X1 U17695 ( .A(n20446), .ZN(n19543) );
  NOR2_X1 U17696 ( .A1(n18106), .A2(n20496), .ZN(n15606) );
  AOI21_X1 U17697 ( .B1(n18106), .B2(n20496), .A(n15606), .ZN(n20498) );
  INV_X1 U17698 ( .A(n20498), .ZN(n15604) );
  OR2_X1 U17699 ( .A1(n15602), .A2(n15601), .ZN(n15603) );
  NAND2_X1 U17700 ( .A1(n12250), .A2(n15603), .ZN(n20547) );
  NOR2_X1 U17701 ( .A1(n18098), .A2(n20547), .ZN(n20550) );
  NOR2_X1 U17702 ( .A1(n15604), .A2(n20550), .ZN(n15605) );
  NOR2_X1 U17703 ( .A1(n15606), .A2(n15605), .ZN(n15607) );
  XNOR2_X1 U17704 ( .A(n19543), .B(n15607), .ZN(n20448) );
  INV_X1 U17705 ( .A(n20448), .ZN(n15609) );
  NAND2_X1 U17706 ( .A1(n15607), .A2(n20446), .ZN(n15608) );
  OAI21_X1 U17707 ( .B1(n15609), .B2(n20447), .A(n15608), .ZN(n20403) );
  XOR2_X1 U17708 ( .A(n20401), .B(n20132), .Z(n20404) );
  NOR2_X1 U17709 ( .A1(n20403), .A2(n20404), .ZN(n20402) );
  INV_X1 U17710 ( .A(n20132), .ZN(n20221) );
  NOR2_X1 U17711 ( .A1(n20221), .A2(n20401), .ZN(n15612) );
  OAI21_X1 U17712 ( .B1(n15554), .B2(n15611), .A(n15610), .ZN(n15613) );
  OAI21_X1 U17713 ( .B1(n20402), .B2(n15612), .A(n15613), .ZN(n20317) );
  XOR2_X1 U17714 ( .A(n20315), .B(n20317), .Z(n15617) );
  INV_X1 U17715 ( .A(n15613), .ZN(n15753) );
  INV_X1 U17716 ( .A(n17404), .ZN(n17344) );
  INV_X1 U17717 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n18137) );
  OAI22_X1 U17718 ( .A1(n20557), .A2(n20361), .B1(n20546), .B2(n18137), .ZN(
        n15615) );
  AOI21_X1 U17719 ( .B1(n15753), .B2(n20497), .A(n15615), .ZN(n15616) );
  OAI21_X1 U17720 ( .B1(n15617), .B2(n20405), .A(n15616), .ZN(P2_U2915) );
  XNOR2_X1 U17721 ( .A(n15618), .B(n15619), .ZN(n18066) );
  INV_X1 U17722 ( .A(n17924), .ZN(n15620) );
  NOR2_X1 U17723 ( .A1(n15620), .A2(n15624), .ZN(n15833) );
  AND2_X1 U17724 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19526), .ZN(n15621) );
  AOI21_X1 U17725 ( .B1(n15834), .B2(n15833), .A(n15621), .ZN(n15622) );
  OAI21_X1 U17726 ( .B1(n18062), .B2(n19514), .A(n15622), .ZN(n15626) );
  AOI21_X1 U17727 ( .B1(n15624), .B2(n17834), .A(n15623), .ZN(n15838) );
  NOR2_X1 U17728 ( .A1(n15838), .A2(n15834), .ZN(n15625) );
  AOI211_X1 U17729 ( .C1(n19527), .C2(n15753), .A(n15626), .B(n15625), .ZN(
        n15631) );
  OR2_X1 U17730 ( .A1(n15627), .A2(n15834), .ZN(n15628) );
  AND2_X1 U17731 ( .A1(n15629), .A2(n15628), .ZN(n18064) );
  OR2_X1 U17732 ( .A1(n18064), .A2(n17944), .ZN(n15630) );
  OAI211_X1 U17733 ( .C1(n18066), .C2(n19546), .A(n15631), .B(n15630), .ZN(
        P2_U3042) );
  INV_X1 U17734 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n15642) );
  OAI211_X1 U17735 ( .C1(n15633), .C2(n15636), .A(n15635), .B(n17303), .ZN(
        n15641) );
  INV_X1 U17736 ( .A(n15846), .ZN(n15637) );
  OAI21_X1 U17737 ( .B1(n15677), .B2(n15638), .A(n15637), .ZN(n17851) );
  INV_X1 U17738 ( .A(n17851), .ZN(n15639) );
  NAND2_X1 U17739 ( .A1(n15639), .A2(n17309), .ZN(n15640) );
  OAI211_X1 U17740 ( .C1(n17309), .C2(n15642), .A(n15641), .B(n15640), .ZN(
        P2_U2874) );
  XNOR2_X1 U17741 ( .A(n15644), .B(n15643), .ZN(n15761) );
  INV_X1 U17742 ( .A(n15645), .ZN(n15787) );
  OAI21_X1 U17743 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17103), .A(
        n15787), .ZN(n15674) );
  NAND2_X1 U17744 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15646), .ZN(
        n15789) );
  AOI21_X1 U17745 ( .B1(n15648), .B2(n15647), .A(n15789), .ZN(n15649) );
  NAND2_X1 U17746 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15790) );
  AOI22_X1 U17747 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15674), .B1(
        n15649), .B2(n15790), .ZN(n15655) );
  INV_X1 U17748 ( .A(n15650), .ZN(n15652) );
  INV_X1 U17749 ( .A(n15690), .ZN(n15651) );
  AOI21_X1 U17750 ( .B1(n15653), .B2(n15652), .A(n15651), .ZN(n22302) );
  NOR2_X1 U17751 ( .A1(n22129), .A2(n20749), .ZN(n15757) );
  AOI21_X1 U17752 ( .B1(n22199), .B2(n22302), .A(n15757), .ZN(n15654) );
  OAI211_X1 U17753 ( .C1(n15761), .C2(n22218), .A(n15655), .B(n15654), .ZN(
        P1_U3023) );
  OAI21_X1 U17754 ( .B1(n15658), .B2(n15657), .A(n15656), .ZN(n20312) );
  NOR2_X1 U17755 ( .A1(n19396), .A2(n15659), .ZN(n15660) );
  XNOR2_X1 U17756 ( .A(n15660), .B(n15827), .ZN(n15661) );
  NAND2_X1 U17757 ( .A1(n15661), .A2(n19484), .ZN(n15669) );
  INV_X1 U17758 ( .A(n15839), .ZN(n15667) );
  OAI21_X1 U17759 ( .B1(n12115), .B2(n19464), .A(n19301), .ZN(n15663) );
  INV_X1 U17760 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15828) );
  NOR2_X1 U17761 ( .A1(n19462), .A2(n15828), .ZN(n15662) );
  AOI211_X1 U17762 ( .C1(n19494), .C2(P2_REIP_REG_5__SCAN_IN), .A(n15663), .B(
        n15662), .ZN(n15664) );
  OAI21_X1 U17763 ( .B1(n15665), .B2(n19393), .A(n15664), .ZN(n15666) );
  AOI21_X1 U17764 ( .B1(n15667), .B2(n19498), .A(n15666), .ZN(n15668) );
  OAI211_X1 U17765 ( .C1(n20312), .C2(n19477), .A(n15669), .B(n15668), .ZN(
        P2_U2850) );
  XOR2_X1 U17766 ( .A(n15671), .B(n15670), .Z(n20839) );
  NAND2_X1 U17767 ( .A1(n20839), .A2(n22200), .ZN(n15676) );
  NAND2_X1 U17768 ( .A1(n22202), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n20840) );
  INV_X1 U17769 ( .A(n20840), .ZN(n15673) );
  NOR2_X1 U17770 ( .A1(n22214), .A2(n22293), .ZN(n15672) );
  AOI211_X1 U17771 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n15674), .A(
        n15673), .B(n15672), .ZN(n15675) );
  OAI211_X1 U17772 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n15789), .A(
        n15676), .B(n15675), .ZN(P1_U3024) );
  AOI21_X1 U17773 ( .B1(n15679), .B2(n15678), .A(n15677), .ZN(n19321) );
  INV_X1 U17774 ( .A(n19321), .ZN(n15681) );
  NOR2_X1 U17775 ( .A1(n15681), .A2(n15680), .ZN(n15685) );
  AOI211_X1 U17776 ( .C1(n15683), .C2(n15682), .A(n17316), .B(n15633), .ZN(
        n15684) );
  AOI211_X1 U17777 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n15680), .A(n15685), .B(
        n15684), .ZN(n15686) );
  INV_X1 U17778 ( .A(n15686), .ZN(P2_U2875) );
  NOR2_X1 U17779 ( .A1(n11326), .A2(n15687), .ZN(n15688) );
  OR2_X1 U17780 ( .A1(n11321), .A2(n15688), .ZN(n16687) );
  NAND2_X1 U17781 ( .A1(n15690), .A2(n15689), .ZN(n15691) );
  NAND2_X1 U17782 ( .A1(n15856), .A2(n15691), .ZN(n16677) );
  OAI222_X1 U17783 ( .A1(n16687), .A2(n20812), .B1(n16682), .B2(n20833), .C1(
        n16677), .C2(n20828), .ZN(P1_U2863) );
  OR2_X1 U17784 ( .A1(n16757), .A2(n20904), .ZN(n15693) );
  NAND2_X1 U17785 ( .A1(n16757), .A2(DATAI_9_), .ZN(n15692) );
  AND2_X1 U17786 ( .A1(n15693), .A2(n15692), .ZN(n22485) );
  INV_X1 U17787 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15694) );
  OAI222_X1 U17788 ( .A1(n16687), .A2(n16837), .B1(n22485), .B2(n16836), .C1(
        n15694), .C2(n16834), .ZN(P1_U2895) );
  NOR2_X1 U17789 ( .A1(n19396), .A2(n19563), .ZN(n19501) );
  INV_X1 U17790 ( .A(n17229), .ZN(n15817) );
  NAND2_X1 U17791 ( .A1(n19484), .A2(n19396), .ZN(n19311) );
  INV_X1 U17792 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15695) );
  AOI21_X1 U17793 ( .B1(n19462), .B2(n19311), .A(n15695), .ZN(n15696) );
  AOI21_X1 U17794 ( .B1(n19501), .B2(n15817), .A(n15696), .ZN(n15702) );
  OAI22_X1 U17795 ( .A1(n19393), .A2(n15697), .B1(n12545), .B2(n19464), .ZN(
        n15699) );
  OAI22_X1 U17796 ( .A1(n19477), .A2(n20547), .B1(n19386), .B2(n18010), .ZN(
        n15698) );
  AOI211_X1 U17797 ( .C1(n15700), .C2(n19498), .A(n15699), .B(n15698), .ZN(
        n15701) );
  OAI211_X1 U17798 ( .C1(n17240), .C2(n18098), .A(n15702), .B(n15701), .ZN(
        P2_U2855) );
  NAND2_X1 U17799 ( .A1(n11252), .A2(n15703), .ZN(n15704) );
  XNOR2_X1 U17800 ( .A(n15705), .B(n15704), .ZN(n15706) );
  NAND2_X1 U17801 ( .A1(n15706), .A2(n19484), .ZN(n15715) );
  OAI22_X1 U17802 ( .A1(n12089), .A2(n19464), .B1(n15707), .B2(n19386), .ZN(
        n15710) );
  NOR2_X1 U17803 ( .A1(n19462), .A2(n15708), .ZN(n15709) );
  AOI211_X1 U17804 ( .C1(n19492), .C2(n15711), .A(n15710), .B(n15709), .ZN(
        n15712) );
  OAI21_X1 U17805 ( .B1(n19543), .B2(n19477), .A(n15712), .ZN(n15713) );
  AOI21_X1 U17806 ( .B1(n19551), .B2(n19498), .A(n15713), .ZN(n15714) );
  OAI211_X1 U17807 ( .C1(n20447), .C2(n17240), .A(n15715), .B(n15714), .ZN(
        P2_U2853) );
  OAI21_X1 U17808 ( .B1(n15718), .B2(n15717), .A(n15716), .ZN(n19525) );
  NAND2_X1 U17809 ( .A1(n11252), .A2(n15719), .ZN(n15720) );
  XNOR2_X1 U17810 ( .A(n18072), .B(n15720), .ZN(n15721) );
  NAND2_X1 U17811 ( .A1(n15721), .A2(n19484), .ZN(n15731) );
  INV_X1 U17812 ( .A(n15722), .ZN(n15729) );
  INV_X1 U17813 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n15727) );
  NAND2_X1 U17814 ( .A1(n19498), .A2(n19531), .ZN(n15726) );
  OAI21_X1 U17815 ( .B1(n15723), .B2(n19464), .A(n19301), .ZN(n15724) );
  AOI21_X1 U17816 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19495), .A(
        n15724), .ZN(n15725) );
  OAI211_X1 U17817 ( .C1(n15727), .C2(n19386), .A(n15726), .B(n15725), .ZN(
        n15728) );
  AOI21_X1 U17818 ( .B1(n15729), .B2(n19492), .A(n15728), .ZN(n15730) );
  OAI211_X1 U17819 ( .C1(n19477), .C2(n19525), .A(n15731), .B(n15730), .ZN(
        P2_U2849) );
  XOR2_X1 U17820 ( .A(n15732), .B(n17221), .Z(n20069) );
  INV_X1 U17821 ( .A(n20069), .ZN(n15744) );
  NAND2_X1 U17822 ( .A1(n11252), .A2(n15733), .ZN(n15734) );
  XNOR2_X1 U17823 ( .A(n18082), .B(n15734), .ZN(n15735) );
  NAND2_X1 U17824 ( .A1(n15735), .A2(n19484), .ZN(n15743) );
  INV_X1 U17825 ( .A(n15736), .ZN(n18087) );
  INV_X1 U17826 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n15738) );
  AOI22_X1 U17827 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19495), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19494), .ZN(n15737) );
  OAI211_X1 U17828 ( .C1(n19464), .C2(n15738), .A(n15737), .B(n19301), .ZN(
        n15741) );
  NOR2_X1 U17829 ( .A1(n15739), .A2(n19393), .ZN(n15740) );
  AOI211_X1 U17830 ( .C1(n18087), .C2(n19498), .A(n15741), .B(n15740), .ZN(
        n15742) );
  OAI211_X1 U17831 ( .C1(n15744), .C2(n19477), .A(n15743), .B(n15742), .ZN(
        P2_U2845) );
  AND2_X1 U17832 ( .A1(n11252), .A2(n15745), .ZN(n15747) );
  AOI21_X1 U17833 ( .B1(n18061), .B2(n15747), .A(n19563), .ZN(n15746) );
  OAI21_X1 U17834 ( .B1(n18061), .B2(n15747), .A(n15746), .ZN(n15755) );
  AOI22_X1 U17835 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19491), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19494), .ZN(n15748) );
  OAI211_X1 U17836 ( .C1(n19462), .C2(n18071), .A(n19301), .B(n15748), .ZN(
        n15749) );
  AOI21_X1 U17837 ( .B1(n19492), .B2(n15750), .A(n15749), .ZN(n15751) );
  OAI21_X1 U17838 ( .B1(n18062), .B2(n19467), .A(n15751), .ZN(n15752) );
  AOI21_X1 U17839 ( .B1(n15753), .B2(n12449), .A(n15752), .ZN(n15754) );
  OAI211_X1 U17840 ( .C1(n17240), .C2(n20315), .A(n15755), .B(n15754), .ZN(
        P2_U2851) );
  XOR2_X1 U17841 ( .A(n15756), .B(n15584), .Z(n22305) );
  AOI21_X1 U17842 ( .B1(n20870), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15757), .ZN(n15758) );
  OAI21_X1 U17843 ( .B1(n20877), .B2(n22303), .A(n15758), .ZN(n15759) );
  AOI21_X1 U17844 ( .B1(n22305), .B2(n20873), .A(n15759), .ZN(n15760) );
  OAI21_X1 U17845 ( .B1(n15761), .B2(n22385), .A(n15760), .ZN(P1_U2991) );
  NAND2_X1 U17846 ( .A1(n20114), .A2(n20203), .ZN(n20412) );
  NOR2_X1 U17847 ( .A1(n20663), .A2(n20668), .ZN(n15762) );
  OAI21_X1 U17848 ( .B1(n15762), .B2(n22410), .A(n20222), .ZN(n15774) );
  INV_X1 U17849 ( .A(n15763), .ZN(n20561) );
  NAND2_X1 U17850 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n17995), .ZN(n19271) );
  NAND2_X1 U17851 ( .A1(n15765), .A2(n19271), .ZN(n19574) );
  INV_X1 U17852 ( .A(n12585), .ZN(n15770) );
  NAND2_X1 U17853 ( .A1(n15767), .A2(n20162), .ZN(n20209) );
  NOR2_X1 U17854 ( .A1(n15770), .A2(n20209), .ZN(n15768) );
  OAI22_X1 U17855 ( .A1(n15774), .A2(n20561), .B1(n20184), .B2(n15768), .ZN(
        n15769) );
  NOR2_X1 U17856 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20246) );
  NAND2_X1 U17857 ( .A1(n20205), .A2(n20246), .ZN(n15779) );
  OAI21_X1 U17858 ( .B1(n15770), .B2(n20235), .A(n15779), .ZN(n15771) );
  NOR2_X1 U17859 ( .A1(n15771), .A2(n20561), .ZN(n15773) );
  INV_X1 U17860 ( .A(n15771), .ZN(n15772) );
  OAI22_X1 U17861 ( .A1(n15774), .A2(n15773), .B1(n15772), .B2(n20235), .ZN(
        n20666) );
  INV_X1 U17862 ( .A(n20668), .ZN(n15781) );
  INV_X1 U17863 ( .A(n20454), .ZN(n20560) );
  INV_X1 U17864 ( .A(n15779), .ZN(n20662) );
  AOI22_X1 U17865 ( .A1(n20442), .A2(n20663), .B1(n20441), .B2(n20662), .ZN(
        n15780) );
  OAI21_X1 U17866 ( .B1(n15781), .B2(n20445), .A(n15780), .ZN(n15782) );
  AOI21_X1 U17867 ( .B1(n20666), .B2(n15775), .A(n15782), .ZN(n15783) );
  OAI21_X1 U17868 ( .B1(n20672), .B2(n15784), .A(n15783), .ZN(P2_U3051) );
  NOR2_X1 U17869 ( .A1(n15786), .A2(n15790), .ZN(n16968) );
  OAI21_X1 U17870 ( .B1(n17103), .B2(n16968), .A(n15787), .ZN(n17147) );
  INV_X1 U17871 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20751) );
  OAI22_X1 U17872 ( .A1(n22214), .A2(n16677), .B1(n20751), .B2(n22129), .ZN(
        n15788) );
  AOI21_X1 U17873 ( .B1(n17147), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15788), .ZN(n15792) );
  NOR2_X1 U17874 ( .A1(n15790), .A2(n15789), .ZN(n17146) );
  NAND2_X1 U17875 ( .A1(n17146), .A2(n17144), .ZN(n15791) );
  OAI211_X1 U17876 ( .C1(n15880), .C2(n22218), .A(n15792), .B(n15791), .ZN(
        P1_U3022) );
  INV_X1 U17877 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n15796) );
  INV_X1 U17878 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20902) );
  INV_X1 U17879 ( .A(DATAI_8_), .ZN(n16153) );
  AOI22_X1 U17880 ( .A1(n15793), .A2(n20902), .B1(n16153), .B2(n16757), .ZN(
        n15794) );
  INV_X1 U17881 ( .A(n15794), .ZN(n22479) );
  INV_X1 U17882 ( .A(n22305), .ZN(n15795) );
  OAI222_X1 U17883 ( .A1(n16834), .A2(n15796), .B1(n22479), .B2(n16836), .C1(
        n16837), .C2(n15795), .ZN(P1_U2896) );
  OAI211_X1 U17884 ( .C1(n15797), .C2(n15798), .A(n11279), .B(n17303), .ZN(
        n15803) );
  AOI21_X1 U17885 ( .B1(n15801), .B2(n15799), .A(n15800), .ZN(n19343) );
  NAND2_X1 U17886 ( .A1(n19343), .A2(n17309), .ZN(n15802) );
  OAI211_X1 U17887 ( .C1(n17309), .C2(n12147), .A(n15803), .B(n15802), .ZN(
        P2_U2872) );
  AOI21_X1 U17888 ( .B1(n15806), .B2(n15804), .A(n15805), .ZN(n20059) );
  INV_X1 U17889 ( .A(n20059), .ZN(n17855) );
  OAI22_X1 U17890 ( .A1(n17851), .A2(n19467), .B1(n19462), .B2(n15807), .ZN(
        n15808) );
  AOI21_X1 U17891 ( .B1(n15809), .B2(n19492), .A(n15808), .ZN(n15813) );
  NAND2_X1 U17892 ( .A1(n11253), .A2(n19325), .ZN(n15810) );
  NOR2_X1 U17893 ( .A1(n19563), .A2(n15810), .ZN(n19333) );
  OAI21_X1 U17894 ( .B1(n15811), .B2(n17588), .A(n19333), .ZN(n15812) );
  OAI211_X1 U17895 ( .C1(n17855), .C2(n19477), .A(n15813), .B(n15812), .ZN(
        n15816) );
  AOI22_X1 U17896 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19491), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19494), .ZN(n15814) );
  OAI211_X1 U17897 ( .C1(n17588), .C2(n19311), .A(n15814), .B(n19301), .ZN(
        n15815) );
  OR2_X1 U17898 ( .A1(n15816), .A2(n15815), .ZN(P2_U2842) );
  NAND2_X1 U17899 ( .A1(n17948), .A2(n20162), .ZN(n19557) );
  INV_X1 U17900 ( .A(n19557), .ZN(n17955) );
  INV_X1 U17901 ( .A(n17961), .ZN(n19572) );
  AOI22_X1 U17902 ( .A1(n19396), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n15817), .B2(n11253), .ZN(n17949) );
  AOI222_X1 U17903 ( .A1(n15818), .A2(n17955), .B1(n19572), .B2(n20554), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n17949), .ZN(n15823) );
  NAND2_X1 U17904 ( .A1(n15819), .A2(n19570), .ZN(n15821) );
  AOI22_X1 U17905 ( .A1(n17995), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19567), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n15820) );
  NAND2_X1 U17906 ( .A1(n15821), .A2(n15820), .ZN(n19510) );
  INV_X1 U17907 ( .A(n19510), .ZN(n19507) );
  NAND2_X1 U17908 ( .A1(n19507), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15822) );
  OAI21_X1 U17909 ( .B1(n15823), .B2(n19507), .A(n15822), .ZN(P2_U3601) );
  XNOR2_X1 U17910 ( .A(n15824), .B(n15837), .ZN(n15844) );
  XOR2_X1 U17911 ( .A(n15826), .B(n15825), .Z(n15842) );
  OAI22_X1 U17912 ( .A1(n15828), .A2(n18093), .B1(n17638), .B2(n15827), .ZN(
        n15829) );
  AOI21_X1 U17913 ( .B1(P2_REIP_REG_5__SCAN_IN), .B2(n19526), .A(n15829), .ZN(
        n15830) );
  OAI21_X1 U17914 ( .B1(n17641), .B2(n15839), .A(n15830), .ZN(n15831) );
  AOI21_X1 U17915 ( .B1(n15842), .B2(n18089), .A(n15831), .ZN(n15832) );
  OAI21_X1 U17916 ( .B1(n18063), .B2(n15844), .A(n15832), .ZN(P2_U3009) );
  OAI221_X1 U17917 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15834), .C2(n15837), .A(
        n15833), .ZN(n15836) );
  NAND2_X1 U17918 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19526), .ZN(n15835) );
  OAI211_X1 U17919 ( .C1(n15838), .C2(n15837), .A(n15836), .B(n15835), .ZN(
        n15841) );
  OAI22_X1 U17920 ( .A1(n20312), .A2(n19542), .B1(n19514), .B2(n15839), .ZN(
        n15840) );
  AOI211_X1 U17921 ( .C1(n15842), .C2(n19530), .A(n15841), .B(n15840), .ZN(
        n15843) );
  OAI21_X1 U17922 ( .B1(n17944), .B2(n15844), .A(n15843), .ZN(P2_U3041) );
  OR2_X1 U17923 ( .A1(n15846), .A2(n15845), .ZN(n15847) );
  AND2_X1 U17924 ( .A1(n15799), .A2(n15847), .ZN(n19331) );
  INV_X1 U17925 ( .A(n19331), .ZN(n15848) );
  NOR2_X1 U17926 ( .A1(n15848), .A2(n15680), .ZN(n15851) );
  AOI211_X1 U17927 ( .C1(n15849), .C2(n15635), .A(n17316), .B(n15797), .ZN(
        n15850) );
  AOI211_X1 U17928 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n15680), .A(n15851), .B(
        n15850), .ZN(n15852) );
  INV_X1 U17929 ( .A(n15852), .ZN(P2_U2873) );
  XOR2_X1 U17930 ( .A(n15853), .B(n11321), .Z(n20844) );
  INV_X1 U17931 ( .A(n20844), .ZN(n15899) );
  OAI21_X1 U17932 ( .B1(n22312), .B2(n22323), .A(n22255), .ZN(n22330) );
  OAI21_X1 U17933 ( .B1(n22323), .B2(n15854), .A(n20753), .ZN(n15864) );
  NAND2_X1 U17934 ( .A1(n15856), .A2(n15855), .ZN(n15857) );
  NAND2_X1 U17935 ( .A1(n17115), .A2(n15857), .ZN(n20816) );
  INV_X1 U17936 ( .A(n15858), .ZN(n20843) );
  NAND2_X1 U17937 ( .A1(n22255), .A2(n15859), .ZN(n22354) );
  OAI21_X1 U17938 ( .B1(n22337), .B2(n13401), .A(n22354), .ZN(n15861) );
  NOR2_X1 U17939 ( .A1(n22374), .A2(n20819), .ZN(n15860) );
  AOI211_X1 U17940 ( .C1(n22353), .C2(n20843), .A(n15861), .B(n15860), .ZN(
        n15862) );
  OAI21_X1 U17941 ( .B1(n22375), .B2(n20816), .A(n15862), .ZN(n15863) );
  AOI21_X1 U17942 ( .B1(n22330), .B2(n15864), .A(n15863), .ZN(n15865) );
  OAI21_X1 U17943 ( .B1(n15899), .B2(n22377), .A(n15865), .ZN(P1_U2830) );
  AOI21_X1 U17944 ( .B1(n15867), .B2(n11279), .A(n15866), .ZN(n15884) );
  AND2_X1 U17945 ( .A1(n17816), .A2(n15868), .ZN(n15869) );
  OR2_X1 U17946 ( .A1(n15869), .A2(n11325), .ZN(n19358) );
  OAI22_X1 U17947 ( .A1(n17404), .A2(n20559), .B1(n15870), .B2(n20546), .ZN(
        n15871) );
  AOI21_X1 U17948 ( .B1(n20048), .B2(BUF2_REG_16__SCAN_IN), .A(n15871), .ZN(
        n15873) );
  NAND2_X1 U17949 ( .A1(n20050), .A2(BUF1_REG_16__SCAN_IN), .ZN(n15872) );
  OAI211_X1 U17950 ( .C1(n19358), .C2(n20548), .A(n15873), .B(n15872), .ZN(
        n15874) );
  AOI21_X1 U17951 ( .B1(n15884), .B2(n20551), .A(n15874), .ZN(n15875) );
  INV_X1 U17952 ( .A(n15875), .ZN(P2_U2903) );
  INV_X1 U17953 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15876) );
  OAI22_X1 U17954 ( .A1(n20842), .A2(n15876), .B1(n22129), .B2(n20751), .ZN(
        n15878) );
  NOR2_X1 U17955 ( .A1(n16687), .A2(n20853), .ZN(n15877) );
  AOI211_X1 U17956 ( .C1(n20862), .C2(n16680), .A(n15878), .B(n15877), .ZN(
        n15879) );
  OAI21_X1 U17957 ( .B1(n22385), .B2(n15880), .A(n15879), .ZN(P1_U2990) );
  NAND2_X1 U17958 ( .A1(n15882), .A2(n15881), .ZN(n15883) );
  NAND2_X1 U17959 ( .A1(n15903), .A2(n15883), .ZN(n17804) );
  NAND2_X1 U17960 ( .A1(n15884), .A2(n17303), .ZN(n15886) );
  NAND2_X1 U17961 ( .A1(n15680), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15885) );
  OAI211_X1 U17962 ( .C1(n17804), .C2(n15680), .A(n15886), .B(n15885), .ZN(
        P2_U2871) );
  OAI21_X1 U17963 ( .B1(n15866), .B2(n15888), .A(n15887), .ZN(n15907) );
  NOR2_X1 U17964 ( .A1(n11325), .A2(n15889), .ZN(n15890) );
  OR2_X1 U17965 ( .A1(n15921), .A2(n15890), .ZN(n17793) );
  OAI22_X1 U17966 ( .A1(n17404), .A2(n20502), .B1(n20546), .B2(n15891), .ZN(
        n15892) );
  AOI21_X1 U17967 ( .B1(n20048), .B2(BUF2_REG_17__SCAN_IN), .A(n15892), .ZN(
        n15894) );
  NAND2_X1 U17968 ( .A1(n20050), .A2(BUF1_REG_17__SCAN_IN), .ZN(n15893) );
  OAI211_X1 U17969 ( .C1(n17793), .C2(n20548), .A(n15894), .B(n15893), .ZN(
        n15895) );
  INV_X1 U17970 ( .A(n15895), .ZN(n15896) );
  OAI21_X1 U17971 ( .B1(n15907), .B2(n20405), .A(n15896), .ZN(P2_U2902) );
  INV_X1 U17972 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15900) );
  OR2_X1 U17973 ( .A1(n16757), .A2(n20906), .ZN(n15898) );
  NAND2_X1 U17974 ( .A1(n16757), .A2(DATAI_10_), .ZN(n15897) );
  AND2_X1 U17975 ( .A1(n15898), .A2(n15897), .ZN(n22492) );
  OAI222_X1 U17976 ( .A1(n16834), .A2(n15900), .B1(n22492), .B2(n16836), .C1(
        n16837), .C2(n15899), .ZN(P1_U2894) );
  AND2_X1 U17977 ( .A1(n15903), .A2(n15902), .ZN(n15904) );
  NOR2_X1 U17978 ( .A1(n15901), .A2(n15904), .ZN(n17790) );
  INV_X1 U17979 ( .A(n17790), .ZN(n17208) );
  NOR2_X1 U17980 ( .A1(n17208), .A2(n15680), .ZN(n15905) );
  AOI21_X1 U17981 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15680), .A(n15905), .ZN(
        n15906) );
  OAI21_X1 U17982 ( .B1(n15907), .B2(n17316), .A(n15906), .ZN(P2_U2870) );
  OR2_X1 U17983 ( .A1(n15909), .A2(n15908), .ZN(n15911) );
  INV_X1 U17984 ( .A(n16660), .ZN(n15912) );
  XNOR2_X1 U17985 ( .A(n16661), .B(n15912), .ZN(n22318) );
  INV_X1 U17986 ( .A(n22318), .ZN(n20852) );
  INV_X1 U17987 ( .A(n16836), .ZN(n15915) );
  OR2_X1 U17988 ( .A1(n16757), .A2(n20908), .ZN(n15914) );
  NAND2_X1 U17989 ( .A1(n16757), .A2(DATAI_11_), .ZN(n15913) );
  NAND2_X1 U17990 ( .A1(n15914), .A2(n15913), .ZN(n22499) );
  INV_X1 U17991 ( .A(n16834), .ZN(n16819) );
  AOI22_X1 U17992 ( .A1(n15915), .A2(n22499), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n16819), .ZN(n15916) );
  OAI21_X1 U17993 ( .B1(n20852), .B2(n16837), .A(n15916), .ZN(P1_U2893) );
  XNOR2_X1 U17994 ( .A(n17115), .B(n17117), .ZN(n22313) );
  AOI22_X1 U17995 ( .A1(n22313), .A2(n20825), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n16714), .ZN(n15917) );
  OAI21_X1 U17996 ( .B1(n20852), .B2(n20812), .A(n15917), .ZN(P1_U2861) );
  AOI21_X1 U17997 ( .B1(n15919), .B2(n15887), .A(n15918), .ZN(n15929) );
  OR2_X1 U17998 ( .A1(n15921), .A2(n15920), .ZN(n15922) );
  NAND2_X1 U17999 ( .A1(n17400), .A2(n15922), .ZN(n19373) );
  OAI22_X1 U18000 ( .A1(n17404), .A2(n20452), .B1(n15923), .B2(n20546), .ZN(
        n15924) );
  AOI21_X1 U18001 ( .B1(n20048), .B2(BUF2_REG_18__SCAN_IN), .A(n15924), .ZN(
        n15926) );
  NAND2_X1 U18002 ( .A1(n20050), .A2(BUF1_REG_18__SCAN_IN), .ZN(n15925) );
  OAI211_X1 U18003 ( .C1(n19373), .C2(n20548), .A(n15926), .B(n15925), .ZN(
        n15927) );
  AOI21_X1 U18004 ( .B1(n15929), .B2(n20551), .A(n15927), .ZN(n15928) );
  INV_X1 U18005 ( .A(n15928), .ZN(P2_U2901) );
  INV_X1 U18006 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15934) );
  NAND2_X1 U18007 ( .A1(n15929), .A2(n17303), .ZN(n15933) );
  OR2_X1 U18008 ( .A1(n15901), .A2(n15930), .ZN(n15931) );
  AND2_X1 U18009 ( .A1(n15931), .A2(n17312), .ZN(n19367) );
  NAND2_X1 U18010 ( .A1(n19367), .A2(n17309), .ZN(n15932) );
  OAI211_X1 U18011 ( .C1(n17309), .C2(n15934), .A(n15933), .B(n15932), .ZN(
        P2_U2869) );
  AOI21_X1 U18012 ( .B1(n15938), .B2(n15936), .A(n11700), .ZN(n16953) );
  NOR2_X1 U18013 ( .A1(n22323), .A2(n16668), .ZN(n15939) );
  AOI21_X1 U18014 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n22339), .A(n15939), 
        .ZN(n15948) );
  NAND2_X1 U18015 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15939), .ZN(n16625) );
  INV_X1 U18016 ( .A(n16625), .ZN(n22338) );
  NAND2_X1 U18017 ( .A1(n22371), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15942) );
  INV_X1 U18018 ( .A(n16951), .ZN(n15940) );
  NAND2_X1 U18019 ( .A1(n22353), .A2(n15940), .ZN(n15941) );
  NAND3_X1 U18020 ( .A1(n15942), .A2(n15941), .A3(n22354), .ZN(n15943) );
  AOI21_X1 U18021 ( .B1(n22358), .B2(P1_EBX_REG_14__SCAN_IN), .A(n15943), .ZN(
        n15947) );
  NAND2_X1 U18022 ( .A1(n16666), .A2(n15944), .ZN(n15945) );
  AND2_X1 U18023 ( .A1(n16735), .A2(n15945), .ZN(n22132) );
  NAND2_X1 U18024 ( .A1(n22327), .A2(n22132), .ZN(n15946) );
  OAI211_X1 U18025 ( .C1(n15948), .C2(n22338), .A(n15947), .B(n15946), .ZN(
        n15949) );
  AOI21_X1 U18026 ( .B1(n16953), .B2(n22362), .A(n15949), .ZN(n15950) );
  INV_X1 U18027 ( .A(n15950), .ZN(P1_U2826) );
  INV_X1 U18028 ( .A(n16953), .ZN(n15955) );
  AOI22_X1 U18029 ( .A1(n22132), .A2(n20825), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n16714), .ZN(n15951) );
  OAI21_X1 U18030 ( .B1(n15955), .B2(n20812), .A(n15951), .ZN(P1_U2858) );
  INV_X1 U18031 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20914) );
  OR2_X1 U18032 ( .A1(n16757), .A2(n20914), .ZN(n15953) );
  NAND2_X1 U18033 ( .A1(n16757), .A2(DATAI_14_), .ZN(n15952) );
  AND2_X1 U18034 ( .A1(n15953), .A2(n15952), .ZN(n22519) );
  INV_X1 U18035 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15954) );
  OAI222_X1 U18036 ( .A1(n15955), .A2(n16837), .B1(n22519), .B2(n16836), .C1(
        n15954), .C2(n16834), .ZN(P1_U2890) );
  INV_X1 U18037 ( .A(n15956), .ZN(n15962) );
  NAND2_X1 U18038 ( .A1(n15967), .A2(n17753), .ZN(n15958) );
  NAND4_X1 U18039 ( .A1(n15958), .A2(n15957), .A3(n17550), .A4(n17534), .ZN(
        n15960) );
  NOR2_X1 U18040 ( .A1(n15960), .A2(n15959), .ZN(n15961) );
  NOR2_X1 U18041 ( .A1(n15965), .A2(n15964), .ZN(n15966) );
  OAI211_X1 U18042 ( .C1(n15967), .C2(n17753), .A(n15966), .B(n17527), .ZN(
        n15969) );
  NAND2_X1 U18043 ( .A1(n15975), .A2(n15974), .ZN(n15976) );
  AND2_X1 U18044 ( .A1(n15979), .A2(n15976), .ZN(n19409) );
  NAND2_X1 U18045 ( .A1(n19409), .A2(n16014), .ZN(n15977) );
  INV_X1 U18046 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17731) );
  NOR2_X1 U18047 ( .A1(n15977), .A2(n17731), .ZN(n17494) );
  XNOR2_X1 U18048 ( .A(n15979), .B(n15978), .ZN(n19416) );
  NAND2_X1 U18049 ( .A1(n19416), .A2(n16014), .ZN(n15980) );
  INV_X1 U18050 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17722) );
  AND2_X1 U18051 ( .A1(n15980), .A2(n17722), .ZN(n17485) );
  INV_X1 U18052 ( .A(n15980), .ZN(n15981) );
  XNOR2_X1 U18053 ( .A(n15983), .B(n15982), .ZN(n19427) );
  NAND2_X1 U18054 ( .A1(n19427), .A2(n16014), .ZN(n15984) );
  NOR2_X1 U18055 ( .A1(n15984), .A2(n17707), .ZN(n17474) );
  NAND2_X1 U18056 ( .A1(n19449), .A2(n16014), .ZN(n15987) );
  XOR2_X1 U18057 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15987), .Z(
        n17453) );
  INV_X1 U18058 ( .A(n15988), .ZN(n15989) );
  XNOR2_X1 U18059 ( .A(n15990), .B(n15989), .ZN(n19436) );
  AOI21_X1 U18060 ( .B1(n19436), .B2(n16014), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17466) );
  NOR2_X2 U18061 ( .A1(n17453), .A2(n17466), .ZN(n15991) );
  INV_X1 U18062 ( .A(n15992), .ZN(n15993) );
  NAND2_X1 U18063 ( .A1(n11313), .A2(n15993), .ZN(n15994) );
  NAND2_X1 U18064 ( .A1(n15997), .A2(n15994), .ZN(n17181) );
  NOR2_X1 U18065 ( .A1(n17181), .A2(n16007), .ZN(n16052) );
  XNOR2_X1 U18066 ( .A(n15997), .B(n15996), .ZN(n19470) );
  NAND2_X1 U18067 ( .A1(n19470), .A2(n16014), .ZN(n16002) );
  NOR2_X1 U18068 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16001) );
  NAND3_X1 U18069 ( .A1(n19449), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n16014), .ZN(n16000) );
  NOR2_X1 U18070 ( .A1(n16007), .A2(n17700), .ZN(n15999) );
  NAND2_X1 U18071 ( .A1(n19436), .A2(n15999), .ZN(n17464) );
  AND2_X1 U18072 ( .A1(n16000), .A2(n17464), .ZN(n16049) );
  OAI21_X1 U18073 ( .B1(n16002), .B2(n16001), .A(n16049), .ZN(n16003) );
  INV_X1 U18074 ( .A(n16003), .ZN(n16004) );
  XNOR2_X1 U18075 ( .A(n16006), .B(n16005), .ZN(n16010) );
  OAI21_X1 U18076 ( .B1(n16010), .B2(n16007), .A(n17659), .ZN(n17431) );
  AOI21_X1 U18077 ( .B1(n16009), .B2(n16014), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17422) );
  INV_X1 U18078 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17645) );
  NOR2_X1 U18079 ( .A1(n16007), .A2(n17645), .ZN(n16008) );
  NAND2_X1 U18080 ( .A1(n16009), .A2(n16008), .ZN(n17420) );
  INV_X1 U18081 ( .A(n16010), .ZN(n19478) );
  NAND3_X1 U18082 ( .A1(n19478), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16014), .ZN(n17432) );
  NOR2_X1 U18083 ( .A1(n16011), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16012) );
  MUX2_X1 U18084 ( .A(n16013), .B(n16012), .S(n20322), .Z(n19493) );
  NAND2_X1 U18085 ( .A1(n19493), .A2(n16014), .ZN(n16015) );
  XNOR2_X1 U18086 ( .A(n16015), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16016) );
  XNOR2_X1 U18087 ( .A(n16017), .B(n16016), .ZN(n17418) );
  AND2_X1 U18088 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16031) );
  INV_X1 U18089 ( .A(n16057), .ZN(n17459) );
  NAND2_X1 U18090 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17646) );
  INV_X1 U18091 ( .A(n17646), .ZN(n17657) );
  AND2_X1 U18092 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16018) );
  NAND2_X1 U18093 ( .A1(n17657), .A2(n16018), .ZN(n16034) );
  INV_X1 U18094 ( .A(n17425), .ZN(n16019) );
  NAND2_X1 U18095 ( .A1(n17425), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16020) );
  AOI22_X1 U18096 ( .A1(n12196), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n16022) );
  OAI21_X1 U18097 ( .B1(n16023), .B2(n17243), .A(n16022), .ZN(n16024) );
  AOI21_X1 U18098 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n16024), .ZN(n16026) );
  INV_X1 U18099 ( .A(n16034), .ZN(n16028) );
  OAI211_X1 U18100 ( .C1(n16031), .C2(n19521), .A(n17732), .B(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17709) );
  INV_X1 U18101 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17689) );
  NOR2_X1 U18102 ( .A1(n17689), .A2(n17700), .ZN(n16033) );
  INV_X1 U18103 ( .A(n16033), .ZN(n17686) );
  OAI21_X1 U18104 ( .B1(n17709), .B2(n17686), .A(n17685), .ZN(n17676) );
  OAI21_X1 U18105 ( .B1(n19521), .B2(n16028), .A(n17676), .ZN(n17648) );
  INV_X1 U18106 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n16029) );
  NOR2_X1 U18107 ( .A1(n19301), .A2(n16029), .ZN(n17413) );
  OR2_X1 U18108 ( .A1(n17794), .A2(n16030), .ZN(n17719) );
  NAND2_X1 U18109 ( .A1(n16031), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16032) );
  NOR2_X1 U18110 ( .A1(n17719), .A2(n16032), .ZN(n17701) );
  NAND2_X1 U18111 ( .A1(n17701), .A2(n16033), .ZN(n17658) );
  NOR3_X1 U18112 ( .A1(n17658), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16034), .ZN(n16035) );
  AOI211_X1 U18113 ( .C1(n17648), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n17413), .B(n16035), .ZN(n16036) );
  OAI21_X1 U18114 ( .B1(n17241), .B2(n19514), .A(n16036), .ZN(n16037) );
  AOI222_X1 U18115 ( .A1(n16041), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n16040), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12262), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16042) );
  INV_X1 U18116 ( .A(n16042), .ZN(n16043) );
  XNOR2_X1 U18117 ( .A(n16044), .B(n16043), .ZN(n19496) );
  NAND2_X1 U18118 ( .A1(n16046), .A2(n16045), .ZN(n16047) );
  OAI21_X1 U18119 ( .B1(n17418), .B2(n19546), .A(n16048), .ZN(P2_U3015) );
  NAND2_X1 U18120 ( .A1(n16054), .A2(n16053), .ZN(n16056) );
  XNOR2_X1 U18121 ( .A(n16056), .B(n16055), .ZN(n16073) );
  XNOR2_X2 U18122 ( .A(n17184), .B(n16058), .ZN(n19468) );
  NOR2_X1 U18123 ( .A1(n19468), .A2(n17641), .ZN(n16061) );
  NAND2_X1 U18124 ( .A1(n19526), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16066) );
  NAND2_X1 U18125 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16059) );
  OAI211_X1 U18126 ( .C1(n17638), .C2(n19473), .A(n16066), .B(n16059), .ZN(
        n16060) );
  AOI211_X1 U18127 ( .C1(n16071), .C2(n18086), .A(n16061), .B(n16060), .ZN(
        n16062) );
  OAI21_X1 U18128 ( .B1(n16073), .B2(n18065), .A(n16062), .ZN(P2_U2986) );
  XNOR2_X1 U18129 ( .A(n16063), .B(n16064), .ZN(n19476) );
  INV_X1 U18130 ( .A(n17658), .ZN(n16065) );
  NAND2_X1 U18131 ( .A1(n16065), .A2(n15995), .ZN(n17675) );
  NAND2_X1 U18132 ( .A1(n17676), .A2(n17675), .ZN(n17664) );
  OR2_X1 U18133 ( .A1(n17658), .A2(n15995), .ZN(n17661) );
  OAI21_X1 U18134 ( .B1(n17661), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16066), .ZN(n16068) );
  NOR2_X1 U18135 ( .A1(n19468), .A2(n19514), .ZN(n16067) );
  AOI211_X1 U18136 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n17664), .A(
        n16068), .B(n16067), .ZN(n16069) );
  OAI21_X1 U18137 ( .B1(n19476), .B2(n19542), .A(n16069), .ZN(n16070) );
  OAI21_X1 U18138 ( .B1(n16073), .B2(n19546), .A(n16072), .ZN(P2_U3018) );
  OAI22_X1 U18139 ( .A1(n17404), .A2(n20056), .B1(n20546), .B2(n16074), .ZN(
        n16075) );
  AOI21_X1 U18140 ( .B1(n20048), .B2(BUF2_REG_30__SCAN_IN), .A(n16075), .ZN(
        n16077) );
  NAND2_X1 U18141 ( .A1(n20050), .A2(BUF1_REG_30__SCAN_IN), .ZN(n16076) );
  OAI211_X1 U18142 ( .C1(n17652), .C2(n20548), .A(n16077), .B(n16076), .ZN(
        n16078) );
  AOI21_X1 U18143 ( .B1(n16079), .B2(n20551), .A(n16078), .ZN(n16080) );
  INV_X1 U18144 ( .A(n16080), .ZN(P2_U2889) );
  NOR2_X1 U18145 ( .A1(n19396), .A2(n16081), .ZN(n16083) );
  XNOR2_X1 U18146 ( .A(n16083), .B(n16082), .ZN(n16084) );
  NAND2_X1 U18147 ( .A1(n16084), .A2(n19484), .ZN(n16093) );
  NAND2_X1 U18148 ( .A1(n12449), .A2(n20401), .ZN(n16089) );
  OAI22_X1 U18149 ( .A1(n16086), .A2(n19464), .B1(n16085), .B2(n19386), .ZN(
        n16087) );
  AOI21_X1 U18150 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19495), .A(
        n16087), .ZN(n16088) );
  OAI211_X1 U18151 ( .C1(n19393), .C2(n16090), .A(n16089), .B(n16088), .ZN(
        n16091) );
  AOI21_X1 U18152 ( .B1(n11260), .B2(n19498), .A(n16091), .ZN(n16092) );
  OAI211_X1 U18153 ( .C1(n20132), .C2(n17240), .A(n16093), .B(n16092), .ZN(
        P2_U2852) );
  INV_X1 U18154 ( .A(n16106), .ZN(n16094) );
  OAI21_X1 U18155 ( .B1(n16094), .B2(n22402), .A(P1_MEMORYFETCH_REG_SCAN_IN), 
        .ZN(n16095) );
  NAND3_X1 U18156 ( .A1(n16096), .A2(n20881), .A3(n16095), .ZN(P1_U2801) );
  INV_X1 U18157 ( .A(n16097), .ZN(n16099) );
  NOR2_X1 U18158 ( .A1(n16099), .A2(n16098), .ZN(n16100) );
  AOI21_X1 U18159 ( .B1(n16108), .B2(n14191), .A(n16100), .ZN(n16104) );
  INV_X1 U18160 ( .A(n16101), .ZN(n16102) );
  NAND2_X1 U18161 ( .A1(n16108), .A2(n16102), .ZN(n16103) );
  OAI211_X1 U18162 ( .C1(n16105), .C2(n16108), .A(n16104), .B(n16103), .ZN(
        n18032) );
  NOR2_X1 U18163 ( .A1(n16106), .A2(n14191), .ZN(n16107) );
  AOI21_X1 U18164 ( .B1(n16108), .B2(n16688), .A(n16107), .ZN(n20878) );
  OR2_X1 U18165 ( .A1(n16109), .A2(n18044), .ZN(n16110) );
  NAND2_X1 U18166 ( .A1(n16110), .A2(n22424), .ZN(n22107) );
  AND2_X1 U18167 ( .A1(n20878), .A2(n22107), .ZN(n18030) );
  NOR2_X1 U18168 ( .A1(n18030), .A2(n22402), .ZN(n22387) );
  MUX2_X1 U18169 ( .A(P1_MORE_REG_SCAN_IN), .B(n18032), .S(n22387), .Z(
        P1_U3484) );
  INV_X1 U18170 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20799) );
  AOI21_X1 U18171 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n16111) );
  INV_X1 U18172 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n22247) );
  AOI22_X1 U18173 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n16111), .B2(n22247), .ZN(n16122) );
  NOR4_X1 U18174 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16115) );
  AOI211_X1 U18175 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16114) );
  NOR4_X1 U18176 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16113) );
  NOR4_X1 U18177 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16112) );
  NAND4_X1 U18178 ( .A1(n16115), .A2(n16114), .A3(n16113), .A4(n16112), .ZN(
        n16121) );
  NOR4_X1 U18179 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16119) );
  NOR4_X1 U18180 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16118) );
  NOR4_X1 U18181 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16117) );
  NOR4_X1 U18182 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16116) );
  NAND4_X1 U18183 ( .A1(n16119), .A2(n16118), .A3(n16117), .A4(n16116), .ZN(
        n16120) );
  NOR2_X1 U18184 ( .A1(n16121), .A2(n16120), .ZN(n20804) );
  MUX2_X1 U18185 ( .A(n20799), .B(n16122), .S(n20804), .Z(n16493) );
  XNOR2_X1 U18186 ( .A(DATAI_31_), .B(keyinput_1), .ZN(n16126) );
  XNOR2_X1 U18187 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_0), .ZN(n16125) );
  XNOR2_X1 U18188 ( .A(DATAI_28_), .B(keyinput_4), .ZN(n16124) );
  XNOR2_X1 U18189 ( .A(DATAI_30_), .B(keyinput_2), .ZN(n16123) );
  OAI211_X1 U18190 ( .C1(n16126), .C2(n16125), .A(n16124), .B(n16123), .ZN(
        n16129) );
  XOR2_X1 U18191 ( .A(DATAI_27_), .B(keyinput_5), .Z(n16128) );
  XNOR2_X1 U18192 ( .A(DATAI_29_), .B(keyinput_3), .ZN(n16127) );
  NOR3_X1 U18193 ( .A1(n16129), .A2(n16128), .A3(n16127), .ZN(n16133) );
  XNOR2_X1 U18194 ( .A(DATAI_26_), .B(keyinput_6), .ZN(n16132) );
  XNOR2_X1 U18195 ( .A(DATAI_24_), .B(keyinput_8), .ZN(n16131) );
  XNOR2_X1 U18196 ( .A(DATAI_25_), .B(keyinput_7), .ZN(n16130) );
  OAI211_X1 U18197 ( .C1(n16133), .C2(n16132), .A(n16131), .B(n16130), .ZN(
        n16137) );
  XNOR2_X1 U18198 ( .A(DATAI_23_), .B(keyinput_9), .ZN(n16136) );
  XOR2_X1 U18199 ( .A(DATAI_22_), .B(keyinput_10), .Z(n16135) );
  XNOR2_X1 U18200 ( .A(DATAI_21_), .B(keyinput_11), .ZN(n16134) );
  AOI211_X1 U18201 ( .C1(n16137), .C2(n16136), .A(n16135), .B(n16134), .ZN(
        n16143) );
  XOR2_X1 U18202 ( .A(DATAI_20_), .B(keyinput_12), .Z(n16142) );
  XOR2_X1 U18203 ( .A(DATAI_19_), .B(keyinput_13), .Z(n16140) );
  XOR2_X1 U18204 ( .A(DATAI_17_), .B(keyinput_15), .Z(n16139) );
  XNOR2_X1 U18205 ( .A(DATAI_18_), .B(keyinput_14), .ZN(n16138) );
  NOR3_X1 U18206 ( .A1(n16140), .A2(n16139), .A3(n16138), .ZN(n16141) );
  OAI21_X1 U18207 ( .B1(n16143), .B2(n16142), .A(n16141), .ZN(n16149) );
  XNOR2_X1 U18208 ( .A(DATAI_16_), .B(keyinput_16), .ZN(n16148) );
  XOR2_X1 U18209 ( .A(DATAI_13_), .B(keyinput_19), .Z(n16146) );
  XOR2_X1 U18210 ( .A(DATAI_14_), .B(keyinput_18), .Z(n16145) );
  XNOR2_X1 U18211 ( .A(DATAI_15_), .B(keyinput_17), .ZN(n16144) );
  NAND3_X1 U18212 ( .A1(n16146), .A2(n16145), .A3(n16144), .ZN(n16147) );
  AOI21_X1 U18213 ( .B1(n16149), .B2(n16148), .A(n16147), .ZN(n16152) );
  XOR2_X1 U18214 ( .A(DATAI_11_), .B(keyinput_21), .Z(n16151) );
  XNOR2_X1 U18215 ( .A(DATAI_12_), .B(keyinput_20), .ZN(n16150) );
  NOR3_X1 U18216 ( .A1(n16152), .A2(n16151), .A3(n16150), .ZN(n16157) );
  XOR2_X1 U18217 ( .A(DATAI_10_), .B(keyinput_22), .Z(n16156) );
  XNOR2_X1 U18218 ( .A(n16153), .B(keyinput_24), .ZN(n16155) );
  XNOR2_X1 U18219 ( .A(DATAI_9_), .B(keyinput_23), .ZN(n16154) );
  NOR4_X1 U18220 ( .A1(n16157), .A2(n16156), .A3(n16155), .A4(n16154), .ZN(
        n16160) );
  XNOR2_X1 U18221 ( .A(DATAI_7_), .B(keyinput_25), .ZN(n16159) );
  XNOR2_X1 U18222 ( .A(DATAI_6_), .B(keyinput_26), .ZN(n16158) );
  OAI21_X1 U18223 ( .B1(n16160), .B2(n16159), .A(n16158), .ZN(n16163) );
  XNOR2_X1 U18224 ( .A(n16339), .B(keyinput_27), .ZN(n16162) );
  XOR2_X1 U18225 ( .A(DATAI_4_), .B(keyinput_28), .Z(n16161) );
  NAND3_X1 U18226 ( .A1(n16163), .A2(n16162), .A3(n16161), .ZN(n16166) );
  XNOR2_X1 U18227 ( .A(DATAI_3_), .B(keyinput_29), .ZN(n16165) );
  XNOR2_X1 U18228 ( .A(DATAI_2_), .B(keyinput_30), .ZN(n16164) );
  AOI21_X1 U18229 ( .B1(n16166), .B2(n16165), .A(n16164), .ZN(n16169) );
  XNOR2_X1 U18230 ( .A(n16348), .B(keyinput_31), .ZN(n16168) );
  XNOR2_X1 U18231 ( .A(DATAI_0_), .B(keyinput_32), .ZN(n16167) );
  NOR3_X1 U18232 ( .A1(n16169), .A2(n16168), .A3(n16167), .ZN(n16179) );
  XNOR2_X1 U18233 ( .A(READY2), .B(keyinput_37), .ZN(n16171) );
  XNOR2_X1 U18234 ( .A(READY1), .B(keyinput_36), .ZN(n16170) );
  NOR2_X1 U18235 ( .A1(n16171), .A2(n16170), .ZN(n16176) );
  INV_X1 U18236 ( .A(keyinput_35), .ZN(n16172) );
  XNOR2_X1 U18237 ( .A(n16172), .B(BS16), .ZN(n16175) );
  XNOR2_X1 U18238 ( .A(HOLD), .B(keyinput_33), .ZN(n16174) );
  XNOR2_X1 U18239 ( .A(NA), .B(keyinput_34), .ZN(n16173) );
  NAND4_X1 U18240 ( .A1(n16176), .A2(n16175), .A3(n16174), .A4(n16173), .ZN(
        n16178) );
  XNOR2_X1 U18241 ( .A(P1_READREQUEST_REG_SCAN_IN), .B(keyinput_38), .ZN(
        n16177) );
  OAI21_X1 U18242 ( .B1(n16179), .B2(n16178), .A(n16177), .ZN(n16183) );
  INV_X1 U18243 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n18058) );
  XNOR2_X1 U18244 ( .A(n18058), .B(keyinput_39), .ZN(n16182) );
  XOR2_X1 U18245 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_40), .Z(n16181)
         );
  XNOR2_X1 U18246 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_41), .ZN(n16180) );
  AOI211_X1 U18247 ( .C1(n16183), .C2(n16182), .A(n16181), .B(n16180), .ZN(
        n16186) );
  XNOR2_X1 U18248 ( .A(P1_D_C_N_REG_SCAN_IN), .B(keyinput_42), .ZN(n16185) );
  XNOR2_X1 U18249 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_43), .ZN(
        n16184) );
  NOR3_X1 U18250 ( .A1(n16186), .A2(n16185), .A3(n16184), .ZN(n16189) );
  XNOR2_X1 U18251 ( .A(n22405), .B(keyinput_44), .ZN(n16188) );
  XNOR2_X1 U18252 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_45), .ZN(n16187) );
  OAI21_X1 U18253 ( .B1(n16189), .B2(n16188), .A(n16187), .ZN(n16195) );
  XOR2_X1 U18254 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_46), .Z(n16194) );
  XOR2_X1 U18255 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_48), .Z(
        n16192) );
  XOR2_X1 U18256 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_49), .Z(
        n16191) );
  XNOR2_X1 U18257 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_47), .ZN(n16190) );
  NAND3_X1 U18258 ( .A1(n16192), .A2(n16191), .A3(n16190), .ZN(n16193) );
  AOI21_X1 U18259 ( .B1(n16195), .B2(n16194), .A(n16193), .ZN(n16199) );
  XOR2_X1 U18260 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_52), .Z(n16198) );
  XOR2_X1 U18261 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_51), .Z(
        n16197) );
  XNOR2_X1 U18262 ( .A(n20799), .B(keyinput_50), .ZN(n16196) );
  NOR4_X1 U18263 ( .A1(n16199), .A2(n16198), .A3(n16197), .A4(n16196), .ZN(
        n16203) );
  XNOR2_X1 U18264 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_53), .ZN(n16202)
         );
  XNOR2_X1 U18265 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_55), .ZN(n16201)
         );
  XNOR2_X1 U18266 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_54), .ZN(n16200)
         );
  OAI211_X1 U18267 ( .C1(n16203), .C2(n16202), .A(n16201), .B(n16200), .ZN(
        n16206) );
  XOR2_X1 U18268 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_56), .Z(n16205) );
  XNOR2_X1 U18269 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_57), .ZN(n16204)
         );
  NAND3_X1 U18270 ( .A1(n16206), .A2(n16205), .A3(n16204), .ZN(n16219) );
  AOI22_X1 U18271 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_65), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_58), .ZN(n16207) );
  OAI221_X1 U18272 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_65), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_58), .A(n16207), .ZN(n16216) );
  INV_X1 U18273 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U18274 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_61), .B1(n20778), .B2(keyinput_59), .ZN(n16208) );
  OAI221_X1 U18275 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_61), .C1(
        n20778), .C2(keyinput_59), .A(n16208), .ZN(n16212) );
  XOR2_X1 U18276 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_63), .Z(n16211) );
  XNOR2_X1 U18277 ( .A(n20777), .B(keyinput_60), .ZN(n16210) );
  XNOR2_X1 U18278 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_62), .ZN(n16209)
         );
  OR4_X1 U18279 ( .A1(n16212), .A2(n16211), .A3(n16210), .A4(n16209), .ZN(
        n16215) );
  XNOR2_X1 U18280 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_64), .ZN(n16214)
         );
  XNOR2_X1 U18281 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_66), .ZN(n16213)
         );
  NOR4_X1 U18282 ( .A1(n16216), .A2(n16215), .A3(n16214), .A4(n16213), .ZN(
        n16218) );
  XOR2_X1 U18283 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_67), .Z(n16217) );
  AOI21_X1 U18284 ( .B1(n16219), .B2(n16218), .A(n16217), .ZN(n16223) );
  XNOR2_X1 U18285 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_68), .ZN(n16222)
         );
  XNOR2_X1 U18286 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n16221)
         );
  XNOR2_X1 U18287 ( .A(P1_REIP_REG_13__SCAN_IN), .B(keyinput_70), .ZN(n16220)
         );
  OAI211_X1 U18288 ( .C1(n16223), .C2(n16222), .A(n16221), .B(n16220), .ZN(
        n16227) );
  XNOR2_X1 U18289 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_71), .ZN(n16226)
         );
  XNOR2_X1 U18290 ( .A(P1_REIP_REG_11__SCAN_IN), .B(keyinput_72), .ZN(n16225)
         );
  XNOR2_X1 U18291 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_73), .ZN(n16224)
         );
  AOI211_X1 U18292 ( .C1(n16227), .C2(n16226), .A(n16225), .B(n16224), .ZN(
        n16233) );
  XOR2_X1 U18293 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_74), .Z(n16229) );
  XNOR2_X1 U18294 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_75), .ZN(n16228)
         );
  NAND2_X1 U18295 ( .A1(n16229), .A2(n16228), .ZN(n16232) );
  XOR2_X1 U18296 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_76), .Z(n16231) );
  XNOR2_X1 U18297 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_77), .ZN(n16230)
         );
  OAI211_X1 U18298 ( .C1(n16233), .C2(n16232), .A(n16231), .B(n16230), .ZN(
        n16236) );
  XOR2_X1 U18299 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_79), .Z(n16235) );
  XNOR2_X1 U18300 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_78), .ZN(n16234)
         );
  NAND3_X1 U18301 ( .A1(n16236), .A2(n16235), .A3(n16234), .ZN(n16244) );
  XOR2_X1 U18302 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_80), .Z(n16243) );
  XOR2_X1 U18303 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_82), .Z(n16242) );
  XOR2_X1 U18304 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_81), .Z(n16240) );
  XOR2_X1 U18305 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_84), .Z(n16239) );
  INV_X1 U18306 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n16707) );
  XNOR2_X1 U18307 ( .A(n16707), .B(keyinput_85), .ZN(n16238) );
  XNOR2_X1 U18308 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_83), .ZN(n16237)
         );
  NOR4_X1 U18309 ( .A1(n16240), .A2(n16239), .A3(n16238), .A4(n16237), .ZN(
        n16241) );
  NAND4_X1 U18310 ( .A1(n16244), .A2(n16243), .A3(n16242), .A4(n16241), .ZN(
        n16251) );
  XNOR2_X1 U18311 ( .A(n16427), .B(keyinput_88), .ZN(n16250) );
  XOR2_X1 U18312 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_90), .Z(n16249) );
  XNOR2_X1 U18313 ( .A(n16708), .B(keyinput_86), .ZN(n16247) );
  XNOR2_X1 U18314 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_87), .ZN(n16246)
         );
  XNOR2_X1 U18315 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_89), .ZN(n16245)
         );
  NOR3_X1 U18316 ( .A1(n16247), .A2(n16246), .A3(n16245), .ZN(n16248) );
  NAND4_X1 U18317 ( .A1(n16251), .A2(n16250), .A3(n16249), .A4(n16248), .ZN(
        n16254) );
  XNOR2_X1 U18318 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_91), .ZN(n16253)
         );
  XNOR2_X1 U18319 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_92), .ZN(n16252)
         );
  AOI21_X1 U18320 ( .B1(n16254), .B2(n16253), .A(n16252), .ZN(n16260) );
  INV_X1 U18321 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16728) );
  INV_X1 U18322 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n22373) );
  AOI22_X1 U18323 ( .A1(n16728), .A2(keyinput_96), .B1(keyinput_94), .B2(
        n22373), .ZN(n16255) );
  OAI221_X1 U18324 ( .B1(n16728), .B2(keyinput_96), .C1(n22373), .C2(
        keyinput_94), .A(n16255), .ZN(n16259) );
  INV_X1 U18325 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16717) );
  AOI22_X1 U18326 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(keyinput_97), .B1(n16717), 
        .B2(keyinput_93), .ZN(n16256) );
  OAI221_X1 U18327 ( .B1(P1_EBX_REG_18__SCAN_IN), .B2(keyinput_97), .C1(n16717), .C2(keyinput_93), .A(n16256), .ZN(n16258) );
  XNOR2_X1 U18328 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_95), .ZN(n16257)
         );
  NOR4_X1 U18329 ( .A1(n16260), .A2(n16259), .A3(n16258), .A4(n16257), .ZN(
        n16262) );
  XNOR2_X1 U18330 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_98), .ZN(n16261)
         );
  NOR2_X1 U18331 ( .A1(n16262), .A2(n16261), .ZN(n16266) );
  XNOR2_X1 U18332 ( .A(n16738), .B(keyinput_100), .ZN(n16265) );
  XNOR2_X1 U18333 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n16264)
         );
  XNOR2_X1 U18334 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_99), .ZN(n16263)
         );
  NOR4_X1 U18335 ( .A1(n16266), .A2(n16265), .A3(n16264), .A4(n16263), .ZN(
        n16270) );
  XNOR2_X1 U18336 ( .A(n16739), .B(keyinput_102), .ZN(n16269) );
  XNOR2_X1 U18337 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_104), .ZN(n16268)
         );
  XNOR2_X1 U18338 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_103), .ZN(n16267)
         );
  OAI211_X1 U18339 ( .C1(n16270), .C2(n16269), .A(n16268), .B(n16267), .ZN(
        n16273) );
  XOR2_X1 U18340 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_105), .Z(n16272) );
  XNOR2_X1 U18341 ( .A(n16682), .B(keyinput_106), .ZN(n16271) );
  AOI21_X1 U18342 ( .B1(n16273), .B2(n16272), .A(n16271), .ZN(n16276) );
  XNOR2_X1 U18343 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_107), .ZN(n16275)
         );
  XNOR2_X1 U18344 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_108), .ZN(n16274)
         );
  OAI21_X1 U18345 ( .B1(n16276), .B2(n16275), .A(n16274), .ZN(n16280) );
  XOR2_X1 U18346 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_109), .Z(n16279) );
  XOR2_X1 U18347 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_110), .Z(n16278) );
  XNOR2_X1 U18348 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n16277)
         );
  AOI211_X1 U18349 ( .C1(n16280), .C2(n16279), .A(n16278), .B(n16277), .ZN(
        n16284) );
  XNOR2_X1 U18350 ( .A(n22228), .B(keyinput_113), .ZN(n16283) );
  XOR2_X1 U18351 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_112), .Z(n16282) );
  XNOR2_X1 U18352 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_114), .ZN(n16281)
         );
  NOR4_X1 U18353 ( .A1(n16284), .A2(n16283), .A3(n16282), .A4(n16281), .ZN(
        n16287) );
  XNOR2_X1 U18354 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_115), .ZN(n16286)
         );
  XOR2_X1 U18355 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_116), .Z(n16285) );
  OAI21_X1 U18356 ( .B1(n16287), .B2(n16286), .A(n16285), .ZN(n16291) );
  XOR2_X1 U18357 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_117), .Z(n16290) );
  XOR2_X1 U18358 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_118), .Z(n16289) );
  XNOR2_X1 U18359 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_119), .ZN(n16288)
         );
  NAND4_X1 U18360 ( .A1(n16291), .A2(n16290), .A3(n16289), .A4(n16288), .ZN(
        n16294) );
  XOR2_X1 U18361 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_120), .Z(n16293) );
  XOR2_X1 U18362 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_121), .Z(n16292) );
  NAND3_X1 U18363 ( .A1(n16294), .A2(n16293), .A3(n16292), .ZN(n16297) );
  XOR2_X1 U18364 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_122), .Z(n16296) );
  XOR2_X1 U18365 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_123), .Z(n16295) );
  AOI21_X1 U18366 ( .B1(n16297), .B2(n16296), .A(n16295), .ZN(n16300) );
  XOR2_X1 U18367 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_124), .Z(n16299) );
  XNOR2_X1 U18368 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_125), .ZN(n16298)
         );
  OAI21_X1 U18369 ( .B1(n16300), .B2(n16299), .A(n16298), .ZN(n16491) );
  XOR2_X1 U18370 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_126), .Z(n16490) );
  XOR2_X1 U18371 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_127), .Z(n16489) );
  XOR2_X1 U18372 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_128), .Z(n16304) );
  XNOR2_X1 U18373 ( .A(n15058), .B(keyinput_129), .ZN(n16303) );
  XOR2_X1 U18374 ( .A(DATAI_27_), .B(keyinput_133), .Z(n16302) );
  XOR2_X1 U18375 ( .A(DATAI_29_), .B(keyinput_131), .Z(n16301) );
  AOI211_X1 U18376 ( .C1(n16304), .C2(n16303), .A(n16302), .B(n16301), .ZN(
        n16307) );
  XOR2_X1 U18377 ( .A(DATAI_30_), .B(keyinput_130), .Z(n16306) );
  XOR2_X1 U18378 ( .A(DATAI_28_), .B(keyinput_132), .Z(n16305) );
  NAND3_X1 U18379 ( .A1(n16307), .A2(n16306), .A3(n16305), .ZN(n16311) );
  XOR2_X1 U18380 ( .A(DATAI_26_), .B(keyinput_134), .Z(n16310) );
  XOR2_X1 U18381 ( .A(DATAI_24_), .B(keyinput_136), .Z(n16309) );
  XNOR2_X1 U18382 ( .A(DATAI_25_), .B(keyinput_135), .ZN(n16308) );
  AOI211_X1 U18383 ( .C1(n16311), .C2(n16310), .A(n16309), .B(n16308), .ZN(
        n16315) );
  XNOR2_X1 U18384 ( .A(DATAI_23_), .B(keyinput_137), .ZN(n16314) );
  XOR2_X1 U18385 ( .A(DATAI_22_), .B(keyinput_138), .Z(n16313) );
  XNOR2_X1 U18386 ( .A(DATAI_21_), .B(keyinput_139), .ZN(n16312) );
  OAI211_X1 U18387 ( .C1(n16315), .C2(n16314), .A(n16313), .B(n16312), .ZN(
        n16321) );
  XNOR2_X1 U18388 ( .A(DATAI_20_), .B(keyinput_140), .ZN(n16320) );
  XOR2_X1 U18389 ( .A(DATAI_19_), .B(keyinput_141), .Z(n16318) );
  XOR2_X1 U18390 ( .A(DATAI_17_), .B(keyinput_143), .Z(n16317) );
  XNOR2_X1 U18391 ( .A(DATAI_18_), .B(keyinput_142), .ZN(n16316) );
  NAND3_X1 U18392 ( .A1(n16318), .A2(n16317), .A3(n16316), .ZN(n16319) );
  AOI21_X1 U18393 ( .B1(n16321), .B2(n16320), .A(n16319), .ZN(n16327) );
  XNOR2_X1 U18394 ( .A(DATAI_16_), .B(keyinput_144), .ZN(n16326) );
  XOR2_X1 U18395 ( .A(DATAI_13_), .B(keyinput_147), .Z(n16324) );
  XOR2_X1 U18396 ( .A(DATAI_15_), .B(keyinput_145), .Z(n16323) );
  XOR2_X1 U18397 ( .A(DATAI_14_), .B(keyinput_146), .Z(n16322) );
  NOR3_X1 U18398 ( .A1(n16324), .A2(n16323), .A3(n16322), .ZN(n16325) );
  OAI21_X1 U18399 ( .B1(n16327), .B2(n16326), .A(n16325), .ZN(n16330) );
  XOR2_X1 U18400 ( .A(DATAI_11_), .B(keyinput_149), .Z(n16329) );
  XNOR2_X1 U18401 ( .A(DATAI_12_), .B(keyinput_148), .ZN(n16328) );
  NAND3_X1 U18402 ( .A1(n16330), .A2(n16329), .A3(n16328), .ZN(n16334) );
  XNOR2_X1 U18403 ( .A(DATAI_8_), .B(keyinput_152), .ZN(n16333) );
  XNOR2_X1 U18404 ( .A(DATAI_10_), .B(keyinput_150), .ZN(n16332) );
  XNOR2_X1 U18405 ( .A(DATAI_9_), .B(keyinput_151), .ZN(n16331) );
  NAND4_X1 U18406 ( .A1(n16334), .A2(n16333), .A3(n16332), .A4(n16331), .ZN(
        n16338) );
  XNOR2_X1 U18407 ( .A(DATAI_7_), .B(keyinput_153), .ZN(n16337) );
  XNOR2_X1 U18408 ( .A(n16335), .B(keyinput_154), .ZN(n16336) );
  AOI21_X1 U18409 ( .B1(n16338), .B2(n16337), .A(n16336), .ZN(n16342) );
  XNOR2_X1 U18410 ( .A(n16339), .B(keyinput_155), .ZN(n16341) );
  XNOR2_X1 U18411 ( .A(DATAI_4_), .B(keyinput_156), .ZN(n16340) );
  NOR3_X1 U18412 ( .A1(n16342), .A2(n16341), .A3(n16340), .ZN(n16347) );
  XNOR2_X1 U18413 ( .A(n16343), .B(keyinput_157), .ZN(n16346) );
  XNOR2_X1 U18414 ( .A(n16344), .B(keyinput_158), .ZN(n16345) );
  OAI21_X1 U18415 ( .B1(n16347), .B2(n16346), .A(n16345), .ZN(n16351) );
  XNOR2_X1 U18416 ( .A(n16348), .B(keyinput_159), .ZN(n16350) );
  XOR2_X1 U18417 ( .A(DATAI_0_), .B(keyinput_160), .Z(n16349) );
  NAND3_X1 U18418 ( .A1(n16351), .A2(n16350), .A3(n16349), .ZN(n16358) );
  XOR2_X1 U18419 ( .A(BS16), .B(keyinput_163), .Z(n16357) );
  XOR2_X1 U18420 ( .A(HOLD), .B(keyinput_161), .Z(n16354) );
  XOR2_X1 U18421 ( .A(READY2), .B(keyinput_165), .Z(n16353) );
  XNOR2_X1 U18422 ( .A(READY1), .B(keyinput_164), .ZN(n16352) );
  NOR3_X1 U18423 ( .A1(n16354), .A2(n16353), .A3(n16352), .ZN(n16356) );
  XNOR2_X1 U18424 ( .A(NA), .B(keyinput_162), .ZN(n16355) );
  NAND4_X1 U18425 ( .A1(n16358), .A2(n16357), .A3(n16356), .A4(n16355), .ZN(
        n16361) );
  XOR2_X1 U18426 ( .A(P1_READREQUEST_REG_SCAN_IN), .B(keyinput_166), .Z(n16360) );
  XNOR2_X1 U18427 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_167), .ZN(n16359) );
  AOI21_X1 U18428 ( .B1(n16361), .B2(n16360), .A(n16359), .ZN(n16364) );
  XOR2_X1 U18429 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_169), .Z(n16363) );
  XNOR2_X1 U18430 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_168), .ZN(n16362) );
  NOR3_X1 U18431 ( .A1(n16364), .A2(n16363), .A3(n16362), .ZN(n16367) );
  INV_X1 U18432 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22426) );
  XNOR2_X1 U18433 ( .A(n22426), .B(keyinput_171), .ZN(n16366) );
  XNOR2_X1 U18434 ( .A(P1_D_C_N_REG_SCAN_IN), .B(keyinput_170), .ZN(n16365) );
  NOR3_X1 U18435 ( .A1(n16367), .A2(n16366), .A3(n16365), .ZN(n16370) );
  XNOR2_X1 U18436 ( .A(P1_STATEBS16_REG_SCAN_IN), .B(keyinput_172), .ZN(n16369) );
  XNOR2_X1 U18437 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_173), .ZN(n16368) );
  OAI21_X1 U18438 ( .B1(n16370), .B2(n16369), .A(n16368), .ZN(n16376) );
  XNOR2_X1 U18439 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_174), .ZN(n16375) );
  XOR2_X1 U18440 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_175), .Z(n16373) );
  XOR2_X1 U18441 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_176), .Z(
        n16372) );
  XNOR2_X1 U18442 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_177), .ZN(
        n16371) );
  NAND3_X1 U18443 ( .A1(n16373), .A2(n16372), .A3(n16371), .ZN(n16374) );
  AOI21_X1 U18444 ( .B1(n16376), .B2(n16375), .A(n16374), .ZN(n16380) );
  XOR2_X1 U18445 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_180), .Z(n16379)
         );
  XNOR2_X1 U18446 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_179), .ZN(
        n16378) );
  XNOR2_X1 U18447 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_178), .ZN(
        n16377) );
  NOR4_X1 U18448 ( .A1(n16380), .A2(n16379), .A3(n16378), .A4(n16377), .ZN(
        n16384) );
  XNOR2_X1 U18449 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_181), .ZN(n16383)
         );
  XOR2_X1 U18450 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_183), .Z(n16382)
         );
  XOR2_X1 U18451 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_182), .Z(n16381)
         );
  OAI211_X1 U18452 ( .C1(n16384), .C2(n16383), .A(n16382), .B(n16381), .ZN(
        n16387) );
  XOR2_X1 U18453 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_184), .Z(n16386)
         );
  XOR2_X1 U18454 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_185), .Z(n16385)
         );
  NAND3_X1 U18455 ( .A1(n16387), .A2(n16386), .A3(n16385), .ZN(n16401) );
  OAI22_X1 U18456 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_193), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(keyinput_192), .ZN(n16389) );
  AND2_X1 U18457 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_193), .ZN(n16388) );
  AOI211_X1 U18458 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(keyinput_192), .A(
        n16389), .B(n16388), .ZN(n16393) );
  XOR2_X1 U18459 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_187), .Z(n16392)
         );
  XNOR2_X1 U18460 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_194), .ZN(n16391)
         );
  XNOR2_X1 U18461 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_190), .ZN(n16390)
         );
  NAND4_X1 U18462 ( .A1(n16393), .A2(n16392), .A3(n16391), .A4(n16390), .ZN(
        n16398) );
  INV_X1 U18463 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20774) );
  AOI22_X1 U18464 ( .A1(n20777), .A2(keyinput_188), .B1(n20774), .B2(
        keyinput_189), .ZN(n16394) );
  OAI221_X1 U18465 ( .B1(n20777), .B2(keyinput_188), .C1(n20774), .C2(
        keyinput_189), .A(n16394), .ZN(n16397) );
  XNOR2_X1 U18466 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_191), .ZN(n16396)
         );
  XNOR2_X1 U18467 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_186), .ZN(n16395)
         );
  NOR4_X1 U18468 ( .A1(n16398), .A2(n16397), .A3(n16396), .A4(n16395), .ZN(
        n16400) );
  XOR2_X1 U18469 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_195), .Z(n16399)
         );
  AOI21_X1 U18470 ( .B1(n16401), .B2(n16400), .A(n16399), .ZN(n16405) );
  XOR2_X1 U18471 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_196), .Z(n16404)
         );
  XOR2_X1 U18472 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_197), .Z(n16403)
         );
  XOR2_X1 U18473 ( .A(P1_REIP_REG_13__SCAN_IN), .B(keyinput_198), .Z(n16402)
         );
  OAI211_X1 U18474 ( .C1(n16405), .C2(n16404), .A(n16403), .B(n16402), .ZN(
        n16409) );
  XNOR2_X1 U18475 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_199), .ZN(n16408)
         );
  XOR2_X1 U18476 ( .A(P1_REIP_REG_11__SCAN_IN), .B(keyinput_200), .Z(n16407)
         );
  XNOR2_X1 U18477 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_201), .ZN(n16406)
         );
  AOI211_X1 U18478 ( .C1(n16409), .C2(n16408), .A(n16407), .B(n16406), .ZN(
        n16415) );
  XOR2_X1 U18479 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_202), .Z(n16411) );
  XNOR2_X1 U18480 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_203), .ZN(n16410)
         );
  NAND2_X1 U18481 ( .A1(n16411), .A2(n16410), .ZN(n16414) );
  XOR2_X1 U18482 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_204), .Z(n16413) );
  XOR2_X1 U18483 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_205), .Z(n16412) );
  OAI211_X1 U18484 ( .C1(n16415), .C2(n16414), .A(n16413), .B(n16412), .ZN(
        n16418) );
  XNOR2_X1 U18485 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_206), .ZN(n16417)
         );
  XNOR2_X1 U18486 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_207), .ZN(n16416)
         );
  NAND3_X1 U18487 ( .A1(n16418), .A2(n16417), .A3(n16416), .ZN(n16426) );
  XOR2_X1 U18488 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_211), .Z(n16425) );
  XNOR2_X1 U18489 ( .A(n16707), .B(keyinput_213), .ZN(n16424) );
  XOR2_X1 U18490 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_208), .Z(n16422) );
  XOR2_X1 U18491 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_209), .Z(n16421) );
  XOR2_X1 U18492 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_210), .Z(n16420) );
  XOR2_X1 U18493 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_212), .Z(n16419) );
  NOR4_X1 U18494 ( .A1(n16422), .A2(n16421), .A3(n16420), .A4(n16419), .ZN(
        n16423) );
  NAND4_X1 U18495 ( .A1(n16426), .A2(n16425), .A3(n16424), .A4(n16423), .ZN(
        n16434) );
  XNOR2_X1 U18496 ( .A(n16427), .B(keyinput_216), .ZN(n16433) );
  XNOR2_X1 U18497 ( .A(n16708), .B(keyinput_214), .ZN(n16430) );
  XNOR2_X1 U18498 ( .A(n16709), .B(keyinput_215), .ZN(n16429) );
  XNOR2_X1 U18499 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_218), .ZN(n16428)
         );
  NOR3_X1 U18500 ( .A1(n16430), .A2(n16429), .A3(n16428), .ZN(n16432) );
  XNOR2_X1 U18501 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_217), .ZN(n16431)
         );
  NAND4_X1 U18502 ( .A1(n16434), .A2(n16433), .A3(n16432), .A4(n16431), .ZN(
        n16438) );
  XNOR2_X1 U18503 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_219), .ZN(n16437)
         );
  XNOR2_X1 U18504 ( .A(n16435), .B(keyinput_220), .ZN(n16436) );
  AOI21_X1 U18505 ( .B1(n16438), .B2(n16437), .A(n16436), .ZN(n16444) );
  INV_X1 U18506 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n16723) );
  INV_X1 U18507 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16729) );
  AOI22_X1 U18508 ( .A1(n16723), .A2(keyinput_223), .B1(keyinput_225), .B2(
        n16729), .ZN(n16439) );
  OAI221_X1 U18509 ( .B1(n16723), .B2(keyinput_223), .C1(n16729), .C2(
        keyinput_225), .A(n16439), .ZN(n16443) );
  AOI22_X1 U18510 ( .A1(n22373), .A2(keyinput_222), .B1(n16728), .B2(
        keyinput_224), .ZN(n16440) );
  OAI221_X1 U18511 ( .B1(n22373), .B2(keyinput_222), .C1(n16728), .C2(
        keyinput_224), .A(n16440), .ZN(n16442) );
  XNOR2_X1 U18512 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_221), .ZN(n16441)
         );
  NOR4_X1 U18513 ( .A1(n16444), .A2(n16443), .A3(n16442), .A4(n16441), .ZN(
        n16446) );
  XNOR2_X1 U18514 ( .A(n20824), .B(keyinput_226), .ZN(n16445) );
  NOR2_X1 U18515 ( .A1(n16446), .A2(n16445), .ZN(n16450) );
  XNOR2_X1 U18516 ( .A(n16738), .B(keyinput_228), .ZN(n16449) );
  XNOR2_X1 U18517 ( .A(n16731), .B(keyinput_227), .ZN(n16448) );
  XNOR2_X1 U18518 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_229), .ZN(n16447)
         );
  NOR4_X1 U18519 ( .A1(n16450), .A2(n16449), .A3(n16448), .A4(n16447), .ZN(
        n16454) );
  XNOR2_X1 U18520 ( .A(n16739), .B(keyinput_230), .ZN(n16453) );
  XNOR2_X1 U18521 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_232), .ZN(n16452)
         );
  XNOR2_X1 U18522 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_231), .ZN(n16451)
         );
  OAI211_X1 U18523 ( .C1(n16454), .C2(n16453), .A(n16452), .B(n16451), .ZN(
        n16457) );
  XOR2_X1 U18524 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_233), .Z(n16456) );
  XNOR2_X1 U18525 ( .A(n16682), .B(keyinput_234), .ZN(n16455) );
  AOI21_X1 U18526 ( .B1(n16457), .B2(n16456), .A(n16455), .ZN(n16460) );
  XOR2_X1 U18527 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_235), .Z(n16459) );
  XOR2_X1 U18528 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_236), .Z(n16458) );
  OAI21_X1 U18529 ( .B1(n16460), .B2(n16459), .A(n16458), .ZN(n16464) );
  XNOR2_X1 U18530 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_237), .ZN(n16463)
         );
  XOR2_X1 U18531 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_239), .Z(n16462) );
  XNOR2_X1 U18532 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_238), .ZN(n16461)
         );
  AOI211_X1 U18533 ( .C1(n16464), .C2(n16463), .A(n16462), .B(n16461), .ZN(
        n16468) );
  XOR2_X1 U18534 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_240), .Z(n16467) );
  XNOR2_X1 U18535 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_242), .ZN(n16466)
         );
  XNOR2_X1 U18536 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_241), .ZN(n16465)
         );
  NOR4_X1 U18537 ( .A1(n16468), .A2(n16467), .A3(n16466), .A4(n16465), .ZN(
        n16471) );
  XOR2_X1 U18538 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_243), .Z(n16470) );
  XOR2_X1 U18539 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_244), .Z(n16469) );
  OAI21_X1 U18540 ( .B1(n16471), .B2(n16470), .A(n16469), .ZN(n16475) );
  XOR2_X1 U18541 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_247), .Z(n16474) );
  XNOR2_X1 U18542 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_246), .ZN(n16473)
         );
  XNOR2_X1 U18543 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n16472)
         );
  NAND4_X1 U18544 ( .A1(n16475), .A2(n16474), .A3(n16473), .A4(n16472), .ZN(
        n16478) );
  XOR2_X1 U18545 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_248), .Z(n16477) );
  XNOR2_X1 U18546 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_249), .ZN(n16476)
         );
  NAND3_X1 U18547 ( .A1(n16478), .A2(n16477), .A3(n16476), .ZN(n16481) );
  XOR2_X1 U18548 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_250), .Z(n16480) );
  XNOR2_X1 U18549 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_251), .ZN(n16479)
         );
  AOI21_X1 U18550 ( .B1(n16481), .B2(n16480), .A(n16479), .ZN(n16484) );
  XOR2_X1 U18551 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_252), .Z(n16483) );
  XOR2_X1 U18552 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_253), .Z(n16482) );
  OAI21_X1 U18553 ( .B1(n16484), .B2(n16483), .A(n16482), .ZN(n16487) );
  XOR2_X1 U18554 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_255), .Z(n16486) );
  XNOR2_X1 U18555 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_254), .ZN(n16485)
         );
  NAND3_X1 U18556 ( .A1(n16487), .A2(n16486), .A3(n16485), .ZN(n16488) );
  NAND4_X1 U18557 ( .A1(n16491), .A2(n16490), .A3(n16489), .A4(n16488), .ZN(
        n16492) );
  XOR2_X1 U18558 ( .A(n16493), .B(n16492), .Z(P1_U3481) );
  AOI22_X1 U18559 ( .A1(n16495), .A2(n16995), .B1(n11155), .B2(n16707), .ZN(
        n16513) );
  MUX2_X1 U18560 ( .A(n16513), .B(n16496), .S(n16497), .Z(n16502) );
  INV_X1 U18561 ( .A(n16497), .ZN(n16512) );
  NAND2_X1 U18562 ( .A1(n16512), .A2(n16513), .ZN(n16501) );
  AOI22_X1 U18563 ( .A1(n16499), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n16498), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16500) );
  NAND2_X1 U18564 ( .A1(n16743), .A2(n22362), .ZN(n16509) );
  NAND2_X1 U18565 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n16503) );
  NOR2_X1 U18566 ( .A1(n16534), .A2(n16503), .ZN(n16504) );
  NOR2_X1 U18567 ( .A1(n16504), .A2(n16675), .ZN(n16521) );
  INV_X1 U18568 ( .A(n16504), .ZN(n16506) );
  AOI22_X1 U18569 ( .A1(n22358), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n22371), .ZN(n16505) );
  OAI21_X1 U18570 ( .B1(n16506), .B2(P1_REIP_REG_31__SCAN_IN), .A(n16505), 
        .ZN(n16507) );
  AOI21_X1 U18571 ( .B1(n16521), .B2(P1_REIP_REG_31__SCAN_IN), .A(n16507), 
        .ZN(n16508) );
  OAI211_X1 U18572 ( .C1(n16967), .C2(n22375), .A(n16509), .B(n16508), .ZN(
        P1_U2809) );
  INV_X1 U18573 ( .A(n16530), .ZN(n16510) );
  OAI22_X1 U18574 ( .A1(n16512), .A2(n14293), .B1(n16511), .B2(n16510), .ZN(
        n16514) );
  XNOR2_X1 U18575 ( .A(n16514), .B(n16513), .ZN(n16992) );
  INV_X1 U18576 ( .A(n16515), .ZN(n16516) );
  XNOR2_X1 U18577 ( .A(n16517), .B(n16516), .ZN(n16847) );
  NAND2_X1 U18578 ( .A1(n16847), .A2(n22362), .ZN(n16523) );
  INV_X1 U18579 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20790) );
  INV_X1 U18580 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20793) );
  OAI21_X1 U18581 ( .B1(n16534), .B2(n20790), .A(n20793), .ZN(n16520) );
  AOI22_X1 U18582 ( .A1(n16843), .A2(n22353), .B1(n22371), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16518) );
  OAI21_X1 U18583 ( .B1(n22374), .B2(n16707), .A(n16518), .ZN(n16519) );
  AOI21_X1 U18584 ( .B1(n16521), .B2(n16520), .A(n16519), .ZN(n16522) );
  OAI211_X1 U18585 ( .C1(n16992), .C2(n22375), .A(n16523), .B(n16522), .ZN(
        P1_U2810) );
  OAI21_X1 U18586 ( .B1(n16675), .B2(n20787), .A(n16541), .ZN(n16533) );
  AOI22_X1 U18587 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n22371), .B1(
        n22353), .B2(n16863), .ZN(n16527) );
  OAI21_X1 U18588 ( .B1(n22374), .B2(n16709), .A(n16527), .ZN(n16532) );
  NOR2_X1 U18589 ( .A1(n16539), .A2(n16528), .ZN(n16529) );
  OR2_X1 U18590 ( .A1(n16530), .A2(n16529), .ZN(n17013) );
  NOR2_X1 U18591 ( .A1(n17013), .A2(n22375), .ZN(n16531) );
  AOI211_X1 U18592 ( .C1(n16534), .C2(n16533), .A(n16532), .B(n16531), .ZN(
        n16535) );
  OAI21_X1 U18593 ( .B1(n16861), .B2(n22377), .A(n16535), .ZN(P1_U2812) );
  AOI21_X1 U18594 ( .B1(n16538), .B2(n16537), .A(n16536), .ZN(n16869) );
  INV_X1 U18595 ( .A(n16869), .ZN(n16767) );
  AOI21_X1 U18596 ( .B1(n16540), .B2(n16557), .A(n16539), .ZN(n17028) );
  AOI21_X1 U18597 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n22339), .A(n16553), 
        .ZN(n16546) );
  INV_X1 U18598 ( .A(n16541), .ZN(n16545) );
  OAI22_X1 U18599 ( .A1(n16542), .A2(n22337), .B1(n22383), .B2(n16867), .ZN(
        n16543) );
  AOI21_X1 U18600 ( .B1(n22358), .B2(P1_EBX_REG_27__SCAN_IN), .A(n16543), .ZN(
        n16544) );
  OAI21_X1 U18601 ( .B1(n16546), .B2(n16545), .A(n16544), .ZN(n16547) );
  AOI21_X1 U18602 ( .B1(n17028), .B2(n22327), .A(n16547), .ZN(n16548) );
  OAI21_X1 U18603 ( .B1(n16767), .B2(n22377), .A(n16548), .ZN(P1_U2813) );
  XOR2_X1 U18604 ( .A(n16550), .B(n16549), .Z(n16876) );
  INV_X1 U18605 ( .A(n16876), .ZN(n16771) );
  INV_X1 U18606 ( .A(n16551), .ZN(n16874) );
  OAI22_X1 U18607 ( .A1(n16552), .A2(n22337), .B1(n22383), .B2(n16874), .ZN(
        n16556) );
  NAND2_X1 U18608 ( .A1(n22339), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16554) );
  AOI21_X1 U18609 ( .B1(n16569), .B2(n16554), .A(n16553), .ZN(n16555) );
  AOI211_X1 U18610 ( .C1(n22358), .C2(P1_EBX_REG_26__SCAN_IN), .A(n16556), .B(
        n16555), .ZN(n16560) );
  AOI21_X1 U18611 ( .B1(n16558), .B2(n16561), .A(n11567), .ZN(n17037) );
  NAND2_X1 U18612 ( .A1(n17037), .A2(n22327), .ZN(n16559) );
  OAI211_X1 U18613 ( .C1(n16771), .C2(n22377), .A(n16560), .B(n16559), .ZN(
        P1_U2814) );
  OAI21_X1 U18614 ( .B1(n16580), .B2(n16562), .A(n16561), .ZN(n17041) );
  AOI21_X1 U18615 ( .B1(n16565), .B2(n16564), .A(n16549), .ZN(n16885) );
  NAND2_X1 U18616 ( .A1(n16885), .A2(n22362), .ZN(n16572) );
  INV_X1 U18617 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20782) );
  OAI22_X1 U18618 ( .A1(n16675), .A2(n20782), .B1(n16578), .B2(n20778), .ZN(
        n16570) );
  AND2_X1 U18619 ( .A1(n22358), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n16568) );
  OAI22_X1 U18620 ( .A1(n16566), .A2(n22337), .B1(n22383), .B2(n16883), .ZN(
        n16567) );
  AOI211_X1 U18621 ( .C1(n16570), .C2(n16569), .A(n16568), .B(n16567), .ZN(
        n16571) );
  OAI211_X1 U18622 ( .C1(n22375), .C2(n17041), .A(n16572), .B(n16571), .ZN(
        P1_U2815) );
  OAI21_X1 U18623 ( .B1(n16573), .B2(n16574), .A(n16564), .ZN(n16891) );
  INV_X1 U18624 ( .A(n16578), .ZN(n16575) );
  NOR2_X1 U18625 ( .A1(n16575), .A2(n16675), .ZN(n16588) );
  AOI22_X1 U18626 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n22371), .B1(
        n22353), .B2(n16894), .ZN(n16577) );
  NAND2_X1 U18627 ( .A1(n22358), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n16576) );
  OAI211_X1 U18628 ( .C1(n16578), .C2(P1_REIP_REG_24__SCAN_IN), .A(n16577), 
        .B(n16576), .ZN(n16579) );
  AOI21_X1 U18629 ( .B1(n16588), .B2(P1_REIP_REG_24__SCAN_IN), .A(n16579), 
        .ZN(n16583) );
  AOI21_X1 U18630 ( .B1(n16581), .B2(n16593), .A(n16580), .ZN(n17057) );
  NAND2_X1 U18631 ( .A1(n17057), .A2(n22327), .ZN(n16582) );
  OAI211_X1 U18632 ( .C1(n16891), .C2(n22377), .A(n16583), .B(n16582), .ZN(
        P1_U2816) );
  AOI21_X1 U18633 ( .B1(n16586), .B2(n16585), .A(n16573), .ZN(n16902) );
  INV_X1 U18634 ( .A(n16902), .ZN(n16784) );
  INV_X1 U18635 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16587) );
  OAI22_X1 U18636 ( .A1(n16587), .A2(n22337), .B1(n22383), .B2(n16900), .ZN(
        n16592) );
  INV_X1 U18637 ( .A(n16588), .ZN(n16589) );
  AOI21_X1 U18638 ( .B1(n20777), .B2(n16590), .A(n16589), .ZN(n16591) );
  AOI211_X1 U18639 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n22358), .A(n16592), .B(
        n16591), .ZN(n16597) );
  INV_X1 U18640 ( .A(n16593), .ZN(n16594) );
  AOI21_X1 U18641 ( .B1(n16595), .B2(n16603), .A(n16594), .ZN(n17065) );
  NAND2_X1 U18642 ( .A1(n17065), .A2(n22327), .ZN(n16596) );
  OAI211_X1 U18643 ( .C1(n16784), .C2(n22377), .A(n16597), .B(n16596), .ZN(
        P1_U2817) );
  OAI21_X1 U18644 ( .B1(n16599), .B2(n16600), .A(n16585), .ZN(n16907) );
  NAND2_X1 U18645 ( .A1(n16718), .A2(n16601), .ZN(n16602) );
  NAND2_X1 U18646 ( .A1(n16603), .A2(n16602), .ZN(n16716) );
  INV_X1 U18647 ( .A(n16716), .ZN(n22198) );
  NOR2_X1 U18648 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22323), .ZN(n22369) );
  OAI21_X1 U18649 ( .B1(n22370), .B2(n22323), .A(n22255), .ZN(n22381) );
  OAI21_X1 U18650 ( .B1(n22369), .B2(n22381), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n16605) );
  AOI22_X1 U18651 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n22371), .B1(
        n22353), .B2(n16908), .ZN(n16604) );
  OAI211_X1 U18652 ( .C1(n16717), .C2(n22374), .A(n16605), .B(n16604), .ZN(
        n16608) );
  INV_X1 U18653 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20773) );
  OR3_X1 U18654 ( .A1(n22323), .A2(n16668), .A3(n16606), .ZN(n16613) );
  NOR4_X1 U18655 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n20773), .A3(n20771), 
        .A4(n16613), .ZN(n16607) );
  AOI211_X1 U18656 ( .C1(n22198), .C2(n22327), .A(n16608), .B(n16607), .ZN(
        n16609) );
  OAI21_X1 U18657 ( .B1(n16907), .B2(n22377), .A(n16609), .ZN(P1_U2818) );
  OAI21_X1 U18658 ( .B1(n16610), .B2(n16612), .A(n16611), .ZN(n16924) );
  NAND2_X1 U18659 ( .A1(n20771), .A2(n16613), .ZN(n16618) );
  AOI21_X1 U18660 ( .B1(n16614), .B2(n11292), .A(n16720), .ZN(n22191) );
  NAND2_X1 U18661 ( .A1(n22191), .A2(n22327), .ZN(n16616) );
  AOI22_X1 U18662 ( .A1(n22371), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n22353), .B2(n16921), .ZN(n16615) );
  OAI211_X1 U18663 ( .C1(n16723), .C2(n22374), .A(n16616), .B(n16615), .ZN(
        n16617) );
  AOI21_X1 U18664 ( .B1(n22381), .B2(n16618), .A(n16617), .ZN(n16619) );
  OAI21_X1 U18665 ( .B1(n16924), .B2(n22377), .A(n16619), .ZN(P1_U2820) );
  INV_X1 U18666 ( .A(n16622), .ZN(n16623) );
  AOI21_X1 U18667 ( .B1(n16624), .B2(n16621), .A(n16623), .ZN(n16930) );
  INV_X1 U18668 ( .A(n16930), .ZN(n16813) );
  NOR2_X1 U18669 ( .A1(n20762), .A2(n16625), .ZN(n22341) );
  NAND2_X1 U18670 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n22341), .ZN(n16653) );
  NOR2_X1 U18671 ( .A1(n20765), .A2(n16653), .ZN(n22350) );
  NOR2_X1 U18672 ( .A1(n16675), .A2(n22350), .ZN(n22365) );
  INV_X1 U18673 ( .A(n16649), .ZN(n16637) );
  OAI21_X1 U18674 ( .B1(n16637), .B2(n16636), .A(n16626), .ZN(n16627) );
  NAND2_X1 U18675 ( .A1(n16627), .A2(n11333), .ZN(n22172) );
  INV_X1 U18676 ( .A(n16628), .ZN(n16928) );
  OAI21_X1 U18677 ( .B1(n22383), .B2(n16928), .A(n22354), .ZN(n16630) );
  NOR2_X1 U18678 ( .A1(n22374), .A2(n16729), .ZN(n16629) );
  AOI211_X1 U18679 ( .C1(n22371), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16630), .B(n16629), .ZN(n16631) );
  OAI21_X1 U18680 ( .B1(n22375), .B2(n22172), .A(n16631), .ZN(n16632) );
  INV_X1 U18681 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20767) );
  AND2_X1 U18682 ( .A1(n20767), .A2(n22350), .ZN(n22364) );
  AOI211_X1 U18683 ( .C1(n22365), .C2(P1_REIP_REG_18__SCAN_IN), .A(n16632), 
        .B(n22364), .ZN(n16633) );
  OAI21_X1 U18684 ( .B1(n16813), .B2(n22377), .A(n16633), .ZN(P1_U2822) );
  OAI21_X1 U18685 ( .B1(n16634), .B2(n16635), .A(n16621), .ZN(n20820) );
  NAND2_X1 U18686 ( .A1(n20765), .A2(n16653), .ZN(n16643) );
  XNOR2_X1 U18687 ( .A(n16637), .B(n16636), .ZN(n20821) );
  NAND2_X1 U18688 ( .A1(n22353), .A2(n20861), .ZN(n16638) );
  OAI211_X1 U18689 ( .C1(n22337), .C2(n16639), .A(n16638), .B(n22354), .ZN(
        n16640) );
  AOI21_X1 U18690 ( .B1(n22358), .B2(P1_EBX_REG_17__SCAN_IN), .A(n16640), .ZN(
        n16641) );
  OAI21_X1 U18691 ( .B1(n20821), .B2(n22375), .A(n16641), .ZN(n16642) );
  AOI21_X1 U18692 ( .B1(n22365), .B2(n16643), .A(n16642), .ZN(n16644) );
  OAI21_X1 U18693 ( .B1(n20820), .B2(n22377), .A(n16644), .ZN(P1_U2823) );
  AOI21_X1 U18694 ( .B1(n16645), .B2(n16646), .A(n16634), .ZN(n16940) );
  INV_X1 U18695 ( .A(n16940), .ZN(n16827) );
  NOR2_X1 U18696 ( .A1(n16736), .A2(n16647), .ZN(n16648) );
  OR2_X1 U18697 ( .A1(n16649), .A2(n16648), .ZN(n16730) );
  INV_X1 U18698 ( .A(n16730), .ZN(n22181) );
  INV_X1 U18699 ( .A(n22354), .ZN(n22325) );
  INV_X1 U18700 ( .A(n16650), .ZN(n16938) );
  NOR2_X1 U18701 ( .A1(n22383), .A2(n16938), .ZN(n16651) );
  AOI211_X1 U18702 ( .C1(n22371), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n22325), .B(n16651), .ZN(n16652) );
  OAI21_X1 U18703 ( .B1(n22374), .B2(n16731), .A(n16652), .ZN(n16657) );
  AOI21_X1 U18704 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n22339), .A(n22341), 
        .ZN(n16655) );
  INV_X1 U18705 ( .A(n16653), .ZN(n16654) );
  NOR2_X1 U18706 ( .A1(n16655), .A2(n16654), .ZN(n16656) );
  AOI211_X1 U18707 ( .C1(n22181), .C2(n22327), .A(n16657), .B(n16656), .ZN(
        n16658) );
  OAI21_X1 U18708 ( .B1(n16827), .B2(n22377), .A(n16658), .ZN(P1_U2824) );
  INV_X1 U18709 ( .A(n15910), .ZN(n16659) );
  AOI21_X1 U18710 ( .B1(n16661), .B2(n16660), .A(n16659), .ZN(n16833) );
  INV_X1 U18711 ( .A(n16662), .ZN(n16832) );
  NOR2_X1 U18712 ( .A1(n16833), .A2(n16832), .ZN(n16831) );
  OAI21_X1 U18713 ( .B1(n16831), .B2(n16663), .A(n15936), .ZN(n16962) );
  OR2_X1 U18714 ( .A1(n17119), .A2(n16664), .ZN(n16665) );
  NAND2_X1 U18715 ( .A1(n16666), .A2(n16665), .ZN(n22125) );
  INV_X1 U18716 ( .A(n22125), .ZN(n16673) );
  AOI22_X1 U18717 ( .A1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n22371), .B1(
        n22353), .B2(n16965), .ZN(n16667) );
  OAI21_X1 U18718 ( .B1(n22374), .B2(n16739), .A(n16667), .ZN(n16672) );
  INV_X1 U18719 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n22130) );
  OAI211_X1 U18720 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n16669), .A(n22248), 
        .B(n16668), .ZN(n16670) );
  OAI211_X1 U18721 ( .C1(n22255), .C2(n22130), .A(n22354), .B(n16670), .ZN(
        n16671) );
  AOI211_X1 U18722 ( .C1(n16673), .C2(n22327), .A(n16672), .B(n16671), .ZN(
        n16674) );
  OAI21_X1 U18723 ( .B1(n16962), .B2(n22377), .A(n16674), .ZN(P1_U2827) );
  AOI21_X1 U18724 ( .B1(n16678), .B2(n22248), .A(n16675), .ZN(n22306) );
  AOI22_X1 U18725 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n22306), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n22371), .ZN(n16676) );
  OAI211_X1 U18726 ( .C1(n16677), .C2(n22375), .A(n16676), .B(n22354), .ZN(
        n16685) );
  INV_X1 U18727 ( .A(n16678), .ZN(n16679) );
  NOR3_X1 U18728 ( .A1(n22323), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n16679), .ZN(
        n16684) );
  INV_X1 U18729 ( .A(n16680), .ZN(n16681) );
  OAI22_X1 U18730 ( .A1(n22374), .A2(n16682), .B1(n22383), .B2(n16681), .ZN(
        n16683) );
  NOR3_X1 U18731 ( .A1(n16685), .A2(n16684), .A3(n16683), .ZN(n16686) );
  OAI21_X1 U18732 ( .B1(n16687), .B2(n22377), .A(n16686), .ZN(P1_U2831) );
  NOR2_X1 U18733 ( .A1(n16691), .A2(n16688), .ZN(n16689) );
  OR2_X1 U18734 ( .A1(n16689), .A2(n22362), .ZN(n22275) );
  OR2_X1 U18735 ( .A1(n16691), .A2(n16690), .ZN(n22265) );
  NOR2_X1 U18736 ( .A1(n22265), .A2(n22611), .ZN(n16694) );
  AOI22_X1 U18737 ( .A1(n22371), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n22238), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n16692) );
  OAI21_X1 U18738 ( .B1(n22383), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16692), .ZN(n16693) );
  AOI211_X1 U18739 ( .C1(n22327), .C2(n16695), .A(n16694), .B(n16693), .ZN(
        n16697) );
  AOI22_X1 U18740 ( .A1(n22248), .A2(n22247), .B1(n22358), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n16696) );
  OAI211_X1 U18741 ( .C1(n22259), .C2(n16698), .A(n16697), .B(n16696), .ZN(
        P1_U2839) );
  OAI21_X1 U18742 ( .B1(n22371), .B2(n22353), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16699) );
  OAI21_X1 U18743 ( .B1(n22265), .B2(n16700), .A(n16699), .ZN(n16701) );
  AOI21_X1 U18744 ( .B1(n22358), .B2(P1_EBX_REG_0__SCAN_IN), .A(n16701), .ZN(
        n16702) );
  OAI21_X1 U18745 ( .B1(n22375), .B2(n22213), .A(n16702), .ZN(n16703) );
  AOI21_X1 U18746 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n22339), .A(n16703), .ZN(
        n16704) );
  OAI21_X1 U18747 ( .B1(n22259), .B2(n16705), .A(n16704), .ZN(P1_U2840) );
  INV_X1 U18748 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16706) );
  OAI22_X1 U18749 ( .A1(n16967), .A2(n20828), .B1(n20833), .B2(n16706), .ZN(
        P1_U2841) );
  INV_X1 U18750 ( .A(n16847), .ZN(n16750) );
  OAI222_X1 U18751 ( .A1(n16750), .A2(n20812), .B1(n16707), .B2(n20833), .C1(
        n20828), .C2(n16992), .ZN(P1_U2842) );
  OAI222_X1 U18752 ( .A1(n20812), .A2(n16756), .B1(n16708), .B2(n20833), .C1(
        n17008), .C2(n20828), .ZN(P1_U2843) );
  OAI222_X1 U18753 ( .A1(n20812), .A2(n16861), .B1(n16709), .B2(n20833), .C1(
        n17013), .C2(n20828), .ZN(P1_U2844) );
  AOI22_X1 U18754 ( .A1(n17028), .A2(n20825), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n16714), .ZN(n16710) );
  OAI21_X1 U18755 ( .B1(n16767), .B2(n20812), .A(n16710), .ZN(P1_U2845) );
  AOI22_X1 U18756 ( .A1(n17037), .A2(n20825), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n16714), .ZN(n16711) );
  OAI21_X1 U18757 ( .B1(n16771), .B2(n20812), .A(n16711), .ZN(P1_U2846) );
  INV_X1 U18758 ( .A(n16885), .ZN(n16775) );
  INV_X1 U18759 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n16712) );
  OAI222_X1 U18760 ( .A1(n20812), .A2(n16775), .B1(n16712), .B2(n20833), .C1(
        n17041), .C2(n20828), .ZN(P1_U2847) );
  AOI22_X1 U18761 ( .A1(n17057), .A2(n20825), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n16714), .ZN(n16713) );
  OAI21_X1 U18762 ( .B1(n16891), .B2(n20812), .A(n16713), .ZN(P1_U2848) );
  AOI22_X1 U18763 ( .A1(n17065), .A2(n20825), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n16714), .ZN(n16715) );
  OAI21_X1 U18764 ( .B1(n16784), .B2(n20812), .A(n16715), .ZN(P1_U2849) );
  OAI222_X1 U18765 ( .A1(n16907), .A2(n20812), .B1(n20833), .B2(n16717), .C1(
        n16716), .C2(n20828), .ZN(P1_U2850) );
  OAI21_X1 U18766 ( .B1(n16720), .B2(n16719), .A(n16718), .ZN(n22376) );
  AOI21_X1 U18767 ( .B1(n16721), .B2(n16611), .A(n16599), .ZN(n20874) );
  INV_X1 U18768 ( .A(n20874), .ZN(n22378) );
  OAI222_X1 U18769 ( .A1(n20828), .A2(n22376), .B1(n20833), .B2(n22373), .C1(
        n22378), .C2(n20812), .ZN(P1_U2851) );
  INV_X1 U18770 ( .A(n22191), .ZN(n16722) );
  OAI222_X1 U18771 ( .A1(n20812), .A2(n16924), .B1(n20833), .B2(n16723), .C1(
        n16722), .C2(n20828), .ZN(P1_U2852) );
  NAND2_X1 U18772 ( .A1(n11333), .A2(n16724), .ZN(n16725) );
  NAND2_X1 U18773 ( .A1(n11292), .A2(n16725), .ZN(n22368) );
  AND2_X1 U18774 ( .A1(n16622), .A2(n16726), .ZN(n16727) );
  NOR2_X1 U18775 ( .A1(n16610), .A2(n16727), .ZN(n22363) );
  INV_X1 U18776 ( .A(n22363), .ZN(n16807) );
  OAI222_X1 U18777 ( .A1(n22368), .A2(n20828), .B1(n20833), .B2(n16728), .C1(
        n16807), .C2(n20812), .ZN(P1_U2853) );
  OAI222_X1 U18778 ( .A1(n22172), .A2(n20828), .B1(n20833), .B2(n16729), .C1(
        n16813), .C2(n20812), .ZN(P1_U2854) );
  OAI222_X1 U18779 ( .A1(n16827), .A2(n20812), .B1(n16731), .B2(n20833), .C1(
        n16730), .C2(n20828), .ZN(P1_U2856) );
  INV_X1 U18780 ( .A(n16645), .ZN(n16732) );
  AOI21_X1 U18781 ( .B1(n16733), .B2(n15937), .A(n16732), .ZN(n22345) );
  INV_X1 U18782 ( .A(n22345), .ZN(n16829) );
  AND2_X1 U18783 ( .A1(n16735), .A2(n16734), .ZN(n16737) );
  OR2_X1 U18784 ( .A1(n16737), .A2(n16736), .ZN(n22348) );
  OAI222_X1 U18785 ( .A1(n16829), .A2(n20812), .B1(n16738), .B2(n20833), .C1(
        n22348), .C2(n20828), .ZN(P1_U2857) );
  OAI222_X1 U18786 ( .A1(n16962), .A2(n20812), .B1(n16739), .B2(n20833), .C1(
        n22125), .C2(n20828), .ZN(P1_U2859) );
  INV_X1 U18787 ( .A(n16744), .ZN(n16740) );
  NAND2_X1 U18788 ( .A1(n16743), .A2(n16742), .ZN(n16746) );
  AOI22_X1 U18789 ( .A1(n16825), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n16819), .ZN(n16745) );
  OAI211_X1 U18790 ( .C1(n15058), .C2(n16823), .A(n16746), .B(n16745), .ZN(
        P1_U2873) );
  OAI22_X1 U18791 ( .A1(n16792), .A2(n22519), .B1(n22526), .B2(n16834), .ZN(
        n16747) );
  AOI21_X1 U18792 ( .B1(n16794), .B2(DATAI_30_), .A(n16747), .ZN(n16749) );
  NAND2_X1 U18793 ( .A1(n16825), .A2(BUF1_REG_30__SCAN_IN), .ZN(n16748) );
  OAI211_X1 U18794 ( .C1(n16750), .C2(n16837), .A(n16749), .B(n16748), .ZN(
        P1_U2874) );
  INV_X1 U18795 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20912) );
  OR2_X1 U18796 ( .A1(n16757), .A2(n20912), .ZN(n16752) );
  NAND2_X1 U18797 ( .A1(n16757), .A2(DATAI_13_), .ZN(n16751) );
  AND2_X1 U18798 ( .A1(n16752), .A2(n16751), .ZN(n22512) );
  OAI22_X1 U18799 ( .A1(n16792), .A2(n22512), .B1(n22516), .B2(n16834), .ZN(
        n16753) );
  AOI21_X1 U18800 ( .B1(n16794), .B2(DATAI_29_), .A(n16753), .ZN(n16755) );
  NAND2_X1 U18801 ( .A1(n16825), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16754) );
  OAI211_X1 U18802 ( .C1(n16756), .C2(n16837), .A(n16755), .B(n16754), .ZN(
        P1_U2875) );
  OR2_X1 U18803 ( .A1(n16757), .A2(n20910), .ZN(n16759) );
  NAND2_X1 U18804 ( .A1(n16757), .A2(DATAI_12_), .ZN(n16758) );
  AND2_X1 U18805 ( .A1(n16759), .A2(n16758), .ZN(n22505) );
  OAI22_X1 U18806 ( .A1(n16792), .A2(n22505), .B1(n22509), .B2(n16834), .ZN(
        n16760) );
  AOI21_X1 U18807 ( .B1(n16794), .B2(DATAI_28_), .A(n16760), .ZN(n16762) );
  NAND2_X1 U18808 ( .A1(n16825), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16761) );
  OAI211_X1 U18809 ( .C1(n16861), .C2(n16837), .A(n16762), .B(n16761), .ZN(
        P1_U2876) );
  INV_X1 U18810 ( .A(n16792), .ZN(n16821) );
  AOI22_X1 U18811 ( .A1(n16821), .A2(n22499), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16819), .ZN(n16763) );
  OAI21_X1 U18812 ( .B1(n16823), .B2(n16764), .A(n16763), .ZN(n16765) );
  AOI21_X1 U18813 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n16825), .A(n16765), .ZN(
        n16766) );
  OAI21_X1 U18814 ( .B1(n16767), .B2(n16837), .A(n16766), .ZN(P1_U2877) );
  OAI22_X1 U18815 ( .A1(n16792), .A2(n22492), .B1(n22496), .B2(n16834), .ZN(
        n16768) );
  AOI21_X1 U18816 ( .B1(n16794), .B2(DATAI_26_), .A(n16768), .ZN(n16770) );
  NAND2_X1 U18817 ( .A1(n16825), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16769) );
  OAI211_X1 U18818 ( .C1(n16771), .C2(n16837), .A(n16770), .B(n16769), .ZN(
        P1_U2878) );
  OAI22_X1 U18819 ( .A1(n16792), .A2(n22485), .B1(n22489), .B2(n16834), .ZN(
        n16772) );
  AOI21_X1 U18820 ( .B1(n16794), .B2(DATAI_25_), .A(n16772), .ZN(n16774) );
  NAND2_X1 U18821 ( .A1(n16825), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16773) );
  OAI211_X1 U18822 ( .C1(n16775), .C2(n16837), .A(n16774), .B(n16773), .ZN(
        P1_U2879) );
  OAI22_X1 U18823 ( .A1(n16792), .A2(n22479), .B1(n22482), .B2(n16834), .ZN(
        n16776) );
  AOI21_X1 U18824 ( .B1(n16794), .B2(DATAI_24_), .A(n16776), .ZN(n16778) );
  NAND2_X1 U18825 ( .A1(n16825), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16777) );
  OAI211_X1 U18826 ( .C1(n16891), .C2(n16837), .A(n16778), .B(n16777), .ZN(
        P1_U2880) );
  AOI22_X1 U18827 ( .A1(n16821), .A2(n16779), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16819), .ZN(n16780) );
  OAI21_X1 U18828 ( .B1(n16823), .B2(n16781), .A(n16780), .ZN(n16782) );
  AOI21_X1 U18829 ( .B1(n16825), .B2(BUF1_REG_23__SCAN_IN), .A(n16782), .ZN(
        n16783) );
  OAI21_X1 U18830 ( .B1(n16784), .B2(n16837), .A(n16783), .ZN(P1_U2881) );
  AOI22_X1 U18831 ( .A1(n16821), .A2(n16785), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n16819), .ZN(n16786) );
  OAI21_X1 U18832 ( .B1(n16823), .B2(n16787), .A(n16786), .ZN(n16788) );
  AOI21_X1 U18833 ( .B1(n16825), .B2(BUF1_REG_22__SCAN_IN), .A(n16788), .ZN(
        n16789) );
  OAI21_X1 U18834 ( .B1(n16907), .B2(n16837), .A(n16789), .ZN(P1_U2882) );
  OAI22_X1 U18835 ( .A1(n16792), .A2(n16791), .B1(n16790), .B2(n16834), .ZN(
        n16793) );
  AOI21_X1 U18836 ( .B1(n16794), .B2(DATAI_21_), .A(n16793), .ZN(n16796) );
  NAND2_X1 U18837 ( .A1(n16825), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16795) );
  OAI211_X1 U18838 ( .C1(n22378), .C2(n16837), .A(n16796), .B(n16795), .ZN(
        P1_U2883) );
  AOI22_X1 U18839 ( .A1(n16821), .A2(n16797), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16819), .ZN(n16798) );
  OAI21_X1 U18840 ( .B1(n16823), .B2(n16799), .A(n16798), .ZN(n16800) );
  AOI21_X1 U18841 ( .B1(n16825), .B2(BUF1_REG_20__SCAN_IN), .A(n16800), .ZN(
        n16801) );
  OAI21_X1 U18842 ( .B1(n16924), .B2(n16837), .A(n16801), .ZN(P1_U2884) );
  AOI22_X1 U18843 ( .A1(n16821), .A2(n16802), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16819), .ZN(n16803) );
  OAI21_X1 U18844 ( .B1(n16823), .B2(n16804), .A(n16803), .ZN(n16805) );
  AOI21_X1 U18845 ( .B1(n16825), .B2(BUF1_REG_19__SCAN_IN), .A(n16805), .ZN(
        n16806) );
  OAI21_X1 U18846 ( .B1(n16807), .B2(n16837), .A(n16806), .ZN(P1_U2885) );
  AOI22_X1 U18847 ( .A1(n16821), .A2(n16808), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16819), .ZN(n16809) );
  OAI21_X1 U18848 ( .B1(n16823), .B2(n16810), .A(n16809), .ZN(n16811) );
  AOI21_X1 U18849 ( .B1(n16825), .B2(BUF1_REG_18__SCAN_IN), .A(n16811), .ZN(
        n16812) );
  OAI21_X1 U18850 ( .B1(n16813), .B2(n16837), .A(n16812), .ZN(P1_U2886) );
  AOI22_X1 U18851 ( .A1(n16821), .A2(n16814), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16819), .ZN(n16815) );
  OAI21_X1 U18852 ( .B1(n16823), .B2(n16816), .A(n16815), .ZN(n16817) );
  AOI21_X1 U18853 ( .B1(n16825), .B2(BUF1_REG_17__SCAN_IN), .A(n16817), .ZN(
        n16818) );
  OAI21_X1 U18854 ( .B1(n20820), .B2(n16837), .A(n16818), .ZN(P1_U2887) );
  AOI22_X1 U18855 ( .A1(n16821), .A2(n16820), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16819), .ZN(n16822) );
  OAI21_X1 U18856 ( .B1(n16823), .B2(n14998), .A(n16822), .ZN(n16824) );
  AOI21_X1 U18857 ( .B1(n16825), .B2(BUF1_REG_16__SCAN_IN), .A(n16824), .ZN(
        n16826) );
  OAI21_X1 U18858 ( .B1(n16827), .B2(n16837), .A(n16826), .ZN(P1_U2888) );
  INV_X1 U18859 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20737) );
  OAI222_X1 U18860 ( .A1(n16829), .A2(n16837), .B1(n16836), .B2(n16828), .C1(
        n16834), .C2(n20737), .ZN(P1_U2889) );
  INV_X1 U18861 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n16830) );
  OAI222_X1 U18862 ( .A1(n16962), .A2(n16837), .B1(n22512), .B2(n16836), .C1(
        n16830), .C2(n16834), .ZN(P1_U2891) );
  AOI21_X1 U18863 ( .B1(n16833), .B2(n16832), .A(n16831), .ZN(n22328) );
  INV_X1 U18864 ( .A(n22328), .ZN(n16838) );
  OAI222_X1 U18865 ( .A1(n16838), .A2(n16837), .B1(n22505), .B2(n16836), .C1(
        n16835), .C2(n16834), .ZN(P1_U2892) );
  INV_X1 U18866 ( .A(n16839), .ZN(n16841) );
  XNOR2_X1 U18867 ( .A(n11160), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16850) );
  XNOR2_X1 U18868 ( .A(n16842), .B(n16995), .ZN(n17002) );
  NAND2_X1 U18869 ( .A1(n20862), .A2(n16843), .ZN(n16844) );
  NAND2_X1 U18870 ( .A1(n22202), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16996) );
  OAI211_X1 U18871 ( .C1(n20842), .C2(n16845), .A(n16844), .B(n16996), .ZN(
        n16846) );
  AOI21_X1 U18872 ( .B1(n16847), .B2(n20873), .A(n16846), .ZN(n16848) );
  OAI21_X1 U18873 ( .B1(n17002), .B2(n22385), .A(n16848), .ZN(P1_U2969) );
  XOR2_X1 U18874 ( .A(n16850), .B(n16849), .Z(n17012) );
  NOR2_X1 U18875 ( .A1(n22129), .A2(n20790), .ZN(n17006) );
  AOI21_X1 U18876 ( .B1(n20870), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n17006), .ZN(n16851) );
  OAI21_X1 U18877 ( .B1(n20877), .B2(n16852), .A(n16851), .ZN(n16853) );
  AOI21_X1 U18878 ( .B1(n16854), .B2(n20873), .A(n16853), .ZN(n16855) );
  OAI21_X1 U18879 ( .B1(n22385), .B2(n17012), .A(n16855), .ZN(P1_U2970) );
  NAND2_X1 U18880 ( .A1(n17134), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16857) );
  OAI21_X1 U18881 ( .B1(n17134), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16857), .ZN(n16859) );
  INV_X1 U18882 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17034) );
  INV_X1 U18883 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16860) );
  NAND2_X1 U18884 ( .A1(n22202), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n17015) );
  OAI21_X1 U18885 ( .B1(n20842), .B2(n16860), .A(n17015), .ZN(n16862) );
  NAND2_X1 U18886 ( .A1(n16871), .A2(n11294), .ZN(n16865) );
  XNOR2_X1 U18887 ( .A(n11160), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16864) );
  XNOR2_X1 U18888 ( .A(n16865), .B(n16864), .ZN(n17030) );
  NAND2_X1 U18889 ( .A1(n22202), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n17023) );
  NAND2_X1 U18890 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16866) );
  OAI211_X1 U18891 ( .C1(n20877), .C2(n16867), .A(n17023), .B(n16866), .ZN(
        n16868) );
  AOI21_X1 U18892 ( .B1(n16869), .B2(n20873), .A(n16868), .ZN(n16870) );
  OAI21_X1 U18893 ( .B1(n17030), .B2(n22385), .A(n16870), .ZN(P1_U2972) );
  OAI21_X1 U18894 ( .B1(n16872), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16871), .ZN(n17040) );
  NOR2_X1 U18895 ( .A1(n22129), .A2(n20784), .ZN(n17036) );
  AOI21_X1 U18896 ( .B1(n20870), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17036), .ZN(n16873) );
  OAI21_X1 U18897 ( .B1(n20877), .B2(n16874), .A(n16873), .ZN(n16875) );
  AOI21_X1 U18898 ( .B1(n16876), .B2(n20873), .A(n16875), .ZN(n16877) );
  OAI21_X1 U18899 ( .B1(n22385), .B2(n17040), .A(n16877), .ZN(P1_U2973) );
  INV_X1 U18900 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16878) );
  AOI21_X1 U18901 ( .B1(n16897), .B2(n16878), .A(n16984), .ZN(n16880) );
  NOR2_X1 U18902 ( .A1(n11160), .A2(n17052), .ZN(n16896) );
  NOR3_X1 U18903 ( .A1(n16880), .A2(n16879), .A3(n16896), .ZN(n16881) );
  XNOR2_X1 U18904 ( .A(n16881), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17049) );
  NOR2_X1 U18905 ( .A1(n22129), .A2(n20782), .ZN(n17042) );
  AOI21_X1 U18906 ( .B1(n20870), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17042), .ZN(n16882) );
  OAI21_X1 U18907 ( .B1(n20877), .B2(n16883), .A(n16882), .ZN(n16884) );
  AOI21_X1 U18908 ( .B1(n16885), .B2(n20873), .A(n16884), .ZN(n16886) );
  OAI21_X1 U18909 ( .B1(n22385), .B2(n17049), .A(n16886), .ZN(P1_U2974) );
  NAND2_X1 U18910 ( .A1(n13229), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16888) );
  NAND3_X1 U18911 ( .A1(n16897), .A2(n17134), .A3(n17052), .ZN(n16887) );
  OAI21_X1 U18912 ( .B1(n16897), .B2(n16888), .A(n16887), .ZN(n16889) );
  XNOR2_X1 U18913 ( .A(n16889), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17060) );
  NAND2_X1 U18914 ( .A1(n22202), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n17051) );
  OAI21_X1 U18915 ( .B1(n20842), .B2(n16890), .A(n17051), .ZN(n16893) );
  NOR2_X1 U18916 ( .A1(n16891), .A2(n20853), .ZN(n16892) );
  AOI211_X1 U18917 ( .C1(n20862), .C2(n16894), .A(n16893), .B(n16892), .ZN(
        n16895) );
  OAI21_X1 U18918 ( .B1(n17060), .B2(n22385), .A(n16895), .ZN(P1_U2975) );
  AOI21_X1 U18919 ( .B1(n13229), .B2(n17052), .A(n16896), .ZN(n16898) );
  XOR2_X1 U18920 ( .A(n16898), .B(n16897), .Z(n17068) );
  NOR2_X1 U18921 ( .A1(n22129), .A2(n20777), .ZN(n17062) );
  AOI21_X1 U18922 ( .B1(n20870), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17062), .ZN(n16899) );
  OAI21_X1 U18923 ( .B1(n20877), .B2(n16900), .A(n16899), .ZN(n16901) );
  AOI21_X1 U18924 ( .B1(n16902), .B2(n20873), .A(n16901), .ZN(n16903) );
  OAI21_X1 U18925 ( .B1(n17068), .B2(n22385), .A(n16903), .ZN(P1_U2976) );
  NOR2_X1 U18926 ( .A1(n16905), .A2(n16904), .ZN(n16906) );
  XNOR2_X1 U18927 ( .A(n16906), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n22197) );
  INV_X1 U18928 ( .A(n16907), .ZN(n16912) );
  INV_X1 U18929 ( .A(n16908), .ZN(n16910) );
  AOI22_X1 U18930 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n22202), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16909) );
  OAI21_X1 U18931 ( .B1(n20877), .B2(n16910), .A(n16909), .ZN(n16911) );
  AOI21_X1 U18932 ( .B1(n16912), .B2(n20873), .A(n16911), .ZN(n16913) );
  OAI21_X1 U18933 ( .B1(n22385), .B2(n22197), .A(n16913), .ZN(P1_U2977) );
  INV_X1 U18934 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n22196) );
  INV_X1 U18935 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17081) );
  MUX2_X1 U18936 ( .A(n16915), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .S(
        n13229), .Z(n16926) );
  NAND2_X1 U18937 ( .A1(n16914), .A2(n16926), .ZN(n16925) );
  OR2_X1 U18938 ( .A1(n13229), .A2(n16915), .ZN(n16916) );
  INV_X1 U18939 ( .A(n17083), .ZN(n16917) );
  MUX2_X1 U18940 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17083), .S(
        n17134), .Z(n17070) );
  OAI21_X1 U18941 ( .B1(n17081), .B2(n16917), .A(n17070), .ZN(n16918) );
  XOR2_X1 U18942 ( .A(n22196), .B(n16918), .Z(n22192) );
  NAND2_X1 U18943 ( .A1(n22192), .A2(n20872), .ZN(n16923) );
  OAI22_X1 U18944 ( .A1(n20842), .A2(n16919), .B1(n22129), .B2(n20771), .ZN(
        n16920) );
  AOI21_X1 U18945 ( .B1(n20862), .B2(n16921), .A(n16920), .ZN(n16922) );
  OAI211_X1 U18946 ( .C1(n20853), .C2(n16924), .A(n16923), .B(n16922), .ZN(
        P1_U2979) );
  OAI21_X1 U18947 ( .B1(n16914), .B2(n16926), .A(n16925), .ZN(n22169) );
  AOI22_X1 U18948 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n22202), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n16927) );
  OAI21_X1 U18949 ( .B1(n20877), .B2(n16928), .A(n16927), .ZN(n16929) );
  AOI21_X1 U18950 ( .B1(n16930), .B2(n20873), .A(n16929), .ZN(n16931) );
  OAI21_X1 U18951 ( .B1(n22385), .B2(n22169), .A(n16931), .ZN(P1_U2981) );
  NOR2_X1 U18952 ( .A1(n11305), .A2(n16932), .ZN(n16933) );
  INV_X1 U18953 ( .A(n16933), .ZN(n20858) );
  NOR2_X1 U18954 ( .A1(n20858), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16935) );
  NOR2_X1 U18955 ( .A1(n16933), .A2(n14256), .ZN(n16934) );
  MUX2_X1 U18956 ( .A(n16935), .B(n16934), .S(n13229), .Z(n16936) );
  XNOR2_X1 U18957 ( .A(n16936), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n22180) );
  AOI22_X1 U18958 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n22202), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16937) );
  OAI21_X1 U18959 ( .B1(n20877), .B2(n16938), .A(n16937), .ZN(n16939) );
  AOI21_X1 U18960 ( .B1(n16940), .B2(n20873), .A(n16939), .ZN(n16941) );
  OAI21_X1 U18961 ( .B1(n22180), .B2(n22385), .A(n16941), .ZN(P1_U2983) );
  NOR2_X1 U18962 ( .A1(n17137), .A2(n16943), .ZN(n17091) );
  AOI21_X1 U18963 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17134), .ZN(n16956) );
  NOR3_X1 U18964 ( .A1(n17091), .A2(n16956), .A3(n16944), .ZN(n16947) );
  INV_X1 U18965 ( .A(n16945), .ZN(n16946) );
  NOR2_X1 U18966 ( .A1(n16947), .A2(n16946), .ZN(n16949) );
  XNOR2_X1 U18967 ( .A(n17134), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16948) );
  XNOR2_X1 U18968 ( .A(n16949), .B(n16948), .ZN(n22131) );
  AOI22_X1 U18969 ( .A1(n20870), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n22202), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16950) );
  OAI21_X1 U18970 ( .B1(n20877), .B2(n16951), .A(n16950), .ZN(n16952) );
  AOI21_X1 U18971 ( .B1(n16953), .B2(n20873), .A(n16952), .ZN(n16954) );
  OAI21_X1 U18972 ( .B1(n22131), .B2(n22385), .A(n16954), .ZN(P1_U2985) );
  OAI22_X1 U18973 ( .A1(n11414), .A2(n16956), .B1(n16955), .B2(n11160), .ZN(
        n17114) );
  INV_X1 U18974 ( .A(n16958), .ZN(n16957) );
  OAI21_X1 U18975 ( .B1(n13229), .B2(n16970), .A(n16957), .ZN(n17113) );
  NOR2_X1 U18976 ( .A1(n17114), .A2(n17113), .ZN(n17112) );
  NOR2_X1 U18977 ( .A1(n17112), .A2(n16958), .ZN(n16959) );
  XOR2_X1 U18978 ( .A(n16960), .B(n16959), .Z(n22124) );
  INV_X1 U18979 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16961) );
  OAI22_X1 U18980 ( .A1(n20842), .A2(n16961), .B1(n22129), .B2(n22130), .ZN(
        n16964) );
  NOR2_X1 U18981 ( .A1(n16962), .A2(n20853), .ZN(n16963) );
  AOI211_X1 U18982 ( .C1(n20862), .C2(n16965), .A(n16964), .B(n16963), .ZN(
        n16966) );
  OAI21_X1 U18983 ( .B1(n22124), .B2(n22385), .A(n16966), .ZN(P1_U2986) );
  NAND2_X1 U18984 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17100) );
  NOR3_X1 U18985 ( .A1(n16915), .A2(n22168), .A3(n17100), .ZN(n16974) );
  NAND3_X1 U18986 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n16968), .ZN(n16972) );
  NOR2_X1 U18987 ( .A1(n16972), .A2(n16969), .ZN(n17072) );
  NAND2_X1 U18988 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17072), .ZN(
        n17124) );
  NOR2_X1 U18989 ( .A1(n16970), .A2(n17124), .ZN(n22120) );
  NAND2_X1 U18990 ( .A1(n16974), .A2(n22120), .ZN(n17084) );
  INV_X1 U18991 ( .A(n16975), .ZN(n22207) );
  NAND2_X1 U18992 ( .A1(n22207), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16971) );
  NOR2_X1 U18993 ( .A1(n17084), .A2(n16971), .ZN(n16981) );
  INV_X1 U18994 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n22205) );
  NOR2_X1 U18995 ( .A1(n16973), .A2(n16972), .ZN(n17121) );
  NAND3_X1 U18996 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n17121), .ZN(n22122) );
  INV_X1 U18997 ( .A(n22122), .ZN(n22116) );
  NAND2_X1 U18998 ( .A1(n22116), .A2(n16974), .ZN(n17073) );
  NOR3_X1 U18999 ( .A1(n22205), .A2(n16975), .A3(n17073), .ZN(n16980) );
  OR2_X1 U19000 ( .A1(n17122), .A2(n16980), .ZN(n16976) );
  OAI21_X1 U19001 ( .B1(n22119), .B2(n16981), .A(n16976), .ZN(n16977) );
  NOR2_X1 U19002 ( .A1(n17102), .A2(n16977), .ZN(n17061) );
  OAI21_X1 U19003 ( .B1(n17103), .B2(n16984), .A(n17061), .ZN(n17043) );
  NAND2_X1 U19004 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16986) );
  NAND2_X1 U19005 ( .A1(n17103), .A2(n22118), .ZN(n17075) );
  OAI21_X1 U19006 ( .B1(n17043), .B2(n16986), .A(n17075), .ZN(n17025) );
  NAND2_X1 U19007 ( .A1(n17025), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16978) );
  AOI21_X1 U19008 ( .B1(n16978), .B2(n17075), .A(n16995), .ZN(n16993) );
  INV_X1 U19009 ( .A(n17075), .ZN(n17003) );
  AOI211_X1 U19010 ( .C1(n16993), .C2(n11437), .A(n17003), .B(n16979), .ZN(
        n16990) );
  NAND2_X1 U19011 ( .A1(n17105), .A2(n16980), .ZN(n16983) );
  NAND2_X1 U19012 ( .A1(n17125), .A2(n16981), .ZN(n16982) );
  INV_X1 U19013 ( .A(n16984), .ZN(n16985) );
  NOR2_X1 U19014 ( .A1(n17053), .A2(n16985), .ZN(n17031) );
  INV_X1 U19015 ( .A(n16986), .ZN(n17032) );
  NAND2_X1 U19016 ( .A1(n17031), .A2(n17032), .ZN(n17022) );
  OR3_X1 U19017 ( .A1(n17022), .A2(n17004), .A3(n16987), .ZN(n16994) );
  NOR3_X1 U19018 ( .A1(n16994), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16995), .ZN(n16988) );
  INV_X1 U19019 ( .A(n16992), .ZN(n17000) );
  AOI21_X1 U19020 ( .B1(n16995), .B2(n16994), .A(n16993), .ZN(n16999) );
  NAND3_X1 U19021 ( .A1(n17075), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n17004), .ZN(n16997) );
  NAND2_X1 U19022 ( .A1(n16997), .A2(n16996), .ZN(n16998) );
  AOI211_X1 U19023 ( .C1(n17000), .C2(n22199), .A(n16999), .B(n16998), .ZN(
        n17001) );
  OAI21_X1 U19024 ( .B1(n17002), .B2(n22218), .A(n17001), .ZN(P1_U3001) );
  OAI21_X1 U19025 ( .B1(n11437), .B2(n17003), .A(n17025), .ZN(n17007) );
  NOR3_X1 U19026 ( .A1(n17022), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n17004), .ZN(n17005) );
  AOI211_X1 U19027 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n17007), .A(
        n17006), .B(n17005), .ZN(n17011) );
  INV_X1 U19028 ( .A(n17008), .ZN(n17009) );
  NAND2_X1 U19029 ( .A1(n17009), .A2(n22199), .ZN(n17010) );
  OAI211_X1 U19030 ( .C1(n17012), .C2(n22218), .A(n17011), .B(n17010), .ZN(
        P1_U3002) );
  INV_X1 U19031 ( .A(n17013), .ZN(n17019) );
  NOR3_X1 U19032 ( .A1(n17022), .A2(n17014), .A3(n11437), .ZN(n17018) );
  INV_X1 U19033 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17016) );
  OAI21_X1 U19034 ( .B1(n17025), .B2(n17016), .A(n17015), .ZN(n17017) );
  AOI211_X1 U19035 ( .C1(n17019), .C2(n22199), .A(n17018), .B(n17017), .ZN(
        n17020) );
  OAI21_X1 U19036 ( .B1(n17021), .B2(n22218), .A(n17020), .ZN(P1_U3003) );
  NOR2_X1 U19037 ( .A1(n17022), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17027) );
  OAI21_X1 U19038 ( .B1(n17025), .B2(n17024), .A(n17023), .ZN(n17026) );
  AOI211_X1 U19039 ( .C1(n17028), .C2(n22199), .A(n17027), .B(n17026), .ZN(
        n17029) );
  OAI21_X1 U19040 ( .B1(n17030), .B2(n22218), .A(n17029), .ZN(P1_U3004) );
  INV_X1 U19041 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17033) );
  INV_X1 U19042 ( .A(n17031), .ZN(n17045) );
  AOI211_X1 U19043 ( .C1(n17034), .C2(n17033), .A(n17032), .B(n17045), .ZN(
        n17035) );
  AOI211_X1 U19044 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17043), .A(
        n17036), .B(n17035), .ZN(n17039) );
  NAND2_X1 U19045 ( .A1(n17037), .A2(n22199), .ZN(n17038) );
  OAI211_X1 U19046 ( .C1(n17040), .C2(n22218), .A(n17039), .B(n17038), .ZN(
        P1_U3005) );
  INV_X1 U19047 ( .A(n17041), .ZN(n17047) );
  AOI21_X1 U19048 ( .B1(n17043), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17042), .ZN(n17044) );
  OAI21_X1 U19049 ( .B1(n17045), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17044), .ZN(n17046) );
  AOI21_X1 U19050 ( .B1(n17047), .B2(n22199), .A(n17046), .ZN(n17048) );
  OAI21_X1 U19051 ( .B1(n17049), .B2(n22218), .A(n17048), .ZN(P1_U3006) );
  NOR2_X1 U19052 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17053), .ZN(
        n17063) );
  INV_X1 U19053 ( .A(n17063), .ZN(n17050) );
  NAND2_X1 U19054 ( .A1(n17061), .A2(n17050), .ZN(n17056) );
  INV_X1 U19055 ( .A(n17051), .ZN(n17055) );
  NOR3_X1 U19056 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17053), .A3(
        n17052), .ZN(n17054) );
  AOI211_X1 U19057 ( .C1(n17056), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n17055), .B(n17054), .ZN(n17059) );
  NAND2_X1 U19058 ( .A1(n17057), .A2(n22199), .ZN(n17058) );
  OAI211_X1 U19059 ( .C1(n17060), .C2(n22218), .A(n17059), .B(n17058), .ZN(
        P1_U3007) );
  INV_X1 U19060 ( .A(n17061), .ZN(n17064) );
  AOI211_X1 U19061 ( .C1(n17064), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17063), .B(n17062), .ZN(n17067) );
  NAND2_X1 U19062 ( .A1(n17065), .A2(n22199), .ZN(n17066) );
  OAI211_X1 U19063 ( .C1(n17068), .C2(n22218), .A(n17067), .B(n17066), .ZN(
        P1_U3008) );
  AOI22_X1 U19064 ( .A1(n17083), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n22196), .ZN(n17069) );
  NAND2_X1 U19065 ( .A1(n17070), .A2(n17069), .ZN(n17071) );
  XNOR2_X1 U19066 ( .A(n17071), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n20871) );
  AOI22_X1 U19067 ( .A1(n17125), .A2(n17072), .B1(n17121), .B2(n17105), .ZN(
        n22139) );
  OR3_X1 U19068 ( .A1(n22196), .A2(n17081), .A3(n17084), .ZN(n17076) );
  NOR3_X1 U19069 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n22139), .A3(
        n17076), .ZN(n22203) );
  AOI22_X1 U19070 ( .A1(n17125), .A2(n17084), .B1(n22147), .B2(n17073), .ZN(
        n17074) );
  NAND2_X1 U19071 ( .A1(n22118), .A2(n17074), .ZN(n22186) );
  OAI21_X1 U19072 ( .B1(n22186), .B2(n17076), .A(n17075), .ZN(n17077) );
  INV_X1 U19073 ( .A(n17077), .ZN(n22204) );
  AOI22_X1 U19074 ( .A1(n22204), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n22202), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n17078) );
  OAI21_X1 U19075 ( .B1(n22376), .B2(n22214), .A(n17078), .ZN(n17079) );
  AOI211_X1 U19076 ( .C1(n20871), .C2(n22200), .A(n22203), .B(n17079), .ZN(
        n17080) );
  INV_X1 U19077 ( .A(n17080), .ZN(P1_U3010) );
  MUX2_X1 U19078 ( .A(n17081), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .S(
        n13229), .Z(n17082) );
  XNOR2_X1 U19079 ( .A(n17083), .B(n17082), .ZN(n20867) );
  NOR2_X1 U19080 ( .A1(n22139), .A2(n17084), .ZN(n22206) );
  AOI22_X1 U19081 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n22186), .B1(
        n22206), .B2(n17081), .ZN(n17086) );
  NAND2_X1 U19082 ( .A1(n22202), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n17085) );
  OAI211_X1 U19083 ( .C1(n22214), .C2(n22368), .A(n17086), .B(n17085), .ZN(
        n17087) );
  AOI21_X1 U19084 ( .B1(n20867), .B2(n22200), .A(n17087), .ZN(n17088) );
  INV_X1 U19085 ( .A(n17088), .ZN(P1_U3012) );
  INV_X1 U19086 ( .A(n17089), .ZN(n17090) );
  NOR2_X1 U19087 ( .A1(n17091), .A2(n17090), .ZN(n17092) );
  AOI211_X1 U19088 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n17134), .A(
        n17093), .B(n17092), .ZN(n17094) );
  INV_X1 U19089 ( .A(n17094), .ZN(n17097) );
  AOI21_X1 U19090 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11160), .A(
        n17094), .ZN(n17095) );
  AOI21_X1 U19091 ( .B1(n13229), .B2(n17098), .A(n17095), .ZN(n17096) );
  OAI21_X1 U19092 ( .B1(n17098), .B2(n17097), .A(n17096), .ZN(n17099) );
  XNOR2_X1 U19093 ( .A(n17099), .B(n17108), .ZN(n20866) );
  INV_X1 U19094 ( .A(n22168), .ZN(n17104) );
  NOR2_X1 U19095 ( .A1(n22122), .A2(n17100), .ZN(n17106) );
  INV_X1 U19096 ( .A(n22120), .ZN(n22115) );
  NOR2_X1 U19097 ( .A1(n17100), .A2(n22115), .ZN(n17107) );
  OAI22_X1 U19098 ( .A1(n17122), .A2(n17106), .B1(n17107), .B2(n22119), .ZN(
        n17101) );
  NOR2_X1 U19099 ( .A1(n17102), .A2(n17101), .ZN(n22185) );
  OAI21_X1 U19100 ( .B1(n17104), .B2(n17103), .A(n22185), .ZN(n22173) );
  AOI22_X1 U19101 ( .A1(n17125), .A2(n17107), .B1(n17106), .B2(n17105), .ZN(
        n22177) );
  OAI21_X1 U19102 ( .B1(n22177), .B2(n22178), .A(n17108), .ZN(n17110) );
  OAI22_X1 U19103 ( .A1(n20821), .A2(n22214), .B1(n22129), .B2(n20765), .ZN(
        n17109) );
  AOI21_X1 U19104 ( .B1(n22173), .B2(n17110), .A(n17109), .ZN(n17111) );
  OAI21_X1 U19105 ( .B1(n20866), .B2(n22218), .A(n17111), .ZN(P1_U3014) );
  AOI21_X1 U19106 ( .B1(n17114), .B2(n17113), .A(n17112), .ZN(n20856) );
  NOR2_X1 U19107 ( .A1(n20856), .A2(n22218), .ZN(n17133) );
  INV_X1 U19108 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17126) );
  NOR3_X1 U19109 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n22139), .A3(
        n17126), .ZN(n17132) );
  INV_X1 U19110 ( .A(n17115), .ZN(n17118) );
  AOI21_X1 U19111 ( .B1(n17118), .B2(n17117), .A(n17116), .ZN(n17120) );
  OR2_X1 U19112 ( .A1(n17120), .A2(n17119), .ZN(n20813) );
  OAI21_X1 U19113 ( .B1(n17122), .B2(n17121), .A(n22118), .ZN(n17123) );
  AOI21_X1 U19114 ( .B1(n17125), .B2(n17124), .A(n17123), .ZN(n17127) );
  AOI22_X1 U19115 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17127), .B1(
        n22139), .B2(n17126), .ZN(n17138) );
  INV_X1 U19116 ( .A(n17127), .ZN(n17128) );
  OAI21_X1 U19117 ( .B1(n17138), .B2(n17128), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17130) );
  NAND2_X1 U19118 ( .A1(n22202), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n17129) );
  OAI211_X1 U19119 ( .C1(n20813), .C2(n22214), .A(n17130), .B(n17129), .ZN(
        n17131) );
  OR3_X1 U19120 ( .A1(n17133), .A2(n17132), .A3(n17131), .ZN(P1_U3019) );
  MUX2_X1 U19121 ( .A(n17135), .B(n17137), .S(n17134), .Z(n17140) );
  INV_X1 U19122 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17136) );
  NOR2_X1 U19123 ( .A1(n17140), .A2(n17136), .ZN(n17141) );
  INV_X1 U19124 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20755) );
  NOR2_X1 U19125 ( .A1(n22129), .A2(n20755), .ZN(n20850) );
  AOI211_X1 U19126 ( .C1(n22199), .C2(n22313), .A(n20850), .B(n17138), .ZN(
        n17139) );
  OAI21_X1 U19127 ( .B1(n20848), .B2(n22218), .A(n17139), .ZN(P1_U3020) );
  INV_X1 U19128 ( .A(n17140), .ZN(n17143) );
  INV_X1 U19129 ( .A(n17141), .ZN(n17142) );
  OAI21_X1 U19130 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17143), .A(
        n17142), .ZN(n20847) );
  AOI22_X1 U19131 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(n17136), .B2(n17144), .ZN(
        n17145) );
  AOI22_X1 U19132 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17147), .B1(
        n17146), .B2(n17145), .ZN(n17150) );
  OAI22_X1 U19133 ( .A1(n22214), .A2(n20816), .B1(n22129), .B2(n20753), .ZN(
        n17148) );
  INV_X1 U19134 ( .A(n17148), .ZN(n17149) );
  OAI211_X1 U19135 ( .C1(n20847), .C2(n22218), .A(n17150), .B(n17149), .ZN(
        P1_U3021) );
  NAND2_X1 U19136 ( .A1(n17152), .A2(n17151), .ZN(n22563) );
  NOR2_X1 U19137 ( .A1(n11254), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n17154) );
  INV_X1 U19138 ( .A(n17153), .ZN(n17160) );
  OAI22_X1 U19139 ( .A1(n22563), .A2(n17154), .B1(n22611), .B2(n17160), .ZN(
        n17156) );
  MUX2_X1 U19140 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n17156), .S(
        n17155), .Z(P1_U3477) );
  MUX2_X1 U19141 ( .A(n22563), .B(n17157), .S(n13301), .Z(n17158) );
  OAI21_X1 U19142 ( .B1(n17160), .B2(n17159), .A(n17158), .ZN(n17161) );
  MUX2_X1 U19143 ( .A(n17161), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n18057), .Z(P1_U3476) );
  INV_X1 U19144 ( .A(n17162), .ZN(n17172) );
  NAND3_X1 U19145 ( .A1(n17163), .A2(n17171), .A3(n17172), .ZN(n17164) );
  OAI21_X1 U19146 ( .B1(n17165), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n17164), .ZN(n17166) );
  AOI21_X1 U19147 ( .B1(n22629), .B2(n17167), .A(n17166), .ZN(n18016) );
  INV_X1 U19148 ( .A(n17168), .ZN(n17169) );
  NAND2_X1 U19149 ( .A1(n17170), .A2(n17169), .ZN(n17174) );
  NAND3_X1 U19150 ( .A1(n17172), .A2(n22396), .A3(n17171), .ZN(n17173) );
  OAI211_X1 U19151 ( .C1(n18016), .C2(n17175), .A(n17174), .B(n17173), .ZN(
        n17176) );
  MUX2_X1 U19152 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n17176), .S(
        n17979), .Z(P1_U3473) );
  AND2_X1 U19153 ( .A1(n11264), .A2(n17177), .ZN(n17178) );
  OR2_X1 U19154 ( .A1(n17178), .A2(n16063), .ZN(n17680) );
  OAI211_X1 U19155 ( .C1(n17180), .C2(n17446), .A(n19484), .B(n17179), .ZN(
        n17192) );
  NOR2_X1 U19156 ( .A1(n17181), .A2(n19393), .ZN(n17190) );
  NAND2_X1 U19157 ( .A1(n17262), .A2(n17182), .ZN(n17183) );
  NAND2_X1 U19158 ( .A1(n17184), .A2(n17183), .ZN(n17672) );
  NOR2_X1 U19159 ( .A1(n17672), .A2(n19467), .ZN(n17189) );
  INV_X1 U19160 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17185) );
  INV_X1 U19161 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17445) );
  OAI22_X1 U19162 ( .A1(n17185), .A2(n19462), .B1(n17445), .B2(n19386), .ZN(
        n17188) );
  INV_X1 U19163 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n17186) );
  NOR2_X1 U19164 ( .A1(n19464), .A2(n17186), .ZN(n17187) );
  NOR4_X1 U19165 ( .A1(n17190), .A2(n17189), .A3(n17188), .A4(n17187), .ZN(
        n17191) );
  OAI211_X1 U19166 ( .C1(n17680), .C2(n19477), .A(n17192), .B(n17191), .ZN(
        P2_U2828) );
  AOI21_X1 U19167 ( .B1(n17194), .B2(n17193), .A(n19563), .ZN(n17195) );
  NAND2_X1 U19168 ( .A1(n17196), .A2(n17195), .ZN(n17202) );
  AOI22_X1 U19169 ( .A1(n19491), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19495), .ZN(n17198) );
  NAND2_X1 U19170 ( .A1(n19494), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n17197) );
  OAI211_X1 U19171 ( .C1(n17297), .C2(n19467), .A(n17198), .B(n17197), .ZN(
        n17199) );
  AOI21_X1 U19172 ( .B1(n17200), .B2(n19492), .A(n17199), .ZN(n17201) );
  OAI211_X1 U19173 ( .C1(n19477), .C2(n17385), .A(n17202), .B(n17201), .ZN(
        P2_U2834) );
  AOI211_X1 U19174 ( .C1(n17540), .C2(n17204), .A(n17203), .B(n19563), .ZN(
        n17205) );
  INV_X1 U19175 ( .A(n17205), .ZN(n17213) );
  AOI22_X1 U19176 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19495), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19494), .ZN(n17206) );
  OAI211_X1 U19177 ( .C1(n19464), .C2(n17207), .A(n17206), .B(n19301), .ZN(
        n17210) );
  NOR2_X1 U19178 ( .A1(n17208), .A2(n19467), .ZN(n17209) );
  AOI211_X1 U19179 ( .C1(n19492), .C2(n17211), .A(n17210), .B(n17209), .ZN(
        n17212) );
  OAI211_X1 U19180 ( .C1(n19477), .C2(n17793), .A(n17213), .B(n17212), .ZN(
        P2_U2838) );
  NOR2_X1 U19181 ( .A1(n19396), .A2(n17214), .ZN(n17215) );
  XNOR2_X1 U19182 ( .A(n17215), .B(n17614), .ZN(n17216) );
  NAND2_X1 U19183 ( .A1(n17216), .A2(n19484), .ZN(n17227) );
  AOI22_X1 U19184 ( .A1(n17217), .A2(n19492), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19495), .ZN(n17218) );
  OAI211_X1 U19185 ( .C1(n12129), .C2(n19464), .A(n17218), .B(n19301), .ZN(
        n17219) );
  AOI21_X1 U19186 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n19494), .A(n17219), .ZN(
        n17226) );
  INV_X1 U19187 ( .A(n17221), .ZN(n17222) );
  AOI21_X1 U19188 ( .B1(n17223), .B2(n17220), .A(n17222), .ZN(n20074) );
  NAND2_X1 U19189 ( .A1(n20074), .A2(n12449), .ZN(n17225) );
  NAND2_X1 U19190 ( .A1(n17906), .A2(n19498), .ZN(n17224) );
  NAND4_X1 U19191 ( .A1(n17227), .A2(n17226), .A3(n17225), .A4(n17224), .ZN(
        P2_U2846) );
  INV_X1 U19192 ( .A(n20496), .ZN(n17236) );
  NAND2_X1 U19193 ( .A1(n19492), .A2(n17228), .ZN(n17235) );
  XOR2_X1 U19194 ( .A(n17230), .B(n17229), .Z(n17946) );
  NAND2_X1 U19195 ( .A1(n17946), .A2(n19501), .ZN(n17232) );
  AOI22_X1 U19196 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19495), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19494), .ZN(n17231) );
  OAI211_X1 U19197 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19311), .A(
        n17232), .B(n17231), .ZN(n17233) );
  AOI21_X1 U19198 ( .B1(n19491), .B2(P2_EBX_REG_1__SCAN_IN), .A(n17233), .ZN(
        n17234) );
  OAI211_X1 U19199 ( .C1(n17236), .C2(n19477), .A(n17235), .B(n17234), .ZN(
        n17237) );
  AOI21_X1 U19200 ( .B1(n19498), .B2(n17238), .A(n17237), .ZN(n17239) );
  OAI21_X1 U19201 ( .B1(n20108), .B2(n17240), .A(n17239), .ZN(P2_U2854) );
  INV_X1 U19202 ( .A(n17241), .ZN(n19497) );
  NAND2_X1 U19203 ( .A1(n19497), .A2(n17309), .ZN(n17242) );
  OAI21_X1 U19204 ( .B1(n17309), .B2(n17243), .A(n17242), .ZN(P2_U2856) );
  INV_X1 U19205 ( .A(n17244), .ZN(n17251) );
  NOR2_X1 U19206 ( .A1(n17251), .A2(n17245), .ZN(n17247) );
  XNOR2_X1 U19207 ( .A(n17247), .B(n17246), .ZN(n17322) );
  NAND2_X1 U19208 ( .A1(n17322), .A2(n17303), .ZN(n17249) );
  NAND2_X1 U19209 ( .A1(n15680), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n17248) );
  OAI211_X1 U19210 ( .C1(n19468), .C2(n15680), .A(n17249), .B(n17248), .ZN(
        P2_U2859) );
  NOR2_X1 U19211 ( .A1(n17250), .A2(n17251), .ZN(n17253) );
  XNOR2_X1 U19212 ( .A(n17253), .B(n17252), .ZN(n17324) );
  NAND2_X1 U19213 ( .A1(n17324), .A2(n17303), .ZN(n17255) );
  NAND2_X1 U19214 ( .A1(n15680), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n17254) );
  OAI211_X1 U19215 ( .C1(n15680), .C2(n17672), .A(n17255), .B(n17254), .ZN(
        P2_U2860) );
  OAI21_X1 U19216 ( .B1(n17256), .B2(n17258), .A(n17257), .ZN(n17339) );
  NAND2_X1 U19217 ( .A1(n15680), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n17264) );
  NAND2_X1 U19218 ( .A1(n17259), .A2(n17260), .ZN(n17261) );
  NAND2_X1 U19219 ( .A1(n19450), .A2(n17309), .ZN(n17263) );
  OAI211_X1 U19220 ( .C1(n17339), .C2(n17316), .A(n17264), .B(n17263), .ZN(
        P2_U2861) );
  OAI21_X1 U19221 ( .B1(n17273), .B2(n17265), .A(n17259), .ZN(n19437) );
  AOI21_X1 U19222 ( .B1(n17266), .B2(n17268), .A(n17267), .ZN(n17343) );
  NAND2_X1 U19223 ( .A1(n17343), .A2(n17303), .ZN(n17270) );
  NAND2_X1 U19224 ( .A1(n15680), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n17269) );
  OAI211_X1 U19225 ( .C1(n19437), .C2(n15680), .A(n17270), .B(n17269), .ZN(
        P2_U2862) );
  NOR2_X1 U19226 ( .A1(n17282), .A2(n17271), .ZN(n17272) );
  OR2_X1 U19227 ( .A1(n17273), .A2(n17272), .ZN(n17712) );
  AOI21_X1 U19228 ( .B1(n17274), .B2(n17276), .A(n17275), .ZN(n17352) );
  NAND2_X1 U19229 ( .A1(n17352), .A2(n17303), .ZN(n17278) );
  NAND2_X1 U19230 ( .A1(n15680), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n17277) );
  OAI211_X1 U19231 ( .C1(n17712), .C2(n15680), .A(n17278), .B(n17277), .ZN(
        P2_U2863) );
  XNOR2_X1 U19232 ( .A(n17279), .B(n17280), .ZN(n17361) );
  AND2_X1 U19233 ( .A1(n17292), .A2(n17281), .ZN(n17283) );
  OR2_X1 U19234 ( .A1(n17283), .A2(n17282), .ZN(n19417) );
  NOR2_X1 U19235 ( .A1(n19417), .A2(n15680), .ZN(n17284) );
  AOI21_X1 U19236 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n15680), .A(n17284), .ZN(
        n17285) );
  OAI21_X1 U19237 ( .B1(n17361), .B2(n17316), .A(n17285), .ZN(P2_U2864) );
  AOI21_X1 U19238 ( .B1(n17288), .B2(n17287), .A(n17279), .ZN(n17379) );
  NAND2_X1 U19239 ( .A1(n17379), .A2(n17303), .ZN(n17294) );
  NAND2_X1 U19240 ( .A1(n17290), .A2(n17289), .ZN(n17291) );
  NAND2_X1 U19241 ( .A1(n19404), .A2(n17309), .ZN(n17293) );
  OAI211_X1 U19242 ( .C1(n17309), .C2(n12172), .A(n17294), .B(n17293), .ZN(
        P2_U2865) );
  OAI21_X1 U19243 ( .B1(n17295), .B2(n17296), .A(n17287), .ZN(n17388) );
  NOR2_X1 U19244 ( .A1(n17297), .A2(n15680), .ZN(n17298) );
  AOI21_X1 U19245 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n15680), .A(n17298), .ZN(
        n17299) );
  OAI21_X1 U19246 ( .B1(n17388), .B2(n17316), .A(n17299), .ZN(P2_U2866) );
  INV_X1 U19247 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n19388) );
  AOI21_X1 U19248 ( .B1(n17302), .B2(n17301), .A(n17295), .ZN(n17397) );
  NAND2_X1 U19249 ( .A1(n17397), .A2(n17303), .ZN(n17308) );
  AOI21_X1 U19250 ( .B1(n17306), .B2(n17304), .A(n17305), .ZN(n19391) );
  NAND2_X1 U19251 ( .A1(n19391), .A2(n17309), .ZN(n17307) );
  OAI211_X1 U19252 ( .C1(n17309), .C2(n19388), .A(n17308), .B(n17307), .ZN(
        P2_U2867) );
  OAI21_X1 U19253 ( .B1(n15918), .B2(n17310), .A(n17301), .ZN(n17410) );
  NAND2_X1 U19254 ( .A1(n17312), .A2(n17311), .ZN(n17313) );
  NAND2_X1 U19255 ( .A1(n17304), .A2(n17313), .ZN(n19378) );
  NOR2_X1 U19256 ( .A1(n19378), .A2(n15680), .ZN(n17314) );
  AOI21_X1 U19257 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15680), .A(n17314), .ZN(
        n17315) );
  OAI21_X1 U19258 ( .B1(n17410), .B2(n17316), .A(n17315), .ZN(P2_U2868) );
  OAI22_X1 U19259 ( .A1(n17404), .A2(n20062), .B1(n20546), .B2(n17317), .ZN(
        n17318) );
  AOI21_X1 U19260 ( .B1(n20048), .B2(BUF2_REG_28__SCAN_IN), .A(n17318), .ZN(
        n17320) );
  NAND2_X1 U19261 ( .A1(n20050), .A2(BUF1_REG_28__SCAN_IN), .ZN(n17319) );
  OAI211_X1 U19262 ( .C1(n19476), .C2(n20548), .A(n17320), .B(n17319), .ZN(
        n17321) );
  AOI21_X1 U19263 ( .B1(n17322), .B2(n20551), .A(n17321), .ZN(n17323) );
  INV_X1 U19264 ( .A(n17323), .ZN(P2_U2891) );
  NAND2_X1 U19265 ( .A1(n17324), .A2(n20551), .ZN(n17329) );
  INV_X1 U19266 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n17326) );
  INV_X1 U19267 ( .A(n20546), .ZN(n20495) );
  AOI22_X1 U19268 ( .A1(n17344), .A2(n20065), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n20495), .ZN(n17325) );
  OAI21_X1 U19269 ( .B1(n17355), .B2(n17326), .A(n17325), .ZN(n17327) );
  AOI21_X1 U19270 ( .B1(n20050), .B2(BUF1_REG_27__SCAN_IN), .A(n17327), .ZN(
        n17328) );
  OAI211_X1 U19271 ( .C1(n20548), .C2(n17680), .A(n17329), .B(n17328), .ZN(
        P2_U2892) );
  NAND2_X1 U19272 ( .A1(n17330), .A2(n17331), .ZN(n17332) );
  NAND2_X1 U19273 ( .A1(n11264), .A2(n17332), .ZN(n19452) );
  OAI22_X1 U19274 ( .A1(n17404), .A2(n20071), .B1(n20546), .B2(n17333), .ZN(
        n17334) );
  AOI21_X1 U19275 ( .B1(n20048), .B2(BUF2_REG_26__SCAN_IN), .A(n17334), .ZN(
        n17336) );
  NAND2_X1 U19276 ( .A1(n20050), .A2(BUF1_REG_26__SCAN_IN), .ZN(n17335) );
  OAI211_X1 U19277 ( .C1(n19452), .C2(n20548), .A(n17336), .B(n17335), .ZN(
        n17337) );
  INV_X1 U19278 ( .A(n17337), .ZN(n17338) );
  OAI21_X1 U19279 ( .B1(n17339), .B2(n20405), .A(n17338), .ZN(P2_U2893) );
  OR2_X1 U19280 ( .A1(n17341), .A2(n17340), .ZN(n17342) );
  AND2_X1 U19281 ( .A1(n17330), .A2(n17342), .ZN(n19439) );
  INV_X1 U19282 ( .A(n19439), .ZN(n17350) );
  NAND2_X1 U19283 ( .A1(n17343), .A2(n20551), .ZN(n17349) );
  INV_X1 U19284 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U19285 ( .A1(n17344), .A2(n20073), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n20495), .ZN(n17345) );
  OAI21_X1 U19286 ( .B1(n17355), .B2(n17346), .A(n17345), .ZN(n17347) );
  AOI21_X1 U19287 ( .B1(n20050), .B2(BUF1_REG_25__SCAN_IN), .A(n17347), .ZN(
        n17348) );
  OAI211_X1 U19288 ( .C1(n17350), .C2(n20548), .A(n17349), .B(n17348), .ZN(
        P2_U2894) );
  XOR2_X1 U19289 ( .A(n17351), .B(n11265), .Z(n19429) );
  INV_X1 U19290 ( .A(n19429), .ZN(n17360) );
  NAND2_X1 U19291 ( .A1(n17352), .A2(n20551), .ZN(n17359) );
  OAI22_X1 U19292 ( .A1(n17404), .A2(n20077), .B1(n17353), .B2(n20546), .ZN(
        n17357) );
  INV_X1 U19293 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17354) );
  NOR2_X1 U19294 ( .A1(n17355), .A2(n17354), .ZN(n17356) );
  AOI211_X1 U19295 ( .C1(BUF1_REG_24__SCAN_IN), .C2(n20050), .A(n17357), .B(
        n17356), .ZN(n17358) );
  OAI211_X1 U19296 ( .C1(n17360), .C2(n20548), .A(n17359), .B(n17358), .ZN(
        P2_U2895) );
  OR2_X1 U19297 ( .A1(n17361), .A2(n20405), .ZN(n17370) );
  OAI22_X1 U19298 ( .A1(n17404), .A2(n20085), .B1(n20546), .B2(n17362), .ZN(
        n17363) );
  AOI21_X1 U19299 ( .B1(n20048), .B2(BUF2_REG_23__SCAN_IN), .A(n17363), .ZN(
        n17369) );
  NAND2_X1 U19300 ( .A1(n17364), .A2(n17365), .ZN(n17366) );
  AND2_X1 U19301 ( .A1(n11265), .A2(n17366), .ZN(n19419) );
  NAND2_X1 U19302 ( .A1(n19419), .A2(n20497), .ZN(n17368) );
  NAND2_X1 U19303 ( .A1(n20050), .A2(BUF1_REG_23__SCAN_IN), .ZN(n17367) );
  NAND4_X1 U19304 ( .A1(n17370), .A2(n17369), .A3(n17368), .A4(n17367), .ZN(
        P2_U2896) );
  OR2_X1 U19305 ( .A1(n17372), .A2(n17371), .ZN(n17373) );
  NAND2_X1 U19306 ( .A1(n17364), .A2(n17373), .ZN(n19415) );
  OAI22_X1 U19307 ( .A1(n17404), .A2(n20271), .B1(n17374), .B2(n20546), .ZN(
        n17375) );
  AOI21_X1 U19308 ( .B1(n20048), .B2(BUF2_REG_22__SCAN_IN), .A(n17375), .ZN(
        n17377) );
  NAND2_X1 U19309 ( .A1(n20050), .A2(BUF1_REG_22__SCAN_IN), .ZN(n17376) );
  OAI211_X1 U19310 ( .C1(n19415), .C2(n20548), .A(n17377), .B(n17376), .ZN(
        n17378) );
  AOI21_X1 U19311 ( .B1(n17379), .B2(n20551), .A(n17378), .ZN(n17380) );
  INV_X1 U19312 ( .A(n17380), .ZN(P2_U2897) );
  OAI22_X1 U19313 ( .A1(n17404), .A2(n20320), .B1(n20546), .B2(n17381), .ZN(
        n17382) );
  AOI21_X1 U19314 ( .B1(n20048), .B2(BUF2_REG_21__SCAN_IN), .A(n17382), .ZN(
        n17384) );
  NAND2_X1 U19315 ( .A1(n20050), .A2(BUF1_REG_21__SCAN_IN), .ZN(n17383) );
  OAI211_X1 U19316 ( .C1(n17385), .C2(n20548), .A(n17384), .B(n17383), .ZN(
        n17386) );
  INV_X1 U19317 ( .A(n17386), .ZN(n17387) );
  OAI21_X1 U19318 ( .B1(n17388), .B2(n20405), .A(n17387), .ZN(P2_U2898) );
  NAND2_X1 U19319 ( .A1(n17402), .A2(n17389), .ZN(n17390) );
  NAND2_X1 U19320 ( .A1(n17391), .A2(n17390), .ZN(n19403) );
  OAI22_X1 U19321 ( .A1(n17404), .A2(n20361), .B1(n20546), .B2(n17392), .ZN(
        n17393) );
  AOI21_X1 U19322 ( .B1(n20048), .B2(BUF2_REG_20__SCAN_IN), .A(n17393), .ZN(
        n17395) );
  NAND2_X1 U19323 ( .A1(n20050), .A2(BUF1_REG_20__SCAN_IN), .ZN(n17394) );
  OAI211_X1 U19324 ( .C1(n19403), .C2(n20548), .A(n17395), .B(n17394), .ZN(
        n17396) );
  AOI21_X1 U19325 ( .B1(n17397), .B2(n20551), .A(n17396), .ZN(n17398) );
  INV_X1 U19326 ( .A(n17398), .ZN(P2_U2899) );
  NAND2_X1 U19327 ( .A1(n17400), .A2(n17399), .ZN(n17401) );
  NAND2_X1 U19328 ( .A1(n17402), .A2(n17401), .ZN(n19385) );
  OAI22_X1 U19329 ( .A1(n17404), .A2(n20409), .B1(n20546), .B2(n17403), .ZN(
        n17405) );
  AOI21_X1 U19330 ( .B1(n20048), .B2(BUF2_REG_19__SCAN_IN), .A(n17405), .ZN(
        n17407) );
  NAND2_X1 U19331 ( .A1(n20050), .A2(BUF1_REG_19__SCAN_IN), .ZN(n17406) );
  OAI211_X1 U19332 ( .C1(n19385), .C2(n20548), .A(n17407), .B(n17406), .ZN(
        n17408) );
  INV_X1 U19333 ( .A(n17408), .ZN(n17409) );
  OAI21_X1 U19334 ( .B1(n17410), .B2(n20405), .A(n17409), .ZN(P2_U2900) );
  NOR2_X1 U19335 ( .A1(n17638), .A2(n17411), .ZN(n17412) );
  AOI211_X1 U19336 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n17612), .A(
        n17413), .B(n17412), .ZN(n17414) );
  OAI21_X1 U19337 ( .B1(n17241), .B2(n17641), .A(n17414), .ZN(n17415) );
  AOI21_X1 U19338 ( .B1(n17416), .B2(n18086), .A(n17415), .ZN(n17417) );
  OAI21_X1 U19339 ( .B1(n17418), .B2(n18065), .A(n17417), .ZN(P2_U2983) );
  NAND2_X1 U19340 ( .A1(n17419), .A2(n17432), .ZN(n17424) );
  INV_X1 U19341 ( .A(n17420), .ZN(n17421) );
  NOR2_X1 U19342 ( .A1(n17422), .A2(n17421), .ZN(n17423) );
  INV_X1 U19343 ( .A(n17435), .ZN(n17426) );
  AOI21_X1 U19344 ( .B1(n17426), .B2(n17645), .A(n17425), .ZN(n17655) );
  NOR2_X1 U19345 ( .A1(n17651), .A2(n17641), .ZN(n17429) );
  NAND2_X1 U19346 ( .A1(n19526), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n17650) );
  NAND2_X1 U19347 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17427) );
  OAI211_X1 U19348 ( .C1(n17638), .C2(n19500), .A(n17650), .B(n17427), .ZN(
        n17428) );
  AOI211_X1 U19349 ( .C1(n17655), .C2(n18086), .A(n17429), .B(n17428), .ZN(
        n17430) );
  NAND2_X1 U19350 ( .A1(n17432), .A2(n17431), .ZN(n17434) );
  XOR2_X1 U19351 ( .A(n17434), .B(n17433), .Z(n17671) );
  AOI21_X1 U19352 ( .B1(n17444), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17436) );
  NAND2_X1 U19353 ( .A1(n19526), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n17666) );
  OAI21_X1 U19354 ( .B1(n18093), .B2(n17437), .A(n17666), .ZN(n17438) );
  AOI21_X1 U19355 ( .B1(n18083), .B2(n17439), .A(n17438), .ZN(n17440) );
  OAI21_X1 U19356 ( .B1(n19480), .B2(n17641), .A(n17440), .ZN(n17441) );
  AOI21_X1 U19357 ( .B1(n17669), .B2(n18086), .A(n17441), .ZN(n17442) );
  OAI21_X1 U19358 ( .B1(n17671), .B2(n18065), .A(n17442), .ZN(P2_U2985) );
  XNOR2_X1 U19359 ( .A(n17443), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17684) );
  AOI21_X1 U19360 ( .B1(n15995), .B2(n17459), .A(n17444), .ZN(n17682) );
  NOR2_X1 U19361 ( .A1(n19301), .A2(n17445), .ZN(n17673) );
  NOR2_X1 U19362 ( .A1(n17638), .A2(n17446), .ZN(n17447) );
  AOI211_X1 U19363 ( .C1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17612), .A(
        n17673), .B(n17447), .ZN(n17448) );
  OAI21_X1 U19364 ( .B1(n17672), .B2(n17641), .A(n17448), .ZN(n17449) );
  AOI21_X1 U19365 ( .B1(n17682), .B2(n18086), .A(n17449), .ZN(n17450) );
  OAI21_X1 U19366 ( .B1(n17684), .B2(n18065), .A(n17450), .ZN(P2_U2987) );
  AOI21_X1 U19368 ( .B1(n17452), .B2(n17464), .A(n17466), .ZN(n17454) );
  MUX2_X1 U19369 ( .A(n17464), .B(n17454), .S(n17453), .Z(n17455) );
  NAND2_X1 U19370 ( .A1(n17456), .A2(n17455), .ZN(n17695) );
  NAND2_X1 U19371 ( .A1(n19526), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n17687) );
  NAND2_X1 U19372 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17457) );
  OAI211_X1 U19373 ( .C1(n17638), .C2(n19455), .A(n17687), .B(n17457), .ZN(
        n17461) );
  OAI21_X1 U19374 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17458), .A(
        n17459), .ZN(n17692) );
  NOR2_X1 U19375 ( .A1(n17692), .A2(n18063), .ZN(n17460) );
  OAI21_X1 U19376 ( .B1(n17695), .B2(n18065), .A(n17462), .ZN(P2_U2988) );
  INV_X1 U19377 ( .A(n17458), .ZN(n17463) );
  OAI21_X1 U19378 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17477), .A(
        n17463), .ZN(n17706) );
  INV_X1 U19379 ( .A(n17464), .ZN(n17465) );
  NOR2_X1 U19380 ( .A1(n17466), .A2(n17465), .ZN(n17467) );
  XNOR2_X1 U19381 ( .A(n17452), .B(n17467), .ZN(n17696) );
  NAND2_X1 U19382 ( .A1(n17696), .A2(n18089), .ZN(n17472) );
  NAND2_X1 U19383 ( .A1(n19526), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17697) );
  OAI21_X1 U19384 ( .B1(n18093), .B2(n17468), .A(n17697), .ZN(n17470) );
  NOR2_X1 U19385 ( .A1(n19437), .A2(n17641), .ZN(n17469) );
  AOI211_X1 U19386 ( .C1(n18083), .C2(n19440), .A(n17470), .B(n17469), .ZN(
        n17471) );
  OAI211_X1 U19387 ( .C1(n18063), .C2(n17706), .A(n17472), .B(n17471), .ZN(
        P2_U2989) );
  NOR2_X1 U19388 ( .A1(n17474), .A2(n11330), .ZN(n17475) );
  XNOR2_X1 U19389 ( .A(n17473), .B(n17475), .ZN(n17717) );
  INV_X1 U19390 ( .A(n17712), .ZN(n19428) );
  NAND2_X1 U19391 ( .A1(n19526), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n17711) );
  NAND2_X1 U19392 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17476) );
  OAI211_X1 U19393 ( .C1(n17638), .C2(n19431), .A(n17711), .B(n17476), .ZN(
        n17482) );
  INV_X1 U19394 ( .A(n17477), .ZN(n17480) );
  NAND2_X1 U19395 ( .A1(n17478), .A2(n17707), .ZN(n17479) );
  NAND2_X1 U19396 ( .A1(n17480), .A2(n17479), .ZN(n17713) );
  NOR2_X1 U19397 ( .A1(n17713), .A2(n18063), .ZN(n17481) );
  AOI211_X1 U19398 ( .C1(n19428), .C2(n18088), .A(n17482), .B(n17481), .ZN(
        n17483) );
  OAI21_X1 U19399 ( .B1(n17717), .B2(n18065), .A(n17483), .ZN(P2_U2990) );
  NOR2_X1 U19400 ( .A1(n17500), .A2(n17731), .ZN(n17499) );
  OAI21_X1 U19401 ( .B1(n17499), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17478), .ZN(n17727) );
  NOR2_X1 U19402 ( .A1(n11327), .A2(n17485), .ZN(n17486) );
  XNOR2_X1 U19403 ( .A(n17484), .B(n17486), .ZN(n17718) );
  NAND2_X1 U19404 ( .A1(n17718), .A2(n18089), .ZN(n17492) );
  NAND2_X1 U19405 ( .A1(n19526), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17721) );
  OAI21_X1 U19406 ( .B1(n18093), .B2(n17487), .A(n17721), .ZN(n17489) );
  NOR2_X1 U19407 ( .A1(n19417), .A2(n17641), .ZN(n17488) );
  AOI211_X1 U19408 ( .C1(n18083), .C2(n17490), .A(n17489), .B(n17488), .ZN(
        n17491) );
  OAI211_X1 U19409 ( .C1(n18063), .C2(n17727), .A(n17492), .B(n17491), .ZN(
        P2_U2991) );
  NOR2_X1 U19410 ( .A1(n17494), .A2(n11331), .ZN(n17495) );
  XNOR2_X1 U19411 ( .A(n17493), .B(n17495), .ZN(n17740) );
  NOR2_X1 U19412 ( .A1(n19301), .A2(n17496), .ZN(n17728) );
  AOI21_X1 U19413 ( .B1(n17612), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17728), .ZN(n17497) );
  OAI21_X1 U19414 ( .B1(n17638), .B2(n19412), .A(n17497), .ZN(n17498) );
  AOI21_X1 U19415 ( .B1(n19404), .B2(n18088), .A(n17498), .ZN(n17502) );
  INV_X1 U19416 ( .A(n17499), .ZN(n17737) );
  NAND2_X1 U19417 ( .A1(n17500), .A2(n17731), .ZN(n17736) );
  NAND3_X1 U19418 ( .A1(n17737), .A2(n18086), .A3(n17736), .ZN(n17501) );
  OAI211_X1 U19419 ( .C1(n17740), .C2(n18065), .A(n17502), .B(n17501), .ZN(
        P2_U2992) );
  XNOR2_X1 U19420 ( .A(n17503), .B(n17753), .ZN(n17759) );
  NAND2_X1 U19421 ( .A1(n19526), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n17752) );
  NAND2_X1 U19422 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17504) );
  OAI211_X1 U19423 ( .C1(n19397), .C2(n17638), .A(n17752), .B(n17504), .ZN(
        n17505) );
  AOI21_X1 U19424 ( .B1(n19391), .B2(n18088), .A(n17505), .ZN(n17509) );
  INV_X1 U19425 ( .A(n17749), .ZN(n17506) );
  NAND2_X1 U19426 ( .A1(n17543), .A2(n17506), .ZN(n17516) );
  AOI21_X1 U19427 ( .B1(n17516), .B2(n17753), .A(n17507), .ZN(n17757) );
  NAND2_X1 U19428 ( .A1(n17757), .A2(n18086), .ZN(n17508) );
  OAI211_X1 U19429 ( .C1(n17759), .C2(n18065), .A(n17509), .B(n17508), .ZN(
        P2_U2994) );
  NAND2_X1 U19430 ( .A1(n17511), .A2(n17510), .ZN(n17515) );
  INV_X1 U19431 ( .A(n17529), .ZN(n17513) );
  NOR2_X1 U19432 ( .A1(n17512), .A2(n17513), .ZN(n17514) );
  XOR2_X1 U19433 ( .A(n17515), .B(n17514), .Z(n17772) );
  INV_X1 U19434 ( .A(n17516), .ZN(n17518) );
  AOI21_X1 U19435 ( .B1(n17543), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17517) );
  NOR2_X1 U19436 ( .A1(n17518), .A2(n17517), .ZN(n17769) );
  INV_X1 U19437 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n17519) );
  NOR2_X1 U19438 ( .A1(n19301), .A2(n17519), .ZN(n17761) );
  NOR2_X1 U19439 ( .A1(n18093), .A2(n19375), .ZN(n17520) );
  AOI211_X1 U19440 ( .C1(n19379), .C2(n18083), .A(n17761), .B(n17520), .ZN(
        n17521) );
  OAI21_X1 U19441 ( .B1(n19378), .B2(n17641), .A(n17521), .ZN(n17522) );
  AOI21_X1 U19442 ( .B1(n17769), .B2(n18086), .A(n17522), .ZN(n17523) );
  OAI21_X1 U19443 ( .B1(n17772), .B2(n18065), .A(n17523), .ZN(P2_U2995) );
  XNOR2_X1 U19444 ( .A(n17543), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17782) );
  NOR2_X1 U19445 ( .A1(n19301), .A2(n19365), .ZN(n17774) );
  AOI21_X1 U19446 ( .B1(n17612), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17774), .ZN(n17524) );
  OAI21_X1 U19447 ( .B1(n17638), .B2(n17525), .A(n17524), .ZN(n17531) );
  AOI21_X1 U19448 ( .B1(n17529), .B2(n17527), .A(n17526), .ZN(n17528) );
  AOI21_X1 U19449 ( .B1(n17512), .B2(n17529), .A(n17528), .ZN(n17773) );
  NOR2_X1 U19450 ( .A1(n17773), .A2(n18065), .ZN(n17530) );
  AOI211_X1 U19451 ( .C1(n18088), .C2(n19367), .A(n17531), .B(n17530), .ZN(
        n17532) );
  OAI21_X1 U19452 ( .B1(n18063), .B2(n17782), .A(n17532), .ZN(P2_U2996) );
  NAND2_X1 U19453 ( .A1(n17534), .A2(n17533), .ZN(n17539) );
  INV_X1 U19454 ( .A(n17535), .ZN(n17537) );
  NAND2_X1 U19455 ( .A1(n17537), .A2(n17536), .ZN(n17538) );
  XOR2_X1 U19456 ( .A(n17539), .B(n17538), .Z(n17802) );
  NAND2_X1 U19457 ( .A1(n17540), .A2(n18083), .ZN(n17541) );
  NAND2_X1 U19458 ( .A1(n19526), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17792) );
  OAI211_X1 U19459 ( .C1(n17542), .C2(n18093), .A(n17541), .B(n17792), .ZN(
        n17546) );
  AOI211_X1 U19460 ( .C1(n17544), .C2(n11229), .A(n18063), .B(n17543), .ZN(
        n17545) );
  OAI21_X1 U19461 ( .B1(n17802), .B2(n18065), .A(n17547), .ZN(P2_U2997) );
  INV_X1 U19462 ( .A(n17804), .ZN(n19356) );
  INV_X1 U19463 ( .A(n19352), .ZN(n17549) );
  NAND2_X1 U19464 ( .A1(n19526), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17803) );
  NAND2_X1 U19465 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17548) );
  OAI211_X1 U19466 ( .C1(n17638), .C2(n17549), .A(n17803), .B(n17548), .ZN(
        n17553) );
  NOR2_X1 U19467 ( .A1(n17551), .A2(n17550), .ZN(n17805) );
  NOR3_X1 U19468 ( .A1(n17805), .A2(n17535), .A3(n18065), .ZN(n17552) );
  AOI211_X1 U19469 ( .C1(n19356), .C2(n18088), .A(n17553), .B(n17552), .ZN(
        n17555) );
  OAI211_X1 U19470 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17826), .A(
        n11229), .B(n18086), .ZN(n17554) );
  NAND2_X1 U19471 ( .A1(n17555), .A2(n17554), .ZN(P2_U2998) );
  INV_X1 U19472 ( .A(n17595), .ZN(n17557) );
  NOR2_X1 U19473 ( .A1(n17556), .A2(n17557), .ZN(n17586) );
  INV_X1 U19474 ( .A(n17583), .ZN(n17558) );
  OAI21_X1 U19475 ( .B1(n17586), .B2(n17558), .A(n17584), .ZN(n17575) );
  AND2_X1 U19476 ( .A1(n17560), .A2(n17559), .ZN(n17574) );
  NAND2_X1 U19477 ( .A1(n17575), .A2(n17574), .ZN(n17573) );
  NAND2_X1 U19478 ( .A1(n17573), .A2(n17560), .ZN(n17564) );
  NAND2_X1 U19479 ( .A1(n17562), .A2(n17561), .ZN(n17563) );
  XNOR2_X1 U19480 ( .A(n17564), .B(n17563), .ZN(n17831) );
  NAND2_X1 U19481 ( .A1(n19526), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n17819) );
  NAND2_X1 U19482 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17565) );
  OAI211_X1 U19483 ( .C1(n17638), .C2(n17566), .A(n17819), .B(n17565), .ZN(
        n17569) );
  NOR2_X1 U19484 ( .A1(n17567), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17827) );
  NOR3_X1 U19485 ( .A1(n17827), .A2(n17826), .A3(n18063), .ZN(n17568) );
  AOI211_X1 U19486 ( .C1(n18088), .C2(n19343), .A(n17569), .B(n17568), .ZN(
        n17570) );
  OAI21_X1 U19487 ( .B1(n17831), .B2(n18065), .A(n17570), .ZN(P2_U2999) );
  INV_X1 U19488 ( .A(n17581), .ZN(n17572) );
  OAI21_X1 U19489 ( .B1(n17572), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17795), .ZN(n17846) );
  OAI21_X1 U19490 ( .B1(n17575), .B2(n17574), .A(n17573), .ZN(n17832) );
  NAND2_X1 U19491 ( .A1(n17832), .A2(n18089), .ZN(n17579) );
  NAND2_X1 U19492 ( .A1(n19526), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n17838) );
  NAND2_X1 U19493 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17576) );
  OAI211_X1 U19494 ( .C1(n17638), .C2(n19332), .A(n17838), .B(n17576), .ZN(
        n17577) );
  AOI21_X1 U19495 ( .B1(n19331), .B2(n18088), .A(n17577), .ZN(n17578) );
  OAI211_X1 U19496 ( .C1(n18063), .C2(n17846), .A(n17579), .B(n17578), .ZN(
        P2_U3000) );
  NAND2_X1 U19497 ( .A1(n17580), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17902) );
  NAND2_X1 U19498 ( .A1(n17893), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17600) );
  OAI21_X1 U19499 ( .B1(n17600), .B2(n17865), .A(n17847), .ZN(n17582) );
  NAND2_X1 U19500 ( .A1(n17582), .A2(n17581), .ZN(n17859) );
  NAND2_X1 U19501 ( .A1(n17584), .A2(n17583), .ZN(n17585) );
  XNOR2_X1 U19502 ( .A(n17586), .B(n17585), .ZN(n17857) );
  NOR2_X1 U19503 ( .A1(n17851), .A2(n17641), .ZN(n17590) );
  NAND2_X1 U19504 ( .A1(n19526), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n17850) );
  NAND2_X1 U19505 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17587) );
  OAI211_X1 U19506 ( .C1(n17638), .C2(n17588), .A(n17850), .B(n17587), .ZN(
        n17589) );
  AOI211_X1 U19507 ( .C1(n17857), .C2(n18089), .A(n17590), .B(n17589), .ZN(
        n17591) );
  OAI21_X1 U19508 ( .B1(n18063), .B2(n17859), .A(n17591), .ZN(P2_U3001) );
  XNOR2_X1 U19509 ( .A(n17600), .B(n17865), .ZN(n17872) );
  NAND2_X1 U19510 ( .A1(n18083), .A2(n19319), .ZN(n17592) );
  NAND2_X1 U19511 ( .A1(n19526), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17861) );
  OAI211_X1 U19512 ( .C1(n19313), .C2(n18093), .A(n17592), .B(n17861), .ZN(
        n17598) );
  NAND2_X1 U19513 ( .A1(n17595), .A2(n17594), .ZN(n17596) );
  XNOR2_X1 U19514 ( .A(n17593), .B(n17596), .ZN(n17867) );
  NOR2_X1 U19515 ( .A1(n17867), .A2(n18065), .ZN(n17597) );
  AOI211_X1 U19516 ( .C1(n18088), .C2(n19321), .A(n17598), .B(n17597), .ZN(
        n17599) );
  OAI21_X1 U19517 ( .B1(n18063), .B2(n17872), .A(n17599), .ZN(P2_U3002) );
  OAI21_X1 U19518 ( .B1(n17893), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17600), .ZN(n17885) );
  XOR2_X1 U19519 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17602), .Z(
        n17603) );
  XNOR2_X1 U19520 ( .A(n17601), .B(n17603), .ZN(n17883) );
  NOR2_X1 U19521 ( .A1(n17641), .A2(n19306), .ZN(n17606) );
  NAND2_X1 U19522 ( .A1(n19526), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n17876) );
  NAND2_X1 U19523 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17604) );
  OAI211_X1 U19524 ( .C1(n17638), .C2(n19312), .A(n17876), .B(n17604), .ZN(
        n17605) );
  AOI211_X1 U19525 ( .C1(n17883), .C2(n18089), .A(n17606), .B(n17605), .ZN(
        n17607) );
  OAI21_X1 U19526 ( .B1(n17885), .B2(n18063), .A(n17607), .ZN(P2_U3003) );
  INV_X1 U19527 ( .A(n17886), .ZN(n17608) );
  NOR2_X1 U19528 ( .A1(n17609), .A2(n17608), .ZN(n17611) );
  XOR2_X1 U19529 ( .A(n17611), .B(n17610), .Z(n17914) );
  OR2_X1 U19530 ( .A1(n17580), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17903) );
  NAND3_X1 U19531 ( .A1(n17903), .A2(n17902), .A3(n18086), .ZN(n17617) );
  NAND2_X1 U19532 ( .A1(n19526), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n17907) );
  NAND2_X1 U19533 ( .A1(n17612), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17613) );
  OAI211_X1 U19534 ( .C1(n17638), .C2(n17614), .A(n17907), .B(n17613), .ZN(
        n17615) );
  AOI21_X1 U19535 ( .B1(n18088), .B2(n17906), .A(n17615), .ZN(n17616) );
  OAI211_X1 U19536 ( .C1(n18065), .C2(n17914), .A(n17617), .B(n17616), .ZN(
        P2_U3005) );
  NAND2_X1 U19537 ( .A1(n17620), .A2(n17619), .ZN(n17621) );
  XNOR2_X1 U19538 ( .A(n17618), .B(n17621), .ZN(n17932) );
  OR2_X1 U19539 ( .A1(n17623), .A2(n17622), .ZN(n17915) );
  NAND3_X1 U19540 ( .A1(n17915), .A2(n17624), .A3(n18086), .ZN(n17630) );
  NOR2_X1 U19541 ( .A1(n17641), .A2(n19294), .ZN(n17628) );
  INV_X1 U19542 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n17625) );
  OAI22_X1 U19543 ( .A1(n17626), .A2(n18093), .B1(n17625), .B2(n19301), .ZN(
        n17627) );
  AOI211_X1 U19544 ( .C1(n18083), .C2(n19293), .A(n17628), .B(n17627), .ZN(
        n17629) );
  OAI211_X1 U19545 ( .C1(n18065), .C2(n17932), .A(n17630), .B(n17629), .ZN(
        P2_U3006) );
  NAND2_X1 U19546 ( .A1(n17632), .A2(n17631), .ZN(n17634) );
  XOR2_X1 U19547 ( .A(n17634), .B(n11230), .Z(n17945) );
  NAND2_X1 U19548 ( .A1(n11352), .A2(n17636), .ZN(n17637) );
  XNOR2_X1 U19549 ( .A(n17635), .B(n17637), .ZN(n17942) );
  INV_X1 U19550 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17639) );
  OAI22_X1 U19551 ( .A1(n17639), .A2(n18093), .B1(n17638), .B2(n19280), .ZN(
        n17643) );
  OAI22_X1 U19552 ( .A1(n17641), .A2(n19283), .B1(n17640), .B2(n19301), .ZN(
        n17642) );
  AOI211_X1 U19553 ( .C1(n17942), .C2(n18089), .A(n17643), .B(n17642), .ZN(
        n17644) );
  OAI21_X1 U19554 ( .B1(n17945), .B2(n18063), .A(n17644), .ZN(P2_U3007) );
  OAI21_X1 U19555 ( .B1(n17661), .B2(n17646), .A(n17645), .ZN(n17647) );
  NAND2_X1 U19556 ( .A1(n17648), .A2(n17647), .ZN(n17649) );
  OAI211_X1 U19557 ( .C1(n17651), .C2(n19514), .A(n17650), .B(n17649), .ZN(
        n17654) );
  NOR2_X1 U19558 ( .A1(n17652), .A2(n19542), .ZN(n17653) );
  AOI211_X1 U19559 ( .C1(n17655), .C2(n19537), .A(n17654), .B(n17653), .ZN(
        n17656) );
  NOR2_X1 U19560 ( .A1(n19479), .A2(n19542), .ZN(n17668) );
  NOR2_X1 U19561 ( .A1(n17658), .A2(n17657), .ZN(n17663) );
  INV_X1 U19562 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17660) );
  OAI21_X1 U19563 ( .B1(n17661), .B2(n17660), .A(n17659), .ZN(n17662) );
  OAI21_X1 U19564 ( .B1(n17664), .B2(n17663), .A(n17662), .ZN(n17665) );
  OAI211_X1 U19565 ( .C1(n19480), .C2(n19514), .A(n17666), .B(n17665), .ZN(
        n17667) );
  OAI21_X1 U19566 ( .B1(n17671), .B2(n19546), .A(n17670), .ZN(P2_U3017) );
  INV_X1 U19567 ( .A(n17672), .ZN(n17678) );
  INV_X1 U19568 ( .A(n17673), .ZN(n17674) );
  OAI211_X1 U19569 ( .C1(n17676), .C2(n15995), .A(n17675), .B(n17674), .ZN(
        n17677) );
  AOI21_X1 U19570 ( .B1(n17678), .B2(n19550), .A(n17677), .ZN(n17679) );
  OAI21_X1 U19571 ( .B1(n17680), .B2(n19542), .A(n17679), .ZN(n17681) );
  AOI21_X1 U19572 ( .B1(n17682), .B2(n19537), .A(n17681), .ZN(n17683) );
  OAI21_X1 U19573 ( .B1(n17684), .B2(n19546), .A(n17683), .ZN(P2_U3019) );
  NAND2_X1 U19574 ( .A1(n17685), .A2(n17709), .ZN(n17698) );
  OAI211_X1 U19575 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17701), .B(n17686), .ZN(
        n17688) );
  OAI211_X1 U19576 ( .C1(n17698), .C2(n17689), .A(n17688), .B(n17687), .ZN(
        n17691) );
  NOR2_X1 U19577 ( .A1(n19452), .A2(n19542), .ZN(n17690) );
  AOI211_X1 U19578 ( .C1(n19450), .C2(n19550), .A(n17691), .B(n17690), .ZN(
        n17694) );
  OR2_X1 U19579 ( .A1(n17692), .A2(n17944), .ZN(n17693) );
  OAI211_X1 U19580 ( .C1(n17695), .C2(n19546), .A(n17694), .B(n17693), .ZN(
        P2_U3020) );
  NAND2_X1 U19581 ( .A1(n17696), .A2(n19530), .ZN(n17705) );
  OAI21_X1 U19582 ( .B1(n17698), .B2(n17700), .A(n17697), .ZN(n17699) );
  AOI21_X1 U19583 ( .B1(n17701), .B2(n17700), .A(n17699), .ZN(n17702) );
  OAI21_X1 U19584 ( .B1(n19437), .B2(n19514), .A(n17702), .ZN(n17703) );
  AOI21_X1 U19585 ( .B1(n19439), .B2(n19527), .A(n17703), .ZN(n17704) );
  OAI211_X1 U19586 ( .C1(n17706), .C2(n17944), .A(n17705), .B(n17704), .ZN(
        P2_U3021) );
  OAI21_X1 U19587 ( .B1(n17719), .B2(n11593), .A(n17707), .ZN(n17708) );
  NAND2_X1 U19588 ( .A1(n17709), .A2(n17708), .ZN(n17710) );
  OAI211_X1 U19589 ( .C1(n17712), .C2(n19514), .A(n17711), .B(n17710), .ZN(
        n17715) );
  NOR2_X1 U19590 ( .A1(n17713), .A2(n17944), .ZN(n17714) );
  AOI211_X1 U19591 ( .C1(n19527), .C2(n19429), .A(n17715), .B(n17714), .ZN(
        n17716) );
  OAI21_X1 U19592 ( .B1(n17717), .B2(n19546), .A(n17716), .ZN(P2_U3022) );
  NAND2_X1 U19593 ( .A1(n17718), .A2(n19530), .ZN(n17726) );
  NOR2_X1 U19594 ( .A1(n19417), .A2(n19514), .ZN(n17724) );
  INV_X1 U19595 ( .A(n17719), .ZN(n17729) );
  OAI211_X1 U19596 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17729), .B(n11593), .ZN(
        n17720) );
  OAI211_X1 U19597 ( .C1(n17732), .C2(n17722), .A(n17721), .B(n17720), .ZN(
        n17723) );
  AOI211_X1 U19598 ( .C1(n19419), .C2(n19527), .A(n17724), .B(n17723), .ZN(
        n17725) );
  OAI211_X1 U19599 ( .C1(n17727), .C2(n17944), .A(n17726), .B(n17725), .ZN(
        P2_U3023) );
  AOI21_X1 U19600 ( .B1(n17729), .B2(n17731), .A(n17728), .ZN(n17730) );
  OAI21_X1 U19601 ( .B1(n17732), .B2(n17731), .A(n17730), .ZN(n17733) );
  AOI21_X1 U19602 ( .B1(n19404), .B2(n19550), .A(n17733), .ZN(n17734) );
  OAI21_X1 U19603 ( .B1(n19415), .B2(n19542), .A(n17734), .ZN(n17735) );
  INV_X1 U19604 ( .A(n17735), .ZN(n17739) );
  NAND3_X1 U19605 ( .A1(n17737), .A2(n19537), .A3(n17736), .ZN(n17738) );
  OAI211_X1 U19606 ( .C1(n17740), .C2(n19546), .A(n17739), .B(n17738), .ZN(
        P2_U3024) );
  INV_X1 U19607 ( .A(n17747), .ZN(n17741) );
  OR2_X1 U19608 ( .A1(n17794), .A2(n17741), .ZN(n17748) );
  NOR2_X1 U19609 ( .A1(n17748), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17776) );
  INV_X1 U19610 ( .A(n17784), .ZN(n17742) );
  AND2_X1 U19611 ( .A1(n19539), .A2(n17742), .ZN(n17743) );
  NOR2_X1 U19612 ( .A1(n17744), .A2(n17743), .ZN(n17788) );
  NAND2_X1 U19613 ( .A1(n17785), .A2(n17784), .ZN(n17745) );
  NAND2_X1 U19614 ( .A1(n17919), .A2(n17745), .ZN(n17746) );
  OAI211_X1 U19615 ( .C1(n19521), .C2(n17747), .A(n17788), .B(n17746), .ZN(
        n17775) );
  NOR2_X1 U19616 ( .A1(n17776), .A2(n17775), .ZN(n17760) );
  INV_X1 U19617 ( .A(n17748), .ZN(n17763) );
  NAND2_X1 U19618 ( .A1(n17749), .A2(n17753), .ZN(n17750) );
  OAI211_X1 U19619 ( .C1(n17753), .C2(n17762), .A(n17763), .B(n17750), .ZN(
        n17751) );
  OAI211_X1 U19620 ( .C1(n17760), .C2(n17753), .A(n17752), .B(n17751), .ZN(
        n17754) );
  AOI21_X1 U19621 ( .B1(n19391), .B2(n19550), .A(n17754), .ZN(n17755) );
  OAI21_X1 U19622 ( .B1(n19403), .B2(n19542), .A(n17755), .ZN(n17756) );
  AOI21_X1 U19623 ( .B1(n17757), .B2(n19537), .A(n17756), .ZN(n17758) );
  OAI21_X1 U19624 ( .B1(n17759), .B2(n19546), .A(n17758), .ZN(P2_U3026) );
  INV_X1 U19625 ( .A(n19385), .ZN(n17768) );
  NOR2_X1 U19626 ( .A1(n17760), .A2(n17762), .ZN(n17767) );
  INV_X1 U19627 ( .A(n17761), .ZN(n17765) );
  NAND3_X1 U19628 ( .A1(n17763), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17762), .ZN(n17764) );
  OAI211_X1 U19629 ( .C1(n19378), .C2(n19514), .A(n17765), .B(n17764), .ZN(
        n17766) );
  AOI211_X1 U19630 ( .C1(n17768), .C2(n19527), .A(n17767), .B(n17766), .ZN(
        n17771) );
  NAND2_X1 U19631 ( .A1(n17769), .A2(n19537), .ZN(n17770) );
  OAI211_X1 U19632 ( .C1(n17772), .C2(n19546), .A(n17771), .B(n17770), .ZN(
        P2_U3027) );
  INV_X1 U19633 ( .A(n17773), .ZN(n17780) );
  AOI21_X1 U19634 ( .B1(n17775), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17774), .ZN(n17778) );
  AOI21_X1 U19635 ( .B1(n19367), .B2(n19550), .A(n17776), .ZN(n17777) );
  OAI211_X1 U19636 ( .C1(n19373), .C2(n19542), .A(n17778), .B(n17777), .ZN(
        n17779) );
  AOI21_X1 U19637 ( .B1(n17780), .B2(n19530), .A(n17779), .ZN(n17781) );
  OAI21_X1 U19638 ( .B1(n17944), .B2(n17782), .A(n17781), .ZN(P2_U3028) );
  INV_X1 U19639 ( .A(n19539), .ZN(n19523) );
  NAND2_X1 U19640 ( .A1(n19523), .A2(n17944), .ZN(n17809) );
  NAND2_X1 U19641 ( .A1(n11229), .A2(n17809), .ZN(n17789) );
  NAND3_X1 U19642 ( .A1(n17785), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n17784), .ZN(n17786) );
  NAND2_X1 U19643 ( .A1(n17919), .A2(n17786), .ZN(n17787) );
  AND2_X1 U19644 ( .A1(n17788), .A2(n17787), .ZN(n17825) );
  OAI211_X1 U19645 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n19521), .A(
        n17789), .B(n17825), .ZN(n17800) );
  NAND2_X1 U19646 ( .A1(n17790), .A2(n19550), .ZN(n17791) );
  OAI211_X1 U19647 ( .C1(n17793), .C2(n19542), .A(n17792), .B(n17791), .ZN(
        n17799) );
  OAI21_X1 U19648 ( .B1(n17795), .B2(n17944), .A(n17794), .ZN(n17796) );
  NAND2_X1 U19649 ( .A1(n17796), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17814) );
  NOR3_X1 U19650 ( .A1(n17814), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n17797), .ZN(n17798) );
  AOI211_X1 U19651 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17800), .A(
        n17799), .B(n17798), .ZN(n17801) );
  OAI21_X1 U19652 ( .B1(n17802), .B2(n19546), .A(n17801), .ZN(P2_U3029) );
  INV_X1 U19653 ( .A(n19358), .ZN(n17808) );
  OAI21_X1 U19654 ( .B1(n17804), .B2(n19514), .A(n17803), .ZN(n17807) );
  NOR3_X1 U19655 ( .A1(n17805), .A2(n17535), .A3(n19546), .ZN(n17806) );
  AOI211_X1 U19656 ( .C1(n19527), .C2(n17808), .A(n17807), .B(n17806), .ZN(
        n17813) );
  INV_X1 U19657 ( .A(n17809), .ZN(n17810) );
  OAI21_X1 U19658 ( .B1(n17826), .B2(n17810), .A(n17825), .ZN(n17811) );
  NAND2_X1 U19659 ( .A1(n17811), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17812) );
  OAI211_X1 U19660 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17814), .A(
        n17813), .B(n17812), .ZN(P2_U3030) );
  INV_X1 U19661 ( .A(n17816), .ZN(n17817) );
  AOI21_X1 U19662 ( .B1(n17818), .B2(n17815), .A(n17817), .ZN(n20053) );
  INV_X1 U19663 ( .A(n19343), .ZN(n17820) );
  OAI21_X1 U19664 ( .B1(n17820), .B2(n19514), .A(n17819), .ZN(n17821) );
  AOI21_X1 U19665 ( .B1(n17822), .B2(n17824), .A(n17821), .ZN(n17823) );
  OAI21_X1 U19666 ( .B1(n17825), .B2(n17824), .A(n17823), .ZN(n17829) );
  NOR3_X1 U19667 ( .A1(n17827), .A2(n17826), .A3(n17944), .ZN(n17828) );
  AOI211_X1 U19668 ( .C1(n19527), .C2(n20053), .A(n17829), .B(n17828), .ZN(
        n17830) );
  OAI21_X1 U19669 ( .B1(n17831), .B2(n19546), .A(n17830), .ZN(P2_U3031) );
  NAND2_X1 U19670 ( .A1(n17832), .A2(n19530), .ZN(n17845) );
  INV_X1 U19671 ( .A(n17836), .ZN(n17833) );
  AOI21_X1 U19672 ( .B1(n17834), .B2(n17833), .A(n17875), .ZN(n17866) );
  AND2_X1 U19673 ( .A1(n17836), .A2(n17865), .ZN(n17835) );
  NAND2_X1 U19674 ( .A1(n17877), .A2(n17835), .ZN(n17863) );
  NAND2_X1 U19675 ( .A1(n17866), .A2(n17863), .ZN(n17853) );
  INV_X1 U19676 ( .A(n17877), .ZN(n17909) );
  OAI21_X1 U19677 ( .B1(n17865), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17837) );
  OAI211_X1 U19678 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n17837), .B(n17836), .ZN(
        n17840) );
  NAND2_X1 U19679 ( .A1(n19331), .A2(n19550), .ZN(n17839) );
  OAI211_X1 U19680 ( .C1(n17909), .C2(n17840), .A(n17839), .B(n17838), .ZN(
        n17843) );
  OAI21_X1 U19681 ( .B1(n15805), .B2(n17841), .A(n17815), .ZN(n20058) );
  NOR2_X1 U19682 ( .A1(n20058), .A2(n19542), .ZN(n17842) );
  AOI211_X1 U19683 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17853), .A(
        n17843), .B(n17842), .ZN(n17844) );
  OAI211_X1 U19684 ( .C1(n17846), .C2(n17944), .A(n17845), .B(n17844), .ZN(
        P2_U3032) );
  NAND3_X1 U19685 ( .A1(n17877), .A2(n17848), .A3(n17847), .ZN(n17849) );
  OAI211_X1 U19686 ( .C1(n17851), .C2(n19514), .A(n17850), .B(n17849), .ZN(
        n17852) );
  AOI21_X1 U19687 ( .B1(n17853), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n17852), .ZN(n17854) );
  OAI21_X1 U19688 ( .B1(n17855), .B2(n19542), .A(n17854), .ZN(n17856) );
  AOI21_X1 U19689 ( .B1(n17857), .B2(n19530), .A(n17856), .ZN(n17858) );
  OAI21_X1 U19690 ( .B1(n17944), .B2(n17859), .A(n17858), .ZN(P2_U3033) );
  OAI21_X1 U19691 ( .B1(n11594), .B2(n11363), .A(n15804), .ZN(n20064) );
  INV_X1 U19692 ( .A(n20064), .ZN(n17870) );
  INV_X1 U19693 ( .A(n17861), .ZN(n17862) );
  AOI21_X1 U19694 ( .B1(n19321), .B2(n19550), .A(n17862), .ZN(n17864) );
  OAI211_X1 U19695 ( .C1(n17866), .C2(n17865), .A(n17864), .B(n17863), .ZN(
        n17869) );
  NOR2_X1 U19696 ( .A1(n17867), .A2(n19546), .ZN(n17868) );
  AOI211_X1 U19697 ( .C1(n19527), .C2(n17870), .A(n17869), .B(n17868), .ZN(
        n17871) );
  OAI21_X1 U19698 ( .B1(n17944), .B2(n17872), .A(n17871), .ZN(P2_U3034) );
  OAI21_X1 U19699 ( .B1(n17874), .B2(n17873), .A(n17860), .ZN(n19299) );
  INV_X1 U19700 ( .A(n17875), .ZN(n17905) );
  OAI21_X1 U19701 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19521), .A(
        n17905), .ZN(n17895) );
  OAI21_X1 U19702 ( .B1(n19306), .B2(n19514), .A(n17876), .ZN(n17880) );
  NAND2_X1 U19703 ( .A1(n17877), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17898) );
  XNOR2_X1 U19704 ( .A(n12661), .B(n17894), .ZN(n17878) );
  NOR2_X1 U19705 ( .A1(n17898), .A2(n17878), .ZN(n17879) );
  AOI211_X1 U19706 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n17895), .A(
        n17880), .B(n17879), .ZN(n17881) );
  OAI21_X1 U19707 ( .B1(n19299), .B2(n19542), .A(n17881), .ZN(n17882) );
  AOI21_X1 U19708 ( .B1(n17883), .B2(n19530), .A(n17882), .ZN(n17884) );
  OAI21_X1 U19709 ( .B1(n17885), .B2(n17944), .A(n17884), .ZN(P2_U3035) );
  NAND2_X1 U19710 ( .A1(n17887), .A2(n17886), .ZN(n17892) );
  INV_X1 U19711 ( .A(n17888), .ZN(n17890) );
  NOR2_X1 U19712 ( .A1(n17890), .A2(n17889), .ZN(n17891) );
  XNOR2_X1 U19713 ( .A(n17892), .B(n17891), .ZN(n18084) );
  AOI21_X1 U19714 ( .B1(n17894), .B2(n17902), .A(n17893), .ZN(n18085) );
  NAND2_X1 U19715 ( .A1(n18085), .A2(n19537), .ZN(n17901) );
  NAND2_X1 U19716 ( .A1(n17895), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17897) );
  AOI22_X1 U19717 ( .A1(n19550), .A2(n18087), .B1(P2_REIP_REG_10__SCAN_IN), 
        .B2(n19526), .ZN(n17896) );
  OAI211_X1 U19718 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17898), .A(
        n17897), .B(n17896), .ZN(n17899) );
  AOI21_X1 U19719 ( .B1(n20069), .B2(n19527), .A(n17899), .ZN(n17900) );
  OAI211_X1 U19720 ( .C1(n18084), .C2(n19546), .A(n17901), .B(n17900), .ZN(
        P2_U3036) );
  NAND3_X1 U19721 ( .A1(n17903), .A2(n17902), .A3(n19537), .ZN(n17913) );
  NOR2_X1 U19722 ( .A1(n17905), .A2(n17904), .ZN(n17911) );
  NAND2_X1 U19723 ( .A1(n19550), .A2(n17906), .ZN(n17908) );
  OAI211_X1 U19724 ( .C1(n17909), .C2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17908), .B(n17907), .ZN(n17910) );
  AOI211_X1 U19725 ( .C1(n20074), .C2(n19527), .A(n17911), .B(n17910), .ZN(
        n17912) );
  OAI211_X1 U19726 ( .C1(n17914), .C2(n19546), .A(n17913), .B(n17912), .ZN(
        P2_U3037) );
  NAND3_X1 U19727 ( .A1(n17915), .A2(n17624), .A3(n19537), .ZN(n17931) );
  INV_X1 U19728 ( .A(n17916), .ZN(n17920) );
  AOI21_X1 U19729 ( .B1(n17919), .B2(n17918), .A(n17917), .ZN(n19522) );
  OAI21_X1 U19730 ( .B1(n17920), .B2(n19523), .A(n19522), .ZN(n17934) );
  NAND2_X1 U19731 ( .A1(n17922), .A2(n17921), .ZN(n17923) );
  NAND2_X1 U19732 ( .A1(n17220), .A2(n17923), .ZN(n20079) );
  NAND2_X1 U19733 ( .A1(n19524), .A2(n17924), .ZN(n19535) );
  NOR2_X1 U19734 ( .A1(n18074), .A2(n19535), .ZN(n17936) );
  OAI211_X1 U19735 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n17936), .B(n17925), .ZN(n17928) );
  OAI22_X1 U19736 ( .A1(n19514), .A2(n19294), .B1(n17625), .B2(n19301), .ZN(
        n17926) );
  INV_X1 U19737 ( .A(n17926), .ZN(n17927) );
  OAI211_X1 U19738 ( .C1(n20079), .C2(n19542), .A(n17928), .B(n17927), .ZN(
        n17929) );
  AOI21_X1 U19739 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17934), .A(
        n17929), .ZN(n17930) );
  OAI211_X1 U19740 ( .C1(n17932), .C2(n19546), .A(n17931), .B(n17930), .ZN(
        P2_U3038) );
  AND2_X1 U19741 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19526), .ZN(n17933) );
  AOI221_X1 U19742 ( .B1(n17936), .B2(n17935), .C1(n17934), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n17933), .ZN(n17937) );
  INV_X1 U19743 ( .A(n17937), .ZN(n17941) );
  XNOR2_X1 U19744 ( .A(n17938), .B(n17939), .ZN(n20082) );
  OAI22_X1 U19745 ( .A1(n20082), .A2(n19542), .B1(n19514), .B2(n19283), .ZN(
        n17940) );
  AOI211_X1 U19746 ( .C1(n17942), .C2(n19530), .A(n17941), .B(n17940), .ZN(
        n17943) );
  OAI21_X1 U19747 ( .B1(n17945), .B2(n17944), .A(n17943), .ZN(P2_U3039) );
  AOI22_X1 U19748 ( .A1(n19396), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n17946), .B2(n11253), .ZN(n17947) );
  INV_X1 U19749 ( .A(n17947), .ZN(n17954) );
  NOR2_X1 U19750 ( .A1(n17949), .A2(n17948), .ZN(n17953) );
  INV_X1 U19751 ( .A(n17953), .ZN(n17951) );
  OAI222_X1 U19752 ( .A1(n17954), .A2(n17951), .B1(n19557), .B2(n17950), .C1(
        n17961), .C2(n20108), .ZN(n17952) );
  MUX2_X1 U19753 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n17952), .S(
        n19510), .Z(P2_U3600) );
  AOI222_X1 U19754 ( .A1(n17956), .A2(n17955), .B1(n18109), .B2(n19572), .C1(
        n17954), .C2(n17953), .ZN(n17959) );
  NAND2_X1 U19755 ( .A1(n19507), .A2(n17957), .ZN(n17958) );
  OAI21_X1 U19756 ( .B1(n17959), .B2(n19507), .A(n17958), .ZN(P2_U3599) );
  OAI22_X1 U19757 ( .A1(n20132), .A2(n17961), .B1(n17960), .B2(n19557), .ZN(
        n17962) );
  MUX2_X1 U19758 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17962), .S(
        n19510), .Z(P2_U3596) );
  NOR2_X1 U19759 ( .A1(n21619), .A2(n21998), .ZN(n18578) );
  NOR2_X1 U19760 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18578), .ZN(n20957) );
  NAND2_X1 U19761 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19105) );
  NAND2_X1 U19762 ( .A1(n20957), .A2(n19105), .ZN(n17967) );
  NOR2_X1 U19763 ( .A1(n19636), .A2(n19609), .ZN(n19632) );
  AOI21_X1 U19764 ( .B1(n17967), .B2(n22084), .A(n19632), .ZN(n17966) );
  NAND2_X1 U19765 ( .A1(n19653), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19627) );
  NAND2_X1 U19766 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18578), .ZN(n22083) );
  NAND2_X1 U19767 ( .A1(n17963), .A2(n17972), .ZN(n17964) );
  NOR2_X1 U19768 ( .A1(n18616), .A2(n17964), .ZN(n18579) );
  INV_X1 U19769 ( .A(n22087), .ZN(n17965) );
  OAI221_X1 U19770 ( .B1(n22083), .B2(n18579), .C1(n22083), .C2(n22102), .A(
        n19863), .ZN(n19153) );
  NAND2_X1 U19771 ( .A1(n19627), .A2(n19153), .ZN(n19154) );
  NOR2_X1 U19772 ( .A1(n17966), .A2(n19154), .ZN(n19151) );
  NOR3_X2 U19773 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n22414), .ZN(n19648) );
  OAI21_X1 U19774 ( .B1(n19653), .B2(n22084), .A(n17967), .ZN(n19152) );
  OAI221_X1 U19775 ( .B1(n19648), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19648), .C2(n19152), .A(n19153), .ZN(n19149) );
  AOI22_X1 U19776 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19151), .B1(
        n19149), .B2(n19609), .ZN(P3_U2865) );
  NOR2_X1 U19777 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n22084), .ZN(n19613) );
  NOR2_X1 U19778 ( .A1(n22102), .A2(n22083), .ZN(n17968) );
  INV_X1 U19779 ( .A(n21639), .ZN(n21636) );
  NOR2_X1 U19780 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21634) );
  NAND3_X1 U19781 ( .A1(n21636), .A2(n21634), .A3(n17970), .ZN(n17971) );
  OAI21_X1 U19782 ( .B1(n21636), .B2(n17972), .A(n17971), .ZN(P3_U3284) );
  NOR2_X1 U19783 ( .A1(n17974), .A2(n17973), .ZN(n17975) );
  XNOR2_X1 U19784 ( .A(n17975), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n22266) );
  NAND3_X1 U19785 ( .A1(n11207), .A2(n17977), .A3(n17976), .ZN(n17978) );
  OAI21_X1 U19786 ( .B1(n17979), .B2(n18038), .A(n17978), .ZN(P1_U3468) );
  INV_X1 U19787 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17982) );
  INV_X2 U19788 ( .A(n22421), .ZN(n22469) );
  OAI21_X1 U19789 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n17980), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n19219) );
  INV_X1 U19790 ( .A(n22417), .ZN(n17983) );
  NOR2_X1 U19791 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n19180) );
  OAI21_X1 U19792 ( .B1(BS16), .B2(n19180), .A(n22417), .ZN(n22415) );
  INV_X1 U19793 ( .A(n22415), .ZN(n17981) );
  AOI21_X1 U19794 ( .B1(n17982), .B2(n17983), .A(n17981), .ZN(P3_U3280) );
  AND2_X1 U19795 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17983), .ZN(P3_U3028) );
  AND2_X1 U19796 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17983), .ZN(P3_U3027) );
  AND2_X1 U19797 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17983), .ZN(P3_U3026) );
  AND2_X1 U19798 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17983), .ZN(P3_U3025) );
  AND2_X1 U19799 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17983), .ZN(P3_U3024) );
  AND2_X1 U19800 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17983), .ZN(P3_U3023) );
  AND2_X1 U19801 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17983), .ZN(P3_U3022) );
  AND2_X1 U19802 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17983), .ZN(P3_U3021) );
  AND2_X1 U19803 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17983), .ZN(
        P3_U3020) );
  AND2_X1 U19804 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17983), .ZN(
        P3_U3019) );
  AND2_X1 U19805 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17983), .ZN(
        P3_U3018) );
  AND2_X1 U19806 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17983), .ZN(
        P3_U3017) );
  AND2_X1 U19807 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17983), .ZN(
        P3_U3016) );
  AND2_X1 U19808 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17983), .ZN(
        P3_U3015) );
  AND2_X1 U19809 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17983), .ZN(
        P3_U3014) );
  AND2_X1 U19810 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17983), .ZN(
        P3_U3013) );
  AND2_X1 U19811 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17983), .ZN(
        P3_U3012) );
  AND2_X1 U19812 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17983), .ZN(
        P3_U3011) );
  AND2_X1 U19813 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17983), .ZN(
        P3_U3010) );
  AND2_X1 U19814 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17983), .ZN(
        P3_U3009) );
  AND2_X1 U19815 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17983), .ZN(
        P3_U3008) );
  AND2_X1 U19816 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17983), .ZN(
        P3_U3007) );
  AND2_X1 U19817 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17983), .ZN(
        P3_U3006) );
  AND2_X1 U19818 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17983), .ZN(
        P3_U3005) );
  AND2_X1 U19819 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17983), .ZN(
        P3_U3004) );
  AND2_X1 U19820 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17983), .ZN(
        P3_U3003) );
  AND2_X1 U19821 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17983), .ZN(
        P3_U3002) );
  AND2_X1 U19822 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17983), .ZN(
        P3_U3001) );
  AND2_X1 U19823 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17983), .ZN(
        P3_U3000) );
  AND2_X1 U19824 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17983), .ZN(
        P3_U2999) );
  AOI21_X1 U19825 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17986)
         );
  INV_X1 U19826 ( .A(n22083), .ZN(n17985) );
  AOI211_X1 U19827 ( .C1(n19105), .C2(n17986), .A(n17985), .B(n17984), .ZN(
        P3_U2998) );
  NOR2_X1 U19828 ( .A1(n17987), .A2(n19153), .ZN(P3_U2867) );
  AND2_X1 U19829 ( .A1(n19208), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U19830 ( .A1(n18577), .A2(n20954), .ZN(n17991) );
  OAI22_X1 U19831 ( .A1(P3_READREQUEST_REG_SCAN_IN), .A2(n17991), .B1(n20961), 
        .B2(n20954), .ZN(n17990) );
  INV_X1 U19832 ( .A(n17990), .ZN(P3_U3298) );
  NOR2_X1 U19833 ( .A1(P3_MEMORYFETCH_REG_SCAN_IN), .A2(n17991), .ZN(n17992)
         );
  NOR2_X1 U19834 ( .A1(n21421), .A2(n17992), .ZN(P3_U3299) );
  NOR2_X1 U19835 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n22444), .ZN(n22450) );
  AOI21_X1 U19836 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n22450), .A(n17993), 
        .ZN(n17994) );
  INV_X1 U19837 ( .A(n17994), .ZN(n22413) );
  INV_X1 U19838 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18009) );
  INV_X1 U19839 ( .A(BS16), .ZN(n18011) );
  INV_X1 U19840 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22461) );
  NAND2_X1 U19841 ( .A1(n22444), .A2(n22461), .ZN(n22443) );
  AOI21_X1 U19842 ( .B1(n18011), .B2(n22443), .A(n18125), .ZN(n22409) );
  AOI21_X1 U19843 ( .B1(n18125), .B2(n18009), .A(n22409), .ZN(P2_U3591) );
  AND2_X1 U19844 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n18125), .ZN(P2_U3208) );
  AND2_X1 U19845 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17994), .ZN(P2_U3207) );
  AND2_X1 U19846 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n18125), .ZN(P2_U3206) );
  AND2_X1 U19847 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n18125), .ZN(P2_U3205) );
  AND2_X1 U19848 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n18125), .ZN(P2_U3204) );
  AND2_X1 U19849 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n18125), .ZN(P2_U3203) );
  AND2_X1 U19850 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17994), .ZN(P2_U3202) );
  AND2_X1 U19851 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17994), .ZN(P2_U3201) );
  AND2_X1 U19852 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17994), .ZN(
        P2_U3200) );
  AND2_X1 U19853 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17994), .ZN(
        P2_U3199) );
  AND2_X1 U19854 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17994), .ZN(
        P2_U3198) );
  AND2_X1 U19855 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17994), .ZN(
        P2_U3197) );
  AND2_X1 U19856 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17994), .ZN(
        P2_U3196) );
  AND2_X1 U19857 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17994), .ZN(
        P2_U3195) );
  AND2_X1 U19858 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17994), .ZN(
        P2_U3194) );
  AND2_X1 U19859 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17994), .ZN(
        P2_U3193) );
  AND2_X1 U19860 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17994), .ZN(
        P2_U3192) );
  AND2_X1 U19861 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17994), .ZN(
        P2_U3191) );
  AND2_X1 U19862 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n18125), .ZN(
        P2_U3190) );
  AND2_X1 U19863 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n18125), .ZN(
        P2_U3189) );
  AND2_X1 U19864 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n18125), .ZN(
        P2_U3188) );
  AND2_X1 U19865 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n18125), .ZN(
        P2_U3187) );
  AND2_X1 U19866 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17994), .ZN(
        P2_U3186) );
  AND2_X1 U19867 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n18125), .ZN(
        P2_U3185) );
  AND2_X1 U19868 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n18125), .ZN(
        P2_U3184) );
  AND2_X1 U19869 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n18125), .ZN(
        P2_U3183) );
  AND2_X1 U19870 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n18125), .ZN(
        P2_U3182) );
  AND2_X1 U19871 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n18125), .ZN(
        P2_U3181) );
  AND2_X1 U19872 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n18125), .ZN(
        P2_U3180) );
  AND2_X1 U19873 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n18125), .ZN(
        P2_U3179) );
  OAI221_X1 U19874 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(
        P2_STATEBS16_REG_SCAN_IN), .C1(n17995), .C2(n22445), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17996) );
  AOI21_X1 U19875 ( .B1(n17996), .B2(n20235), .A(n19567), .ZN(P2_U3178) );
  INV_X1 U19876 ( .A(n19568), .ZN(n17997) );
  AOI221_X1 U19877 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n19567), .C1(n17997), .C2(
        n19567), .A(n20257), .ZN(n18115) );
  INV_X1 U19878 ( .A(n18115), .ZN(n18113) );
  NOR2_X1 U19879 ( .A1(n17998), .A2(n18113), .ZN(P2_U3047) );
  AND2_X1 U19880 ( .A1(n18145), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19881 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18002) );
  NOR4_X1 U19882 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18001) );
  NOR4_X1 U19883 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18000) );
  NOR4_X1 U19884 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17999) );
  NAND4_X1 U19885 ( .A1(n18002), .A2(n18001), .A3(n18000), .A4(n17999), .ZN(
        n18008) );
  NOR4_X1 U19886 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18006) );
  AOI211_X1 U19887 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18005) );
  NOR4_X1 U19888 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18004) );
  NOR4_X1 U19889 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18003) );
  NAND4_X1 U19890 ( .A1(n18006), .A2(n18005), .A3(n18004), .A4(n18003), .ZN(
        n18007) );
  NOR2_X1 U19891 ( .A1(n18008), .A2(n18007), .ZN(n18123) );
  INV_X1 U19892 ( .A(n18123), .ZN(n18122) );
  NOR2_X1 U19893 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18122), .ZN(n18116) );
  INV_X1 U19894 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22412) );
  NAND3_X1 U19895 ( .A1(n18010), .A2(n22412), .A3(n18009), .ZN(n18121) );
  INV_X1 U19896 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18197) );
  AOI22_X1 U19897 ( .A1(n18116), .A2(n18121), .B1(n18122), .B2(n18197), .ZN(
        P2_U2821) );
  INV_X1 U19898 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18195) );
  AOI22_X1 U19899 ( .A1(n18116), .A2(n18010), .B1(n18122), .B2(n18195), .ZN(
        P2_U2820) );
  INV_X1 U19900 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18012) );
  INV_X2 U19901 ( .A(n22852), .ZN(n22855) );
  INV_X1 U19902 ( .A(n22408), .ZN(n18013) );
  INV_X1 U19903 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n22440) );
  NAND2_X1 U19904 ( .A1(n22433), .A2(n22440), .ZN(n20883) );
  AOI21_X1 U19905 ( .B1(n18011), .B2(n20883), .A(n18013), .ZN(n22404) );
  AOI21_X1 U19906 ( .B1(n18012), .B2(n18013), .A(n22404), .ZN(P1_U3464) );
  AND2_X1 U19907 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n18013), .ZN(P1_U3193) );
  AND2_X1 U19908 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n18013), .ZN(P1_U3192) );
  AND2_X1 U19909 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n18013), .ZN(P1_U3191) );
  AND2_X1 U19910 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n18013), .ZN(P1_U3190) );
  AND2_X1 U19911 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n18013), .ZN(P1_U3189) );
  AND2_X1 U19912 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n18013), .ZN(P1_U3188) );
  AND2_X1 U19913 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n18013), .ZN(P1_U3187) );
  AND2_X1 U19914 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n18013), .ZN(P1_U3186) );
  AND2_X1 U19915 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n18013), .ZN(
        P1_U3185) );
  AND2_X1 U19916 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n18013), .ZN(
        P1_U3184) );
  AND2_X1 U19917 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n18013), .ZN(
        P1_U3183) );
  AND2_X1 U19918 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n18013), .ZN(
        P1_U3182) );
  AND2_X1 U19919 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n18013), .ZN(
        P1_U3181) );
  AND2_X1 U19920 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n18013), .ZN(
        P1_U3180) );
  AND2_X1 U19921 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n18013), .ZN(
        P1_U3179) );
  AND2_X1 U19922 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n18013), .ZN(
        P1_U3178) );
  AND2_X1 U19923 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n18013), .ZN(
        P1_U3177) );
  AND2_X1 U19924 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n18013), .ZN(
        P1_U3176) );
  AND2_X1 U19925 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n18013), .ZN(
        P1_U3175) );
  AND2_X1 U19926 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n18013), .ZN(
        P1_U3174) );
  AND2_X1 U19927 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n18013), .ZN(
        P1_U3173) );
  AND2_X1 U19928 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n18013), .ZN(
        P1_U3172) );
  AND2_X1 U19929 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n18013), .ZN(
        P1_U3171) );
  AND2_X1 U19930 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n18013), .ZN(
        P1_U3170) );
  AND2_X1 U19931 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n18013), .ZN(
        P1_U3169) );
  AND2_X1 U19932 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n18013), .ZN(
        P1_U3168) );
  AND2_X1 U19933 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n18013), .ZN(
        P1_U3167) );
  AND2_X1 U19934 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n18013), .ZN(
        P1_U3166) );
  AND2_X1 U19935 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n18013), .ZN(
        P1_U3165) );
  AND2_X1 U19936 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n18013), .ZN(
        P1_U3164) );
  MUX2_X1 U19937 ( .A(n18014), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n18017), .Z(n18042) );
  MUX2_X1 U19938 ( .A(n18015), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n18017), .Z(n18041) );
  OR2_X1 U19939 ( .A1(n18017), .A2(n18016), .ZN(n18023) );
  AOI21_X1 U19940 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18019), .A(
        n18018), .ZN(n18020) );
  AOI22_X1 U19941 ( .A1(n18023), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18020), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18021) );
  INV_X1 U19942 ( .A(n18021), .ZN(n18022) );
  OAI21_X1 U19943 ( .B1(n18023), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n18022), .ZN(n18024) );
  AOI222_X1 U19944 ( .A1(n18042), .A2(n22552), .B1(n18042), .B2(n18024), .C1(
        n22552), .C2(n18024), .ZN(n18027) );
  NAND2_X1 U19945 ( .A1(n22553), .A2(n18041), .ZN(n18026) );
  INV_X1 U19946 ( .A(n18041), .ZN(n18025) );
  AOI221_X1 U19947 ( .B1(n18027), .B2(n18026), .C1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n18025), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18040) );
  INV_X1 U19948 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n18028) );
  NAND2_X1 U19949 ( .A1(n18028), .A2(n22386), .ZN(n18029) );
  NAND2_X1 U19950 ( .A1(n18030), .A2(n18029), .ZN(n18034) );
  NOR2_X1 U19951 ( .A1(n18032), .A2(n18031), .ZN(n18033) );
  AND2_X1 U19952 ( .A1(n18034), .A2(n18033), .ZN(n18036) );
  INV_X1 U19953 ( .A(n11207), .ZN(n18035) );
  OAI211_X1 U19954 ( .C1(n18038), .C2(n18037), .A(n18036), .B(n18035), .ZN(
        n18039) );
  AOI211_X1 U19955 ( .C1(n18042), .C2(n18041), .A(n18040), .B(n18039), .ZN(
        n22403) );
  INV_X1 U19956 ( .A(n22403), .ZN(n18050) );
  NAND3_X1 U19957 ( .A1(n18045), .A2(n18044), .A3(n18043), .ZN(n18049) );
  OAI21_X1 U19958 ( .B1(n22424), .B2(n18047), .A(n18046), .ZN(n18048) );
  NAND2_X1 U19959 ( .A1(n18049), .A2(n18048), .ZN(n18056) );
  AOI221_X1 U19960 ( .B1(n22392), .B2(n22388), .C1(n18050), .C2(n22388), .A(
        n18056), .ZN(n22395) );
  NOR2_X1 U19961 ( .A1(n22395), .A2(n22392), .ZN(n22394) );
  INV_X1 U19962 ( .A(n18051), .ZN(n22397) );
  NAND2_X1 U19963 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22397), .ZN(n18052) );
  OAI211_X1 U19964 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n22424), .A(n22394), 
        .B(n18052), .ZN(n22399) );
  NAND4_X1 U19965 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n22556), .A4(n22424), .ZN(n18053) );
  AND2_X1 U19966 ( .A1(n18054), .A2(n18053), .ZN(n22389) );
  NAND2_X1 U19967 ( .A1(n22389), .A2(n22391), .ZN(n18055) );
  AOI22_X1 U19968 ( .A1(n22388), .A2(n22399), .B1(n18056), .B2(n18055), .ZN(
        P1_U3162) );
  AND2_X1 U19969 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18057), .ZN(
        P1_U3032) );
  AND2_X1 U19970 ( .A1(n20722), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI21_X1 U19971 ( .B1(n18059), .B2(n18058), .A(n22855), .ZN(P1_U2802) );
  INV_X1 U19972 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18060) );
  INV_X1 U19973 ( .A(n19565), .ZN(n19560) );
  OAI22_X1 U19974 ( .A1(n19275), .A2(n18060), .B1(n19560), .B2(n19557), .ZN(
        P2_U2816) );
  AOI22_X1 U19975 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19526), .B1(n18083), 
        .B2(n18061), .ZN(n18070) );
  INV_X1 U19976 ( .A(n18062), .ZN(n18068) );
  OAI22_X1 U19977 ( .A1(n18066), .A2(n18065), .B1(n18064), .B2(n18063), .ZN(
        n18067) );
  AOI21_X1 U19978 ( .B1(n18088), .B2(n18068), .A(n18067), .ZN(n18069) );
  OAI211_X1 U19979 ( .C1(n18071), .C2(n18093), .A(n18070), .B(n18069), .ZN(
        P2_U3010) );
  AOI22_X1 U19980 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19526), .B1(n18083), 
        .B2(n18072), .ZN(n18080) );
  XNOR2_X1 U19981 ( .A(n11239), .B(n18074), .ZN(n19532) );
  XOR2_X1 U19982 ( .A(n18076), .B(n18075), .Z(n19529) );
  AOI22_X1 U19983 ( .A1(n19532), .A2(n18086), .B1(n18089), .B2(n19529), .ZN(
        n18077) );
  INV_X1 U19984 ( .A(n18077), .ZN(n18078) );
  AOI21_X1 U19985 ( .B1(n18088), .B2(n19531), .A(n18078), .ZN(n18079) );
  OAI211_X1 U19986 ( .C1(n18081), .C2(n18093), .A(n18080), .B(n18079), .ZN(
        P2_U3008) );
  AOI22_X1 U19987 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19526), .B1(n18083), 
        .B2(n18082), .ZN(n18092) );
  INV_X1 U19988 ( .A(n18084), .ZN(n18090) );
  AOI222_X1 U19989 ( .A1(n18090), .A2(n18089), .B1(n18088), .B2(n18087), .C1(
        n18086), .C2(n18085), .ZN(n18091) );
  OAI211_X1 U19990 ( .C1(n18094), .C2(n18093), .A(n18092), .B(n18091), .ZN(
        P2_U3004) );
  INV_X1 U19991 ( .A(n18095), .ZN(n18097) );
  OAI22_X1 U19992 ( .A1(n18098), .A2(n19273), .B1(n18097), .B2(n18096), .ZN(
        n18099) );
  AOI21_X1 U19993 ( .B1(n20247), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n18099), 
        .ZN(n18100) );
  OAI22_X1 U19994 ( .A1(n20247), .A2(n18113), .B1(n18115), .B2(n18100), .ZN(
        P2_U3605) );
  OR2_X1 U19995 ( .A1(n20108), .A2(n22410), .ZN(n20173) );
  INV_X1 U19996 ( .A(n20173), .ZN(n18101) );
  NAND2_X1 U19997 ( .A1(n20447), .A2(n18101), .ZN(n20220) );
  AOI21_X1 U19998 ( .B1(n18101), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n19273), 
        .ZN(n18110) );
  NAND2_X1 U19999 ( .A1(n18110), .A2(n18109), .ZN(n18103) );
  NAND2_X1 U20000 ( .A1(n20446), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18102) );
  OAI211_X1 U20001 ( .C1(n20220), .C2(n20254), .A(n18103), .B(n18102), .ZN(
        n18104) );
  INV_X1 U20002 ( .A(n18104), .ZN(n18105) );
  AOI22_X1 U20003 ( .A1(n18115), .A2(n20161), .B1(n18105), .B2(n18113), .ZN(
        P2_U3603) );
  AND2_X1 U20004 ( .A1(n20222), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n18111) );
  OR2_X1 U20005 ( .A1(n18106), .A2(n18111), .ZN(n18107) );
  AOI22_X1 U20006 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20496), .B1(n18110), 
        .B2(n18107), .ZN(n18108) );
  AOI22_X1 U20007 ( .A1(n18115), .A2(n20245), .B1(n18108), .B2(n18113), .ZN(
        P2_U3604) );
  INV_X1 U20008 ( .A(n20192), .ZN(n20193) );
  OAI21_X1 U20009 ( .B1(n20193), .B2(n20108), .A(n20150), .ZN(n18112) );
  AOI222_X1 U20010 ( .A1(n18112), .A2(n18111), .B1(n20221), .B2(n18110), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n20401), .ZN(n18114) );
  AOI22_X1 U20011 ( .A1(n18115), .A2(n20140), .B1(n18114), .B2(n18113), .ZN(
        P2_U3602) );
  NAND2_X1 U20012 ( .A1(n18116), .A2(n22412), .ZN(n18120) );
  AOI21_X1 U20013 ( .B1(P2_REIP_REG_1__SCAN_IN), .B2(P2_REIP_REG_0__SCAN_IN), 
        .A(n18122), .ZN(n18117) );
  INV_X1 U20014 ( .A(n18117), .ZN(n18118) );
  OAI21_X1 U20015 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18123), .A(n18118), 
        .ZN(n18119) );
  OAI221_X1 U20016 ( .B1(n18120), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18120), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18119), .ZN(P2_U2822) );
  INV_X1 U20017 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18199) );
  OAI221_X1 U20018 ( .B1(n18123), .B2(n18199), .C1(n18122), .C2(n18121), .A(
        n18120), .ZN(P2_U2823) );
  MUX2_X1 U20019 ( .A(P2_M_IO_N_REG_SCAN_IN), .B(P2_MEMORYFETCH_REG_SCAN_IN), 
        .S(n22449), .Z(P2_U3611) );
  INV_X1 U20020 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n18124) );
  AOI22_X1 U20021 ( .A1(n22449), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n18124), 
        .B2(n18186), .ZN(P2_U3608) );
  INV_X1 U20022 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n22455) );
  INV_X1 U20023 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18126) );
  OAI21_X1 U20024 ( .B1(n22455), .B2(n18126), .A(n18125), .ZN(P2_U2815) );
  INV_X1 U20025 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n18129) );
  AOI22_X1 U20026 ( .A1(n18154), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18128) );
  OAI21_X1 U20027 ( .B1(n18129), .B2(n18156), .A(n18128), .ZN(P2_U2951) );
  INV_X1 U20028 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18131) );
  AOI22_X1 U20029 ( .A1(n18154), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18130) );
  OAI21_X1 U20030 ( .B1(n18131), .B2(n18156), .A(n18130), .ZN(P2_U2950) );
  INV_X1 U20031 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18133) );
  AOI22_X1 U20032 ( .A1(n18154), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18132) );
  OAI21_X1 U20033 ( .B1(n18133), .B2(n18156), .A(n18132), .ZN(P2_U2949) );
  INV_X1 U20034 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18135) );
  AOI22_X1 U20035 ( .A1(n18146), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18134) );
  OAI21_X1 U20036 ( .B1(n18135), .B2(n18156), .A(n18134), .ZN(P2_U2948) );
  AOI22_X1 U20037 ( .A1(n18154), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18136) );
  OAI21_X1 U20038 ( .B1(n18137), .B2(n18156), .A(n18136), .ZN(P2_U2947) );
  INV_X1 U20039 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18139) );
  AOI22_X1 U20040 ( .A1(n18146), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18138) );
  OAI21_X1 U20041 ( .B1(n18139), .B2(n18156), .A(n18138), .ZN(P2_U2946) );
  INV_X1 U20042 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18141) );
  AOI22_X1 U20043 ( .A1(n18146), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18140) );
  OAI21_X1 U20044 ( .B1(n18141), .B2(n18156), .A(n18140), .ZN(P2_U2945) );
  INV_X1 U20045 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20080) );
  AOI22_X1 U20046 ( .A1(n18146), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18142) );
  OAI21_X1 U20047 ( .B1(n20080), .B2(n18156), .A(n18142), .ZN(P2_U2944) );
  INV_X1 U20048 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20078) );
  AOI22_X1 U20049 ( .A1(n18146), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18143) );
  OAI21_X1 U20050 ( .B1(n20078), .B2(n18156), .A(n18143), .ZN(P2_U2943) );
  AOI22_X1 U20051 ( .A1(n18154), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18144) );
  OAI21_X1 U20052 ( .B1(n20076), .B2(n18156), .A(n18144), .ZN(P2_U2942) );
  INV_X1 U20053 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n18148) );
  AOI22_X1 U20054 ( .A1(n18146), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18147) );
  OAI21_X1 U20055 ( .B1(n18148), .B2(n18156), .A(n18147), .ZN(P2_U2941) );
  AOI22_X1 U20056 ( .A1(n18154), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18149) );
  OAI21_X1 U20057 ( .B1(n20068), .B2(n18156), .A(n18149), .ZN(P2_U2940) );
  INV_X1 U20058 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20063) );
  AOI22_X1 U20059 ( .A1(n18154), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18150) );
  OAI21_X1 U20060 ( .B1(n20063), .B2(n18156), .A(n18150), .ZN(P2_U2939) );
  INV_X1 U20061 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18152) );
  AOI22_X1 U20062 ( .A1(n18154), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18151) );
  OAI21_X1 U20063 ( .B1(n18152), .B2(n18156), .A(n18151), .ZN(P2_U2938) );
  INV_X1 U20064 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U20065 ( .A1(n18154), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18153) );
  OAI21_X1 U20066 ( .B1(n20057), .B2(n18156), .A(n18153), .ZN(P2_U2937) );
  AOI22_X1 U20067 ( .A1(n18154), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18145), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18155) );
  OAI21_X1 U20068 ( .B1(n18157), .B2(n18156), .A(n18155), .ZN(P2_U2936) );
  AOI21_X1 U20069 ( .B1(n22455), .B2(n18158), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18159) );
  AOI21_X1 U20070 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n22449), .A(n18159), 
        .ZN(P2_U2817) );
  NOR2_X1 U20071 ( .A1(n18186), .A2(n22461), .ZN(n18191) );
  CLKBUF_X1 U20072 ( .A(n18191), .Z(n22446) );
  AOI222_X1 U20073 ( .A1(n18192), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_1__SCAN_IN), 
        .C2(n22446), .ZN(n18160) );
  INV_X1 U20074 ( .A(n18160), .ZN(P2_U3212) );
  AOI222_X1 U20075 ( .A1(n18192), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_2__SCAN_IN), 
        .C2(n18191), .ZN(n18161) );
  INV_X1 U20076 ( .A(n18161), .ZN(P2_U3213) );
  AOI222_X1 U20077 ( .A1(n18184), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_3__SCAN_IN), 
        .C2(n18191), .ZN(n18162) );
  INV_X1 U20078 ( .A(n18162), .ZN(P2_U3214) );
  AOI222_X1 U20079 ( .A1(n18192), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_4__SCAN_IN), 
        .C2(n18191), .ZN(n18163) );
  INV_X1 U20080 ( .A(n18163), .ZN(P2_U3215) );
  AOI222_X1 U20081 ( .A1(n18184), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_5__SCAN_IN), 
        .C2(n22446), .ZN(n18164) );
  INV_X1 U20082 ( .A(n18164), .ZN(P2_U3216) );
  AOI222_X1 U20083 ( .A1(n18192), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_6__SCAN_IN), 
        .C2(n22446), .ZN(n18165) );
  INV_X1 U20084 ( .A(n18165), .ZN(P2_U3217) );
  AOI222_X1 U20085 ( .A1(n18192), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_7__SCAN_IN), 
        .C2(n22446), .ZN(n18166) );
  INV_X1 U20086 ( .A(n18166), .ZN(P2_U3218) );
  AOI222_X1 U20087 ( .A1(n18192), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_8__SCAN_IN), 
        .C2(n22446), .ZN(n18167) );
  INV_X1 U20088 ( .A(n18167), .ZN(P2_U3219) );
  AOI222_X1 U20089 ( .A1(n22446), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_ADDRESS_REG_8__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_10__SCAN_IN), 
        .C2(n18184), .ZN(n18168) );
  INV_X1 U20090 ( .A(n18168), .ZN(P2_U3220) );
  AOI222_X1 U20091 ( .A1(n22446), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_ADDRESS_REG_9__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_11__SCAN_IN), 
        .C2(n18192), .ZN(n18169) );
  INV_X1 U20092 ( .A(n18169), .ZN(P2_U3221) );
  AOI222_X1 U20093 ( .A1(n18191), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_ADDRESS_REG_10__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_12__SCAN_IN), 
        .C2(n18184), .ZN(n18170) );
  INV_X1 U20094 ( .A(n18170), .ZN(P2_U3222) );
  AOI222_X1 U20095 ( .A1(n18191), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_ADDRESS_REG_11__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_13__SCAN_IN), 
        .C2(n18192), .ZN(n18171) );
  INV_X1 U20096 ( .A(n18171), .ZN(P2_U3223) );
  AOI222_X1 U20097 ( .A1(n18191), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_ADDRESS_REG_12__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_14__SCAN_IN), 
        .C2(n18184), .ZN(n18172) );
  INV_X1 U20098 ( .A(n18172), .ZN(P2_U3224) );
  AOI222_X1 U20099 ( .A1(n18191), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_ADDRESS_REG_13__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_15__SCAN_IN), 
        .C2(n18184), .ZN(n18173) );
  INV_X1 U20100 ( .A(n18173), .ZN(P2_U3225) );
  AOI222_X1 U20101 ( .A1(n22446), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_ADDRESS_REG_14__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_16__SCAN_IN), 
        .C2(n18184), .ZN(n18174) );
  INV_X1 U20102 ( .A(n18174), .ZN(P2_U3226) );
  AOI222_X1 U20103 ( .A1(n18191), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_ADDRESS_REG_15__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_17__SCAN_IN), 
        .C2(n18184), .ZN(n18175) );
  INV_X1 U20104 ( .A(n18175), .ZN(P2_U3227) );
  AOI222_X1 U20105 ( .A1(n22446), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_ADDRESS_REG_16__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_18__SCAN_IN), 
        .C2(n18184), .ZN(n18176) );
  INV_X1 U20106 ( .A(n18176), .ZN(P2_U3228) );
  AOI222_X1 U20107 ( .A1(n18192), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_ADDRESS_REG_17__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_18__SCAN_IN), 
        .C2(n22446), .ZN(n18177) );
  INV_X1 U20108 ( .A(n18177), .ZN(P2_U3229) );
  AOI222_X1 U20109 ( .A1(n22446), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_ADDRESS_REG_18__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_20__SCAN_IN), 
        .C2(n18184), .ZN(n18178) );
  INV_X1 U20110 ( .A(n18178), .ZN(P2_U3230) );
  AOI222_X1 U20111 ( .A1(n18192), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_20__SCAN_IN), 
        .C2(n22446), .ZN(n18179) );
  INV_X1 U20112 ( .A(n18179), .ZN(P2_U3231) );
  AOI222_X1 U20113 ( .A1(n18192), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_ADDRESS_REG_20__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_21__SCAN_IN), 
        .C2(n22446), .ZN(n18180) );
  INV_X1 U20114 ( .A(n18180), .ZN(P2_U3232) );
  AOI222_X1 U20115 ( .A1(n18192), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_ADDRESS_REG_21__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_22__SCAN_IN), 
        .C2(n22446), .ZN(n18181) );
  INV_X1 U20116 ( .A(n18181), .ZN(P2_U3233) );
  AOI222_X1 U20117 ( .A1(n18192), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_ADDRESS_REG_22__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_23__SCAN_IN), 
        .C2(n22446), .ZN(n18182) );
  INV_X1 U20118 ( .A(n18182), .ZN(P2_U3234) );
  AOI222_X1 U20119 ( .A1(n18192), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_ADDRESS_REG_23__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_24__SCAN_IN), 
        .C2(n22446), .ZN(n18183) );
  INV_X1 U20120 ( .A(n18183), .ZN(P2_U3235) );
  AOI222_X1 U20121 ( .A1(n22446), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_ADDRESS_REG_24__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_26__SCAN_IN), 
        .C2(n18184), .ZN(n18185) );
  INV_X1 U20122 ( .A(n18185), .ZN(P2_U3236) );
  AOI222_X1 U20123 ( .A1(n18192), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_ADDRESS_REG_25__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_26__SCAN_IN), 
        .C2(n18191), .ZN(n18187) );
  INV_X1 U20124 ( .A(n18187), .ZN(P2_U3237) );
  AOI222_X1 U20125 ( .A1(n22446), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_ADDRESS_REG_26__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_28__SCAN_IN), 
        .C2(n18192), .ZN(n18188) );
  INV_X1 U20126 ( .A(n18188), .ZN(P2_U3238) );
  AOI222_X1 U20127 ( .A1(n18192), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_27__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_28__SCAN_IN), 
        .C2(n18191), .ZN(n18189) );
  INV_X1 U20128 ( .A(n18189), .ZN(P2_U3239) );
  AOI222_X1 U20129 ( .A1(n22446), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_28__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_30__SCAN_IN), 
        .C2(n18192), .ZN(n18190) );
  INV_X1 U20130 ( .A(n18190), .ZN(P2_U3240) );
  AOI222_X1 U20131 ( .A1(n18192), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n18186), .C1(P2_REIP_REG_30__SCAN_IN), 
        .C2(n18191), .ZN(n18193) );
  INV_X1 U20132 ( .A(n18193), .ZN(P2_U3241) );
  INV_X1 U20133 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n18194) );
  AOI22_X1 U20134 ( .A1(n22449), .A2(n18195), .B1(n18194), .B2(n18186), .ZN(
        P2_U3588) );
  INV_X1 U20135 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n18196) );
  AOI22_X1 U20136 ( .A1(n22449), .A2(n18197), .B1(n18196), .B2(n18186), .ZN(
        P2_U3587) );
  MUX2_X1 U20137 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n22449), .Z(P2_U3586) );
  INV_X1 U20138 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U20139 ( .A1(n22449), .A2(n18199), .B1(n18198), .B2(n18186), .ZN(
        P2_U3585) );
  NAND3_X1 U20140 ( .A1(n21435), .A2(n21656), .A3(n18200), .ZN(n18201) );
  NAND3_X1 U20141 ( .A1(n21431), .A2(n21641), .A3(n21428), .ZN(n18562) );
  NAND2_X1 U20142 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18564) );
  NOR2_X1 U20143 ( .A1(n18203), .A2(n18564), .ZN(n18204) );
  NAND3_X1 U20144 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n18204), .ZN(n18342) );
  NOR2_X1 U20145 ( .A1(n18562), .A2(n18342), .ZN(n18230) );
  INV_X1 U20146 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n21037) );
  NOR2_X1 U20147 ( .A1(n21533), .A2(n18562), .ZN(n18568) );
  NAND2_X1 U20148 ( .A1(n18204), .A2(n18568), .ZN(n18210) );
  NOR2_X1 U20149 ( .A1(n21037), .A2(n18210), .ZN(n18209) );
  AOI21_X1 U20150 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18565), .A(n18209), .ZN(
        n18205) );
  INV_X1 U20151 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18646) );
  OAI22_X1 U20152 ( .A1(n18230), .A2(n18205), .B1(n18646), .B2(n18565), .ZN(
        P3_U2699) );
  INV_X1 U20153 ( .A(n18210), .ZN(n18206) );
  AOI21_X1 U20154 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18565), .A(n18206), .ZN(
        n18208) );
  INV_X1 U20155 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18207) );
  OAI22_X1 U20156 ( .A1(n18209), .A2(n18208), .B1(n18207), .B2(n18565), .ZN(
        P3_U2700) );
  INV_X1 U20157 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18614) );
  INV_X1 U20158 ( .A(n18564), .ZN(n18211) );
  OAI221_X1 U20159 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n18572), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n18211), .A(n18210), .ZN(n18212) );
  AOI22_X1 U20160 ( .A1(n18569), .A2(n18614), .B1(n18212), .B2(n18565), .ZN(
        P3_U2701) );
  AOI22_X1 U20161 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U20162 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18215) );
  AOI22_X1 U20163 ( .A1(n18665), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18214) );
  AOI22_X1 U20164 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18213) );
  NAND4_X1 U20165 ( .A1(n18216), .A2(n18215), .A3(n18214), .A4(n18213), .ZN(
        n18222) );
  AOI22_X1 U20166 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18220) );
  AOI22_X1 U20167 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18219) );
  AOI22_X1 U20168 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U20169 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18217) );
  NAND4_X1 U20170 ( .A1(n18220), .A2(n18219), .A3(n18218), .A4(n18217), .ZN(
        n18221) );
  NOR2_X1 U20171 ( .A1(n18222), .A2(n18221), .ZN(n21604) );
  NAND3_X1 U20172 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n18341) );
  INV_X1 U20173 ( .A(n18230), .ZN(n18225) );
  NOR2_X1 U20174 ( .A1(n18341), .A2(n18225), .ZN(n18223) );
  NAND2_X1 U20175 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18223), .ZN(n18261) );
  OAI21_X1 U20176 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n18223), .A(n18261), .ZN(
        n18224) );
  AOI22_X1 U20177 ( .A1(n18569), .A2(n21604), .B1(n18224), .B2(n18565), .ZN(
        P3_U2695) );
  NOR2_X1 U20178 ( .A1(n21068), .A2(n18225), .ZN(n18233) );
  NAND2_X1 U20179 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18233), .ZN(n18228) );
  INV_X1 U20180 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n21090) );
  OAI21_X1 U20181 ( .B1(n18569), .B2(n21090), .A(n18228), .ZN(n18226) );
  OAI221_X1 U20182 ( .B1(n21435), .B2(n18228), .C1(n18228), .C2(n21090), .A(
        n18226), .ZN(n18227) );
  OAI21_X1 U20183 ( .B1(n18402), .B2(n18565), .A(n18227), .ZN(P3_U2696) );
  OAI211_X1 U20184 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18233), .A(n18228), .B(
        n18565), .ZN(n18229) );
  OAI21_X1 U20185 ( .B1(n18565), .B2(n18662), .A(n18229), .ZN(P3_U2697) );
  OAI21_X1 U20186 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18230), .A(n18565), .ZN(
        n18232) );
  INV_X1 U20187 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18231) );
  OAI22_X1 U20188 ( .A1(n18233), .A2(n18232), .B1(n18231), .B2(n18565), .ZN(
        P3_U2698) );
  AOI22_X1 U20189 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U20190 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18236) );
  AOI22_X1 U20191 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18235) );
  AOI22_X1 U20192 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18234) );
  NAND4_X1 U20193 ( .A1(n18237), .A2(n18236), .A3(n18235), .A4(n18234), .ZN(
        n18244) );
  AOI22_X1 U20194 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U20195 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18241) );
  BUF_X2 U20196 ( .A(n18238), .Z(n18658) );
  AOI22_X1 U20197 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18240) );
  AOI22_X1 U20198 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18239) );
  NAND4_X1 U20199 ( .A1(n18242), .A2(n18241), .A3(n18240), .A4(n18239), .ZN(
        n18243) );
  NOR2_X1 U20200 ( .A1(n18244), .A2(n18243), .ZN(n21584) );
  INV_X1 U20201 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n21194) );
  INV_X1 U20202 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n21177) );
  NAND3_X1 U20203 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .ZN(n18262) );
  NOR4_X1 U20204 ( .A1(n21194), .A2(n21177), .A3(n21117), .A4(n18262), .ZN(
        n18259) );
  NAND2_X1 U20205 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n18259), .ZN(n18343) );
  NOR2_X1 U20206 ( .A1(n18343), .A2(n18261), .ZN(n18245) );
  NOR2_X1 U20207 ( .A1(n18569), .A2(n18245), .ZN(n18258) );
  NOR4_X1 U20208 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n21533), .A3(n18343), .A4(
        n18261), .ZN(n18246) );
  AOI21_X1 U20209 ( .B1(n18258), .B2(P3_EBX_REG_16__SCAN_IN), .A(n18246), .ZN(
        n18247) );
  OAI21_X1 U20210 ( .B1(n21584), .B2(n18565), .A(n18247), .ZN(P3_U2687) );
  AOI22_X1 U20211 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18251) );
  AOI22_X1 U20212 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18250) );
  AOI22_X1 U20213 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18249) );
  AOI22_X1 U20214 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18248) );
  NAND4_X1 U20215 ( .A1(n18251), .A2(n18250), .A3(n18249), .A4(n18248), .ZN(
        n18257) );
  AOI22_X1 U20216 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18255) );
  AOI22_X1 U20217 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18254) );
  AOI22_X1 U20218 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18253) );
  AOI22_X1 U20219 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18252) );
  NAND4_X1 U20220 ( .A1(n18255), .A2(n18254), .A3(n18253), .A4(n18252), .ZN(
        n18256) );
  NOR2_X1 U20221 ( .A1(n18257), .A2(n18256), .ZN(n21596) );
  INV_X1 U20222 ( .A(n18261), .ZN(n18338) );
  OAI221_X1 U20223 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n18259), .C1(
        P3_EBX_REG_15__SCAN_IN), .C2(n18338), .A(n18258), .ZN(n18260) );
  OAI21_X1 U20224 ( .B1(n21596), .B2(n18565), .A(n18260), .ZN(P3_U2688) );
  NOR2_X1 U20225 ( .A1(n21117), .A2(n18261), .ZN(n18340) );
  NAND2_X1 U20226 ( .A1(n21435), .A2(n18340), .ZN(n18324) );
  NOR2_X1 U20227 ( .A1(n18262), .A2(n18324), .ZN(n18284) );
  INV_X1 U20228 ( .A(n18284), .ZN(n18297) );
  AOI22_X1 U20229 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18266) );
  AOI22_X1 U20230 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18265) );
  AOI22_X1 U20231 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18264) );
  AOI22_X1 U20232 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18263) );
  NAND4_X1 U20233 ( .A1(n18266), .A2(n18265), .A3(n18264), .A4(n18263), .ZN(
        n18272) );
  AOI22_X1 U20234 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U20235 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18269) );
  AOI22_X1 U20236 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18268) );
  AOI22_X1 U20237 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18267) );
  NAND4_X1 U20238 ( .A1(n18270), .A2(n18269), .A3(n18268), .A4(n18267), .ZN(
        n18271) );
  NOR2_X1 U20239 ( .A1(n18272), .A2(n18271), .ZN(n21440) );
  NAND3_X1 U20240 ( .A1(n18297), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n18565), 
        .ZN(n18273) );
  OAI221_X1 U20241 ( .B1(n18297), .B2(P3_EBX_REG_13__SCAN_IN), .C1(n18565), 
        .C2(n21440), .A(n18273), .ZN(P3_U2690) );
  AOI22_X1 U20242 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18277) );
  AOI22_X1 U20243 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18276) );
  AOI22_X1 U20244 ( .A1(n18665), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U20245 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18274) );
  NAND4_X1 U20246 ( .A1(n18277), .A2(n18276), .A3(n18275), .A4(n18274), .ZN(
        n18283) );
  AOI22_X1 U20247 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18644), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18281) );
  AOI22_X1 U20248 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18280) );
  AOI22_X1 U20249 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18279) );
  AOI22_X1 U20250 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18278) );
  NAND4_X1 U20251 ( .A1(n18281), .A2(n18280), .A3(n18279), .A4(n18278), .ZN(
        n18282) );
  NOR2_X1 U20252 ( .A1(n18283), .A2(n18282), .ZN(n21589) );
  OAI211_X1 U20253 ( .C1(n21177), .C2(n18297), .A(P3_EBX_REG_14__SCAN_IN), .B(
        n18565), .ZN(n18286) );
  NAND3_X1 U20254 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18284), .A3(n21194), 
        .ZN(n18285) );
  OAI211_X1 U20255 ( .C1(n21589), .C2(n18565), .A(n18286), .B(n18285), .ZN(
        P3_U2689) );
  AOI22_X1 U20256 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18290) );
  AOI22_X1 U20257 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18289) );
  AOI22_X1 U20258 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18288) );
  AOI22_X1 U20259 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18287) );
  NAND4_X1 U20260 ( .A1(n18290), .A2(n18289), .A3(n18288), .A4(n18287), .ZN(
        n18296) );
  AOI22_X1 U20261 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18294) );
  AOI22_X1 U20262 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18664), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18293) );
  AOI22_X1 U20263 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18292) );
  AOI22_X1 U20264 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18291) );
  NAND4_X1 U20265 ( .A1(n18294), .A2(n18293), .A3(n18292), .A4(n18291), .ZN(
        n18295) );
  NOR2_X1 U20266 ( .A1(n18296), .A2(n18295), .ZN(n21444) );
  INV_X1 U20267 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n21153) );
  NAND2_X1 U20268 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18340), .ZN(n18325) );
  NOR2_X1 U20269 ( .A1(n21153), .A2(n18325), .ZN(n18312) );
  OAI211_X1 U20270 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n18312), .A(n18297), .B(
        n18565), .ZN(n18298) );
  OAI21_X1 U20271 ( .B1(n21444), .B2(n18565), .A(n18298), .ZN(P3_U2691) );
  AOI22_X1 U20272 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18309) );
  AOI22_X1 U20273 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18308) );
  INV_X1 U20274 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18300) );
  AOI22_X1 U20275 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18299) );
  OAI21_X1 U20276 ( .B1(n18496), .B2(n18300), .A(n18299), .ZN(n18306) );
  AOI22_X1 U20277 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18304) );
  AOI22_X1 U20278 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18303) );
  AOI22_X1 U20279 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18302) );
  AOI22_X1 U20280 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18301) );
  NAND4_X1 U20281 ( .A1(n18304), .A2(n18303), .A3(n18302), .A4(n18301), .ZN(
        n18305) );
  AOI211_X1 U20282 ( .C1(n11158), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n18306), .B(n18305), .ZN(n18307) );
  NAND3_X1 U20283 ( .A1(n18309), .A2(n18308), .A3(n18307), .ZN(n21448) );
  INV_X1 U20284 ( .A(n21448), .ZN(n18313) );
  AOI21_X1 U20285 ( .B1(n21153), .B2(n18325), .A(n18569), .ZN(n18310) );
  INV_X1 U20286 ( .A(n18310), .ZN(n18311) );
  OAI22_X1 U20287 ( .A1(n18313), .A2(n18565), .B1(n18312), .B2(n18311), .ZN(
        P3_U2692) );
  AOI22_X1 U20288 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U20289 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18316) );
  AOI22_X1 U20290 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18315) );
  AOI22_X1 U20291 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18314) );
  NAND4_X1 U20292 ( .A1(n18317), .A2(n18316), .A3(n18315), .A4(n18314), .ZN(
        n18323) );
  AOI22_X1 U20293 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18321) );
  AOI22_X1 U20294 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18320) );
  AOI22_X1 U20295 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18644), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18319) );
  AOI22_X1 U20296 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18318) );
  NAND4_X1 U20297 ( .A1(n18321), .A2(n18320), .A3(n18319), .A4(n18318), .ZN(
        n18322) );
  NOR2_X1 U20298 ( .A1(n18323), .A2(n18322), .ZN(n21452) );
  INV_X1 U20299 ( .A(n18324), .ZN(n18326) );
  OAI21_X1 U20300 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18326), .A(n18325), .ZN(
        n18327) );
  AOI22_X1 U20301 ( .A1(n18569), .A2(n21452), .B1(n18327), .B2(n18565), .ZN(
        P3_U2693) );
  AOI22_X1 U20302 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18331) );
  AOI22_X1 U20303 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18330) );
  AOI22_X1 U20304 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18660), .ZN(n18329) );
  AOI22_X1 U20305 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21043), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18328) );
  NAND4_X1 U20306 ( .A1(n18331), .A2(n18330), .A3(n18329), .A4(n18328), .ZN(
        n18337) );
  AOI22_X1 U20307 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18335) );
  AOI22_X1 U20308 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14377), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n18665), .ZN(n18334) );
  AOI22_X1 U20309 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11163), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n18616), .ZN(n18333) );
  AOI22_X1 U20310 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18658), .ZN(n18332) );
  NAND4_X1 U20311 ( .A1(n18335), .A2(n18334), .A3(n18333), .A4(n18332), .ZN(
        n18336) );
  NOR2_X1 U20312 ( .A1(n18337), .A2(n18336), .ZN(n21459) );
  OAI21_X1 U20313 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18338), .A(n18565), .ZN(
        n18339) );
  OAI22_X1 U20314 ( .A1(n21459), .A2(n18565), .B1(n18340), .B2(n18339), .ZN(
        P3_U2694) );
  INV_X1 U20315 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21405) );
  INV_X1 U20316 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n21240) );
  INV_X1 U20317 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21232) );
  NOR3_X1 U20318 ( .A1(n18343), .A2(n18342), .A3(n18341), .ZN(n18344) );
  NAND3_X1 U20319 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n18344), .ZN(n18560) );
  NOR2_X1 U20320 ( .A1(n21232), .A2(n18560), .ZN(n18559) );
  NAND2_X1 U20321 ( .A1(n18572), .A2(n18559), .ZN(n18533) );
  NAND2_X1 U20322 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18547), .ZN(n18546) );
  INV_X1 U20323 ( .A(n18546), .ZN(n18520) );
  INV_X1 U20324 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21383) );
  INV_X1 U20325 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n18464) );
  INV_X1 U20326 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21283) );
  NAND4_X1 U20327 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n18345)
         );
  NOR4_X1 U20328 ( .A1(n21383), .A2(n18464), .A3(n21283), .A4(n18345), .ZN(
        n18346) );
  NAND4_X1 U20329 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n18446), .A4(n18346), .ZN(n18349) );
  NOR2_X1 U20330 ( .A1(n21405), .A2(n18349), .ZN(n18445) );
  NAND2_X1 U20331 ( .A1(n18565), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18348) );
  NAND2_X1 U20332 ( .A1(n18445), .A2(n21435), .ZN(n18347) );
  OAI22_X1 U20333 ( .A1(n18445), .A2(n18348), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18347), .ZN(P3_U2672) );
  NAND2_X1 U20334 ( .A1(n21405), .A2(n18349), .ZN(n18350) );
  NAND2_X1 U20335 ( .A1(n18350), .A2(n18565), .ZN(n18444) );
  AOI22_X1 U20336 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18354) );
  AOI22_X1 U20337 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18353) );
  AOI22_X1 U20338 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18352) );
  AOI22_X1 U20339 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18351) );
  NAND4_X1 U20340 ( .A1(n18354), .A2(n18353), .A3(n18352), .A4(n18351), .ZN(
        n18360) );
  AOI22_X1 U20341 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18644), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18358) );
  AOI22_X1 U20342 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18357) );
  AOI22_X1 U20343 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18356) );
  AOI22_X1 U20344 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18355) );
  NAND4_X1 U20345 ( .A1(n18358), .A2(n18357), .A3(n18356), .A4(n18355), .ZN(
        n18359) );
  NOR2_X1 U20346 ( .A1(n18360), .A2(n18359), .ZN(n18443) );
  AOI22_X1 U20347 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18364) );
  AOI22_X1 U20348 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18363) );
  AOI22_X1 U20349 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18362) );
  AOI22_X1 U20350 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18361) );
  NAND4_X1 U20351 ( .A1(n18364), .A2(n18363), .A3(n18362), .A4(n18361), .ZN(
        n18370) );
  AOI22_X1 U20352 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18368) );
  AOI22_X1 U20353 ( .A1(n18658), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18367) );
  AOI22_X1 U20354 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18366) );
  AOI22_X1 U20355 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18644), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18365) );
  NAND4_X1 U20356 ( .A1(n18368), .A2(n18367), .A3(n18366), .A4(n18365), .ZN(
        n18369) );
  NOR2_X1 U20357 ( .A1(n18370), .A2(n18369), .ZN(n18470) );
  AOI22_X1 U20358 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18374) );
  AOI22_X1 U20359 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U20360 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18372) );
  AOI22_X1 U20361 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18371) );
  NAND4_X1 U20362 ( .A1(n18374), .A2(n18373), .A3(n18372), .A4(n18371), .ZN(
        n18380) );
  AOI22_X1 U20363 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18378) );
  AOI22_X1 U20364 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18377) );
  AOI22_X1 U20365 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18376) );
  AOI22_X1 U20366 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18375) );
  NAND4_X1 U20367 ( .A1(n18378), .A2(n18377), .A3(n18376), .A4(n18375), .ZN(
        n18379) );
  NOR2_X1 U20368 ( .A1(n18380), .A2(n18379), .ZN(n18475) );
  AOI22_X1 U20369 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18665), .ZN(n18384) );
  AOI22_X1 U20370 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14377), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18663), .ZN(n18383) );
  AOI22_X1 U20371 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18382) );
  AOI22_X1 U20372 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18660), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18381) );
  NAND4_X1 U20373 ( .A1(n18384), .A2(n18383), .A3(n18382), .A4(n18381), .ZN(
        n18390) );
  AOI22_X1 U20374 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11163), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18388) );
  AOI22_X1 U20375 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18644), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18387) );
  AOI22_X1 U20376 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18616), .ZN(n18386) );
  AOI22_X1 U20377 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18385) );
  NAND4_X1 U20378 ( .A1(n18388), .A2(n18387), .A3(n18386), .A4(n18385), .ZN(
        n18389) );
  NOR2_X1 U20379 ( .A1(n18390), .A2(n18389), .ZN(n18485) );
  AOI22_X1 U20380 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18400) );
  AOI22_X1 U20381 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18399) );
  INV_X1 U20382 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18681) );
  AOI22_X1 U20383 ( .A1(n14377), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18391) );
  OAI21_X1 U20384 ( .B1(n18433), .B2(n18681), .A(n18391), .ZN(n18397) );
  AOI22_X1 U20385 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18395) );
  AOI22_X1 U20386 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18394) );
  AOI22_X1 U20387 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18393) );
  AOI22_X1 U20388 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18392) );
  NAND4_X1 U20389 ( .A1(n18395), .A2(n18394), .A3(n18393), .A4(n18392), .ZN(
        n18396) );
  AOI211_X1 U20390 ( .C1(n18648), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n18397), .B(n18396), .ZN(n18398) );
  NAND3_X1 U20391 ( .A1(n18400), .A2(n18399), .A3(n18398), .ZN(n18490) );
  AOI22_X1 U20392 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18664), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18411) );
  AOI22_X1 U20393 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18410) );
  AOI22_X1 U20394 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18401) );
  OAI21_X1 U20395 ( .B1(n18496), .B2(n18402), .A(n18401), .ZN(n18408) );
  AOI22_X1 U20396 ( .A1(n14377), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18406) );
  AOI22_X1 U20397 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18405) );
  AOI22_X1 U20398 ( .A1(n18665), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18404) );
  AOI22_X1 U20399 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18403) );
  NAND4_X1 U20400 ( .A1(n18406), .A2(n18405), .A3(n18404), .A4(n18403), .ZN(
        n18407) );
  AOI211_X1 U20401 ( .C1(n11163), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n18408), .B(n18407), .ZN(n18409) );
  NAND3_X1 U20402 ( .A1(n18411), .A2(n18410), .A3(n18409), .ZN(n18491) );
  NAND2_X1 U20403 ( .A1(n18490), .A2(n18491), .ZN(n18489) );
  NOR2_X1 U20404 ( .A1(n18485), .A2(n18489), .ZN(n18484) );
  AOI22_X1 U20405 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18421) );
  AOI22_X1 U20406 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18420) );
  AOI22_X1 U20407 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18412) );
  OAI21_X1 U20408 ( .B1(n18433), .B2(n18614), .A(n18412), .ZN(n18418) );
  AOI22_X1 U20409 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18416) );
  AOI22_X1 U20410 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18415) );
  AOI22_X1 U20411 ( .A1(n14377), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18414) );
  AOI22_X1 U20412 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18413) );
  NAND4_X1 U20413 ( .A1(n18416), .A2(n18415), .A3(n18414), .A4(n18413), .ZN(
        n18417) );
  AOI211_X1 U20414 ( .C1(n11164), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n18418), .B(n18417), .ZN(n18419) );
  NAND3_X1 U20415 ( .A1(n18421), .A2(n18420), .A3(n18419), .ZN(n18481) );
  NAND2_X1 U20416 ( .A1(n18484), .A2(n18481), .ZN(n18480) );
  NOR2_X1 U20417 ( .A1(n18475), .A2(n18480), .ZN(n18474) );
  AOI22_X1 U20418 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18431) );
  AOI22_X1 U20419 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U20420 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18422) );
  OAI21_X1 U20421 ( .B1(n18433), .B2(n18646), .A(n18422), .ZN(n18428) );
  AOI22_X1 U20422 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18426) );
  AOI22_X1 U20423 ( .A1(n18658), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18425) );
  AOI22_X1 U20424 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18424) );
  AOI22_X1 U20425 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18423) );
  NAND4_X1 U20426 ( .A1(n18426), .A2(n18425), .A3(n18424), .A4(n18423), .ZN(
        n18427) );
  AOI211_X1 U20427 ( .C1(n11158), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n18428), .B(n18427), .ZN(n18429) );
  NAND3_X1 U20428 ( .A1(n18431), .A2(n18430), .A3(n18429), .ZN(n18460) );
  NAND2_X1 U20429 ( .A1(n18474), .A2(n18460), .ZN(n18469) );
  NOR2_X1 U20430 ( .A1(n18470), .A2(n18469), .ZN(n18468) );
  AOI22_X1 U20431 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18442) );
  AOI22_X1 U20432 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18441) );
  AOI22_X1 U20433 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18432) );
  OAI21_X1 U20434 ( .B1(n18433), .B2(n18662), .A(n18432), .ZN(n18439) );
  AOI22_X1 U20435 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18437) );
  AOI22_X1 U20436 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18436) );
  AOI22_X1 U20437 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18679), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18435) );
  AOI22_X1 U20438 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18434) );
  NAND4_X1 U20439 ( .A1(n18437), .A2(n18436), .A3(n18435), .A4(n18434), .ZN(
        n18438) );
  AOI211_X1 U20440 ( .C1(n11164), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n18439), .B(n18438), .ZN(n18440) );
  NAND3_X1 U20441 ( .A1(n18442), .A2(n18441), .A3(n18440), .ZN(n18463) );
  NAND2_X1 U20442 ( .A1(n18468), .A2(n18463), .ZN(n18462) );
  XNOR2_X1 U20443 ( .A(n18443), .B(n18462), .ZN(n21551) );
  OAI22_X1 U20444 ( .A1(n18445), .A2(n18444), .B1(n21551), .B2(n18565), .ZN(
        P3_U2673) );
  NAND2_X1 U20445 ( .A1(n21435), .A2(n18446), .ZN(n18459) );
  NOR2_X1 U20446 ( .A1(n18569), .A2(n18446), .ZN(n18519) );
  AOI22_X1 U20447 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18450) );
  AOI22_X1 U20448 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18449) );
  AOI22_X1 U20449 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18448) );
  AOI22_X1 U20450 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18447) );
  NAND4_X1 U20451 ( .A1(n18450), .A2(n18449), .A3(n18448), .A4(n18447), .ZN(
        n18456) );
  AOI22_X1 U20452 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14377), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18454) );
  AOI22_X1 U20453 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18453) );
  AOI22_X1 U20454 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18452) );
  AOI22_X1 U20455 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18451) );
  NAND4_X1 U20456 ( .A1(n18454), .A2(n18453), .A3(n18452), .A4(n18451), .ZN(
        n18455) );
  NOR2_X1 U20457 ( .A1(n18456), .A2(n18455), .ZN(n21499) );
  INV_X1 U20458 ( .A(n21499), .ZN(n18457) );
  AOI22_X1 U20459 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18519), .B1(n18569), 
        .B2(n18457), .ZN(n18458) );
  OAI21_X1 U20460 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18459), .A(n18458), .ZN(
        P3_U2682) );
  INV_X1 U20461 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21331) );
  NOR2_X1 U20462 ( .A1(n21283), .A2(n18459), .ZN(n18494) );
  NAND2_X1 U20463 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18493), .ZN(n18479) );
  NAND2_X1 U20464 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n18478), .ZN(n18473) );
  AOI21_X1 U20465 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18565), .A(n18478), .ZN(
        n18461) );
  OAI21_X1 U20466 ( .B1(n18474), .B2(n18460), .A(n18469), .ZN(n21567) );
  OAI22_X1 U20467 ( .A1(n18465), .A2(n18461), .B1(n21567), .B2(n18565), .ZN(
        P3_U2676) );
  OAI21_X1 U20468 ( .B1(n18468), .B2(n18463), .A(n18462), .ZN(n21555) );
  NOR2_X1 U20469 ( .A1(n18569), .A2(n18465), .ZN(n18471) );
  OAI221_X1 U20470 ( .B1(n18471), .B2(n18568), .C1(n18471), .C2(n18464), .A(
        P3_EBX_REG_29__SCAN_IN), .ZN(n18467) );
  NAND3_X1 U20471 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18465), .A3(n21383), 
        .ZN(n18466) );
  OAI211_X1 U20472 ( .C1(n18565), .C2(n21555), .A(n18467), .B(n18466), .ZN(
        P3_U2674) );
  AOI21_X1 U20473 ( .B1(n18470), .B2(n18469), .A(n18468), .ZN(n21556) );
  AOI22_X1 U20474 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18471), .B1(n21556), 
        .B2(n18569), .ZN(n18472) );
  OAI21_X1 U20475 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n18473), .A(n18472), .ZN(
        P3_U2675) );
  AOI21_X1 U20476 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18565), .A(n18483), .ZN(
        n18477) );
  AOI21_X1 U20477 ( .B1(n18475), .B2(n18480), .A(n18474), .ZN(n21538) );
  INV_X1 U20478 ( .A(n21538), .ZN(n18476) );
  OAI22_X1 U20479 ( .A1(n18478), .A2(n18477), .B1(n18476), .B2(n18565), .ZN(
        P3_U2677) );
  INV_X1 U20480 ( .A(n18479), .ZN(n18488) );
  AOI21_X1 U20481 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18565), .A(n18488), .ZN(
        n18482) );
  OAI21_X1 U20482 ( .B1(n18484), .B2(n18481), .A(n18480), .ZN(n21537) );
  OAI22_X1 U20483 ( .A1(n18483), .A2(n18482), .B1(n18565), .B2(n21537), .ZN(
        P3_U2678) );
  AOI21_X1 U20484 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18565), .A(n18493), .ZN(
        n18487) );
  AOI21_X1 U20485 ( .B1(n18485), .B2(n18489), .A(n18484), .ZN(n21568) );
  INV_X1 U20486 ( .A(n21568), .ZN(n18486) );
  OAI22_X1 U20487 ( .A1(n18488), .A2(n18487), .B1(n18565), .B2(n18486), .ZN(
        P3_U2679) );
  AOI21_X1 U20488 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18565), .A(n18508), .ZN(
        n18492) );
  OAI21_X1 U20489 ( .B1(n18491), .B2(n18490), .A(n18489), .ZN(n21578) );
  OAI22_X1 U20490 ( .A1(n18493), .A2(n18492), .B1(n18565), .B2(n21578), .ZN(
        P3_U2680) );
  AOI21_X1 U20491 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18565), .A(n18494), .ZN(
        n18507) );
  AOI22_X1 U20492 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18505) );
  AOI22_X1 U20493 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18504) );
  AOI22_X1 U20494 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18495) );
  OAI21_X1 U20495 ( .B1(n18496), .B2(n18662), .A(n18495), .ZN(n18502) );
  AOI22_X1 U20496 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18500) );
  AOI22_X1 U20497 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18499) );
  AOI22_X1 U20498 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18498) );
  AOI22_X1 U20499 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18497) );
  NAND4_X1 U20500 ( .A1(n18500), .A2(n18499), .A3(n18498), .A4(n18497), .ZN(
        n18501) );
  AOI211_X1 U20501 ( .C1(n18678), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n18502), .B(n18501), .ZN(n18503) );
  NAND3_X1 U20502 ( .A1(n18505), .A2(n18504), .A3(n18503), .ZN(n21510) );
  INV_X1 U20503 ( .A(n21510), .ZN(n18506) );
  OAI22_X1 U20504 ( .A1(n18508), .A2(n18507), .B1(n18506), .B2(n18565), .ZN(
        P3_U2681) );
  AOI22_X1 U20505 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18512) );
  AOI22_X1 U20506 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18511) );
  AOI22_X1 U20507 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18510) );
  AOI22_X1 U20508 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18509) );
  NAND4_X1 U20509 ( .A1(n18512), .A2(n18511), .A3(n18510), .A4(n18509), .ZN(
        n18518) );
  AOI22_X1 U20510 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18516) );
  AOI22_X1 U20511 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18515) );
  AOI22_X1 U20512 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18514) );
  AOI22_X1 U20513 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18513) );
  NAND4_X1 U20514 ( .A1(n18516), .A2(n18515), .A3(n18514), .A4(n18513), .ZN(
        n18517) );
  NOR2_X1 U20515 ( .A1(n18518), .A2(n18517), .ZN(n21505) );
  OAI21_X1 U20516 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18520), .A(n18519), .ZN(
        n18521) );
  OAI21_X1 U20517 ( .B1(n21505), .B2(n18565), .A(n18521), .ZN(P3_U2683) );
  AOI22_X1 U20518 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18525) );
  AOI22_X1 U20519 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14377), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18524) );
  AOI22_X1 U20520 ( .A1(n18665), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18523) );
  AOI22_X1 U20521 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18522) );
  NAND4_X1 U20522 ( .A1(n18525), .A2(n18524), .A3(n18523), .A4(n18522), .ZN(
        n18531) );
  AOI22_X1 U20523 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18529) );
  AOI22_X1 U20524 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18528) );
  AOI22_X1 U20525 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18527) );
  AOI22_X1 U20526 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18526) );
  NAND4_X1 U20527 ( .A1(n18529), .A2(n18528), .A3(n18527), .A4(n18526), .ZN(
        n18530) );
  NOR2_X1 U20528 ( .A1(n18531), .A2(n18530), .ZN(n21525) );
  INV_X1 U20529 ( .A(n18533), .ZN(n18532) );
  OAI33_X1 U20530 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n21533), .A3(n18533), 
        .B1(n21240), .B2(n18569), .B3(n18532), .ZN(n18534) );
  INV_X1 U20531 ( .A(n18534), .ZN(n18535) );
  OAI21_X1 U20532 ( .B1(n21525), .B2(n18565), .A(n18535), .ZN(P3_U2685) );
  AOI22_X1 U20533 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18539) );
  AOI22_X1 U20534 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18538) );
  AOI22_X1 U20535 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18537) );
  AOI22_X1 U20536 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18536) );
  NAND4_X1 U20537 ( .A1(n18539), .A2(n18538), .A3(n18537), .A4(n18536), .ZN(
        n18545) );
  AOI22_X1 U20538 ( .A1(n18658), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18543) );
  AOI22_X1 U20539 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18542) );
  AOI22_X1 U20540 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18541) );
  AOI22_X1 U20541 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18540) );
  NAND4_X1 U20542 ( .A1(n18543), .A2(n18542), .A3(n18541), .A4(n18540), .ZN(
        n18544) );
  NOR2_X1 U20543 ( .A1(n18545), .A2(n18544), .ZN(n21519) );
  OAI21_X1 U20544 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18547), .A(n18546), .ZN(
        n18548) );
  AOI22_X1 U20545 ( .A1(n18569), .A2(n21519), .B1(n18548), .B2(n18565), .ZN(
        P3_U2684) );
  AOI22_X1 U20546 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n18616), .ZN(n18552) );
  AOI22_X1 U20547 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18665), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18551) );
  AOI22_X1 U20548 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18660), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18550) );
  AOI22_X1 U20549 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n21043), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n18679), .ZN(n18549) );
  NAND4_X1 U20550 ( .A1(n18552), .A2(n18551), .A3(n18550), .A4(n18549), .ZN(
        n18558) );
  AOI22_X1 U20551 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11164), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n18658), .ZN(n18556) );
  AOI22_X1 U20552 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n18659), .ZN(n18555) );
  AOI22_X1 U20553 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18663), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18554) );
  AOI22_X1 U20554 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18553) );
  NAND4_X1 U20555 ( .A1(n18556), .A2(n18555), .A3(n18554), .A4(n18553), .ZN(
        n18557) );
  NOR2_X1 U20556 ( .A1(n18558), .A2(n18557), .ZN(n21530) );
  AOI21_X1 U20557 ( .B1(n21232), .B2(n18560), .A(n18559), .ZN(n18561) );
  AOI22_X1 U20558 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18562), .B1(n18568), 
        .B2(n18561), .ZN(n18563) );
  OAI21_X1 U20559 ( .B1(n21530), .B2(n18565), .A(n18563), .ZN(P3_U2686) );
  OAI21_X1 U20560 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18564), .ZN(n21024) );
  INV_X1 U20561 ( .A(n18568), .ZN(n18567) );
  OAI222_X1 U20562 ( .A1(n21024), .A2(n18567), .B1(n18566), .B2(n18572), .C1(
        n18629), .C2(n18565), .ZN(P3_U2702) );
  AOI22_X1 U20563 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18569), .B1(
        n18568), .B2(n18571), .ZN(n18570) );
  OAI21_X1 U20564 ( .B1(n18572), .B2(n18571), .A(n18570), .ZN(P3_U2703) );
  INV_X1 U20565 ( .A(n18573), .ZN(n18575) );
  OAI21_X1 U20566 ( .B1(n18575), .B2(n18574), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18576) );
  OAI21_X1 U20567 ( .B1(n18577), .B2(n22095), .A(n18576), .ZN(P3_U2634) );
  INV_X1 U20568 ( .A(n19153), .ZN(n18581) );
  OAI21_X1 U20569 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18579), .A(n18578), .ZN(
        n22093) );
  OAI21_X1 U20570 ( .B1(n20957), .B2(n18581), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18580) );
  OAI221_X1 U20571 ( .B1(n18581), .B2(n22093), .C1(n18581), .C2(n19627), .A(
        n18580), .ZN(P3_U2863) );
  AOI22_X1 U20572 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11164), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18585) );
  AOI22_X1 U20573 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18584) );
  AOI22_X1 U20574 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18583) );
  AOI22_X1 U20575 ( .A1(n21043), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18582) );
  NAND4_X1 U20576 ( .A1(n18585), .A2(n18584), .A3(n18583), .A4(n18582), .ZN(
        n18591) );
  AOI22_X1 U20577 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18589) );
  AOI22_X1 U20578 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18588) );
  AOI22_X1 U20579 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18587) );
  AOI22_X1 U20580 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18586) );
  NAND4_X1 U20581 ( .A1(n18589), .A2(n18588), .A3(n18587), .A4(n18586), .ZN(
        n18590) );
  AOI22_X1 U20582 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18595) );
  AOI22_X1 U20583 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18594) );
  AOI22_X1 U20584 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18593) );
  AOI22_X1 U20585 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18592) );
  NAND4_X1 U20586 ( .A1(n18595), .A2(n18594), .A3(n18593), .A4(n18592), .ZN(
        n18601) );
  AOI22_X1 U20587 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18599) );
  AOI22_X1 U20588 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18598) );
  AOI22_X1 U20589 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18597) );
  AOI22_X1 U20590 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18596) );
  NAND4_X1 U20591 ( .A1(n18599), .A2(n18598), .A3(n18597), .A4(n18596), .ZN(
        n18600) );
  AOI22_X1 U20592 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18605) );
  AOI22_X1 U20593 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18604) );
  AOI22_X1 U20594 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18603) );
  AOI22_X1 U20595 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n21043), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18602) );
  NAND4_X1 U20596 ( .A1(n18605), .A2(n18604), .A3(n18603), .A4(n18602), .ZN(
        n18611) );
  AOI22_X1 U20597 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18648), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18609) );
  AOI22_X1 U20598 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18608) );
  AOI22_X1 U20599 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18607) );
  AOI22_X1 U20600 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18606) );
  NAND4_X1 U20601 ( .A1(n18609), .A2(n18608), .A3(n18607), .A4(n18606), .ZN(
        n18610) );
  AOI22_X1 U20602 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18678), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18626) );
  AOI22_X1 U20603 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18625) );
  AOI22_X1 U20604 ( .A1(n18627), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18613) );
  OAI21_X1 U20605 ( .B1(n11293), .B2(n18614), .A(n18613), .ZN(n18623) );
  AOI22_X1 U20606 ( .A1(n18615), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18621) );
  AOI22_X1 U20607 ( .A1(n18634), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18620) );
  AOI22_X1 U20608 ( .A1(n14404), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18631), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18619) );
  AOI22_X1 U20609 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18630), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18618) );
  NAND4_X1 U20610 ( .A1(n18621), .A2(n18620), .A3(n18619), .A4(n18618), .ZN(
        n18622) );
  NAND3_X1 U20611 ( .A1(n18626), .A2(n18625), .A3(n18624), .ZN(n18706) );
  AOI22_X1 U20612 ( .A1(n14404), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n18647), .ZN(n18643) );
  AOI22_X1 U20613 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18663), .ZN(n18642) );
  AOI22_X1 U20614 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18627), .B1(
        n14377), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18628) );
  OAI21_X1 U20615 ( .B1(n18629), .B2(n11293), .A(n18628), .ZN(n18640) );
  AOI22_X1 U20616 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18677), .B1(
        n18630), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18638) );
  AOI22_X1 U20617 ( .A1(n18632), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18631), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18637) );
  AOI22_X1 U20618 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18238), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n18633), .ZN(n18636) );
  AOI22_X1 U20619 ( .A1(n18634), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14372), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18635) );
  NAND4_X1 U20620 ( .A1(n18638), .A2(n18637), .A3(n18636), .A4(n18635), .ZN(
        n18639) );
  AOI211_X1 U20621 ( .C1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .C2(n18660), .A(
        n18640), .B(n18639), .ZN(n18641) );
  NAND3_X1 U20622 ( .A1(n18643), .A2(n18642), .A3(n18641), .ZN(n21606) );
  NAND2_X1 U20623 ( .A1(n18706), .A2(n21606), .ZN(n18715) );
  AOI22_X1 U20624 ( .A1(n18644), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18657) );
  AOI22_X1 U20625 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18659), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18656) );
  AOI22_X1 U20626 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18645) );
  OAI21_X1 U20627 ( .B1(n11293), .B2(n18646), .A(n18645), .ZN(n18654) );
  AOI22_X1 U20628 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18652) );
  AOI22_X1 U20629 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11163), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18651) );
  AOI22_X1 U20630 ( .A1(n18682), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18650) );
  AOI22_X1 U20631 ( .A1(n18648), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18649) );
  NAND4_X1 U20632 ( .A1(n18652), .A2(n18651), .A3(n18650), .A4(n18649), .ZN(
        n18653) );
  AOI211_X1 U20633 ( .C1(n18664), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n18654), .B(n18653), .ZN(n18655) );
  NAND3_X1 U20634 ( .A1(n18657), .A2(n18656), .A3(n18655), .ZN(n18707) );
  NAND2_X1 U20635 ( .A1(n18676), .A2(n18707), .ZN(n18696) );
  AOI22_X1 U20636 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18682), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18675) );
  AOI22_X1 U20637 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18658), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18674) );
  AOI22_X1 U20638 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18661) );
  OAI21_X1 U20639 ( .B1(n11293), .B2(n18662), .A(n18661), .ZN(n18672) );
  AOI22_X1 U20640 ( .A1(n18664), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18670) );
  AOI22_X1 U20641 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18669) );
  AOI22_X1 U20642 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18665), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18668) );
  AOI22_X1 U20643 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18666), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18667) );
  NAND4_X1 U20644 ( .A1(n18670), .A2(n18669), .A3(n18668), .A4(n18667), .ZN(
        n18671) );
  AOI211_X1 U20645 ( .C1(n18648), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n18672), .B(n18671), .ZN(n18673) );
  NAND3_X1 U20646 ( .A1(n18675), .A2(n18674), .A3(n18673), .ZN(n18708) );
  INV_X1 U20647 ( .A(n18707), .ZN(n21475) );
  XNOR2_X1 U20648 ( .A(n21475), .B(n18676), .ZN(n18694) );
  AND2_X1 U20649 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18694), .ZN(
        n18695) );
  INV_X1 U20650 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21699) );
  INV_X1 U20651 ( .A(n18706), .ZN(n21484) );
  INV_X1 U20652 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21691) );
  INV_X1 U20653 ( .A(n21606), .ZN(n18719) );
  XNOR2_X1 U20654 ( .A(n18719), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19133) );
  AOI22_X1 U20655 ( .A1(n11164), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18677), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18689) );
  AOI22_X1 U20656 ( .A1(n18678), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18647), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18688) );
  AOI22_X1 U20657 ( .A1(n18679), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18680) );
  OAI21_X1 U20658 ( .B1(n11293), .B2(n18681), .A(n18680), .ZN(n18686) );
  AOI22_X1 U20659 ( .A1(n18659), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18685) );
  AOI22_X1 U20660 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18632), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18684) );
  AOI22_X1 U20661 ( .A1(n11163), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18663), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18683) );
  NAND3_X1 U20662 ( .A1(n18689), .A2(n18688), .A3(n18687), .ZN(n21610) );
  NAND2_X1 U20663 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21610), .ZN(
        n19142) );
  INV_X1 U20664 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21712) );
  NOR2_X1 U20665 ( .A1(n18691), .A2(n21712), .ZN(n18693) );
  XNOR2_X1 U20666 ( .A(n21712), .B(n18691), .ZN(n19111) );
  XNOR2_X1 U20667 ( .A(n21479), .B(n18715), .ZN(n19110) );
  NOR2_X1 U20668 ( .A1(n19111), .A2(n19110), .ZN(n18692) );
  NOR2_X1 U20669 ( .A1(n18693), .A2(n18692), .ZN(n19102) );
  XNOR2_X1 U20670 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n18694), .ZN(
        n19101) );
  NOR2_X1 U20671 ( .A1(n19102), .A2(n19101), .ZN(n19100) );
  XNOR2_X1 U20672 ( .A(n21470), .B(n18696), .ZN(n18698) );
  NOR2_X1 U20673 ( .A1(n18697), .A2(n18698), .ZN(n18699) );
  INV_X1 U20674 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21730) );
  XNOR2_X1 U20675 ( .A(n18698), .B(n18697), .ZN(n19087) );
  INV_X1 U20676 ( .A(n18708), .ZN(n21466) );
  XNOR2_X1 U20677 ( .A(n21466), .B(n18700), .ZN(n18701) );
  XNOR2_X1 U20678 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n18701), .ZN(
        n19081) );
  OAI21_X1 U20679 ( .B1(n18702), .B2(n21935), .A(n19019), .ZN(n18703) );
  NOR2_X1 U20680 ( .A1(n18767), .A2(n18703), .ZN(n18704) );
  INV_X1 U20681 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21756) );
  INV_X2 U20682 ( .A(n19052), .ZN(n19000) );
  NOR2_X2 U20683 ( .A1(n21641), .A2(n22101), .ZN(n19072) );
  INV_X1 U20684 ( .A(n21610), .ZN(n18717) );
  NOR2_X1 U20685 ( .A1(n18719), .A2(n18717), .ZN(n18718) );
  NOR2_X1 U20686 ( .A1(n21479), .A2(n18714), .ZN(n18723) );
  NAND2_X1 U20687 ( .A1(n18723), .A2(n18707), .ZN(n18711) );
  NOR2_X1 U20688 ( .A1(n21470), .A2(n18711), .ZN(n18710) );
  NAND2_X1 U20689 ( .A1(n18710), .A2(n18708), .ZN(n18709) );
  NOR2_X1 U20690 ( .A1(n21661), .A2(n18709), .ZN(n18733) );
  XNOR2_X1 U20691 ( .A(n21935), .B(n18709), .ZN(n19070) );
  XNOR2_X1 U20692 ( .A(n21466), .B(n18710), .ZN(n18726) );
  XOR2_X1 U20693 ( .A(n21470), .B(n18711), .Z(n18712) );
  NAND2_X1 U20694 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18712), .ZN(
        n18725) );
  XNOR2_X1 U20695 ( .A(n21730), .B(n18712), .ZN(n19092) );
  XOR2_X1 U20696 ( .A(n21479), .B(n18714), .Z(n18713) );
  NAND2_X1 U20697 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18713), .ZN(
        n18721) );
  XOR2_X1 U20698 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18713), .Z(
        n19117) );
  NAND2_X1 U20699 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18716), .ZN(
        n18720) );
  INV_X1 U20700 ( .A(n19133), .ZN(n19135) );
  INV_X1 U20701 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21834) );
  NAND2_X1 U20702 ( .A1(n18717), .A2(n21834), .ZN(n19141) );
  NOR2_X1 U20703 ( .A1(n19135), .A2(n19141), .ZN(n19134) );
  AOI211_X1 U20704 ( .C1(n18719), .C2(n21691), .A(n18718), .B(n19134), .ZN(
        n19125) );
  NAND2_X1 U20705 ( .A1(n19126), .A2(n19125), .ZN(n19124) );
  NAND2_X1 U20706 ( .A1(n18720), .A2(n19124), .ZN(n19116) );
  NAND2_X1 U20707 ( .A1(n19117), .A2(n19116), .ZN(n19115) );
  NAND2_X1 U20708 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18722), .ZN(
        n18724) );
  XNOR2_X1 U20709 ( .A(n21475), .B(n18723), .ZN(n19098) );
  NAND2_X1 U20710 ( .A1(n19092), .A2(n19091), .ZN(n19090) );
  NAND2_X1 U20711 ( .A1(n18726), .A2(n18727), .ZN(n18728) );
  NAND2_X1 U20712 ( .A1(n18733), .A2(n18729), .ZN(n18734) );
  INV_X1 U20713 ( .A(n18729), .ZN(n18732) );
  NAND2_X1 U20714 ( .A1(n19070), .A2(n19069), .ZN(n18731) );
  NAND2_X1 U20715 ( .A1(n18733), .A2(n18732), .ZN(n18730) );
  OAI211_X1 U20716 ( .C1(n18733), .C2(n18732), .A(n18731), .B(n18730), .ZN(
        n19051) );
  NAND2_X1 U20717 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19051), .ZN(
        n19050) );
  INV_X1 U20718 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n22072) );
  NOR2_X1 U20719 ( .A1(n22072), .A2(n22055), .ZN(n21779) );
  NAND2_X1 U20720 ( .A1(n21779), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19013) );
  NAND2_X1 U20721 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21783), .ZN(
        n21798) );
  NOR2_X1 U20722 ( .A1(n21811), .A2(n21798), .ZN(n21822) );
  NAND2_X1 U20723 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21822), .ZN(
        n22022) );
  NOR2_X2 U20724 ( .A1(n19031), .A2(n22022), .ZN(n18988) );
  NOR2_X1 U20725 ( .A1(n22039), .A2(n22028), .ZN(n21658) );
  INV_X1 U20726 ( .A(n21658), .ZN(n22009) );
  INV_X1 U20727 ( .A(n21798), .ZN(n18768) );
  NAND2_X1 U20728 ( .A1(n21766), .A2(n18768), .ZN(n18992) );
  NAND2_X1 U20729 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21820), .ZN(
        n18755) );
  NAND2_X1 U20730 ( .A1(n18768), .A2(n21769), .ZN(n19002) );
  OAI22_X1 U20731 ( .A1(n21812), .A2(n19052), .B1(n18812), .B2(n19148), .ZN(
        n18786) );
  AOI21_X1 U20732 ( .B1(n18988), .B2(n22009), .A(n18786), .ZN(n18991) );
  INV_X1 U20733 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21659) );
  NOR2_X1 U20734 ( .A1(n18736), .A2(n21027), .ZN(n18981) );
  INV_X1 U20735 ( .A(n20957), .ZN(n18735) );
  NAND2_X1 U20736 ( .A1(n19144), .A2(n19105), .ZN(n19078) );
  OAI21_X1 U20737 ( .B1(n19112), .B2(n18736), .A(n19078), .ZN(n18985) );
  OAI21_X1 U20738 ( .B1(n18981), .B2(n19143), .A(n18985), .ZN(n18761) );
  NOR3_X1 U20739 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18889), .A3(
        n18736), .ZN(n18762) );
  INV_X1 U20740 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n22026) );
  INV_X1 U20741 ( .A(n18737), .ZN(n18759) );
  NOR2_X1 U20742 ( .A1(n18759), .A2(n21027), .ZN(n18758) );
  INV_X1 U20743 ( .A(n18758), .ZN(n18738) );
  OAI21_X1 U20744 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18981), .A(
        n18738), .ZN(n21244) );
  OAI22_X1 U20745 ( .A1(n22049), .A2(n22026), .B1(n21244), .B2(n18921), .ZN(
        n18739) );
  AOI211_X1 U20746 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18761), .A(
        n18762), .B(n18739), .ZN(n18751) );
  NOR2_X1 U20747 ( .A1(n21946), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18832) );
  AOI21_X1 U20748 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n21946), .A(
        n18832), .ZN(n18749) );
  NAND2_X1 U20749 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19019), .ZN(
        n18800) );
  NAND2_X1 U20750 ( .A1(n22072), .A2(n22055), .ZN(n19011) );
  NOR4_X1 U20751 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(n19011), .ZN(n18770) );
  NOR2_X1 U20752 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18740) );
  NAND2_X1 U20753 ( .A1(n22013), .A2(n19021), .ZN(n18747) );
  NAND2_X1 U20754 ( .A1(n21946), .A2(n22039), .ZN(n18743) );
  INV_X1 U20755 ( .A(n18746), .ZN(n18748) );
  XNOR2_X1 U20756 ( .A(n18749), .B(n18813), .ZN(n22024) );
  NOR2_X1 U20757 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n22009), .ZN(
        n22023) );
  AOI22_X1 U20758 ( .A1(n19054), .A2(n22024), .B1(n18988), .B2(n22023), .ZN(
        n18750) );
  OAI211_X1 U20759 ( .C1(n18991), .C2(n21659), .A(n18751), .B(n18750), .ZN(
        P3_U2812) );
  INV_X1 U20760 ( .A(n18832), .ZN(n18752) );
  NOR2_X1 U20761 ( .A1(n18752), .A2(n18813), .ZN(n18825) );
  NOR3_X1 U20762 ( .A1(n19019), .A2(n21659), .A3(n18753), .ZN(n18831) );
  NOR2_X1 U20763 ( .A1(n18825), .A2(n18831), .ZN(n18754) );
  INV_X1 U20764 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18842) );
  XNOR2_X1 U20765 ( .A(n18754), .B(n18842), .ZN(n21996) );
  NAND3_X1 U20766 ( .A1(n21658), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18756) );
  NOR2_X1 U20767 ( .A1(n18755), .A2(n18756), .ZN(n21988) );
  NOR2_X1 U20768 ( .A1(n22008), .A2(n18756), .ZN(n21986) );
  OAI22_X1 U20769 ( .A1(n21988), .A2(n19052), .B1(n21986), .B2(n19148), .ZN(
        n18841) );
  NOR2_X1 U20770 ( .A1(n18836), .A2(n21027), .ZN(n18838) );
  INV_X1 U20771 ( .A(n18838), .ZN(n18757) );
  OAI21_X1 U20772 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18758), .A(
        n18757), .ZN(n21251) );
  NOR3_X1 U20773 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18889), .A3(
        n18759), .ZN(n18760) );
  AOI221_X1 U20774 ( .B1(n18762), .B2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(
        n18761), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18760), .ZN(
        n18763) );
  NAND2_X1 U20775 ( .A1(n21869), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21994) );
  OAI211_X1 U20776 ( .C1(n18921), .C2(n21251), .A(n18763), .B(n21994), .ZN(
        n18764) );
  AOI221_X1 U20777 ( .B1(n18885), .B2(n18842), .C1(n18841), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n18764), .ZN(n18765) );
  OAI21_X1 U20778 ( .B1(n21996), .B2(n18961), .A(n18765), .ZN(P3_U2811) );
  INV_X1 U20779 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21829) );
  NAND2_X1 U20780 ( .A1(n19001), .A2(n21829), .ZN(n21824) );
  NAND2_X1 U20781 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18766) );
  NOR3_X1 U20782 ( .A1(n18767), .A2(n19019), .A3(n18766), .ZN(n19039) );
  NAND2_X1 U20783 ( .A1(n18768), .A2(n19039), .ZN(n19003) );
  NAND2_X1 U20784 ( .A1(n18769), .A2(n21756), .ZN(n18791) );
  NAND2_X1 U20785 ( .A1(n18770), .A2(n19040), .ZN(n19004) );
  AOI22_X1 U20786 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19003), .B1(
        n19004), .B2(n21811), .ZN(n18771) );
  XOR2_X1 U20787 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18771), .Z(
        n21825) );
  INV_X1 U20788 ( .A(n18772), .ZN(n21196) );
  NAND2_X1 U20789 ( .A1(n21196), .A2(n18936), .ZN(n18784) );
  NOR2_X1 U20790 ( .A1(n18772), .A2(n21027), .ZN(n18778) );
  OAI21_X1 U20791 ( .B1(n19112), .B2(n18772), .A(n19078), .ZN(n18994) );
  OAI21_X1 U20792 ( .B1(n18778), .B2(n19143), .A(n18994), .ZN(n18781) );
  INV_X1 U20793 ( .A(n18778), .ZN(n18996) );
  XNOR2_X1 U20794 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n18996), .ZN(
        n21197) );
  AOI22_X1 U20795 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18781), .B1(
        n18964), .B2(n21197), .ZN(n18773) );
  NAND2_X1 U20796 ( .A1(n22073), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n21827) );
  OAI211_X1 U20797 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18784), .A(
        n18773), .B(n21827), .ZN(n18774) );
  AOI21_X1 U20798 ( .B1(n19054), .B2(n21825), .A(n18774), .ZN(n18776) );
  OAI21_X1 U20799 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21820), .A(
        n18786), .ZN(n18775) );
  OAI211_X1 U20800 ( .C1(n21824), .C2(n19148), .A(n18776), .B(n18775), .ZN(
        P3_U2815) );
  AOI22_X1 U20801 ( .A1(n21946), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n22039), .B2(n19019), .ZN(n18777) );
  XOR2_X1 U20802 ( .A(n18868), .B(n18777), .Z(n22045) );
  OAI21_X1 U20803 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n21229), .ZN(n18783) );
  INV_X1 U20804 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18780) );
  NAND2_X1 U20805 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18778), .ZN(
        n18779) );
  AND2_X1 U20806 ( .A1(n18984), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18983) );
  AOI21_X1 U20807 ( .B1(n18780), .B2(n18779), .A(n18983), .ZN(n21218) );
  AOI22_X1 U20808 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18781), .B1(
        n18964), .B2(n21218), .ZN(n18782) );
  NAND2_X1 U20809 ( .A1(n22073), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n22042) );
  OAI211_X1 U20810 ( .C1(n18784), .C2(n18783), .A(n18782), .B(n22042), .ZN(
        n18785) );
  AOI221_X1 U20811 ( .B1(n18988), .B2(n22039), .C1(n18786), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n18785), .ZN(n18787) );
  OAI21_X1 U20812 ( .B1(n18961), .B2(n22045), .A(n18787), .ZN(P3_U2814) );
  NOR2_X1 U20813 ( .A1(n21154), .A2(n21027), .ZN(n19008) );
  NAND2_X1 U20814 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19008), .ZN(
        n21173) );
  OAI21_X1 U20815 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19008), .A(
        n21173), .ZN(n21156) );
  NOR2_X1 U20816 ( .A1(n18889), .A2(n21154), .ZN(n18807) );
  INV_X1 U20817 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18790) );
  OAI21_X1 U20818 ( .B1(n19112), .B2(n21154), .A(n19078), .ZN(n18788) );
  OAI21_X1 U20819 ( .B1(n19008), .B2(n19143), .A(n18788), .ZN(n18799) );
  NAND2_X1 U20820 ( .A1(n22073), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21792) );
  INV_X1 U20821 ( .A(n21792), .ZN(n18789) );
  AOI221_X1 U20822 ( .B1(n18807), .B2(n18790), .C1(n18799), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18789), .ZN(n18797) );
  INV_X1 U20823 ( .A(n19013), .ZN(n21790) );
  NOR3_X1 U20824 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n19011), .A3(
        n18791), .ZN(n18802) );
  AOI21_X1 U20825 ( .B1(n19039), .B2(n21790), .A(n18802), .ZN(n18792) );
  XNOR2_X1 U20826 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18792), .ZN(
        n21791) );
  NOR2_X1 U20827 ( .A1(n19031), .A2(n19013), .ZN(n18794) );
  NAND2_X1 U20828 ( .A1(n21766), .A2(n21783), .ZN(n18801) );
  NAND2_X1 U20829 ( .A1(n21783), .A2(n21769), .ZN(n21785) );
  AOI22_X1 U20830 ( .A1(n19000), .A2(n18801), .B1(n19072), .B2(n21785), .ZN(
        n18805) );
  INV_X1 U20831 ( .A(n18805), .ZN(n18793) );
  MUX2_X1 U20832 ( .A(n18794), .B(n18793), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n18795) );
  AOI21_X1 U20833 ( .B1(n19054), .B2(n21791), .A(n18795), .ZN(n18796) );
  OAI211_X1 U20834 ( .C1(n18921), .C2(n21156), .A(n18797), .B(n18796), .ZN(
        P3_U2818) );
  INV_X1 U20835 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18798) );
  AOI22_X1 U20836 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n21167), .B1(
        n18798), .B2(n21173), .ZN(n21175) );
  AOI22_X1 U20837 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18799), .B1(
        n18964), .B2(n21175), .ZN(n18811) );
  NAND2_X1 U20838 ( .A1(n11346), .A2(n18800), .ZN(n19049) );
  NOR2_X1 U20839 ( .A1(n11302), .A2(n19049), .ZN(n19048) );
  INV_X1 U20840 ( .A(n18801), .ZN(n21788) );
  AOI22_X1 U20841 ( .A1(n19048), .A2(n21788), .B1(n18802), .B2(n21797), .ZN(
        n18803) );
  XNOR2_X1 U20842 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18803), .ZN(
        n22046) );
  INV_X1 U20843 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18804) );
  NAND2_X1 U20844 ( .A1(n21783), .A2(n18804), .ZN(n22054) );
  OAI22_X1 U20845 ( .A1(n19031), .A2(n22054), .B1(n18805), .B2(n18804), .ZN(
        n18806) );
  AOI21_X1 U20846 ( .B1(n19054), .B2(n22046), .A(n18806), .ZN(n18810) );
  NAND2_X1 U20847 ( .A1(n22073), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18809) );
  OAI211_X1 U20848 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18807), .B(n18995), .ZN(n18808) );
  NAND4_X1 U20849 ( .A1(n18811), .A2(n18810), .A3(n18809), .A4(n18808), .ZN(
        P3_U2817) );
  NAND2_X1 U20850 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21666) );
  INV_X1 U20851 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21667) );
  NOR2_X1 U20852 ( .A1(n21666), .A2(n21667), .ZN(n21842) );
  INV_X1 U20853 ( .A(n21842), .ZN(n21882) );
  NOR3_X1 U20854 ( .A1(n22009), .A2(n21659), .A3(n21882), .ZN(n18866) );
  NAND2_X1 U20855 ( .A1(n18866), .A2(n18988), .ZN(n18929) );
  INV_X1 U20856 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21856) );
  AOI22_X1 U20857 ( .A1(n19000), .A2(n21957), .B1(n19072), .B2(n18947), .ZN(
        n18830) );
  NOR2_X1 U20858 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18826) );
  NAND3_X1 U20859 ( .A1(n18832), .A2(n18826), .A3(n21667), .ZN(n18845) );
  INV_X1 U20860 ( .A(n18873), .ZN(n18814) );
  AOI21_X1 U20861 ( .B1(n18845), .B2(n18874), .A(n18814), .ZN(n18846) );
  XNOR2_X1 U20862 ( .A(n18846), .B(n21856), .ZN(n21830) );
  INV_X1 U20863 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21292) );
  INV_X1 U20864 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21279) );
  NAND2_X1 U20865 ( .A1(n18816), .A2(n18936), .ZN(n18822) );
  AOI221_X1 U20866 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n21292), .C2(n21279), .A(
        n18822), .ZN(n18820) );
  NAND2_X1 U20867 ( .A1(n18816), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18837) );
  NOR2_X1 U20868 ( .A1(n21279), .A2(n18837), .ZN(n18815) );
  NOR2_X1 U20869 ( .A1(n18848), .A2(n21027), .ZN(n18851) );
  INV_X1 U20870 ( .A(n18851), .ZN(n18849) );
  OAI21_X1 U20871 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18815), .A(
        n18849), .ZN(n21287) );
  OAI22_X1 U20872 ( .A1(n18838), .A2(n19143), .B1(n18816), .B2(n19105), .ZN(
        n18817) );
  NOR2_X1 U20873 ( .A1(n19112), .A2(n18817), .ZN(n18834) );
  OAI21_X1 U20874 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18937), .A(
        n18834), .ZN(n18824) );
  AOI22_X1 U20875 ( .A1(n22073), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18824), .ZN(n18818) );
  OAI21_X1 U20876 ( .B1(n21287), .B2(n18921), .A(n18818), .ZN(n18819) );
  AOI211_X1 U20877 ( .C1(n21830), .C2(n19054), .A(n18820), .B(n18819), .ZN(
        n18821) );
  OAI221_X1 U20878 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18929), 
        .C1(n21856), .C2(n18830), .A(n18821), .ZN(P3_U2808) );
  INV_X1 U20879 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21289) );
  NOR2_X1 U20880 ( .A1(n22049), .A2(n21289), .ZN(n21670) );
  XNOR2_X1 U20881 ( .A(n21279), .B(n18837), .ZN(n21275) );
  OAI22_X1 U20882 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18822), .B1(
        n18921), .B2(n21275), .ZN(n18823) );
  AOI211_X1 U20883 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n18824), .A(
        n21670), .B(n18823), .ZN(n18829) );
  INV_X1 U20884 ( .A(n21666), .ZN(n21664) );
  AOI22_X1 U20885 ( .A1(n21664), .A2(n18831), .B1(n18826), .B2(n18825), .ZN(
        n18827) );
  XNOR2_X1 U20886 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18827), .ZN(
        n21671) );
  NOR2_X1 U20887 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21666), .ZN(
        n21640) );
  AOI22_X1 U20888 ( .A1(n19054), .A2(n21671), .B1(n21640), .B2(n18885), .ZN(
        n18828) );
  OAI211_X1 U20889 ( .C1(n18830), .C2(n21667), .A(n18829), .B(n18828), .ZN(
        P3_U2809) );
  OAI221_X1 U20890 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18832), 
        .C1(n18842), .C2(n18831), .A(n18873), .ZN(n18833) );
  XOR2_X1 U20891 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18833), .Z(
        n22007) );
  AOI221_X1 U20892 ( .B1(n18836), .B2(n18835), .C1(n19862), .C2(n18835), .A(
        n18834), .ZN(n18840) );
  OAI21_X1 U20893 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18838), .A(
        n18837), .ZN(n21269) );
  NAND2_X1 U20894 ( .A1(n22073), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n22005) );
  OAI221_X1 U20895 ( .B1(n21269), .B2(n18921), .C1(n21269), .C2(n18937), .A(
        n22005), .ZN(n18839) );
  AOI211_X1 U20896 ( .C1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n18841), .A(
        n18840), .B(n18839), .ZN(n18844) );
  NOR2_X1 U20897 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18842), .ZN(
        n22003) );
  NAND2_X1 U20898 ( .A1(n18885), .A2(n22003), .ZN(n18843) );
  OAI211_X1 U20899 ( .C1(n22007), .C2(n18961), .A(n18844), .B(n18843), .ZN(
        P3_U2810) );
  INV_X1 U20900 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21967) );
  NOR2_X1 U20901 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18845), .ZN(
        n18869) );
  OAI221_X1 U20902 ( .B1(n18869), .B2(n21946), .C1(n18869), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18846), .ZN(n18847) );
  XNOR2_X1 U20903 ( .A(n21967), .B(n18847), .ZN(n21974) );
  NOR2_X1 U20904 ( .A1(n11344), .A2(n19862), .ZN(n18854) );
  INV_X1 U20905 ( .A(n18848), .ZN(n18853) );
  INV_X1 U20906 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n21302) );
  NOR2_X1 U20907 ( .A1(n22049), .A2(n21302), .ZN(n21956) );
  AOI211_X1 U20908 ( .C1(n18850), .C2(n18849), .A(n18854), .B(n19112), .ZN(
        n18861) );
  NOR2_X1 U20909 ( .A1(n18917), .A2(n18964), .ZN(n19140) );
  NAND2_X1 U20910 ( .A1(n11344), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18880) );
  OAI21_X1 U20911 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18851), .A(
        n18880), .ZN(n21309) );
  OAI22_X1 U20912 ( .A1(n18861), .A2(n21312), .B1(n19140), .B2(n21309), .ZN(
        n18852) );
  AOI211_X1 U20913 ( .C1(n18854), .C2(n18853), .A(n21956), .B(n18852), .ZN(
        n18859) );
  NAND2_X1 U20914 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21958) );
  OAI21_X1 U20915 ( .B1(n21958), .B2(n18947), .A(n19072), .ZN(n18856) );
  OAI21_X1 U20916 ( .B1(n21958), .B2(n21957), .A(n19000), .ZN(n18855) );
  OAI22_X1 U20917 ( .A1(n18947), .A2(n18856), .B1(n21957), .B2(n18855), .ZN(
        n18857) );
  NAND2_X1 U20918 ( .A1(n18856), .A2(n18855), .ZN(n18886) );
  AOI22_X1 U20919 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18857), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18886), .ZN(n18858) );
  OAI211_X1 U20920 ( .C1(n18961), .C2(n21974), .A(n18859), .B(n18858), .ZN(
        P3_U2807) );
  INV_X1 U20921 ( .A(n21958), .ZN(n21960) );
  NAND2_X1 U20922 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21960), .ZN(
        n21841) );
  NOR2_X1 U20923 ( .A1(n21957), .A2(n21841), .ZN(n18860) );
  XNOR2_X1 U20924 ( .A(n18860), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n21847) );
  OAI21_X1 U20925 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18937), .A(
        n18861), .ZN(n18884) );
  NAND2_X1 U20926 ( .A1(n11344), .A2(n18936), .ZN(n18881) );
  AOI221_X1 U20927 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n11526), .C2(n11527), .A(
        n18881), .ZN(n18864) );
  INV_X1 U20928 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21340) );
  NOR2_X1 U20929 ( .A1(n11527), .A2(n18880), .ZN(n18862) );
  NOR2_X1 U20930 ( .A1(n18923), .A2(n21027), .ZN(n18891) );
  INV_X1 U20931 ( .A(n18891), .ZN(n18919) );
  OAI21_X1 U20932 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18862), .A(
        n18919), .ZN(n21335) );
  OAI22_X1 U20933 ( .A1(n22049), .A2(n21340), .B1(n21335), .B2(n18921), .ZN(
        n18863) );
  AOI211_X1 U20934 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18884), .A(
        n18864), .B(n18863), .ZN(n18877) );
  NOR2_X1 U20935 ( .A1(n18947), .A2(n21841), .ZN(n18865) );
  INV_X1 U20936 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21861) );
  XNOR2_X1 U20937 ( .A(n18865), .B(n21861), .ZN(n21851) );
  NAND2_X1 U20938 ( .A1(n18869), .A2(n21967), .ZN(n18870) );
  NOR2_X1 U20939 ( .A1(n21946), .A2(n18878), .ZN(n18898) );
  INV_X1 U20940 ( .A(n18898), .ZN(n18926) );
  OAI21_X1 U20941 ( .B1(n19019), .B2(n11152), .A(n18926), .ZN(n18875) );
  XNOR2_X1 U20942 ( .A(n18875), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n21852) );
  AOI22_X1 U20943 ( .A1(n19072), .A2(n21851), .B1(n19054), .B2(n21852), .ZN(
        n18876) );
  OAI211_X1 U20944 ( .C1(n21847), .C2(n19052), .A(n18877), .B(n18876), .ZN(
        P3_U2805) );
  AOI21_X1 U20945 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18879), .A(
        n18878), .ZN(n21982) );
  INV_X1 U20946 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21324) );
  NOR2_X1 U20947 ( .A1(n22049), .A2(n21324), .ZN(n18883) );
  XOR2_X1 U20948 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n18880), .Z(
        n21321) );
  OAI22_X1 U20949 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18881), .B1(
        n18921), .B2(n21321), .ZN(n18882) );
  AOI211_X1 U20950 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n18884), .A(
        n18883), .B(n18882), .ZN(n18888) );
  NOR3_X1 U20951 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21882), .A3(
        n21958), .ZN(n21976) );
  AOI22_X1 U20952 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18886), .B1(
        n18885), .B2(n21976), .ZN(n18887) );
  OAI211_X1 U20953 ( .C1(n21982), .C2(n18961), .A(n18888), .B(n18887), .ZN(
        P3_U2806) );
  NOR3_X1 U20954 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18889), .A3(
        n18909), .ZN(n18912) );
  OAI22_X1 U20955 ( .A1(n18891), .A2(n19143), .B1(n18890), .B2(n19105), .ZN(
        n18892) );
  NOR2_X1 U20956 ( .A1(n19112), .A2(n18892), .ZN(n18922) );
  OAI21_X1 U20957 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18937), .A(
        n18922), .ZN(n18913) );
  NAND2_X1 U20958 ( .A1(n18894), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18910) );
  NOR2_X1 U20959 ( .A1(n18968), .A2(n21027), .ZN(n18966) );
  AOI21_X1 U20960 ( .B1(n11524), .B2(n18910), .A(n18966), .ZN(n18893) );
  INV_X1 U20961 ( .A(n18893), .ZN(n21375) );
  NAND2_X1 U20962 ( .A1(n21869), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n18896) );
  NAND3_X1 U20963 ( .A1(n18894), .A2(n11524), .A3(n18936), .ZN(n18895) );
  OAI211_X1 U20964 ( .C1(n21375), .C2(n18921), .A(n18896), .B(n18895), .ZN(
        n18897) );
  AOI221_X1 U20965 ( .B1(n18912), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(
        n18913), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18897), .ZN(
        n18907) );
  INV_X1 U20966 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21859) );
  NOR3_X1 U20967 ( .A1(n21841), .A2(n21859), .A3(n21861), .ZN(n18934) );
  INV_X1 U20968 ( .A(n18934), .ZN(n21891) );
  OR2_X1 U20969 ( .A1(n21891), .A2(n21957), .ZN(n21873) );
  INV_X1 U20970 ( .A(n18947), .ZN(n21959) );
  NAND2_X1 U20971 ( .A1(n18934), .A2(n21959), .ZN(n21857) );
  AOI22_X1 U20972 ( .A1(n19000), .A2(n21873), .B1(n19072), .B2(n21857), .ZN(
        n18933) );
  NAND2_X1 U20973 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18933), .ZN(
        n18914) );
  OAI211_X1 U20974 ( .C1(n19000), .C2(n19072), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18914), .ZN(n18906) );
  NOR2_X1 U20975 ( .A1(n21891), .A2(n18929), .ZN(n18955) );
  INV_X1 U20976 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21934) );
  NAND3_X1 U20977 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18955), .A3(
        n21934), .ZN(n18905) );
  NOR2_X1 U20978 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n21946), .ZN(
        n18941) );
  AOI21_X1 U20979 ( .B1(n21946), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18941), .ZN(n21951) );
  NOR2_X1 U20980 ( .A1(n21859), .A2(n21861), .ZN(n18900) );
  AOI21_X1 U20981 ( .B1(n21859), .B2(n21861), .A(n21946), .ZN(n18899) );
  INV_X1 U20982 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21874) );
  NAND2_X1 U20983 ( .A1(n21952), .A2(n18902), .ZN(n18903) );
  OAI211_X1 U20984 ( .C1(n21951), .C2(n18903), .A(n19054), .B(n21931), .ZN(
        n18904) );
  NAND4_X1 U20985 ( .A1(n18907), .A2(n18906), .A3(n18905), .A4(n18904), .ZN(
        P3_U2802) );
  XNOR2_X1 U20986 ( .A(n18908), .B(n19019), .ZN(n21881) );
  INV_X1 U20987 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21380) );
  NOR2_X1 U20988 ( .A1(n18909), .A2(n21027), .ZN(n18918) );
  OAI21_X1 U20989 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18918), .A(
        n18910), .ZN(n21365) );
  OAI22_X1 U20990 ( .A1(n22049), .A2(n21380), .B1(n21365), .B2(n18921), .ZN(
        n18911) );
  AOI211_X1 U20991 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n18913), .A(
        n18912), .B(n18911), .ZN(n18916) );
  OAI21_X1 U20992 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18955), .A(
        n18914), .ZN(n18915) );
  OAI211_X1 U20993 ( .C1(n21881), .C2(n18961), .A(n18916), .B(n18915), .ZN(
        P3_U2803) );
  AOI21_X1 U20994 ( .B1(n21344), .B2(n18919), .A(n18918), .ZN(n18920) );
  INV_X1 U20995 ( .A(n18920), .ZN(n21352) );
  AOI21_X1 U20996 ( .B1(n18921), .B2(n18937), .A(n21352), .ZN(n18925) );
  AOI221_X1 U20997 ( .B1(n18923), .B2(n21344), .C1(n19862), .C2(n21344), .A(
        n18922), .ZN(n18924) );
  AOI211_X1 U20998 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n22073), .A(n18925), 
        .B(n18924), .ZN(n18932) );
  OAI221_X1 U20999 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n19019), 
        .C1(n21861), .C2(n11152), .A(n18926), .ZN(n18928) );
  XNOR2_X1 U21000 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18928), .ZN(
        n21865) );
  NOR4_X1 U21001 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21841), .A3(
        n21861), .A4(n18929), .ZN(n18930) );
  AOI21_X1 U21002 ( .B1(n19054), .B2(n21865), .A(n18930), .ZN(n18931) );
  OAI211_X1 U21003 ( .C1(n18933), .C2(n21859), .A(n18932), .B(n18931), .ZN(
        P3_U2804) );
  NAND3_X1 U21004 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18934), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21888) );
  INV_X1 U21005 ( .A(n21885), .ZN(n21941) );
  NAND2_X1 U21006 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21918) );
  NOR2_X1 U21007 ( .A1(n21941), .A2(n21918), .ZN(n18935) );
  XNOR2_X1 U21008 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n18935), .ZN(
        n21925) );
  INV_X1 U21009 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21412) );
  NOR2_X1 U21010 ( .A1(n22049), .A2(n21412), .ZN(n21928) );
  NAND2_X1 U21011 ( .A1(n11360), .A2(n18936), .ZN(n18954) );
  INV_X1 U21012 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18938) );
  XOR2_X1 U21013 ( .A(n18938), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n18939) );
  NOR2_X1 U21014 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18937), .ZN(
        n18963) );
  OR2_X1 U21015 ( .A1(n19862), .A2(n11360), .ZN(n18967) );
  OAI211_X1 U21016 ( .C1(n18966), .C2(n19143), .A(n18967), .B(n19144), .ZN(
        n18971) );
  NOR2_X1 U21017 ( .A1(n18963), .A2(n18971), .ZN(n18952) );
  OAI22_X1 U21018 ( .A1(n18954), .A2(n18939), .B1(n18952), .B2(n18938), .ZN(
        n18940) );
  AOI211_X1 U21019 ( .C1(n21399), .C2(n18964), .A(n21928), .B(n18940), .ZN(
        n18950) );
  NAND2_X1 U21020 ( .A1(n18942), .A2(n18941), .ZN(n18972) );
  INV_X1 U21021 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21898) );
  NOR2_X1 U21022 ( .A1(n21934), .A2(n19019), .ZN(n18943) );
  OAI33_X1 U21023 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n18972), .B1(n21898), .B2(
        n21933), .B3(n11452), .ZN(n18946) );
  XNOR2_X1 U21024 ( .A(n18946), .B(n18945), .ZN(n21926) );
  INV_X1 U21025 ( .A(n18962), .ZN(n21940) );
  NOR2_X1 U21026 ( .A1(n21940), .A2(n21918), .ZN(n18948) );
  XOR2_X1 U21027 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n18948), .Z(
        n21921) );
  AOI22_X1 U21028 ( .A1(n19054), .A2(n21926), .B1(n19072), .B2(n21921), .ZN(
        n18949) );
  OAI211_X1 U21029 ( .C1(n21925), .C2(n19052), .A(n18950), .B(n18949), .ZN(
        P3_U2799) );
  OAI22_X1 U21030 ( .A1(n21898), .A2(n21933), .B1(n18972), .B2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18951) );
  XNOR2_X1 U21031 ( .A(n18951), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n21917) );
  XOR2_X1 U21032 ( .A(n18965), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n21409) );
  INV_X1 U21033 ( .A(n21409), .ZN(n18959) );
  NAND2_X1 U21034 ( .A1(n21869), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21915) );
  OAI221_X1 U21035 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18954), .C1(
        n18953), .C2(n18952), .A(n21915), .ZN(n18958) );
  NAND3_X1 U21036 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21908) );
  INV_X1 U21037 ( .A(n18955), .ZN(n18956) );
  NOR2_X1 U21038 ( .A1(n21908), .A2(n18956), .ZN(n18957) );
  NAND2_X1 U21039 ( .A1(n18962), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21886) );
  AOI21_X1 U21040 ( .B1(n21885), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n19052), .ZN(n18974) );
  OAI21_X1 U21041 ( .B1(n21917), .B2(n18961), .A(n18960), .ZN(P3_U2800) );
  AOI21_X1 U21042 ( .B1(n18962), .B2(n19072), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18977) );
  INV_X1 U21043 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21390) );
  NOR2_X1 U21044 ( .A1(n22049), .A2(n21390), .ZN(n21901) );
  NOR2_X1 U21045 ( .A1(n18964), .A2(n18963), .ZN(n18969) );
  OAI21_X1 U21046 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18966), .A(
        n18965), .ZN(n21389) );
  OAI22_X1 U21047 ( .A1(n18969), .A2(n21389), .B1(n18968), .B2(n18967), .ZN(
        n18970) );
  AOI211_X1 U21048 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18971), .A(
        n21901), .B(n18970), .ZN(n18976) );
  NAND2_X1 U21049 ( .A1(n18972), .A2(n21933), .ZN(n18973) );
  XNOR2_X1 U21050 ( .A(n18973), .B(n21898), .ZN(n21902) );
  AOI22_X1 U21051 ( .A1(n21885), .A2(n18974), .B1(n19054), .B2(n21902), .ZN(
        n18975) );
  OAI211_X1 U21052 ( .C1(n18978), .C2(n18977), .A(n18976), .B(n18975), .ZN(
        P3_U2801) );
  OAI21_X1 U21053 ( .B1(n18980), .B2(n22028), .A(n18979), .ZN(n22030) );
  INV_X1 U21054 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21224) );
  NOR2_X1 U21055 ( .A1(n22049), .A2(n21224), .ZN(n22029) );
  INV_X1 U21056 ( .A(n18981), .ZN(n18982) );
  OAI21_X1 U21057 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18983), .A(
        n18982), .ZN(n21231) );
  INV_X2 U21058 ( .A(n19862), .ZN(n19947) );
  AOI21_X1 U21059 ( .B1(n18984), .B2(n19947), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18986) );
  OAI22_X1 U21060 ( .A1(n19140), .A2(n21231), .B1(n18986), .B2(n18985), .ZN(
        n18987) );
  AOI211_X1 U21061 ( .C1(n19054), .C2(n22030), .A(n22029), .B(n18987), .ZN(
        n18990) );
  NAND3_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18988), .A3(
        n22028), .ZN(n18989) );
  OAI211_X1 U21063 ( .C1(n18991), .C2(n22028), .A(n18990), .B(n18989), .ZN(
        P3_U2813) );
  AOI21_X1 U21064 ( .B1(n21811), .B2(n18992), .A(n21820), .ZN(n21803) );
  NOR3_X1 U21065 ( .A1(n19079), .A2(n21078), .A3(n19862), .ZN(n19064) );
  NAND2_X1 U21066 ( .A1(n18993), .A2(n19064), .ZN(n19010) );
  AOI221_X1 U21067 ( .B1(n18995), .B2(n11537), .C1(n19010), .C2(n11537), .A(
        n18994), .ZN(n18999) );
  AND2_X1 U21068 ( .A1(n21167), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18997) );
  OAI21_X1 U21069 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18997), .A(
        n18996), .ZN(n21187) );
  NAND2_X1 U21070 ( .A1(n21869), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n21809) );
  OAI21_X1 U21071 ( .B1(n19140), .B2(n21187), .A(n21809), .ZN(n18998) );
  AOI211_X1 U21072 ( .C1(n21803), .C2(n19000), .A(n18999), .B(n18998), .ZN(
        n19007) );
  AOI21_X1 U21073 ( .B1(n21811), .B2(n19002), .A(n19001), .ZN(n21802) );
  NAND2_X1 U21074 ( .A1(n19004), .A2(n19003), .ZN(n19005) );
  XNOR2_X1 U21075 ( .A(n19005), .B(n21811), .ZN(n21807) );
  AOI22_X1 U21076 ( .A1(n19072), .A2(n21802), .B1(n19054), .B2(n21807), .ZN(
        n19006) );
  NAND2_X1 U21077 ( .A1(n19007), .A2(n19006), .ZN(P3_U2816) );
  INV_X1 U21078 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19047) );
  NAND3_X1 U21079 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19055), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21104) );
  NOR2_X1 U21080 ( .A1(n19047), .A2(n21104), .ZN(n19046) );
  NAND3_X1 U21081 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(n19046), .ZN(n19026) );
  AOI21_X1 U21082 ( .B1(n21149), .B2(n19026), .A(n19008), .ZN(n21145) );
  INV_X1 U21083 ( .A(n19078), .ZN(n19139) );
  INV_X1 U21084 ( .A(n19064), .ZN(n19024) );
  OAI22_X1 U21085 ( .A1(n19139), .A2(n21149), .B1(n19025), .B2(n19024), .ZN(
        n19009) );
  AOI22_X1 U21086 ( .A1(n21145), .A2(n19107), .B1(n19010), .B2(n19009), .ZN(
        n19017) );
  OAI22_X1 U21087 ( .A1(n21766), .A2(n19052), .B1(n19148), .B2(n21769), .ZN(
        n19018) );
  INV_X1 U21088 ( .A(n19011), .ZN(n19032) );
  AOI22_X1 U21089 ( .A1(n21779), .A2(n19039), .B1(n19032), .B2(n19040), .ZN(
        n19012) );
  XNOR2_X1 U21090 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19012), .ZN(
        n21777) );
  AOI22_X1 U21091 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n19018), .B1(
        n19054), .B2(n21777), .ZN(n19016) );
  NAND2_X1 U21092 ( .A1(n21869), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n19015) );
  INV_X1 U21093 ( .A(n19031), .ZN(n19042) );
  OAI211_X1 U21094 ( .C1(n21779), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n19042), .B(n19013), .ZN(n19014) );
  NAND4_X1 U21095 ( .A1(n19017), .A2(n19016), .A3(n19015), .A4(n19014), .ZN(
        P3_U2819) );
  INV_X1 U21096 ( .A(n19018), .ZN(n19045) );
  AOI21_X1 U21097 ( .B1(n19019), .B2(n22072), .A(n19039), .ZN(n19020) );
  AOI21_X1 U21098 ( .B1(n22072), .B2(n19021), .A(n19020), .ZN(n19023) );
  AOI221_X1 U21099 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19039), .C1(
        n22072), .C2(n19040), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n19022) );
  AOI21_X1 U21100 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19023), .A(
        n19022), .ZN(n22056) );
  INV_X1 U21101 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n21139) );
  NOR2_X1 U21102 ( .A1(n22049), .A2(n21139), .ZN(n19030) );
  NOR2_X1 U21103 ( .A1(n19025), .A2(n19024), .ZN(n19028) );
  INV_X1 U21104 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21121) );
  NAND3_X1 U21105 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(n19064), .ZN(n19037) );
  NOR2_X1 U21106 ( .A1(n21121), .A2(n19037), .ZN(n19036) );
  AOI21_X1 U21107 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19078), .A(
        n19036), .ZN(n19027) );
  NAND2_X1 U21108 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19046), .ZN(
        n21129) );
  INV_X1 U21109 ( .A(n21129), .ZN(n21114) );
  OAI21_X1 U21110 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n21114), .A(
        n19026), .ZN(n21130) );
  OAI22_X1 U21111 ( .A1(n19028), .A2(n19027), .B1(n19140), .B2(n21130), .ZN(
        n19029) );
  AOI211_X1 U21112 ( .C1(n22056), .C2(n19054), .A(n19030), .B(n19029), .ZN(
        n19034) );
  OR3_X1 U21113 ( .A1(n21779), .A2(n19032), .A3(n19031), .ZN(n19033) );
  OAI211_X1 U21114 ( .C1(n19045), .C2(n22055), .A(n19034), .B(n19033), .ZN(
        P3_U2820) );
  OAI21_X1 U21115 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19046), .A(
        n21129), .ZN(n19035) );
  INV_X1 U21116 ( .A(n19035), .ZN(n21116) );
  AOI211_X1 U21117 ( .C1(n19037), .C2(n21121), .A(n19139), .B(n19036), .ZN(
        n19038) );
  NOR2_X1 U21118 ( .A1(n22049), .A2(n21127), .ZN(n22076) );
  AOI211_X1 U21119 ( .C1(n21116), .C2(n19107), .A(n19038), .B(n22076), .ZN(
        n19044) );
  NOR2_X1 U21120 ( .A1(n19040), .A2(n19039), .ZN(n19041) );
  XNOR2_X1 U21121 ( .A(n19041), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n22078) );
  AOI22_X1 U21122 ( .A1(n19054), .A2(n22078), .B1(n22072), .B2(n19042), .ZN(
        n19043) );
  OAI211_X1 U21123 ( .C1(n19045), .C2(n22072), .A(n19044), .B(n19043), .ZN(
        P3_U2821) );
  OAI21_X1 U21124 ( .B1(n19055), .B2(n19105), .A(n19144), .ZN(n19065) );
  AOI21_X1 U21125 ( .B1(n19047), .B2(n21104), .A(n19046), .ZN(n21106) );
  AOI22_X1 U21126 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19065), .B1(
        n21106), .B2(n19107), .ZN(n19060) );
  AOI21_X1 U21127 ( .B1(n11302), .B2(n19049), .A(n19048), .ZN(n21762) );
  OAI21_X1 U21128 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19051), .A(
        n19050), .ZN(n21758) );
  OAI22_X1 U21129 ( .A1(n21762), .A2(n19052), .B1(n19148), .B2(n21758), .ZN(
        n19053) );
  AOI21_X1 U21130 ( .B1(n19054), .B2(n21762), .A(n19053), .ZN(n19059) );
  NAND2_X1 U21131 ( .A1(n21869), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n21763) );
  INV_X1 U21132 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19063) );
  INV_X1 U21133 ( .A(n19055), .ZN(n19061) );
  NOR2_X1 U21134 ( .A1(n19063), .A2(n19061), .ZN(n19057) );
  NAND2_X1 U21135 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19056) );
  OAI211_X1 U21136 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n19057), .A(
        n19947), .B(n19056), .ZN(n19058) );
  NAND4_X1 U21137 ( .A1(n19060), .A2(n19059), .A3(n21763), .A4(n19058), .ZN(
        P3_U2822) );
  NOR2_X1 U21138 ( .A1(n19061), .A2(n21027), .ZN(n21074) );
  OAI21_X1 U21139 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n21074), .A(
        n21104), .ZN(n21085) );
  INV_X1 U21140 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n21099) );
  OAI22_X1 U21141 ( .A1(n19140), .A2(n21085), .B1(n22049), .B2(n21099), .ZN(
        n19062) );
  AOI221_X1 U21142 ( .B1(n19065), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n19064), .C2(n19063), .A(n19062), .ZN(n19074) );
  AOI21_X1 U21143 ( .B1(n21755), .B2(n19067), .A(n19066), .ZN(n21750) );
  AOI21_X1 U21144 ( .B1(n19070), .B2(n19069), .A(n19068), .ZN(n19071) );
  XNOR2_X1 U21145 ( .A(n19071), .B(n21755), .ZN(n21749) );
  AOI22_X1 U21146 ( .A1(n19137), .A2(n21750), .B1(n19072), .B2(n21749), .ZN(
        n19073) );
  NAND2_X1 U21147 ( .A1(n19074), .A2(n19073), .ZN(P3_U2823) );
  OAI21_X1 U21148 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19076), .A(
        n19075), .ZN(n21741) );
  INV_X1 U21149 ( .A(n19079), .ZN(n19077) );
  NAND2_X1 U21150 ( .A1(n19077), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19089) );
  AOI21_X1 U21151 ( .B1(n21078), .B2(n19089), .A(n21074), .ZN(n21077) );
  NAND2_X1 U21152 ( .A1(n19077), .A2(n19947), .ZN(n19083) );
  OAI21_X1 U21153 ( .B1(n19862), .B2(n19079), .A(n19078), .ZN(n19095) );
  AOI21_X1 U21154 ( .B1(n11358), .B2(n19081), .A(n19080), .ZN(n21736) );
  AOI22_X1 U21155 ( .A1(n22073), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n19137), 
        .B2(n21736), .ZN(n19082) );
  OAI221_X1 U21156 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19083), .C1(
        n21078), .C2(n19095), .A(n19082), .ZN(n19084) );
  AOI21_X1 U21157 ( .B1(n21077), .B2(n19107), .A(n19084), .ZN(n19085) );
  OAI21_X1 U21158 ( .B1(n19148), .B2(n21741), .A(n19085), .ZN(P3_U2824) );
  AOI21_X1 U21159 ( .B1(n19088), .B2(n19144), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19096) );
  AOI21_X1 U21160 ( .B1(n21730), .B2(n19087), .A(n19086), .ZN(n21729) );
  INV_X1 U21161 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n21065) );
  NOR2_X1 U21162 ( .A1(n22049), .A2(n21065), .ZN(n21723) );
  AND2_X1 U21163 ( .A1(n19088), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n21058) );
  OAI21_X1 U21164 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n21058), .A(
        n19089), .ZN(n21059) );
  OAI21_X1 U21165 ( .B1(n19092), .B2(n19091), .A(n19090), .ZN(n21722) );
  OAI22_X1 U21166 ( .A1(n19140), .A2(n21059), .B1(n19148), .B2(n21722), .ZN(
        n19093) );
  AOI211_X1 U21167 ( .C1(n19137), .C2(n21729), .A(n21723), .B(n19093), .ZN(
        n19094) );
  OAI21_X1 U21168 ( .B1(n19096), .B2(n19095), .A(n19094), .ZN(P3_U2825) );
  OAI21_X1 U21169 ( .B1(n19099), .B2(n19098), .A(n19097), .ZN(n21721) );
  AOI21_X1 U21170 ( .B1(n19102), .B2(n19101), .A(n19100), .ZN(n21713) );
  INV_X1 U21171 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n21054) );
  NOR2_X1 U21172 ( .A1(n22049), .A2(n21054), .ZN(n21717) );
  NOR3_X1 U21173 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19104), .A3(
        n19862), .ZN(n19103) );
  AOI211_X1 U21174 ( .C1(n19137), .C2(n21713), .A(n21717), .B(n19103), .ZN(
        n19109) );
  INV_X1 U21175 ( .A(n19104), .ZN(n19106) );
  OAI21_X1 U21176 ( .B1(n19106), .B2(n19105), .A(n19144), .ZN(n19119) );
  NAND2_X1 U21177 ( .A1(n19106), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19113) );
  AOI21_X1 U21178 ( .B1(n21051), .B2(n19113), .A(n21058), .ZN(n21048) );
  AOI22_X1 U21179 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19119), .B1(
        n21048), .B2(n19107), .ZN(n19108) );
  OAI211_X1 U21180 ( .C1(n19148), .C2(n21721), .A(n19109), .B(n19108), .ZN(
        P3_U2826) );
  XNOR2_X1 U21181 ( .A(n19111), .B(n19110), .ZN(n21706) );
  NOR2_X1 U21182 ( .A1(n19112), .A2(n19130), .ZN(n19131) );
  OAI21_X1 U21183 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19114), .A(
        n19113), .ZN(n21034) );
  OAI21_X1 U21184 ( .B1(n19117), .B2(n19116), .A(n19115), .ZN(n21705) );
  OAI22_X1 U21185 ( .A1(n19140), .A2(n21034), .B1(n19148), .B2(n21705), .ZN(
        n19118) );
  AOI221_X1 U21186 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19119), .C1(
        n19131), .C2(n19119), .A(n19118), .ZN(n19120) );
  NAND2_X1 U21187 ( .A1(n21869), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21709) );
  OAI211_X1 U21188 ( .C1(n19147), .C2(n21706), .A(n19120), .B(n21709), .ZN(
        P3_U2827) );
  AOI21_X1 U21189 ( .B1(n19123), .B2(n19122), .A(n19121), .ZN(n21689) );
  NOR2_X1 U21190 ( .A1(n22049), .A2(n19223), .ZN(n21688) );
  OAI21_X1 U21191 ( .B1(n19126), .B2(n19125), .A(n19124), .ZN(n21694) );
  OAI22_X1 U21192 ( .A1(n19140), .A2(n19127), .B1(n19148), .B2(n21694), .ZN(
        n19128) );
  AOI211_X1 U21193 ( .C1(n19137), .C2(n21689), .A(n21688), .B(n19128), .ZN(
        n19129) );
  OAI221_X1 U21194 ( .B1(n19131), .B2(n19130), .C1(n19131), .C2(n19862), .A(
        n19129), .ZN(P3_U2828) );
  AOI21_X1 U21195 ( .B1(n19133), .B2(n19142), .A(n19132), .ZN(n21679) );
  AOI21_X1 U21196 ( .B1(n19135), .B2(n19141), .A(n19134), .ZN(n21682) );
  OAI22_X1 U21197 ( .A1(n21682), .A2(n19148), .B1(n22049), .B2(n21687), .ZN(
        n19136) );
  AOI21_X1 U21198 ( .B1(n19137), .B2(n21679), .A(n19136), .ZN(n19138) );
  OAI221_X1 U21199 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19140), .C1(
        n21027), .C2(n19139), .A(n19138), .ZN(P3_U2829) );
  NAND2_X1 U21200 ( .A1(n19142), .A2(n19141), .ZN(n21676) );
  INV_X1 U21201 ( .A(n21676), .ZN(n21675) );
  NAND3_X1 U21202 ( .A1(n21619), .A2(n19144), .A3(n19143), .ZN(n19145) );
  AOI22_X1 U21203 ( .A1(n22073), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19145), .ZN(n19146) );
  OAI221_X1 U21204 ( .B1(n21675), .B2(n19148), .C1(n21676), .C2(n19147), .A(
        n19146), .ZN(P3_U2830) );
  NOR2_X1 U21205 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19609), .ZN(
        n19660) );
  NOR2_X1 U21206 ( .A1(n19639), .A2(n19660), .ZN(n19150) );
  OAI22_X1 U21207 ( .A1(n19151), .A2(n19631), .B1(n19150), .B2(n19149), .ZN(
        P3_U2866) );
  NAND2_X1 U21208 ( .A1(n19153), .A2(n19152), .ZN(n19156) );
  OAI21_X1 U21209 ( .B1(n19154), .B2(n19648), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19155) );
  OAI21_X1 U21210 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19156), .A(
        n19155), .ZN(P3_U2864) );
  NOR4_X1 U21211 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19160) );
  NOR4_X1 U21212 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19159) );
  NOR4_X1 U21213 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19158) );
  NOR4_X1 U21214 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19157) );
  NAND4_X1 U21215 ( .A1(n19160), .A2(n19159), .A3(n19158), .A4(n19157), .ZN(
        n19166) );
  NOR4_X1 U21216 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19164) );
  AOI211_X1 U21217 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19163) );
  NOR4_X1 U21218 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19162) );
  NOR4_X1 U21219 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19161) );
  NAND4_X1 U21220 ( .A1(n19164), .A2(n19163), .A3(n19162), .A4(n19161), .ZN(
        n19165) );
  NOR2_X1 U21221 ( .A1(n19166), .A2(n19165), .ZN(n19177) );
  INV_X1 U21222 ( .A(n19177), .ZN(n19175) );
  NOR2_X1 U21223 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19168) );
  NAND2_X1 U21224 ( .A1(n19175), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19167) );
  OAI21_X1 U21225 ( .B1(n19175), .B2(n19168), .A(n19167), .ZN(P3_U3293) );
  AOI211_X1 U21226 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19169) );
  AOI21_X1 U21227 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19169), .ZN(n19170) );
  INV_X1 U21228 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19258) );
  AOI22_X1 U21229 ( .A1(n19177), .A2(n19170), .B1(n19258), .B2(n19175), .ZN(
        P3_U3292) );
  INV_X1 U21230 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19172) );
  NOR3_X1 U21231 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19174) );
  NOR2_X1 U21232 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n19174), .ZN(n19171) );
  MUX2_X1 U21233 ( .A(n19172), .B(n19171), .S(n19177), .Z(n19173) );
  INV_X1 U21234 ( .A(n19173), .ZN(P3_U2638) );
  INV_X1 U21235 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22416) );
  AOI21_X1 U21236 ( .B1(n21687), .B2(n22416), .A(n19174), .ZN(n19176) );
  INV_X1 U21237 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19260) );
  AOI22_X1 U21238 ( .A1(n19177), .A2(n19176), .B1(n19260), .B2(n19175), .ZN(
        P3_U2639) );
  INV_X1 U21239 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19178) );
  INV_X1 U21240 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19261) );
  AOI22_X1 U21241 ( .A1(n22421), .A2(n19178), .B1(n19261), .B2(n22469), .ZN(
        P3_U3297) );
  INV_X1 U21242 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19179) );
  AOI22_X1 U21243 ( .A1(n22421), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19179), 
        .B2(n22469), .ZN(P3_U3294) );
  OAI21_X1 U21244 ( .B1(n19180), .B2(P3_D_C_N_REG_SCAN_IN), .A(n22469), .ZN(
        n19181) );
  OAI21_X1 U21245 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n22469), .A(n19181), 
        .ZN(P3_U2635) );
  INV_X1 U21246 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21615) );
  AOI22_X1 U21247 ( .A1(n19216), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n19182) );
  OAI21_X1 U21248 ( .B1(n21615), .B2(n19198), .A(n19182), .ZN(P3_U2767) );
  INV_X1 U21249 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20998) );
  AOI22_X1 U21250 ( .A1(n19216), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n19183) );
  OAI21_X1 U21251 ( .B1(n20998), .B2(n19198), .A(n19183), .ZN(P3_U2766) );
  INV_X1 U21252 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n21000) );
  AOI22_X1 U21253 ( .A1(n19216), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n19184) );
  OAI21_X1 U21254 ( .B1(n21000), .B2(n19198), .A(n19184), .ZN(P3_U2765) );
  INV_X1 U21255 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n21002) );
  AOI22_X1 U21256 ( .A1(n19216), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n19185) );
  OAI21_X1 U21257 ( .B1(n21002), .B2(n19198), .A(n19185), .ZN(P3_U2764) );
  INV_X1 U21258 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21465) );
  AOI22_X1 U21259 ( .A1(n19216), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n19186) );
  OAI21_X1 U21260 ( .B1(n21465), .B2(n19198), .A(n19186), .ZN(P3_U2763) );
  INV_X1 U21261 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n21005) );
  AOI22_X1 U21262 ( .A1(n19216), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n19187) );
  OAI21_X1 U21263 ( .B1(n21005), .B2(n19198), .A(n19187), .ZN(P3_U2762) );
  INV_X1 U21264 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n21007) );
  AOI22_X1 U21265 ( .A1(n19216), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n19188) );
  OAI21_X1 U21266 ( .B1(n21007), .B2(n19198), .A(n19188), .ZN(P3_U2761) );
  INV_X1 U21267 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n21010) );
  INV_X2 U21268 ( .A(n20955), .ZN(n19216) );
  AOI22_X1 U21269 ( .A1(n19216), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n19189) );
  OAI21_X1 U21270 ( .B1(n21010), .B2(n19198), .A(n19189), .ZN(P3_U2760) );
  INV_X1 U21271 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21597) );
  AOI22_X1 U21272 ( .A1(n19216), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n19190) );
  OAI21_X1 U21273 ( .B1(n21597), .B2(n19198), .A(n19190), .ZN(P3_U2759) );
  INV_X1 U21274 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21457) );
  AOI22_X1 U21275 ( .A1(n19216), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U21276 ( .B1(n21457), .B2(n19198), .A(n19191), .ZN(P3_U2758) );
  INV_X1 U21277 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n21014) );
  AOI22_X1 U21278 ( .A1(n19216), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n19192) );
  OAI21_X1 U21279 ( .B1(n21014), .B2(n19198), .A(n19192), .ZN(P3_U2757) );
  INV_X1 U21280 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21450) );
  AOI22_X1 U21281 ( .A1(n19216), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n19193) );
  OAI21_X1 U21282 ( .B1(n21450), .B2(n19198), .A(n19193), .ZN(P3_U2756) );
  INV_X1 U21283 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n21437) );
  AOI22_X1 U21284 ( .A1(n19216), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U21285 ( .B1(n21437), .B2(n19198), .A(n19194), .ZN(P3_U2755) );
  INV_X1 U21286 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n21018) );
  AOI22_X1 U21287 ( .A1(n19216), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n19195) );
  OAI21_X1 U21288 ( .B1(n21018), .B2(n19198), .A(n19195), .ZN(P3_U2754) );
  INV_X1 U21289 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21585) );
  AOI22_X1 U21290 ( .A1(n19216), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U21291 ( .B1(n21585), .B2(n19198), .A(n19196), .ZN(P3_U2753) );
  INV_X1 U21292 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21592) );
  AOI22_X1 U21293 ( .A1(n19216), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n19197) );
  OAI21_X1 U21294 ( .B1(n21592), .B2(n19198), .A(n19197), .ZN(P3_U2752) );
  INV_X1 U21295 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20971) );
  AOI22_X1 U21296 ( .A1(n19216), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U21297 ( .B1(n20971), .B2(n19218), .A(n19200), .ZN(P3_U2751) );
  INV_X1 U21298 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20973) );
  AOI22_X1 U21299 ( .A1(n19216), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n19201) );
  OAI21_X1 U21300 ( .B1(n20973), .B2(n19218), .A(n19201), .ZN(P3_U2750) );
  INV_X1 U21301 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20975) );
  AOI22_X1 U21302 ( .A1(n19216), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n19202) );
  OAI21_X1 U21303 ( .B1(n20975), .B2(n19218), .A(n19202), .ZN(P3_U2749) );
  INV_X1 U21304 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21489) );
  AOI22_X1 U21305 ( .A1(n19216), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n19203) );
  OAI21_X1 U21306 ( .B1(n21489), .B2(n19218), .A(n19203), .ZN(P3_U2748) );
  INV_X1 U21307 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n21508) );
  AOI22_X1 U21308 ( .A1(n19216), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U21309 ( .B1(n21508), .B2(n19218), .A(n19204), .ZN(P3_U2747) );
  INV_X1 U21310 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21502) );
  AOI22_X1 U21311 ( .A1(n19216), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n19205) );
  OAI21_X1 U21312 ( .B1(n21502), .B2(n19218), .A(n19205), .ZN(P3_U2746) );
  INV_X1 U21313 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n21531) );
  AOI22_X1 U21314 ( .A1(n19216), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n19206) );
  OAI21_X1 U21315 ( .B1(n21531), .B2(n19218), .A(n19206), .ZN(P3_U2745) );
  INV_X1 U21316 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20982) );
  AOI22_X1 U21317 ( .A1(n19216), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U21318 ( .B1(n20982), .B2(n19218), .A(n19207), .ZN(P3_U2744) );
  INV_X1 U21319 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20984) );
  AOI22_X1 U21320 ( .A1(n19216), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U21321 ( .B1(n20984), .B2(n19218), .A(n19209), .ZN(P3_U2743) );
  INV_X1 U21322 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20986) );
  AOI22_X1 U21323 ( .A1(n19216), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n19210) );
  OAI21_X1 U21324 ( .B1(n20986), .B2(n19218), .A(n19210), .ZN(P3_U2742) );
  INV_X1 U21325 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21540) );
  AOI22_X1 U21326 ( .A1(n19216), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U21327 ( .B1(n21540), .B2(n19218), .A(n19211), .ZN(P3_U2741) );
  INV_X1 U21328 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U21329 ( .A1(n19216), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n19212) );
  OAI21_X1 U21330 ( .B1(n20990), .B2(n19218), .A(n19212), .ZN(P3_U2740) );
  INV_X1 U21331 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n21558) );
  AOI22_X1 U21332 ( .A1(n19216), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U21333 ( .B1(n21558), .B2(n19218), .A(n19213), .ZN(P3_U2739) );
  INV_X1 U21334 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20993) );
  AOI22_X1 U21335 ( .A1(n19216), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n19214) );
  OAI21_X1 U21336 ( .B1(n20993), .B2(n19218), .A(n19214), .ZN(P3_U2738) );
  INV_X1 U21337 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20995) );
  AOI22_X1 U21338 ( .A1(n19216), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n19215), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n19217) );
  OAI21_X1 U21339 ( .B1(n20995), .B2(n19218), .A(n19217), .ZN(P3_U2737) );
  NOR2_X1 U21340 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n19219), .ZN(n19220) );
  NOR2_X1 U21341 ( .A1(n22421), .A2(n19220), .ZN(P3_U2633) );
  NOR2_X2 U21342 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22469), .ZN(n22465) );
  AOI22_X1 U21343 ( .A1(n22465), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n22469), .ZN(n19221) );
  OAI21_X1 U21344 ( .B1(n19253), .B2(n21687), .A(n19221), .ZN(P3_U3032) );
  AOI22_X1 U21345 ( .A1(n22465), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n22469), .ZN(n19222) );
  OAI21_X1 U21346 ( .B1(n19253), .B2(n19223), .A(n19222), .ZN(P3_U3033) );
  INV_X1 U21347 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19225) );
  AOI22_X1 U21348 ( .A1(n22465), .A2(P3_REIP_REG_4__SCAN_IN), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n22469), .ZN(n19224) );
  OAI21_X1 U21349 ( .B1(n19253), .B2(n19225), .A(n19224), .ZN(P3_U3034) );
  AOI22_X1 U21350 ( .A1(n22465), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n22469), .ZN(n19226) );
  OAI21_X1 U21351 ( .B1(n19253), .B2(n21054), .A(n19226), .ZN(P3_U3035) );
  AOI22_X1 U21352 ( .A1(n22465), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n22469), .ZN(n19227) );
  OAI21_X1 U21353 ( .B1(n19253), .B2(n21065), .A(n19227), .ZN(P3_U3036) );
  INV_X1 U21354 ( .A(n22465), .ZN(n19256) );
  AOI22_X1 U21355 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n22469), .ZN(n19228) );
  OAI21_X1 U21356 ( .B1(n21099), .B2(n19256), .A(n19228), .ZN(P3_U3037) );
  AOI22_X1 U21357 ( .A1(n22465), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n22469), .ZN(n19229) );
  OAI21_X1 U21358 ( .B1(n19253), .B2(n21099), .A(n19229), .ZN(P3_U3038) );
  AOI22_X1 U21359 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n22469), .ZN(n19230) );
  OAI21_X1 U21360 ( .B1(n21127), .B2(n19256), .A(n19230), .ZN(P3_U3039) );
  AOI22_X1 U21361 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n22469), .ZN(n19231) );
  OAI21_X1 U21362 ( .B1(n21139), .B2(n19256), .A(n19231), .ZN(P3_U3040) );
  AOI22_X1 U21363 ( .A1(n22465), .A2(P3_REIP_REG_11__SCAN_IN), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n22469), .ZN(n19232) );
  OAI21_X1 U21364 ( .B1(n19253), .B2(n21139), .A(n19232), .ZN(P3_U3041) );
  INV_X1 U21365 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n21781) );
  AOI22_X1 U21366 ( .A1(n22465), .A2(P3_REIP_REG_12__SCAN_IN), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n22469), .ZN(n19233) );
  OAI21_X1 U21367 ( .B1(n19253), .B2(n21781), .A(n19233), .ZN(P3_U3042) );
  INV_X1 U21368 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n21185) );
  AOI22_X1 U21369 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n22469), .ZN(n19234) );
  OAI21_X1 U21370 ( .B1(n21185), .B2(n19256), .A(n19234), .ZN(P3_U3043) );
  AOI22_X1 U21371 ( .A1(n22465), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n22469), .ZN(n19235) );
  OAI21_X1 U21372 ( .B1(n19253), .B2(n21185), .A(n19235), .ZN(P3_U3044) );
  INV_X1 U21373 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n21207) );
  AOI22_X1 U21374 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n22469), .ZN(n19236) );
  OAI21_X1 U21375 ( .B1(n21207), .B2(n19256), .A(n19236), .ZN(P3_U3045) );
  AOI22_X1 U21376 ( .A1(n22465), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n22469), .ZN(n19237) );
  OAI21_X1 U21377 ( .B1(n19253), .B2(n21207), .A(n19237), .ZN(P3_U3046) );
  AOI22_X1 U21378 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n22469), .ZN(n19238) );
  OAI21_X1 U21379 ( .B1(n21224), .B2(n19256), .A(n19238), .ZN(P3_U3047) );
  AOI22_X1 U21380 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n22469), .ZN(n19239) );
  OAI21_X1 U21381 ( .B1(n22026), .B2(n19256), .A(n19239), .ZN(P3_U3048) );
  AOI22_X1 U21382 ( .A1(n22465), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n22469), .ZN(n19240) );
  OAI21_X1 U21383 ( .B1(n19253), .B2(n22026), .A(n19240), .ZN(P3_U3049) );
  INV_X1 U21384 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19242) );
  AOI22_X1 U21385 ( .A1(n22465), .A2(P3_REIP_REG_20__SCAN_IN), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n22469), .ZN(n19241) );
  OAI21_X1 U21386 ( .B1(n19253), .B2(n19242), .A(n19241), .ZN(P3_U3050) );
  AOI22_X1 U21387 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n22469), .ZN(n19243) );
  OAI21_X1 U21388 ( .B1(n21289), .B2(n19256), .A(n19243), .ZN(P3_U3051) );
  INV_X1 U21389 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21298) );
  AOI22_X1 U21390 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n22469), .ZN(n19244) );
  OAI21_X1 U21391 ( .B1(n21298), .B2(n19256), .A(n19244), .ZN(P3_U3052) );
  AOI22_X1 U21392 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n22469), .ZN(n19245) );
  OAI21_X1 U21393 ( .B1(n21302), .B2(n19256), .A(n19245), .ZN(P3_U3053) );
  AOI22_X1 U21394 ( .A1(n22465), .A2(P3_REIP_REG_24__SCAN_IN), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n22469), .ZN(n19246) );
  OAI21_X1 U21395 ( .B1(n19253), .B2(n21302), .A(n19246), .ZN(P3_U3054) );
  AOI22_X1 U21396 ( .A1(n22465), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_ADDRESS_REG_23__SCAN_IN), .B2(n22469), .ZN(n19247) );
  OAI21_X1 U21397 ( .B1(n19253), .B2(n21324), .A(n19247), .ZN(P3_U3055) );
  AOI22_X1 U21398 ( .A1(n22465), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n22469), .ZN(n19248) );
  OAI21_X1 U21399 ( .B1(n19253), .B2(n21340), .A(n19248), .ZN(P3_U3056) );
  INV_X1 U21400 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21355) );
  AOI22_X1 U21401 ( .A1(n22465), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n22469), .ZN(n19249) );
  OAI21_X1 U21402 ( .B1(n19253), .B2(n21355), .A(n19249), .ZN(P3_U3057) );
  INV_X1 U21403 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21954) );
  AOI22_X1 U21404 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n22469), .ZN(n19250) );
  OAI21_X1 U21405 ( .B1(n21954), .B2(n19256), .A(n19250), .ZN(P3_U3058) );
  AOI22_X1 U21406 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n22469), .ZN(n19251) );
  OAI21_X1 U21407 ( .B1(n21390), .B2(n19256), .A(n19251), .ZN(P3_U3059) );
  AOI22_X1 U21408 ( .A1(n22465), .A2(P3_REIP_REG_30__SCAN_IN), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n22469), .ZN(n19252) );
  OAI21_X1 U21409 ( .B1(n19253), .B2(n21390), .A(n19252), .ZN(P3_U3060) );
  AOI22_X1 U21410 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n19254), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n22469), .ZN(n19255) );
  OAI21_X1 U21411 ( .B1(n21412), .B2(n19256), .A(n19255), .ZN(P3_U3061) );
  MUX2_X1 U21412 ( .A(P3_BE_N_REG_0__SCAN_IN), .B(P3_BYTEENABLE_REG_0__SCAN_IN), .S(n22421), .Z(P3_U3277) );
  MUX2_X1 U21413 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n22421), .Z(P3_U3276) );
  INV_X1 U21414 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19257) );
  AOI22_X1 U21415 ( .A1(n22421), .A2(n19258), .B1(n19257), .B2(n22469), .ZN(
        P3_U3275) );
  INV_X1 U21416 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19259) );
  AOI22_X1 U21417 ( .A1(n22421), .A2(n19260), .B1(n19259), .B2(n22469), .ZN(
        P3_U3274) );
  NOR4_X1 U21418 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n19263)
         );
  NOR4_X1 U21419 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n19261), .ZN(n19262) );
  INV_X2 U21420 ( .A(n19945), .ZN(U215) );
  NAND3_X1 U21421 ( .A1(n19263), .A2(n19262), .A3(U215), .ZN(U213) );
  NOR2_X1 U21422 ( .A1(n19566), .A2(n20235), .ZN(n19270) );
  NOR3_X1 U21423 ( .A1(n19266), .A2(n19264), .A3(n12045), .ZN(n19268) );
  AOI21_X1 U21424 ( .B1(n19266), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19265), 
        .ZN(n19267) );
  OAI21_X1 U21425 ( .B1(n19268), .B2(n19267), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19269) );
  OAI21_X1 U21426 ( .B1(n19270), .B2(n19574), .A(n19269), .ZN(n19277) );
  INV_X1 U21427 ( .A(n19270), .ZN(n19272) );
  OAI22_X1 U21428 ( .A1(n19570), .A2(n19273), .B1(n19272), .B2(n19271), .ZN(
        n19274) );
  NOR2_X1 U21429 ( .A1(n19275), .A2(n19274), .ZN(n19276) );
  MUX2_X1 U21430 ( .A(n19277), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19276), 
        .Z(P2_U3610) );
  NOR2_X1 U21431 ( .A1(n19396), .A2(n19278), .ZN(n19279) );
  XOR2_X1 U21432 ( .A(n19280), .B(n19279), .Z(n19287) );
  AOI22_X1 U21433 ( .A1(n19281), .A2(n19492), .B1(n19494), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n19282) );
  OAI211_X1 U21434 ( .C1(n11923), .C2(n19464), .A(n19282), .B(n19301), .ZN(
        n19285) );
  OAI22_X1 U21435 ( .A1(n20082), .A2(n19477), .B1(n19467), .B2(n19283), .ZN(
        n19284) );
  AOI211_X1 U21436 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19495), .A(
        n19285), .B(n19284), .ZN(n19286) );
  OAI21_X1 U21437 ( .B1(n19563), .B2(n19287), .A(n19286), .ZN(P2_U2848) );
  AOI22_X1 U21438 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19495), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19494), .ZN(n19288) );
  OAI21_X1 U21439 ( .B1(n19289), .B2(n19393), .A(n19288), .ZN(n19290) );
  AOI211_X1 U21440 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19491), .A(n19526), .B(
        n19290), .ZN(n19298) );
  NAND2_X1 U21441 ( .A1(n11252), .A2(n19291), .ZN(n19292) );
  XNOR2_X1 U21442 ( .A(n19293), .B(n19292), .ZN(n19296) );
  INV_X1 U21443 ( .A(n19294), .ZN(n19295) );
  AOI22_X1 U21444 ( .A1(n19296), .A2(n19484), .B1(n19498), .B2(n19295), .ZN(
        n19297) );
  OAI211_X1 U21445 ( .C1(n19477), .C2(n20079), .A(n19298), .B(n19297), .ZN(
        P2_U2847) );
  AOI22_X1 U21446 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19491), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19494), .ZN(n19303) );
  INV_X1 U21447 ( .A(n19299), .ZN(n20066) );
  AOI22_X1 U21448 ( .A1(n20066), .A2(n12449), .B1(n19492), .B2(n19300), .ZN(
        n19302) );
  NAND3_X1 U21449 ( .A1(n19303), .A2(n19302), .A3(n19301), .ZN(n19309) );
  NAND2_X1 U21450 ( .A1(n11253), .A2(n19304), .ZN(n19320) );
  OAI21_X1 U21451 ( .B1(n19305), .B2(n19312), .A(n19484), .ZN(n19307) );
  OAI22_X1 U21452 ( .A1(n19320), .A2(n19307), .B1(n19306), .B2(n19467), .ZN(
        n19308) );
  AOI211_X1 U21453 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n19495), .A(
        n19309), .B(n19308), .ZN(n19310) );
  OAI21_X1 U21454 ( .B1(n19312), .B2(n19311), .A(n19310), .ZN(P2_U2844) );
  INV_X1 U21455 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19317) );
  OAI22_X1 U21456 ( .A1(n19314), .A2(n19393), .B1(n19462), .B2(n19313), .ZN(
        n19315) );
  INV_X1 U21457 ( .A(n19315), .ZN(n19316) );
  OAI21_X1 U21458 ( .B1(n19317), .B2(n19386), .A(n19316), .ZN(n19318) );
  AOI211_X1 U21459 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19491), .A(n19526), .B(
        n19318), .ZN(n19324) );
  XNOR2_X1 U21460 ( .A(n19320), .B(n19319), .ZN(n19322) );
  AOI22_X1 U21461 ( .A1(n19322), .A2(n19484), .B1(n19321), .B2(n19498), .ZN(
        n19323) );
  OAI211_X1 U21462 ( .C1(n19477), .C2(n20064), .A(n19324), .B(n19323), .ZN(
        P2_U2843) );
  AOI211_X1 U21463 ( .C1(n11253), .C2(n19325), .A(n19563), .B(n19332), .ZN(
        n19330) );
  AOI21_X1 U21464 ( .B1(n19491), .B2(P2_EBX_REG_14__SCAN_IN), .A(n19526), .ZN(
        n19327) );
  NAND2_X1 U21465 ( .A1(n19494), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n19326) );
  OAI211_X1 U21466 ( .C1(n19328), .C2(n19393), .A(n19327), .B(n19326), .ZN(
        n19329) );
  AOI211_X1 U21467 ( .C1(n19495), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n19330), .B(n19329), .ZN(n19335) );
  AOI22_X1 U21468 ( .A1(n19333), .A2(n19332), .B1(n19331), .B2(n19498), .ZN(
        n19334) );
  OAI211_X1 U21469 ( .C1(n20058), .C2(n19477), .A(n19335), .B(n19334), .ZN(
        P2_U2841) );
  NOR2_X1 U21470 ( .A1(n19396), .A2(n19336), .ZN(n19337) );
  XNOR2_X1 U21471 ( .A(n19338), .B(n19337), .ZN(n19346) );
  OAI21_X1 U21472 ( .B1(n12147), .B2(n19464), .A(n19301), .ZN(n19342) );
  INV_X1 U21473 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19339) );
  OAI22_X1 U21474 ( .A1(n19340), .A2(n19393), .B1(n19462), .B2(n19339), .ZN(
        n19341) );
  AOI211_X1 U21475 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19494), .A(n19342), 
        .B(n19341), .ZN(n19345) );
  AOI22_X1 U21476 ( .A1(n20053), .A2(n12449), .B1(n19343), .B2(n19498), .ZN(
        n19344) );
  OAI211_X1 U21477 ( .C1(n19563), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        P2_U2840) );
  INV_X1 U21478 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19350) );
  OAI22_X1 U21479 ( .A1(n19347), .A2(n19393), .B1(n19462), .B2(n11741), .ZN(
        n19348) );
  AOI211_X1 U21480 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19491), .A(n19526), .B(
        n19348), .ZN(n19349) );
  OAI21_X1 U21481 ( .B1(n19350), .B2(n19386), .A(n19349), .ZN(n19355) );
  AOI211_X1 U21482 ( .C1(n19353), .C2(n19352), .A(n19563), .B(n19351), .ZN(
        n19354) );
  AOI211_X1 U21483 ( .C1(n19498), .C2(n19356), .A(n19355), .B(n19354), .ZN(
        n19357) );
  OAI21_X1 U21484 ( .B1(n19358), .B2(n19477), .A(n19357), .ZN(P2_U2839) );
  AOI211_X1 U21485 ( .C1(n19361), .C2(n19360), .A(n19359), .B(n19563), .ZN(
        n19371) );
  NAND2_X1 U21486 ( .A1(n19362), .A2(n19492), .ZN(n19369) );
  AOI21_X1 U21487 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n19491), .A(n19526), .ZN(
        n19364) );
  NAND2_X1 U21488 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19495), .ZN(
        n19363) );
  OAI211_X1 U21489 ( .C1(n19386), .C2(n19365), .A(n19364), .B(n19363), .ZN(
        n19366) );
  AOI21_X1 U21490 ( .B1(n19367), .B2(n19498), .A(n19366), .ZN(n19368) );
  NAND2_X1 U21491 ( .A1(n19369), .A2(n19368), .ZN(n19370) );
  NOR2_X1 U21492 ( .A1(n19371), .A2(n19370), .ZN(n19372) );
  OAI21_X1 U21493 ( .B1(n19373), .B2(n19477), .A(n19372), .ZN(P2_U2837) );
  AOI21_X1 U21494 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19491), .A(n19526), .ZN(
        n19374) );
  OAI21_X1 U21495 ( .B1(n19375), .B2(n19462), .A(n19374), .ZN(n19376) );
  AOI21_X1 U21496 ( .B1(n19494), .B2(P2_REIP_REG_19__SCAN_IN), .A(n19376), 
        .ZN(n19377) );
  OAI21_X1 U21497 ( .B1(n19378), .B2(n19467), .A(n19377), .ZN(n19382) );
  AOI211_X1 U21498 ( .C1(n19380), .C2(n19379), .A(n19563), .B(n19400), .ZN(
        n19381) );
  AOI211_X1 U21499 ( .C1(n19492), .C2(n19383), .A(n19382), .B(n19381), .ZN(
        n19384) );
  OAI21_X1 U21500 ( .B1(n19385), .B2(n19477), .A(n19384), .ZN(P2_U2836) );
  INV_X1 U21501 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19387) );
  OAI22_X1 U21502 ( .A1(n11501), .A2(n19462), .B1(n19387), .B2(n19386), .ZN(
        n19390) );
  NOR2_X1 U21503 ( .A1(n19464), .A2(n19388), .ZN(n19389) );
  AOI211_X1 U21504 ( .C1(n19391), .C2(n19498), .A(n19390), .B(n19389), .ZN(
        n19392) );
  OAI21_X1 U21505 ( .B1(n19394), .B2(n19393), .A(n19392), .ZN(n19395) );
  INV_X1 U21506 ( .A(n19395), .ZN(n19402) );
  OR2_X1 U21507 ( .A1(n19397), .A2(n19396), .ZN(n19399) );
  OAI21_X1 U21508 ( .B1(n19396), .B2(n19400), .A(n19397), .ZN(n19398) );
  OAI211_X1 U21509 ( .C1(n19400), .C2(n19399), .A(n19484), .B(n19398), .ZN(
        n19401) );
  OAI211_X1 U21510 ( .C1(n19477), .C2(n19403), .A(n19402), .B(n19401), .ZN(
        P2_U2835) );
  NAND2_X1 U21511 ( .A1(n19404), .A2(n19498), .ZN(n19407) );
  OAI22_X1 U21512 ( .A1(n19464), .A2(n12172), .B1(n19462), .B2(n11502), .ZN(
        n19405) );
  AOI21_X1 U21513 ( .B1(n19494), .B2(P2_REIP_REG_22__SCAN_IN), .A(n19405), 
        .ZN(n19406) );
  NAND2_X1 U21514 ( .A1(n19407), .A2(n19406), .ZN(n19408) );
  AOI21_X1 U21515 ( .B1(n19409), .B2(n19492), .A(n19408), .ZN(n19414) );
  OAI211_X1 U21516 ( .C1(n19412), .C2(n19411), .A(n19484), .B(n19410), .ZN(
        n19413) );
  OAI211_X1 U21517 ( .C1(n19477), .C2(n19415), .A(n19414), .B(n19413), .ZN(
        P2_U2833) );
  AOI22_X1 U21518 ( .A1(n19416), .A2(n19492), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n19491), .ZN(n19426) );
  AOI22_X1 U21519 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19495), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19494), .ZN(n19425) );
  NOR2_X1 U21520 ( .A1(n19417), .A2(n19467), .ZN(n19418) );
  AOI21_X1 U21521 ( .B1(n19419), .B2(n12449), .A(n19418), .ZN(n19424) );
  OAI211_X1 U21522 ( .C1(n19422), .C2(n19421), .A(n19484), .B(n19420), .ZN(
        n19423) );
  NAND4_X1 U21523 ( .A1(n19426), .A2(n19425), .A3(n19424), .A4(n19423), .ZN(
        P2_U2832) );
  AOI22_X1 U21524 ( .A1(n19427), .A2(n19492), .B1(n19494), .B2(
        P2_REIP_REG_24__SCAN_IN), .ZN(n19435) );
  AOI22_X1 U21525 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19495), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19491), .ZN(n19434) );
  AOI22_X1 U21526 ( .A1(n19429), .A2(n12449), .B1(n19498), .B2(n19428), .ZN(
        n19433) );
  OAI211_X1 U21527 ( .C1(n19431), .C2(n19430), .A(n19484), .B(n19441), .ZN(
        n19432) );
  NAND4_X1 U21528 ( .A1(n19435), .A2(n19434), .A3(n19433), .A4(n19432), .ZN(
        P2_U2831) );
  AOI22_X1 U21529 ( .A1(n19436), .A2(n19492), .B1(n19494), .B2(
        P2_REIP_REG_25__SCAN_IN), .ZN(n19448) );
  AOI22_X1 U21530 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19495), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19491), .ZN(n19447) );
  INV_X1 U21531 ( .A(n19437), .ZN(n19438) );
  AOI22_X1 U21532 ( .A1(n19439), .A2(n12449), .B1(n19438), .B2(n19498), .ZN(
        n19446) );
  INV_X1 U21533 ( .A(n19440), .ZN(n19444) );
  NAND2_X1 U21534 ( .A1(n19441), .A2(n11252), .ZN(n19443) );
  AOI21_X1 U21535 ( .B1(n19444), .B2(n19443), .A(n19563), .ZN(n19442) );
  OAI21_X1 U21536 ( .B1(n19444), .B2(n19443), .A(n19442), .ZN(n19445) );
  NAND4_X1 U21537 ( .A1(n19448), .A2(n19447), .A3(n19446), .A4(n19445), .ZN(
        P2_U2830) );
  AOI22_X1 U21538 ( .A1(n19449), .A2(n19492), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19491), .ZN(n19460) );
  AOI22_X1 U21539 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19495), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19494), .ZN(n19459) );
  INV_X1 U21540 ( .A(n19450), .ZN(n19451) );
  OAI22_X1 U21541 ( .A1(n19452), .A2(n19477), .B1(n19451), .B2(n19467), .ZN(
        n19453) );
  INV_X1 U21542 ( .A(n19453), .ZN(n19458) );
  OAI211_X1 U21543 ( .C1(n19456), .C2(n19455), .A(n19484), .B(n19454), .ZN(
        n19457) );
  NAND4_X1 U21544 ( .A1(n19460), .A2(n19459), .A3(n19458), .A4(n19457), .ZN(
        P2_U2829) );
  OAI22_X1 U21545 ( .A1(n19464), .A2(n19463), .B1(n19462), .B2(n19461), .ZN(
        n19465) );
  AOI21_X1 U21546 ( .B1(n19494), .B2(P2_REIP_REG_28__SCAN_IN), .A(n19465), 
        .ZN(n19466) );
  OAI21_X1 U21547 ( .B1(n19468), .B2(n19467), .A(n19466), .ZN(n19469) );
  AOI21_X1 U21548 ( .B1(n19470), .B2(n19492), .A(n19469), .ZN(n19475) );
  OAI211_X1 U21549 ( .C1(n19473), .C2(n19472), .A(n19484), .B(n19471), .ZN(
        n19474) );
  OAI211_X1 U21550 ( .C1(n19477), .C2(n19476), .A(n19475), .B(n19474), .ZN(
        P2_U2827) );
  AOI22_X1 U21551 ( .A1(n19478), .A2(n19492), .B1(n19494), .B2(
        P2_REIP_REG_29__SCAN_IN), .ZN(n19490) );
  AOI22_X1 U21552 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19491), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19495), .ZN(n19489) );
  INV_X1 U21553 ( .A(n19479), .ZN(n19482) );
  INV_X1 U21554 ( .A(n19480), .ZN(n19481) );
  AOI22_X1 U21555 ( .A1(n19482), .A2(n12449), .B1(n19481), .B2(n19498), .ZN(
        n19488) );
  OAI211_X1 U21556 ( .C1(n19486), .C2(n19485), .A(n19484), .B(n19483), .ZN(
        n19487) );
  NAND4_X1 U21557 ( .A1(n19490), .A2(n19489), .A3(n19488), .A4(n19487), .ZN(
        P2_U2826) );
  AOI22_X1 U21558 ( .A1(n19493), .A2(n19492), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n19491), .ZN(n19505) );
  AOI22_X1 U21559 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19495), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n19494), .ZN(n19504) );
  INV_X1 U21560 ( .A(n19496), .ZN(n20049) );
  AOI22_X1 U21561 ( .A1(n20049), .A2(n12449), .B1(n19498), .B2(n19497), .ZN(
        n19503) );
  NAND3_X1 U21562 ( .A1(n19501), .A2(n19500), .A3(n19499), .ZN(n19502) );
  NAND4_X1 U21563 ( .A1(n19505), .A2(n19504), .A3(n19503), .A4(n19502), .ZN(
        P2_U2824) );
  OR3_X1 U21564 ( .A1(n19507), .A2(n19557), .A3(n19506), .ZN(n19508) );
  OAI21_X1 U21565 ( .B1(n19510), .B2(n19509), .A(n19508), .ZN(P2_U3595) );
  INV_X1 U21566 ( .A(n20547), .ZN(n20553) );
  AOI22_X1 U21567 ( .A1(n19530), .A2(n19511), .B1(n19527), .B2(n20553), .ZN(
        n19520) );
  OAI22_X1 U21568 ( .A1(n19515), .A2(n19514), .B1(n19513), .B2(n19512), .ZN(
        n19516) );
  AOI211_X1 U21569 ( .C1(n19518), .C2(n19537), .A(n19517), .B(n19516), .ZN(
        n19519) );
  OAI211_X1 U21570 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19521), .A(
        n19520), .B(n19519), .ZN(P2_U3046) );
  OAI21_X1 U21571 ( .B1(n19524), .B2(n19523), .A(n19522), .ZN(n19528) );
  INV_X1 U21572 ( .A(n19525), .ZN(n20269) );
  AOI222_X1 U21573 ( .A1(n19528), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19527), .B2(n20269), .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19526), .ZN(
        n19534) );
  AOI222_X1 U21574 ( .A1(n19532), .A2(n19537), .B1(n19550), .B2(n19531), .C1(
        n19530), .C2(n19529), .ZN(n19533) );
  OAI211_X1 U21575 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n19535), .A(
        n19534), .B(n19533), .ZN(P2_U3040) );
  AOI22_X1 U21576 ( .A1(n19539), .A2(n19538), .B1(n19537), .B2(n19536), .ZN(
        n19541) );
  OAI211_X1 U21577 ( .C1(n19543), .C2(n19542), .A(n19541), .B(n19540), .ZN(
        n19549) );
  OAI22_X1 U21578 ( .A1(n19547), .A2(n19546), .B1(n19545), .B2(n19544), .ZN(
        n19548) );
  OAI211_X1 U21579 ( .C1(n19555), .C2(n19554), .A(n19553), .B(n19552), .ZN(
        P2_U3044) );
  NAND2_X1 U21580 ( .A1(n19571), .A2(n19556), .ZN(n19573) );
  NAND2_X1 U21581 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n22445), .ZN(n19558) );
  OAI21_X1 U21582 ( .B1(n19558), .B2(n19557), .A(n19580), .ZN(n19562) );
  NAND2_X1 U21583 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19566), .ZN(n19559) );
  AOI21_X1 U21584 ( .B1(n19560), .B2(n19573), .A(n19559), .ZN(n19561) );
  AOI21_X1 U21585 ( .B1(n19573), .B2(n19562), .A(n19561), .ZN(n19564) );
  NAND2_X1 U21586 ( .A1(n19564), .A2(n19563), .ZN(P2_U3177) );
  AOI22_X1 U21587 ( .A1(n19568), .A2(n19567), .B1(n19566), .B2(n19565), .ZN(
        n19579) );
  AOI22_X1 U21588 ( .A1(n19571), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19570), 
        .B2(n19569), .ZN(n19578) );
  NOR2_X1 U21589 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19572), .ZN(n19575) );
  OAI22_X1 U21590 ( .A1(n19575), .A2(n19574), .B1(n22445), .B2(n19573), .ZN(
        n19576) );
  NAND4_X1 U21591 ( .A1(n19579), .A2(n19578), .A3(n19577), .A4(n19576), .ZN(
        P2_U3176) );
  NOR2_X1 U21592 ( .A1(n19581), .A2(n19580), .ZN(n19584) );
  MUX2_X1 U21593 ( .A(P2_MORE_REG_SCAN_IN), .B(n19582), .S(n19584), .Z(
        P2_U3609) );
  OAI21_X1 U21594 ( .B1(n19584), .B2(n12741), .A(n19583), .ZN(P2_U2819) );
  INV_X1 U21595 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20950) );
  INV_X1 U21596 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19610) );
  AOI22_X1 U21597 ( .A1(n19945), .A2(n20950), .B1(n19610), .B2(U215), .ZN(U282) );
  OAI22_X1 U21598 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19945), .ZN(n19585) );
  INV_X1 U21599 ( .A(n19585), .ZN(U281) );
  OAI22_X1 U21600 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19945), .ZN(n19586) );
  INV_X1 U21601 ( .A(n19586), .ZN(U280) );
  INV_X1 U21602 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n19587) );
  INV_X1 U21603 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21562) );
  AOI22_X1 U21604 ( .A1(n19945), .A2(n19587), .B1(n21562), .B2(U215), .ZN(U279) );
  OAI22_X1 U21605 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19945), .ZN(n19588) );
  INV_X1 U21606 ( .A(n19588), .ZN(U278) );
  INV_X1 U21607 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n19589) );
  INV_X1 U21608 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n21544) );
  AOI22_X1 U21609 ( .A1(n19945), .A2(n19589), .B1(n21544), .B2(U215), .ZN(U277) );
  OAI22_X1 U21610 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19945), .ZN(n19590) );
  INV_X1 U21611 ( .A(n19590), .ZN(U276) );
  INV_X1 U21612 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n19591) );
  AOI22_X1 U21613 ( .A1(n19738), .A2(n19591), .B1(n17354), .B2(U215), .ZN(U275) );
  INV_X1 U21614 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n19592) );
  INV_X1 U21615 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n20083) );
  AOI22_X1 U21616 ( .A1(n19945), .A2(n19592), .B1(n20083), .B2(U215), .ZN(U274) );
  OAI22_X1 U21617 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19945), .ZN(n19593) );
  INV_X1 U21618 ( .A(n19593), .ZN(U273) );
  INV_X1 U21619 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n19594) );
  INV_X1 U21620 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21498) );
  AOI22_X1 U21621 ( .A1(n19738), .A2(n19594), .B1(n21498), .B2(U215), .ZN(U272) );
  INV_X1 U21622 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n19595) );
  INV_X1 U21623 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n21504) );
  AOI22_X1 U21624 ( .A1(n19738), .A2(n19595), .B1(n21504), .B2(U215), .ZN(U271) );
  OAI22_X1 U21625 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19738), .ZN(n19596) );
  INV_X1 U21626 ( .A(n19596), .ZN(U270) );
  INV_X1 U21627 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n19597) );
  INV_X1 U21628 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n21520) );
  AOI22_X1 U21629 ( .A1(n19738), .A2(n19597), .B1(n21520), .B2(U215), .ZN(U269) );
  OAI22_X1 U21630 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19738), .ZN(n19598) );
  INV_X1 U21631 ( .A(n19598), .ZN(U268) );
  OAI22_X1 U21632 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19738), .ZN(n19599) );
  INV_X1 U21633 ( .A(n19599), .ZN(U267) );
  OAI22_X1 U21634 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19945), .ZN(n19600) );
  INV_X1 U21635 ( .A(n19600), .ZN(U266) );
  OAI22_X1 U21636 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19945), .ZN(n19601) );
  INV_X1 U21637 ( .A(n19601), .ZN(U265) );
  INV_X1 U21638 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n19602) );
  INV_X1 U21639 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n21442) );
  AOI22_X1 U21640 ( .A1(n19945), .A2(n19602), .B1(n21442), .B2(U215), .ZN(U264) );
  INV_X1 U21641 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n19603) );
  INV_X1 U21642 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21447) );
  AOI22_X1 U21643 ( .A1(n19738), .A2(n19603), .B1(n21447), .B2(U215), .ZN(U263) );
  OAI22_X1 U21644 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19945), .ZN(n19604) );
  INV_X1 U21645 ( .A(n19604), .ZN(U262) );
  INV_X1 U21646 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n19605) );
  INV_X1 U21647 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n21455) );
  AOI22_X1 U21648 ( .A1(n19945), .A2(n19605), .B1(n21455), .B2(U215), .ZN(U261) );
  INV_X1 U21649 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n19606) );
  INV_X1 U21650 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21462) );
  AOI22_X1 U21651 ( .A1(n19738), .A2(n19606), .B1(n21462), .B2(U215), .ZN(U260) );
  OAI22_X1 U21652 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19945), .ZN(n19607) );
  INV_X1 U21653 ( .A(n19607), .ZN(U259) );
  INV_X1 U21654 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n19608) );
  INV_X1 U21655 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21464) );
  AOI22_X1 U21656 ( .A1(n19945), .A2(n19608), .B1(n21464), .B2(U215), .ZN(U258) );
  NOR3_X1 U21657 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19609), .A3(
        n19631), .ZN(n19611) );
  NAND2_X1 U21658 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19611), .ZN(
        n19944) );
  NAND2_X1 U21659 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19947), .ZN(n19676) );
  NAND2_X1 U21660 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19632), .ZN(
        n19616) );
  NOR2_X1 U21661 ( .A1(n19670), .A2(n19616), .ZN(n19949) );
  NOR2_X2 U21662 ( .A1(n21464), .A2(n19863), .ZN(n19688) );
  INV_X1 U21663 ( .A(n19611), .ZN(n19620) );
  NOR2_X2 U21664 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19620), .ZN(
        n19967) );
  NOR2_X2 U21665 ( .A1(n19610), .A2(n19862), .ZN(n19693) );
  AOI22_X1 U21666 ( .A1(n19949), .A2(n19688), .B1(n19967), .B2(n19693), .ZN(
        n19615) );
  INV_X1 U21667 ( .A(n19616), .ZN(n19684) );
  NAND2_X1 U21668 ( .A1(n19627), .A2(n19948), .ZN(n19638) );
  INV_X1 U21669 ( .A(n19638), .ZN(n19647) );
  AOI22_X1 U21670 ( .A1(n19947), .A2(n19611), .B1(n19684), .B2(n19647), .ZN(
        n19953) );
  NOR2_X2 U21671 ( .A1(n19653), .A2(n19616), .ZN(n19952) );
  NAND2_X1 U21672 ( .A1(n19613), .A2(n19612), .ZN(n19950) );
  NOR2_X1 U21673 ( .A1(n21435), .A2(n19950), .ZN(n19673) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19953), .B1(
        n19952), .B2(n19673), .ZN(n19614) );
  OAI211_X1 U21675 ( .C1(n19944), .C2(n19676), .A(n19615), .B(n19614), .ZN(
        P3_U2995) );
  NOR2_X1 U21676 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19616), .ZN(
        n19617) );
  INV_X1 U21677 ( .A(n19617), .ZN(n20047) );
  NAND2_X1 U21678 ( .A1(n19944), .A2(n20047), .ZN(n19692) );
  AND2_X1 U21679 ( .A1(n19687), .A2(n19692), .ZN(n19957) );
  NAND2_X1 U21680 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19639), .ZN(
        n19628) );
  NOR2_X2 U21681 ( .A1(n19653), .A2(n19628), .ZN(n19974) );
  AOI22_X1 U21682 ( .A1(n19688), .A2(n19957), .B1(n19693), .B2(n19974), .ZN(
        n19619) );
  NAND2_X1 U21683 ( .A1(n19956), .A2(n19965), .ZN(n19624) );
  AOI21_X1 U21684 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19863), .ZN(n19691) );
  OAI221_X1 U21685 ( .B1(n19692), .B2(n19648), .C1(n19692), .C2(n19624), .A(
        n19691), .ZN(n19958) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19958), .B1(
        n19673), .B2(n20031), .ZN(n19618) );
  OAI211_X1 U21687 ( .C1(n19676), .C2(n19956), .A(n19619), .B(n19618), .ZN(
        P3_U2987) );
  INV_X1 U21688 ( .A(n19673), .ZN(n19696) );
  INV_X1 U21689 ( .A(n19676), .ZN(n19689) );
  NOR2_X1 U21690 ( .A1(n19670), .A2(n19620), .ZN(n19961) );
  AOI22_X1 U21691 ( .A1(n19689), .A2(n19974), .B1(n19688), .B2(n19961), .ZN(
        n19623) );
  OAI22_X1 U21692 ( .A1(n19862), .A2(n19628), .B1(n19620), .B2(n19638), .ZN(
        n19621) );
  INV_X1 U21693 ( .A(n19621), .ZN(n19962) );
  NOR2_X2 U21694 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19628), .ZN(
        n19979) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19962), .B1(
        n19693), .B2(n19979), .ZN(n19622) );
  OAI211_X1 U21696 ( .C1(n19944), .C2(n19696), .A(n19623), .B(n19622), .ZN(
        P3_U2979) );
  AND2_X1 U21697 ( .A1(n19687), .A2(n19624), .ZN(n19966) );
  INV_X1 U21698 ( .A(n19639), .ZN(n19637) );
  NAND2_X1 U21699 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19636), .ZN(
        n19664) );
  NOR2_X2 U21700 ( .A1(n19637), .A2(n19664), .ZN(n19985) );
  AOI22_X1 U21701 ( .A1(n19688), .A2(n19966), .B1(n19693), .B2(n19985), .ZN(
        n19626) );
  NAND2_X1 U21702 ( .A1(n19971), .A2(n19977), .ZN(n19633) );
  AOI22_X1 U21703 ( .A1(n19947), .A2(n19633), .B1(n19691), .B2(n19624), .ZN(
        n19968) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19968), .B1(
        n19689), .B2(n19979), .ZN(n19625) );
  OAI211_X1 U21705 ( .C1(n19696), .C2(n19956), .A(n19626), .B(n19625), .ZN(
        P3_U2971) );
  INV_X1 U21706 ( .A(n19648), .ZN(n19655) );
  AOI21_X1 U21707 ( .B1(n19636), .B2(n19655), .A(n19863), .ZN(n19672) );
  NAND3_X1 U21708 ( .A1(n19639), .A2(n19672), .A3(n19627), .ZN(n19973) );
  NOR2_X1 U21709 ( .A1(n19670), .A2(n19628), .ZN(n19972) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19973), .B1(
        n19688), .B2(n19972), .ZN(n19630) );
  NOR2_X2 U21711 ( .A1(n19671), .A2(n19637), .ZN(n19991) );
  AOI22_X1 U21712 ( .A1(n19673), .A2(n19974), .B1(n19693), .B2(n19991), .ZN(
        n19629) );
  OAI211_X1 U21713 ( .C1(n19676), .C2(n19977), .A(n19630), .B(n19629), .ZN(
        P3_U2963) );
  AND2_X1 U21714 ( .A1(n19687), .A2(n19633), .ZN(n19978) );
  NAND2_X1 U21715 ( .A1(n19632), .A2(n19631), .ZN(n19649) );
  NOR2_X2 U21716 ( .A1(n19653), .A2(n19649), .ZN(n19996) );
  AOI22_X1 U21717 ( .A1(n19688), .A2(n19978), .B1(n19693), .B2(n19996), .ZN(
        n19635) );
  NAND2_X1 U21718 ( .A1(n19983), .A2(n19989), .ZN(n19644) );
  OAI221_X1 U21719 ( .B1(n19633), .B2(n19648), .C1(n19633), .C2(n19644), .A(
        n19691), .ZN(n19980) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19980), .B1(
        n19689), .B2(n19991), .ZN(n19634) );
  OAI211_X1 U21721 ( .C1(n19696), .C2(n19971), .A(n19635), .B(n19634), .ZN(
        P3_U2955) );
  NAND2_X1 U21722 ( .A1(n19636), .A2(n19687), .ZN(n19681) );
  NOR2_X1 U21723 ( .A1(n19637), .A2(n19681), .ZN(n19984) );
  AOI22_X1 U21724 ( .A1(n19689), .A2(n19996), .B1(n19688), .B2(n19984), .ZN(
        n19642) );
  INV_X1 U21725 ( .A(n19649), .ZN(n19640) );
  NOR2_X1 U21726 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19638), .ZN(
        n19683) );
  AOI22_X1 U21727 ( .A1(n19947), .A2(n19640), .B1(n19639), .B2(n19683), .ZN(
        n19986) );
  NOR2_X1 U21728 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19649), .ZN(
        n19918) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19986), .B1(
        n19693), .B2(n20002), .ZN(n19641) );
  OAI211_X1 U21730 ( .C1(n19696), .C2(n19977), .A(n19642), .B(n19641), .ZN(
        P3_U2947) );
  AND2_X1 U21731 ( .A1(n19687), .A2(n19644), .ZN(n19990) );
  AOI22_X1 U21732 ( .A1(n19689), .A2(n20002), .B1(n19688), .B2(n19990), .ZN(
        n19646) );
  INV_X1 U21733 ( .A(n19918), .ZN(n19836) );
  INV_X1 U21734 ( .A(n19664), .ZN(n19643) );
  NAND2_X1 U21735 ( .A1(n19643), .A2(n19660), .ZN(n20000) );
  NAND2_X1 U21736 ( .A1(n19836), .A2(n20000), .ZN(n19652) );
  AOI22_X1 U21737 ( .A1(n19947), .A2(n19652), .B1(n19691), .B2(n19644), .ZN(
        n19992) );
  INV_X1 U21738 ( .A(n20000), .ZN(n20007) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19992), .B1(
        n19693), .B2(n20007), .ZN(n19645) );
  OAI211_X1 U21740 ( .C1(n19696), .C2(n19983), .A(n19646), .B(n19645), .ZN(
        P3_U2939) );
  OAI211_X1 U21741 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19648), .A(
        n19647), .B(n19660), .ZN(n19997) );
  NOR2_X1 U21742 ( .A1(n19670), .A2(n19649), .ZN(n19995) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19997), .B1(
        n19688), .B2(n19995), .ZN(n19651) );
  INV_X1 U21744 ( .A(n19660), .ZN(n19659) );
  NOR2_X2 U21745 ( .A1(n19671), .A2(n19659), .ZN(n20013) );
  AOI22_X1 U21746 ( .A1(n19673), .A2(n19996), .B1(n19693), .B2(n20013), .ZN(
        n19650) );
  OAI211_X1 U21747 ( .C1(n19676), .C2(n20000), .A(n19651), .B(n19650), .ZN(
        P3_U2931) );
  INV_X1 U21748 ( .A(n19652), .ZN(n19654) );
  NOR2_X1 U21749 ( .A1(n19670), .A2(n19654), .ZN(n20001) );
  NOR2_X1 U21750 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19682) );
  NAND2_X1 U21751 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19682), .ZN(
        n19669) );
  NOR2_X2 U21752 ( .A1(n19653), .A2(n19669), .ZN(n20018) );
  AOI22_X1 U21753 ( .A1(n19688), .A2(n20001), .B1(n19693), .B2(n20018), .ZN(
        n19658) );
  NOR2_X1 U21754 ( .A1(n20013), .A2(n20018), .ZN(n19665) );
  OAI21_X1 U21755 ( .B1(n19665), .B2(n19655), .A(n19654), .ZN(n19656) );
  OAI211_X1 U21756 ( .C1(n20002), .C2(n22084), .A(n19948), .B(n19656), .ZN(
        n20003) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20003), .B1(
        n19689), .B2(n20013), .ZN(n19657) );
  OAI211_X1 U21758 ( .C1(n19696), .C2(n19836), .A(n19658), .B(n19657), .ZN(
        P3_U2923) );
  NOR2_X1 U21759 ( .A1(n19681), .A2(n19659), .ZN(n20006) );
  AOI22_X1 U21760 ( .A1(n19689), .A2(n20018), .B1(n19688), .B2(n20006), .ZN(
        n19663) );
  INV_X1 U21761 ( .A(n19669), .ZN(n19661) );
  AOI22_X1 U21762 ( .A1(n19947), .A2(n19661), .B1(n19683), .B2(n19660), .ZN(
        n20008) );
  NOR2_X1 U21763 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19669), .ZN(
        n19884) );
  CLKBUF_X1 U21764 ( .A(n19884), .Z(n20025) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20008), .B1(
        n19693), .B2(n20025), .ZN(n19662) );
  OAI211_X1 U21766 ( .C1(n19696), .C2(n20000), .A(n19663), .B(n19662), .ZN(
        P3_U2915) );
  INV_X1 U21767 ( .A(n19884), .ZN(n19764) );
  NOR2_X1 U21768 ( .A1(n19670), .A2(n19665), .ZN(n20012) );
  INV_X1 U21769 ( .A(n19682), .ZN(n19680) );
  NOR2_X2 U21770 ( .A1(n19664), .A2(n19680), .ZN(n20032) );
  AOI22_X1 U21771 ( .A1(n19688), .A2(n20012), .B1(n19693), .B2(n20032), .ZN(
        n19668) );
  NAND2_X1 U21772 ( .A1(n19764), .A2(n20022), .ZN(n19677) );
  INV_X1 U21773 ( .A(n19665), .ZN(n19666) );
  AOI22_X1 U21774 ( .A1(n19947), .A2(n19677), .B1(n19691), .B2(n19666), .ZN(
        n20014) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20014), .B1(
        n19673), .B2(n20013), .ZN(n19667) );
  OAI211_X1 U21776 ( .C1(n19676), .C2(n19764), .A(n19668), .B(n19667), .ZN(
        P3_U2907) );
  NOR2_X1 U21777 ( .A1(n19670), .A2(n19669), .ZN(n20017) );
  NOR2_X2 U21778 ( .A1(n19671), .A2(n19680), .ZN(n20042) );
  AOI22_X1 U21779 ( .A1(n19688), .A2(n20017), .B1(n19693), .B2(n20042), .ZN(
        n19675) );
  OAI211_X1 U21780 ( .C1(n20018), .C2(n22084), .A(n19682), .B(n19672), .ZN(
        n20019) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20019), .B1(
        n19673), .B2(n20018), .ZN(n19674) );
  OAI211_X1 U21782 ( .C1(n19676), .C2(n20022), .A(n19675), .B(n19674), .ZN(
        P3_U2899) );
  AND2_X1 U21783 ( .A1(n19687), .A2(n19677), .ZN(n20023) );
  AOI22_X1 U21784 ( .A1(n19952), .A2(n19693), .B1(n19688), .B2(n20023), .ZN(
        n19679) );
  NAND2_X1 U21785 ( .A1(n20036), .A2(n19849), .ZN(n19690) );
  AOI22_X1 U21786 ( .A1(n19947), .A2(n19690), .B1(n19691), .B2(n19677), .ZN(
        n20026) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20026), .B1(
        n19689), .B2(n20042), .ZN(n19678) );
  OAI211_X1 U21788 ( .C1(n19696), .C2(n19764), .A(n19679), .B(n19678), .ZN(
        P3_U2891) );
  NOR2_X1 U21789 ( .A1(n19681), .A2(n19680), .ZN(n20030) );
  AOI22_X1 U21790 ( .A1(n19689), .A2(n19952), .B1(n19688), .B2(n20030), .ZN(
        n19686) );
  AOI22_X1 U21791 ( .A1(n19947), .A2(n19684), .B1(n19683), .B2(n19682), .ZN(
        n20033) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20033), .B1(
        n19693), .B2(n20031), .ZN(n19685) );
  OAI211_X1 U21793 ( .C1(n19696), .C2(n20022), .A(n19686), .B(n19685), .ZN(
        P3_U2883) );
  AND2_X1 U21794 ( .A1(n19687), .A2(n19690), .ZN(n20038) );
  AOI22_X1 U21795 ( .A1(n19689), .A2(n20031), .B1(n19688), .B2(n20038), .ZN(
        n19695) );
  AOI22_X1 U21796 ( .A1(n19947), .A2(n19692), .B1(n19691), .B2(n19690), .ZN(
        n20043) );
  INV_X1 U21797 ( .A(n19944), .ZN(n20040) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20043), .B1(
        n20040), .B2(n19693), .ZN(n19694) );
  OAI211_X1 U21799 ( .C1(n19696), .C2(n19849), .A(n19695), .B(n19694), .ZN(
        P3_U2875) );
  INV_X1 U21800 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n19697) );
  INV_X1 U21801 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21469) );
  AOI22_X1 U21802 ( .A1(n19945), .A2(n19697), .B1(n21469), .B2(U215), .ZN(U257) );
  NAND2_X1 U21803 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19947), .ZN(n19736) );
  NAND2_X1 U21804 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19947), .ZN(n19728) );
  INV_X1 U21805 ( .A(n19728), .ZN(n19732) );
  NOR2_X2 U21806 ( .A1(n21469), .A2(n19863), .ZN(n19731) );
  AOI22_X1 U21807 ( .A1(n20040), .A2(n19732), .B1(n19949), .B2(n19731), .ZN(
        n19700) );
  INV_X1 U21808 ( .A(n19698), .ZN(n21645) );
  NOR2_X2 U21809 ( .A1(n21645), .A2(n19950), .ZN(n19733) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19953), .B1(
        n19952), .B2(n19733), .ZN(n19699) );
  OAI211_X1 U21811 ( .C1(n19956), .C2(n19736), .A(n19700), .B(n19699), .ZN(
        P3_U2994) );
  INV_X1 U21812 ( .A(n19736), .ZN(n19725) );
  AOI22_X1 U21813 ( .A1(n19974), .A2(n19725), .B1(n19957), .B2(n19731), .ZN(
        n19702) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19958), .B1(
        n20031), .B2(n19733), .ZN(n19701) );
  OAI211_X1 U21815 ( .C1(n19956), .C2(n19728), .A(n19702), .B(n19701), .ZN(
        P3_U2986) );
  AOI22_X1 U21816 ( .A1(n19979), .A2(n19725), .B1(n19961), .B2(n19731), .ZN(
        n19704) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19962), .B1(
        n20040), .B2(n19733), .ZN(n19703) );
  OAI211_X1 U21818 ( .C1(n19965), .C2(n19728), .A(n19704), .B(n19703), .ZN(
        P3_U2978) );
  AOI22_X1 U21819 ( .A1(n19985), .A2(n19725), .B1(n19966), .B2(n19731), .ZN(
        n19706) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19968), .B1(
        n19967), .B2(n19733), .ZN(n19705) );
  OAI211_X1 U21821 ( .C1(n19971), .C2(n19728), .A(n19706), .B(n19705), .ZN(
        P3_U2970) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19973), .B1(
        n19972), .B2(n19731), .ZN(n19708) );
  AOI22_X1 U21823 ( .A1(n19974), .A2(n19733), .B1(n19985), .B2(n19732), .ZN(
        n19707) );
  OAI211_X1 U21824 ( .C1(n19983), .C2(n19736), .A(n19708), .B(n19707), .ZN(
        P3_U2962) );
  AOI22_X1 U21825 ( .A1(n19991), .A2(n19732), .B1(n19978), .B2(n19731), .ZN(
        n19710) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19980), .B1(
        n19979), .B2(n19733), .ZN(n19709) );
  OAI211_X1 U21827 ( .C1(n19989), .C2(n19736), .A(n19710), .B(n19709), .ZN(
        P3_U2954) );
  AOI22_X1 U21828 ( .A1(n19996), .A2(n19732), .B1(n19984), .B2(n19731), .ZN(
        n19712) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19733), .ZN(n19711) );
  OAI211_X1 U21830 ( .C1(n19836), .C2(n19736), .A(n19712), .B(n19711), .ZN(
        P3_U2946) );
  AOI22_X1 U21831 ( .A1(n20002), .A2(n19732), .B1(n19990), .B2(n19731), .ZN(
        n19714) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19992), .B1(
        n19991), .B2(n19733), .ZN(n19713) );
  OAI211_X1 U21833 ( .C1(n20000), .C2(n19736), .A(n19714), .B(n19713), .ZN(
        P3_U2938) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19997), .B1(
        n19995), .B2(n19731), .ZN(n19716) );
  AOI22_X1 U21835 ( .A1(n19996), .A2(n19733), .B1(n20013), .B2(n19725), .ZN(
        n19715) );
  OAI211_X1 U21836 ( .C1(n20000), .C2(n19728), .A(n19716), .B(n19715), .ZN(
        P3_U2930) );
  INV_X1 U21837 ( .A(n20013), .ZN(n19925) );
  AOI22_X1 U21838 ( .A1(n20018), .A2(n19725), .B1(n20001), .B2(n19731), .ZN(
        n19718) );
  AOI22_X1 U21839 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20003), .B1(
        n20002), .B2(n19733), .ZN(n19717) );
  OAI211_X1 U21840 ( .C1(n19925), .C2(n19728), .A(n19718), .B(n19717), .ZN(
        P3_U2922) );
  INV_X1 U21841 ( .A(n20018), .ZN(n20011) );
  AOI22_X1 U21842 ( .A1(n20025), .A2(n19725), .B1(n20006), .B2(n19731), .ZN(
        n19720) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20008), .B1(
        n20007), .B2(n19733), .ZN(n19719) );
  OAI211_X1 U21844 ( .C1(n20011), .C2(n19728), .A(n19720), .B(n19719), .ZN(
        P3_U2914) );
  AOI22_X1 U21845 ( .A1(n20025), .A2(n19732), .B1(n20012), .B2(n19731), .ZN(
        n19722) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20014), .B1(
        n20013), .B2(n19733), .ZN(n19721) );
  OAI211_X1 U21847 ( .C1(n20022), .C2(n19736), .A(n19722), .B(n19721), .ZN(
        P3_U2906) );
  AOI22_X1 U21848 ( .A1(n20032), .A2(n19732), .B1(n20017), .B2(n19731), .ZN(
        n19724) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n19733), .ZN(n19723) );
  OAI211_X1 U21850 ( .C1(n19849), .C2(n19736), .A(n19724), .B(n19723), .ZN(
        P3_U2898) );
  AOI22_X1 U21851 ( .A1(n19952), .A2(n19725), .B1(n20023), .B2(n19731), .ZN(
        n19727) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n19733), .ZN(n19726) );
  OAI211_X1 U21853 ( .C1(n19849), .C2(n19728), .A(n19727), .B(n19726), .ZN(
        P3_U2890) );
  AOI22_X1 U21854 ( .A1(n19952), .A2(n19732), .B1(n20030), .B2(n19731), .ZN(
        n19730) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n19733), .ZN(n19729) );
  OAI211_X1 U21856 ( .C1(n20047), .C2(n19736), .A(n19730), .B(n19729), .ZN(
        P3_U2882) );
  AOI22_X1 U21857 ( .A1(n20031), .A2(n19732), .B1(n20038), .B2(n19731), .ZN(
        n19735) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20043), .B1(
        n20042), .B2(n19733), .ZN(n19734) );
  OAI211_X1 U21859 ( .C1(n19944), .C2(n19736), .A(n19735), .B(n19734), .ZN(
        P3_U2874) );
  INV_X1 U21860 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n19737) );
  INV_X1 U21861 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21473) );
  AOI22_X1 U21862 ( .A1(n19738), .A2(n19737), .B1(n21473), .B2(U215), .ZN(U256) );
  NAND2_X1 U21863 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n19947), .ZN(n19772) );
  NOR2_X2 U21864 ( .A1(n21473), .A2(n19863), .ZN(n19773) );
  NAND2_X1 U21865 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19947), .ZN(n19778) );
  AOI22_X1 U21866 ( .A1(n19949), .A2(n19773), .B1(n19967), .B2(n19769), .ZN(
        n19741) );
  NOR2_X2 U21867 ( .A1(n19739), .A2(n19950), .ZN(n19775) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19953), .B1(
        n19952), .B2(n19775), .ZN(n19740) );
  OAI211_X1 U21869 ( .C1(n19944), .C2(n19772), .A(n19741), .B(n19740), .ZN(
        P3_U2993) );
  INV_X1 U21870 ( .A(n19772), .ZN(n19774) );
  AOI22_X1 U21871 ( .A1(n19967), .A2(n19774), .B1(n19957), .B2(n19773), .ZN(
        n19743) );
  AOI22_X1 U21872 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19958), .B1(
        n20031), .B2(n19775), .ZN(n19742) );
  OAI211_X1 U21873 ( .C1(n19965), .C2(n19778), .A(n19743), .B(n19742), .ZN(
        P3_U2985) );
  AOI22_X1 U21874 ( .A1(n19979), .A2(n19769), .B1(n19961), .B2(n19773), .ZN(
        n19745) );
  AOI22_X1 U21875 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19962), .B1(
        n20040), .B2(n19775), .ZN(n19744) );
  OAI211_X1 U21876 ( .C1(n19965), .C2(n19772), .A(n19745), .B(n19744), .ZN(
        P3_U2977) );
  AOI22_X1 U21877 ( .A1(n19979), .A2(n19774), .B1(n19966), .B2(n19773), .ZN(
        n19747) );
  AOI22_X1 U21878 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19968), .B1(
        n19967), .B2(n19775), .ZN(n19746) );
  OAI211_X1 U21879 ( .C1(n19977), .C2(n19778), .A(n19747), .B(n19746), .ZN(
        P3_U2969) );
  AOI22_X1 U21880 ( .A1(n19991), .A2(n19769), .B1(n19972), .B2(n19773), .ZN(
        n19749) );
  AOI22_X1 U21881 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19973), .B1(
        n19974), .B2(n19775), .ZN(n19748) );
  OAI211_X1 U21882 ( .C1(n19977), .C2(n19772), .A(n19749), .B(n19748), .ZN(
        P3_U2961) );
  AOI22_X1 U21883 ( .A1(n19996), .A2(n19769), .B1(n19978), .B2(n19773), .ZN(
        n19751) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19980), .B1(
        n19979), .B2(n19775), .ZN(n19750) );
  OAI211_X1 U21885 ( .C1(n19983), .C2(n19772), .A(n19751), .B(n19750), .ZN(
        P3_U2953) );
  AOI22_X1 U21886 ( .A1(n19996), .A2(n19774), .B1(n19984), .B2(n19773), .ZN(
        n19753) );
  AOI22_X1 U21887 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19775), .ZN(n19752) );
  OAI211_X1 U21888 ( .C1(n19836), .C2(n19778), .A(n19753), .B(n19752), .ZN(
        P3_U2945) );
  AOI22_X1 U21889 ( .A1(n19918), .A2(n19774), .B1(n19990), .B2(n19773), .ZN(
        n19755) );
  AOI22_X1 U21890 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19992), .B1(
        n19991), .B2(n19775), .ZN(n19754) );
  OAI211_X1 U21891 ( .C1(n20000), .C2(n19778), .A(n19755), .B(n19754), .ZN(
        P3_U2937) );
  AOI22_X1 U21892 ( .A1(n20013), .A2(n19769), .B1(n19995), .B2(n19773), .ZN(
        n19757) );
  AOI22_X1 U21893 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19997), .B1(
        n19996), .B2(n19775), .ZN(n19756) );
  OAI211_X1 U21894 ( .C1(n20000), .C2(n19772), .A(n19757), .B(n19756), .ZN(
        P3_U2929) );
  AOI22_X1 U21895 ( .A1(n20018), .A2(n19769), .B1(n20001), .B2(n19773), .ZN(
        n19759) );
  AOI22_X1 U21896 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20003), .B1(
        n20002), .B2(n19775), .ZN(n19758) );
  OAI211_X1 U21897 ( .C1(n19925), .C2(n19772), .A(n19759), .B(n19758), .ZN(
        P3_U2921) );
  AOI22_X1 U21898 ( .A1(n20018), .A2(n19774), .B1(n20006), .B2(n19773), .ZN(
        n19761) );
  AOI22_X1 U21899 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20008), .B1(
        n20007), .B2(n19775), .ZN(n19760) );
  OAI211_X1 U21900 ( .C1(n19764), .C2(n19778), .A(n19761), .B(n19760), .ZN(
        P3_U2913) );
  AOI22_X1 U21901 ( .A1(n20032), .A2(n19769), .B1(n20012), .B2(n19773), .ZN(
        n19763) );
  AOI22_X1 U21902 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20014), .B1(
        n20013), .B2(n19775), .ZN(n19762) );
  OAI211_X1 U21903 ( .C1(n19764), .C2(n19772), .A(n19763), .B(n19762), .ZN(
        P3_U2905) );
  AOI22_X1 U21904 ( .A1(n20042), .A2(n19769), .B1(n20017), .B2(n19773), .ZN(
        n19766) );
  AOI22_X1 U21905 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n19775), .ZN(n19765) );
  OAI211_X1 U21906 ( .C1(n20022), .C2(n19772), .A(n19766), .B(n19765), .ZN(
        P3_U2897) );
  AOI22_X1 U21907 ( .A1(n20042), .A2(n19774), .B1(n20023), .B2(n19773), .ZN(
        n19768) );
  AOI22_X1 U21908 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n19775), .ZN(n19767) );
  OAI211_X1 U21909 ( .C1(n20036), .C2(n19778), .A(n19768), .B(n19767), .ZN(
        P3_U2889) );
  AOI22_X1 U21910 ( .A1(n20031), .A2(n19769), .B1(n20030), .B2(n19773), .ZN(
        n19771) );
  AOI22_X1 U21911 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n19775), .ZN(n19770) );
  OAI211_X1 U21912 ( .C1(n20036), .C2(n19772), .A(n19771), .B(n19770), .ZN(
        P3_U2881) );
  AOI22_X1 U21913 ( .A1(n20031), .A2(n19774), .B1(n20038), .B2(n19773), .ZN(
        n19777) );
  AOI22_X1 U21914 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20043), .B1(
        n20042), .B2(n19775), .ZN(n19776) );
  OAI211_X1 U21915 ( .C1(n19944), .C2(n19778), .A(n19777), .B(n19776), .ZN(
        P3_U2873) );
  INV_X1 U21916 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n19779) );
  INV_X1 U21917 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21478) );
  AOI22_X1 U21918 ( .A1(n19945), .A2(n19779), .B1(n21478), .B2(U215), .ZN(U255) );
  NAND2_X1 U21919 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19947), .ZN(n19817) );
  NOR2_X1 U21920 ( .A1(n21504), .A2(n19862), .ZN(n19813) );
  NOR2_X2 U21921 ( .A1(n21478), .A2(n19863), .ZN(n19812) );
  AOI22_X1 U21922 ( .A1(n20040), .A2(n19813), .B1(n19949), .B2(n19812), .ZN(
        n19781) );
  NOR2_X2 U21923 ( .A1(n21656), .A2(n19950), .ZN(n19814) );
  AOI22_X1 U21924 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19953), .B1(
        n19952), .B2(n19814), .ZN(n19780) );
  OAI211_X1 U21925 ( .C1(n19956), .C2(n19817), .A(n19781), .B(n19780), .ZN(
        P3_U2992) );
  INV_X1 U21926 ( .A(n19813), .ZN(n19811) );
  INV_X1 U21927 ( .A(n19817), .ZN(n19808) );
  AOI22_X1 U21928 ( .A1(n19974), .A2(n19808), .B1(n19957), .B2(n19812), .ZN(
        n19783) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19958), .B1(
        n20031), .B2(n19814), .ZN(n19782) );
  OAI211_X1 U21930 ( .C1(n19956), .C2(n19811), .A(n19783), .B(n19782), .ZN(
        P3_U2984) );
  AOI22_X1 U21931 ( .A1(n19974), .A2(n19813), .B1(n19961), .B2(n19812), .ZN(
        n19785) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19962), .B1(
        n20040), .B2(n19814), .ZN(n19784) );
  OAI211_X1 U21933 ( .C1(n19971), .C2(n19817), .A(n19785), .B(n19784), .ZN(
        P3_U2976) );
  AOI22_X1 U21934 ( .A1(n19979), .A2(n19813), .B1(n19966), .B2(n19812), .ZN(
        n19787) );
  AOI22_X1 U21935 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19968), .B1(
        n19967), .B2(n19814), .ZN(n19786) );
  OAI211_X1 U21936 ( .C1(n19977), .C2(n19817), .A(n19787), .B(n19786), .ZN(
        P3_U2968) );
  AOI22_X1 U21937 ( .A1(n19985), .A2(n19813), .B1(n19972), .B2(n19812), .ZN(
        n19789) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19973), .B1(
        n19974), .B2(n19814), .ZN(n19788) );
  OAI211_X1 U21939 ( .C1(n19983), .C2(n19817), .A(n19789), .B(n19788), .ZN(
        P3_U2960) );
  AOI22_X1 U21940 ( .A1(n19996), .A2(n19808), .B1(n19978), .B2(n19812), .ZN(
        n19791) );
  AOI22_X1 U21941 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19980), .B1(
        n19979), .B2(n19814), .ZN(n19790) );
  OAI211_X1 U21942 ( .C1(n19983), .C2(n19811), .A(n19791), .B(n19790), .ZN(
        P3_U2952) );
  AOI22_X1 U21943 ( .A1(n20002), .A2(n19808), .B1(n19984), .B2(n19812), .ZN(
        n19793) );
  AOI22_X1 U21944 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19814), .ZN(n19792) );
  OAI211_X1 U21945 ( .C1(n19989), .C2(n19811), .A(n19793), .B(n19792), .ZN(
        P3_U2944) );
  AOI22_X1 U21946 ( .A1(n20007), .A2(n19808), .B1(n19990), .B2(n19812), .ZN(
        n19795) );
  AOI22_X1 U21947 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19992), .B1(
        n19991), .B2(n19814), .ZN(n19794) );
  OAI211_X1 U21948 ( .C1(n19836), .C2(n19811), .A(n19795), .B(n19794), .ZN(
        P3_U2936) );
  AOI22_X1 U21949 ( .A1(n20013), .A2(n19808), .B1(n19995), .B2(n19812), .ZN(
        n19797) );
  AOI22_X1 U21950 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19997), .B1(
        n19996), .B2(n19814), .ZN(n19796) );
  OAI211_X1 U21951 ( .C1(n20000), .C2(n19811), .A(n19797), .B(n19796), .ZN(
        P3_U2928) );
  AOI22_X1 U21952 ( .A1(n20018), .A2(n19808), .B1(n20001), .B2(n19812), .ZN(
        n19799) );
  AOI22_X1 U21953 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20003), .B1(
        n20002), .B2(n19814), .ZN(n19798) );
  OAI211_X1 U21954 ( .C1(n19925), .C2(n19811), .A(n19799), .B(n19798), .ZN(
        P3_U2920) );
  AOI22_X1 U21955 ( .A1(n20025), .A2(n19808), .B1(n20006), .B2(n19812), .ZN(
        n19801) );
  AOI22_X1 U21956 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20008), .B1(
        n20007), .B2(n19814), .ZN(n19800) );
  OAI211_X1 U21957 ( .C1(n20011), .C2(n19811), .A(n19801), .B(n19800), .ZN(
        P3_U2912) );
  AOI22_X1 U21958 ( .A1(n20025), .A2(n19813), .B1(n20012), .B2(n19812), .ZN(
        n19803) );
  AOI22_X1 U21959 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20014), .B1(
        n20013), .B2(n19814), .ZN(n19802) );
  OAI211_X1 U21960 ( .C1(n20022), .C2(n19817), .A(n19803), .B(n19802), .ZN(
        P3_U2904) );
  AOI22_X1 U21961 ( .A1(n20032), .A2(n19813), .B1(n20017), .B2(n19812), .ZN(
        n19805) );
  AOI22_X1 U21962 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n19814), .ZN(n19804) );
  OAI211_X1 U21963 ( .C1(n19849), .C2(n19817), .A(n19805), .B(n19804), .ZN(
        P3_U2896) );
  AOI22_X1 U21964 ( .A1(n19952), .A2(n19808), .B1(n20023), .B2(n19812), .ZN(
        n19807) );
  AOI22_X1 U21965 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n19814), .ZN(n19806) );
  OAI211_X1 U21966 ( .C1(n19849), .C2(n19811), .A(n19807), .B(n19806), .ZN(
        P3_U2888) );
  AOI22_X1 U21967 ( .A1(n20031), .A2(n19808), .B1(n20030), .B2(n19812), .ZN(
        n19810) );
  AOI22_X1 U21968 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n19814), .ZN(n19809) );
  OAI211_X1 U21969 ( .C1(n20036), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        P3_U2880) );
  AOI22_X1 U21970 ( .A1(n20031), .A2(n19813), .B1(n20038), .B2(n19812), .ZN(
        n19816) );
  AOI22_X1 U21971 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20043), .B1(
        n20042), .B2(n19814), .ZN(n19815) );
  OAI211_X1 U21972 ( .C1(n19944), .C2(n19817), .A(n19816), .B(n19815), .ZN(
        P3_U2872) );
  INV_X1 U21973 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n19818) );
  INV_X1 U21974 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21482) );
  AOI22_X1 U21975 ( .A1(n19945), .A2(n19818), .B1(n21482), .B2(U215), .ZN(U254) );
  NAND2_X1 U21976 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19947), .ZN(n19859) );
  NAND2_X1 U21977 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19947), .ZN(n19853) );
  INV_X1 U21978 ( .A(n19853), .ZN(n19855) );
  NOR2_X2 U21979 ( .A1(n21482), .A2(n19863), .ZN(n19854) );
  AOI22_X1 U21980 ( .A1(n20040), .A2(n19855), .B1(n19949), .B2(n19854), .ZN(
        n19821) );
  NOR2_X2 U21981 ( .A1(n19819), .A2(n19950), .ZN(n19856) );
  AOI22_X1 U21982 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19953), .B1(
        n19952), .B2(n19856), .ZN(n19820) );
  OAI211_X1 U21983 ( .C1(n19956), .C2(n19859), .A(n19821), .B(n19820), .ZN(
        P3_U2991) );
  AOI22_X1 U21984 ( .A1(n19967), .A2(n19855), .B1(n19957), .B2(n19854), .ZN(
        n19823) );
  AOI22_X1 U21985 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19958), .B1(
        n20031), .B2(n19856), .ZN(n19822) );
  OAI211_X1 U21986 ( .C1(n19965), .C2(n19859), .A(n19823), .B(n19822), .ZN(
        P3_U2983) );
  AOI22_X1 U21987 ( .A1(n19974), .A2(n19855), .B1(n19961), .B2(n19854), .ZN(
        n19825) );
  AOI22_X1 U21988 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19962), .B1(
        n20040), .B2(n19856), .ZN(n19824) );
  OAI211_X1 U21989 ( .C1(n19971), .C2(n19859), .A(n19825), .B(n19824), .ZN(
        P3_U2975) );
  AOI22_X1 U21990 ( .A1(n19979), .A2(n19855), .B1(n19966), .B2(n19854), .ZN(
        n19827) );
  AOI22_X1 U21991 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19968), .B1(
        n19967), .B2(n19856), .ZN(n19826) );
  OAI211_X1 U21992 ( .C1(n19977), .C2(n19859), .A(n19827), .B(n19826), .ZN(
        P3_U2967) );
  AOI22_X1 U21993 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19973), .B1(
        n19972), .B2(n19854), .ZN(n19829) );
  AOI22_X1 U21994 ( .A1(n19974), .A2(n19856), .B1(n19985), .B2(n19855), .ZN(
        n19828) );
  OAI211_X1 U21995 ( .C1(n19983), .C2(n19859), .A(n19829), .B(n19828), .ZN(
        P3_U2959) );
  INV_X1 U21996 ( .A(n19859), .ZN(n19850) );
  AOI22_X1 U21997 ( .A1(n19996), .A2(n19850), .B1(n19978), .B2(n19854), .ZN(
        n19831) );
  AOI22_X1 U21998 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19980), .B1(
        n19979), .B2(n19856), .ZN(n19830) );
  OAI211_X1 U21999 ( .C1(n19983), .C2(n19853), .A(n19831), .B(n19830), .ZN(
        P3_U2951) );
  AOI22_X1 U22000 ( .A1(n20002), .A2(n19850), .B1(n19984), .B2(n19854), .ZN(
        n19833) );
  AOI22_X1 U22001 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19856), .ZN(n19832) );
  OAI211_X1 U22002 ( .C1(n19989), .C2(n19853), .A(n19833), .B(n19832), .ZN(
        P3_U2943) );
  AOI22_X1 U22003 ( .A1(n20007), .A2(n19850), .B1(n19990), .B2(n19854), .ZN(
        n19835) );
  AOI22_X1 U22004 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19992), .B1(
        n19991), .B2(n19856), .ZN(n19834) );
  OAI211_X1 U22005 ( .C1(n19836), .C2(n19853), .A(n19835), .B(n19834), .ZN(
        P3_U2935) );
  AOI22_X1 U22006 ( .A1(n20013), .A2(n19850), .B1(n19995), .B2(n19854), .ZN(
        n19838) );
  AOI22_X1 U22007 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19997), .B1(
        n19996), .B2(n19856), .ZN(n19837) );
  OAI211_X1 U22008 ( .C1(n20000), .C2(n19853), .A(n19838), .B(n19837), .ZN(
        P3_U2927) );
  AOI22_X1 U22009 ( .A1(n20018), .A2(n19850), .B1(n20001), .B2(n19854), .ZN(
        n19840) );
  AOI22_X1 U22010 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20003), .B1(
        n20002), .B2(n19856), .ZN(n19839) );
  OAI211_X1 U22011 ( .C1(n19925), .C2(n19853), .A(n19840), .B(n19839), .ZN(
        P3_U2919) );
  AOI22_X1 U22012 ( .A1(n20025), .A2(n19850), .B1(n20006), .B2(n19854), .ZN(
        n19842) );
  AOI22_X1 U22013 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20008), .B1(
        n20007), .B2(n19856), .ZN(n19841) );
  OAI211_X1 U22014 ( .C1(n20011), .C2(n19853), .A(n19842), .B(n19841), .ZN(
        P3_U2911) );
  AOI22_X1 U22015 ( .A1(n20025), .A2(n19855), .B1(n20012), .B2(n19854), .ZN(
        n19844) );
  AOI22_X1 U22016 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20014), .B1(
        n20013), .B2(n19856), .ZN(n19843) );
  OAI211_X1 U22017 ( .C1(n20022), .C2(n19859), .A(n19844), .B(n19843), .ZN(
        P3_U2903) );
  AOI22_X1 U22018 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20019), .B1(
        n20017), .B2(n19854), .ZN(n19846) );
  AOI22_X1 U22019 ( .A1(n20018), .A2(n19856), .B1(n20032), .B2(n19855), .ZN(
        n19845) );
  OAI211_X1 U22020 ( .C1(n19849), .C2(n19859), .A(n19846), .B(n19845), .ZN(
        P3_U2895) );
  AOI22_X1 U22021 ( .A1(n19952), .A2(n19850), .B1(n20023), .B2(n19854), .ZN(
        n19848) );
  AOI22_X1 U22022 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n19856), .ZN(n19847) );
  OAI211_X1 U22023 ( .C1(n19849), .C2(n19853), .A(n19848), .B(n19847), .ZN(
        P3_U2887) );
  AOI22_X1 U22024 ( .A1(n20031), .A2(n19850), .B1(n20030), .B2(n19854), .ZN(
        n19852) );
  AOI22_X1 U22025 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n19856), .ZN(n19851) );
  OAI211_X1 U22026 ( .C1(n20036), .C2(n19853), .A(n19852), .B(n19851), .ZN(
        P3_U2879) );
  AOI22_X1 U22027 ( .A1(n20031), .A2(n19855), .B1(n20038), .B2(n19854), .ZN(
        n19858) );
  AOI22_X1 U22028 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20043), .B1(
        n20042), .B2(n19856), .ZN(n19857) );
  OAI211_X1 U22029 ( .C1(n19944), .C2(n19859), .A(n19858), .B(n19857), .ZN(
        P3_U2871) );
  INV_X1 U22030 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n19861) );
  INV_X1 U22031 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21488) );
  AOI22_X1 U22032 ( .A1(n19945), .A2(n19861), .B1(n21488), .B2(U215), .ZN(U253) );
  NAND2_X1 U22033 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19947), .ZN(n19896) );
  NOR2_X1 U22034 ( .A1(n19862), .A2(n21520), .ZN(n19893) );
  NOR2_X2 U22035 ( .A1(n19863), .A2(n21488), .ZN(n19897) );
  AOI22_X1 U22036 ( .A1(n20040), .A2(n19893), .B1(n19949), .B2(n19897), .ZN(
        n19865) );
  NOR2_X2 U22037 ( .A1(n21652), .A2(n19950), .ZN(n19899) );
  AOI22_X1 U22038 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19953), .B1(
        n19952), .B2(n19899), .ZN(n19864) );
  OAI211_X1 U22039 ( .C1(n19956), .C2(n19896), .A(n19865), .B(n19864), .ZN(
        P3_U2990) );
  INV_X1 U22040 ( .A(n19896), .ZN(n19898) );
  AOI22_X1 U22041 ( .A1(n19974), .A2(n19898), .B1(n19957), .B2(n19897), .ZN(
        n19867) );
  AOI22_X1 U22042 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19958), .B1(
        n20031), .B2(n19899), .ZN(n19866) );
  OAI211_X1 U22043 ( .C1(n19956), .C2(n19902), .A(n19867), .B(n19866), .ZN(
        P3_U2982) );
  AOI22_X1 U22044 ( .A1(n19974), .A2(n19893), .B1(n19961), .B2(n19897), .ZN(
        n19869) );
  AOI22_X1 U22045 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19962), .B1(
        n20040), .B2(n19899), .ZN(n19868) );
  OAI211_X1 U22046 ( .C1(n19971), .C2(n19896), .A(n19869), .B(n19868), .ZN(
        P3_U2974) );
  AOI22_X1 U22047 ( .A1(n19985), .A2(n19898), .B1(n19966), .B2(n19897), .ZN(
        n19871) );
  AOI22_X1 U22048 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19968), .B1(
        n19967), .B2(n19899), .ZN(n19870) );
  OAI211_X1 U22049 ( .C1(n19971), .C2(n19902), .A(n19871), .B(n19870), .ZN(
        P3_U2966) );
  AOI22_X1 U22050 ( .A1(n19991), .A2(n19898), .B1(n19972), .B2(n19897), .ZN(
        n19873) );
  AOI22_X1 U22051 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19973), .B1(
        n19974), .B2(n19899), .ZN(n19872) );
  OAI211_X1 U22052 ( .C1(n19977), .C2(n19902), .A(n19873), .B(n19872), .ZN(
        P3_U2958) );
  AOI22_X1 U22053 ( .A1(n19996), .A2(n19898), .B1(n19978), .B2(n19897), .ZN(
        n19875) );
  AOI22_X1 U22054 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19980), .B1(
        n19979), .B2(n19899), .ZN(n19874) );
  OAI211_X1 U22055 ( .C1(n19983), .C2(n19902), .A(n19875), .B(n19874), .ZN(
        P3_U2950) );
  AOI22_X1 U22056 ( .A1(n20002), .A2(n19898), .B1(n19984), .B2(n19897), .ZN(
        n19877) );
  AOI22_X1 U22057 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19899), .ZN(n19876) );
  OAI211_X1 U22058 ( .C1(n19989), .C2(n19902), .A(n19877), .B(n19876), .ZN(
        P3_U2942) );
  AOI22_X1 U22059 ( .A1(n19918), .A2(n19893), .B1(n19990), .B2(n19897), .ZN(
        n19879) );
  AOI22_X1 U22060 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19992), .B1(
        n19991), .B2(n19899), .ZN(n19878) );
  OAI211_X1 U22061 ( .C1(n20000), .C2(n19896), .A(n19879), .B(n19878), .ZN(
        P3_U2934) );
  AOI22_X1 U22062 ( .A1(n20013), .A2(n19898), .B1(n19995), .B2(n19897), .ZN(
        n19881) );
  AOI22_X1 U22063 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19997), .B1(
        n19996), .B2(n19899), .ZN(n19880) );
  OAI211_X1 U22064 ( .C1(n20000), .C2(n19902), .A(n19881), .B(n19880), .ZN(
        P3_U2926) );
  AOI22_X1 U22065 ( .A1(n20018), .A2(n19898), .B1(n20001), .B2(n19897), .ZN(
        n19883) );
  AOI22_X1 U22066 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20003), .B1(
        n20002), .B2(n19899), .ZN(n19882) );
  OAI211_X1 U22067 ( .C1(n19925), .C2(n19902), .A(n19883), .B(n19882), .ZN(
        P3_U2918) );
  AOI22_X1 U22068 ( .A1(n19884), .A2(n19898), .B1(n20006), .B2(n19897), .ZN(
        n19886) );
  AOI22_X1 U22069 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20008), .B1(
        n20007), .B2(n19899), .ZN(n19885) );
  OAI211_X1 U22070 ( .C1(n20011), .C2(n19902), .A(n19886), .B(n19885), .ZN(
        P3_U2910) );
  AOI22_X1 U22071 ( .A1(n20025), .A2(n19893), .B1(n20012), .B2(n19897), .ZN(
        n19888) );
  AOI22_X1 U22072 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20014), .B1(
        n20013), .B2(n19899), .ZN(n19887) );
  OAI211_X1 U22073 ( .C1(n20022), .C2(n19896), .A(n19888), .B(n19887), .ZN(
        P3_U2902) );
  AOI22_X1 U22074 ( .A1(n20042), .A2(n19898), .B1(n20017), .B2(n19897), .ZN(
        n19890) );
  AOI22_X1 U22075 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n19899), .ZN(n19889) );
  OAI211_X1 U22076 ( .C1(n20022), .C2(n19902), .A(n19890), .B(n19889), .ZN(
        P3_U2894) );
  AOI22_X1 U22077 ( .A1(n20042), .A2(n19893), .B1(n20023), .B2(n19897), .ZN(
        n19892) );
  AOI22_X1 U22078 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n19899), .ZN(n19891) );
  OAI211_X1 U22079 ( .C1(n20036), .C2(n19896), .A(n19892), .B(n19891), .ZN(
        P3_U2886) );
  AOI22_X1 U22080 ( .A1(n19952), .A2(n19893), .B1(n20030), .B2(n19897), .ZN(
        n19895) );
  AOI22_X1 U22081 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n19899), .ZN(n19894) );
  OAI211_X1 U22082 ( .C1(n20047), .C2(n19896), .A(n19895), .B(n19894), .ZN(
        P3_U2878) );
  AOI22_X1 U22083 ( .A1(n20040), .A2(n19898), .B1(n20038), .B2(n19897), .ZN(
        n19901) );
  AOI22_X1 U22084 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20043), .B1(
        n20042), .B2(n19899), .ZN(n19900) );
  OAI211_X1 U22085 ( .C1(n20047), .C2(n19902), .A(n19901), .B(n19900), .ZN(
        P3_U2870) );
  OAI22_X1 U22086 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19945), .ZN(n19903) );
  INV_X1 U22087 ( .A(n19903), .ZN(U252) );
  NAND2_X1 U22088 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19947), .ZN(n19943) );
  NAND2_X1 U22089 ( .A1(n19947), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19937) );
  AND2_X1 U22090 ( .A1(n19948), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19938) );
  AOI22_X1 U22091 ( .A1(n20040), .A2(n19939), .B1(n19949), .B2(n19938), .ZN(
        n19905) );
  NOR2_X2 U22092 ( .A1(n20959), .A2(n19950), .ZN(n19940) );
  AOI22_X1 U22093 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19953), .B1(
        n19952), .B2(n19940), .ZN(n19904) );
  OAI211_X1 U22094 ( .C1(n19956), .C2(n19943), .A(n19905), .B(n19904), .ZN(
        P3_U2989) );
  INV_X1 U22095 ( .A(n19943), .ZN(n19934) );
  AOI22_X1 U22096 ( .A1(n19974), .A2(n19934), .B1(n19957), .B2(n19938), .ZN(
        n19907) );
  AOI22_X1 U22097 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19958), .B1(
        n20031), .B2(n19940), .ZN(n19906) );
  OAI211_X1 U22098 ( .C1(n19956), .C2(n19937), .A(n19907), .B(n19906), .ZN(
        P3_U2981) );
  AOI22_X1 U22099 ( .A1(n19974), .A2(n19939), .B1(n19961), .B2(n19938), .ZN(
        n19909) );
  AOI22_X1 U22100 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19962), .B1(
        n20040), .B2(n19940), .ZN(n19908) );
  OAI211_X1 U22101 ( .C1(n19971), .C2(n19943), .A(n19909), .B(n19908), .ZN(
        P3_U2973) );
  AOI22_X1 U22102 ( .A1(n19985), .A2(n19934), .B1(n19966), .B2(n19938), .ZN(
        n19911) );
  AOI22_X1 U22103 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19968), .B1(
        n19967), .B2(n19940), .ZN(n19910) );
  OAI211_X1 U22104 ( .C1(n19971), .C2(n19937), .A(n19911), .B(n19910), .ZN(
        P3_U2965) );
  AOI22_X1 U22105 ( .A1(n19991), .A2(n19934), .B1(n19972), .B2(n19938), .ZN(
        n19913) );
  AOI22_X1 U22106 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19973), .B1(
        n19974), .B2(n19940), .ZN(n19912) );
  OAI211_X1 U22107 ( .C1(n19977), .C2(n19937), .A(n19913), .B(n19912), .ZN(
        P3_U2957) );
  AOI22_X1 U22108 ( .A1(n19991), .A2(n19939), .B1(n19978), .B2(n19938), .ZN(
        n19915) );
  AOI22_X1 U22109 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19980), .B1(
        n19979), .B2(n19940), .ZN(n19914) );
  OAI211_X1 U22110 ( .C1(n19989), .C2(n19943), .A(n19915), .B(n19914), .ZN(
        P3_U2949) );
  AOI22_X1 U22111 ( .A1(n19918), .A2(n19934), .B1(n19984), .B2(n19938), .ZN(
        n19917) );
  AOI22_X1 U22112 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19940), .ZN(n19916) );
  OAI211_X1 U22113 ( .C1(n19989), .C2(n19937), .A(n19917), .B(n19916), .ZN(
        P3_U2941) );
  AOI22_X1 U22114 ( .A1(n19918), .A2(n19939), .B1(n19990), .B2(n19938), .ZN(
        n19920) );
  AOI22_X1 U22115 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19992), .B1(
        n19991), .B2(n19940), .ZN(n19919) );
  OAI211_X1 U22116 ( .C1(n20000), .C2(n19943), .A(n19920), .B(n19919), .ZN(
        P3_U2933) );
  AOI22_X1 U22117 ( .A1(n20007), .A2(n19939), .B1(n19995), .B2(n19938), .ZN(
        n19922) );
  AOI22_X1 U22118 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19997), .B1(
        n19996), .B2(n19940), .ZN(n19921) );
  OAI211_X1 U22119 ( .C1(n19925), .C2(n19943), .A(n19922), .B(n19921), .ZN(
        P3_U2925) );
  AOI22_X1 U22120 ( .A1(n20018), .A2(n19934), .B1(n20001), .B2(n19938), .ZN(
        n19924) );
  AOI22_X1 U22121 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20003), .B1(
        n20002), .B2(n19940), .ZN(n19923) );
  OAI211_X1 U22122 ( .C1(n19925), .C2(n19937), .A(n19924), .B(n19923), .ZN(
        P3_U2917) );
  AOI22_X1 U22123 ( .A1(n20025), .A2(n19934), .B1(n20006), .B2(n19938), .ZN(
        n19927) );
  AOI22_X1 U22124 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20008), .B1(
        n20007), .B2(n19940), .ZN(n19926) );
  OAI211_X1 U22125 ( .C1(n20011), .C2(n19937), .A(n19927), .B(n19926), .ZN(
        P3_U2909) );
  AOI22_X1 U22126 ( .A1(n20025), .A2(n19939), .B1(n20012), .B2(n19938), .ZN(
        n19929) );
  AOI22_X1 U22127 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20014), .B1(
        n20013), .B2(n19940), .ZN(n19928) );
  OAI211_X1 U22128 ( .C1(n20022), .C2(n19943), .A(n19929), .B(n19928), .ZN(
        P3_U2901) );
  AOI22_X1 U22129 ( .A1(n20042), .A2(n19934), .B1(n20017), .B2(n19938), .ZN(
        n19931) );
  AOI22_X1 U22130 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n19940), .ZN(n19930) );
  OAI211_X1 U22131 ( .C1(n20022), .C2(n19937), .A(n19931), .B(n19930), .ZN(
        P3_U2893) );
  AOI22_X1 U22132 ( .A1(n20042), .A2(n19939), .B1(n20023), .B2(n19938), .ZN(
        n19933) );
  AOI22_X1 U22133 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n19940), .ZN(n19932) );
  OAI211_X1 U22134 ( .C1(n20036), .C2(n19943), .A(n19933), .B(n19932), .ZN(
        P3_U2885) );
  AOI22_X1 U22135 ( .A1(n20031), .A2(n19934), .B1(n20030), .B2(n19938), .ZN(
        n19936) );
  AOI22_X1 U22136 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n19940), .ZN(n19935) );
  OAI211_X1 U22137 ( .C1(n20036), .C2(n19937), .A(n19936), .B(n19935), .ZN(
        P3_U2877) );
  AOI22_X1 U22138 ( .A1(n20031), .A2(n19939), .B1(n20038), .B2(n19938), .ZN(
        n19942) );
  AOI22_X1 U22139 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20043), .B1(
        n20042), .B2(n19940), .ZN(n19941) );
  OAI211_X1 U22140 ( .C1(n19944), .C2(n19943), .A(n19942), .B(n19941), .ZN(
        P3_U2869) );
  OAI22_X1 U22141 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19945), .ZN(n19946) );
  INV_X1 U22142 ( .A(n19946), .ZN(U251) );
  NAND2_X1 U22143 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19947), .ZN(n20029) );
  NAND2_X1 U22144 ( .A1(n19947), .A2(BUF2_REG_16__SCAN_IN), .ZN(n20046) );
  INV_X1 U22145 ( .A(n20046), .ZN(n20024) );
  AND2_X1 U22146 ( .A1(n19948), .A2(BUF2_REG_0__SCAN_IN), .ZN(n20037) );
  AOI22_X1 U22147 ( .A1(n20040), .A2(n20024), .B1(n19949), .B2(n20037), .ZN(
        n19955) );
  NOR2_X2 U22148 ( .A1(n19951), .A2(n19950), .ZN(n20041) );
  AOI22_X1 U22149 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19953), .B1(
        n19952), .B2(n20041), .ZN(n19954) );
  OAI211_X1 U22150 ( .C1(n19956), .C2(n20029), .A(n19955), .B(n19954), .ZN(
        P3_U2988) );
  AOI22_X1 U22151 ( .A1(n19967), .A2(n20024), .B1(n19957), .B2(n20037), .ZN(
        n19960) );
  AOI22_X1 U22152 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19958), .B1(
        n20031), .B2(n20041), .ZN(n19959) );
  OAI211_X1 U22153 ( .C1(n19965), .C2(n20029), .A(n19960), .B(n19959), .ZN(
        P3_U2980) );
  INV_X1 U22154 ( .A(n20029), .ZN(n20039) );
  AOI22_X1 U22155 ( .A1(n19979), .A2(n20039), .B1(n19961), .B2(n20037), .ZN(
        n19964) );
  AOI22_X1 U22156 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19962), .B1(
        n20040), .B2(n20041), .ZN(n19963) );
  OAI211_X1 U22157 ( .C1(n19965), .C2(n20046), .A(n19964), .B(n19963), .ZN(
        P3_U2972) );
  AOI22_X1 U22158 ( .A1(n19985), .A2(n20039), .B1(n19966), .B2(n20037), .ZN(
        n19970) );
  AOI22_X1 U22159 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19968), .B1(
        n19967), .B2(n20041), .ZN(n19969) );
  OAI211_X1 U22160 ( .C1(n19971), .C2(n20046), .A(n19970), .B(n19969), .ZN(
        P3_U2964) );
  AOI22_X1 U22161 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19973), .B1(
        n19972), .B2(n20037), .ZN(n19976) );
  AOI22_X1 U22162 ( .A1(n19974), .A2(n20041), .B1(n19991), .B2(n20039), .ZN(
        n19975) );
  OAI211_X1 U22163 ( .C1(n19977), .C2(n20046), .A(n19976), .B(n19975), .ZN(
        P3_U2956) );
  AOI22_X1 U22164 ( .A1(n19996), .A2(n20039), .B1(n19978), .B2(n20037), .ZN(
        n19982) );
  AOI22_X1 U22165 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19980), .B1(
        n19979), .B2(n20041), .ZN(n19981) );
  OAI211_X1 U22166 ( .C1(n19983), .C2(n20046), .A(n19982), .B(n19981), .ZN(
        P3_U2948) );
  AOI22_X1 U22167 ( .A1(n20002), .A2(n20039), .B1(n19984), .B2(n20037), .ZN(
        n19988) );
  AOI22_X1 U22168 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n20041), .ZN(n19987) );
  OAI211_X1 U22169 ( .C1(n19989), .C2(n20046), .A(n19988), .B(n19987), .ZN(
        P3_U2940) );
  AOI22_X1 U22170 ( .A1(n20002), .A2(n20024), .B1(n19990), .B2(n20037), .ZN(
        n19994) );
  AOI22_X1 U22171 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19992), .B1(
        n19991), .B2(n20041), .ZN(n19993) );
  OAI211_X1 U22172 ( .C1(n20000), .C2(n20029), .A(n19994), .B(n19993), .ZN(
        P3_U2932) );
  AOI22_X1 U22173 ( .A1(n20013), .A2(n20039), .B1(n19995), .B2(n20037), .ZN(
        n19999) );
  AOI22_X1 U22174 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19997), .B1(
        n19996), .B2(n20041), .ZN(n19998) );
  OAI211_X1 U22175 ( .C1(n20000), .C2(n20046), .A(n19999), .B(n19998), .ZN(
        P3_U2924) );
  AOI22_X1 U22176 ( .A1(n20013), .A2(n20024), .B1(n20001), .B2(n20037), .ZN(
        n20005) );
  AOI22_X1 U22177 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20003), .B1(
        n20002), .B2(n20041), .ZN(n20004) );
  OAI211_X1 U22178 ( .C1(n20011), .C2(n20029), .A(n20005), .B(n20004), .ZN(
        P3_U2916) );
  AOI22_X1 U22179 ( .A1(n20025), .A2(n20039), .B1(n20006), .B2(n20037), .ZN(
        n20010) );
  AOI22_X1 U22180 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20008), .B1(
        n20007), .B2(n20041), .ZN(n20009) );
  OAI211_X1 U22181 ( .C1(n20011), .C2(n20046), .A(n20010), .B(n20009), .ZN(
        P3_U2908) );
  AOI22_X1 U22182 ( .A1(n20025), .A2(n20024), .B1(n20012), .B2(n20037), .ZN(
        n20016) );
  AOI22_X1 U22183 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20014), .B1(
        n20013), .B2(n20041), .ZN(n20015) );
  OAI211_X1 U22184 ( .C1(n20022), .C2(n20029), .A(n20016), .B(n20015), .ZN(
        P3_U2900) );
  AOI22_X1 U22185 ( .A1(n20042), .A2(n20039), .B1(n20017), .B2(n20037), .ZN(
        n20021) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20019), .B1(
        n20018), .B2(n20041), .ZN(n20020) );
  OAI211_X1 U22187 ( .C1(n20022), .C2(n20046), .A(n20021), .B(n20020), .ZN(
        P3_U2892) );
  AOI22_X1 U22188 ( .A1(n20042), .A2(n20024), .B1(n20023), .B2(n20037), .ZN(
        n20028) );
  AOI22_X1 U22189 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20041), .ZN(n20027) );
  OAI211_X1 U22190 ( .C1(n20036), .C2(n20029), .A(n20028), .B(n20027), .ZN(
        P3_U2884) );
  AOI22_X1 U22191 ( .A1(n20031), .A2(n20039), .B1(n20030), .B2(n20037), .ZN(
        n20035) );
  AOI22_X1 U22192 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n20041), .ZN(n20034) );
  OAI211_X1 U22193 ( .C1(n20036), .C2(n20046), .A(n20035), .B(n20034), .ZN(
        P3_U2876) );
  AOI22_X1 U22194 ( .A1(n20040), .A2(n20039), .B1(n20038), .B2(n20037), .ZN(
        n20045) );
  AOI22_X1 U22195 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20043), .B1(
        n20042), .B2(n20041), .ZN(n20044) );
  OAI211_X1 U22196 ( .C1(n20047), .C2(n20046), .A(n20045), .B(n20044), .ZN(
        P3_U2868) );
  AOI22_X1 U22197 ( .A1(n20049), .A2(n20497), .B1(BUF2_REG_31__SCAN_IN), .B2(
        n20048), .ZN(n20052) );
  AOI22_X1 U22198 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n20495), .B1(n20050), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n20051) );
  NAND2_X1 U22199 ( .A1(n20052), .A2(n20051), .ZN(P2_U2888) );
  AOI22_X1 U22200 ( .A1(P2_EAX_REG_15__SCAN_IN), .A2(n20495), .B1(n20053), 
        .B2(n20313), .ZN(n20054) );
  OAI21_X1 U22201 ( .B1(n20557), .B2(n20055), .A(n20054), .ZN(P2_U2904) );
  OAI222_X1 U22202 ( .A1(n20058), .A2(n20081), .B1(n20057), .B2(n20546), .C1(
        n20557), .C2(n20056), .ZN(P2_U2905) );
  AOI22_X1 U22203 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(n20495), .B1(n20059), 
        .B2(n20313), .ZN(n20060) );
  OAI21_X1 U22204 ( .B1(n20061), .B2(n20557), .A(n20060), .ZN(P2_U2906) );
  OAI222_X1 U22205 ( .A1(n20064), .A2(n20081), .B1(n20063), .B2(n20546), .C1(
        n20557), .C2(n20062), .ZN(P2_U2907) );
  AOI22_X1 U22206 ( .A1(n20066), .A2(n20313), .B1(n20065), .B2(n20072), .ZN(
        n20067) );
  OAI21_X1 U22207 ( .B1(n20546), .B2(n20068), .A(n20067), .ZN(P2_U2908) );
  AOI22_X1 U22208 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n20495), .B1(n20069), 
        .B2(n20313), .ZN(n20070) );
  OAI21_X1 U22209 ( .B1(n20071), .B2(n20557), .A(n20070), .ZN(P2_U2909) );
  AOI22_X1 U22210 ( .A1(n20074), .A2(n20313), .B1(n20073), .B2(n20072), .ZN(
        n20075) );
  OAI21_X1 U22211 ( .B1(n20546), .B2(n20076), .A(n20075), .ZN(P2_U2910) );
  OAI222_X1 U22212 ( .A1(n20079), .A2(n20081), .B1(n20078), .B2(n20546), .C1(
        n20557), .C2(n20077), .ZN(P2_U2911) );
  OAI222_X1 U22213 ( .A1(n20082), .A2(n20081), .B1(n20080), .B2(n20546), .C1(
        n20557), .C2(n20085), .ZN(P2_U2912) );
  OAI22_X2 U22214 ( .A1(n20083), .A2(n20456), .B1(n20934), .B2(n20455), .ZN(
        n20265) );
  INV_X1 U22215 ( .A(n20265), .ZN(n20262) );
  NAND3_X1 U22216 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20094) );
  OAI21_X1 U22217 ( .B1(n20088), .B2(n20561), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20084) );
  OAI21_X1 U22218 ( .B1(n20094), .B2(n20254), .A(n20084), .ZN(n20562) );
  NOR2_X2 U22219 ( .A1(n20087), .A2(n20454), .ZN(n20263) );
  AOI22_X1 U22220 ( .A1(n20562), .A2(n20086), .B1(n20561), .B2(n20263), .ZN(
        n20093) );
  INV_X1 U22221 ( .A(n20244), .ZN(n20264) );
  INV_X1 U22222 ( .A(n20209), .ZN(n20253) );
  AOI211_X1 U22223 ( .C1(n20088), .C2(n20253), .A(n20561), .B(n20222), .ZN(
        n20089) );
  NOR2_X1 U22224 ( .A1(n20558), .A2(n20089), .ZN(n20091) );
  OAI21_X1 U22225 ( .B1(n20109), .B2(n20173), .A(n20094), .ZN(n20090) );
  NAND2_X1 U22226 ( .A1(n20091), .A2(n20090), .ZN(n20565) );
  AOI22_X1 U22227 ( .A1(n20264), .A2(n20570), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n20565), .ZN(n20092) );
  OAI211_X1 U22228 ( .C1(n20262), .C2(n20412), .A(n20093), .B(n20092), .ZN(
        P2_U3175) );
  NOR2_X1 U22229 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20094), .ZN(
        n20569) );
  AOI22_X1 U22230 ( .A1(n20570), .A2(n20265), .B1(n20263), .B2(n20569), .ZN(
        n20105) );
  INV_X1 U22231 ( .A(n20184), .ZN(n20095) );
  OAI21_X1 U22232 ( .B1(n20096), .B2(n20209), .A(n20095), .ZN(n20099) );
  NOR2_X1 U22233 ( .A1(n20570), .A2(n20507), .ZN(n20097) );
  OAI21_X1 U22234 ( .B1(n20097), .B2(n22410), .A(n20222), .ZN(n20103) );
  NAND3_X1 U22235 ( .A1(n20245), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20118) );
  NOR2_X1 U22236 ( .A1(n20247), .A2(n20118), .ZN(n20575) );
  OR2_X1 U22237 ( .A1(n20103), .A2(n20575), .ZN(n20098) );
  AOI22_X1 U22238 ( .A1(n20099), .A2(n20098), .B1(n20569), .B2(n20257), .ZN(
        n20572) );
  NOR2_X1 U22239 ( .A1(n20575), .A2(n20569), .ZN(n20102) );
  OAI21_X1 U22240 ( .B1(n20100), .B2(n20569), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20101) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20572), .B1(
        n20086), .B2(n20571), .ZN(n20104) );
  OAI211_X1 U22242 ( .C1(n20244), .C2(n20580), .A(n20105), .B(n20104), .ZN(
        P2_U3167) );
  OAI21_X1 U22243 ( .B1(n20106), .B2(n20575), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20107) );
  OAI21_X1 U22244 ( .B1(n20118), .B2(n20254), .A(n20107), .ZN(n20576) );
  AOI22_X1 U22245 ( .A1(n20576), .A2(n20086), .B1(n20263), .B2(n20575), .ZN(
        n20116) );
  NAND2_X1 U22246 ( .A1(n20108), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20251) );
  OAI21_X1 U22247 ( .B1(n20109), .B2(n20251), .A(n20118), .ZN(n20113) );
  AOI21_X1 U22248 ( .B1(n20257), .B2(n20575), .A(n20184), .ZN(n20110) );
  OAI21_X1 U22249 ( .B1(n20111), .B2(n20209), .A(n20110), .ZN(n20112) );
  NAND2_X1 U22250 ( .A1(n20113), .A2(n20112), .ZN(n20577) );
  NAND2_X1 U22251 ( .A1(n20191), .A2(n20114), .ZN(n20510) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20577), .B1(
        n20583), .B2(n20264), .ZN(n20115) );
  OAI211_X1 U22253 ( .C1(n20262), .C2(n20580), .A(n20116), .B(n20115), .ZN(
        P2_U3159) );
  NAND2_X1 U22254 ( .A1(n20117), .A2(n20183), .ZN(n20207) );
  NOR2_X1 U22255 ( .A1(n20140), .A2(n20207), .ZN(n20124) );
  INV_X1 U22256 ( .A(n20124), .ZN(n20120) );
  NOR2_X1 U22257 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20118), .ZN(
        n20581) );
  OAI21_X1 U22258 ( .B1(n20121), .B2(n20581), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20119) );
  OAI21_X1 U22259 ( .B1(n20120), .B2(n20254), .A(n20119), .ZN(n20582) );
  AOI22_X1 U22260 ( .A1(n20582), .A2(n20086), .B1(n20263), .B2(n20581), .ZN(
        n20127) );
  AOI21_X1 U22261 ( .B1(n20593), .B2(n20510), .A(n22410), .ZN(n20125) );
  AOI211_X1 U22262 ( .C1(n20121), .C2(n20253), .A(n20222), .B(n20581), .ZN(
        n20122) );
  NOR2_X1 U22263 ( .A1(n20558), .A2(n20122), .ZN(n20123) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20265), .ZN(n20126) );
  OAI211_X1 U22265 ( .C1(n20244), .C2(n20593), .A(n20127), .B(n20126), .ZN(
        P2_U3151) );
  NAND3_X1 U22266 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20161), .ZN(n20137) );
  INV_X1 U22267 ( .A(n20128), .ZN(n20130) );
  NOR2_X1 U22268 ( .A1(n20247), .A2(n20137), .ZN(n20587) );
  OAI21_X1 U22269 ( .B1(n20130), .B2(n20587), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20129) );
  OAI21_X1 U22270 ( .B1(n20137), .B2(n20254), .A(n20129), .ZN(n20588) );
  AOI22_X1 U22271 ( .A1(n20588), .A2(n20086), .B1(n20263), .B2(n20587), .ZN(
        n20136) );
  AOI211_X1 U22272 ( .C1(n20130), .C2(n20253), .A(n20184), .B(n20587), .ZN(
        n20131) );
  NOR2_X1 U22273 ( .A1(n20558), .A2(n20131), .ZN(n20134) );
  OAI21_X1 U22274 ( .B1(n20132), .B2(n20220), .A(n20137), .ZN(n20133) );
  NAND2_X1 U22275 ( .A1(n20134), .A2(n20133), .ZN(n20590) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20264), .ZN(n20135) );
  OAI211_X1 U22277 ( .C1(n20262), .C2(n20593), .A(n20136), .B(n20135), .ZN(
        P2_U3143) );
  AOI22_X1 U22278 ( .A1(n20589), .A2(n20265), .B1(n20263), .B2(n20594), .ZN(
        n20148) );
  INV_X1 U22279 ( .A(n20138), .ZN(n20143) );
  NOR3_X1 U22280 ( .A1(n20143), .A2(n20594), .A3(n20235), .ZN(n20142) );
  NOR2_X1 U22281 ( .A1(n20595), .A2(n20589), .ZN(n20139) );
  OAI21_X1 U22282 ( .B1(n20139), .B2(n22410), .A(n20222), .ZN(n20146) );
  NOR3_X1 U22283 ( .A1(n20140), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20153) );
  INV_X1 U22284 ( .A(n20153), .ZN(n20159) );
  NOR2_X1 U22285 ( .A1(n20601), .A2(n20594), .ZN(n20145) );
  OAI21_X1 U22286 ( .B1(n20143), .B2(n20594), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20144) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20597), .B1(
        n20086), .B2(n20596), .ZN(n20147) );
  OAI211_X1 U22288 ( .C1(n20244), .C2(n20606), .A(n20148), .B(n20147), .ZN(
        P2_U3135) );
  AOI22_X1 U22289 ( .A1(n20595), .A2(n20265), .B1(n20263), .B2(n20601), .ZN(
        n20158) );
  OAI21_X1 U22290 ( .B1(n20150), .B2(n20251), .A(n20222), .ZN(n20156) );
  NOR2_X1 U22291 ( .A1(n20558), .A2(n20151), .ZN(n20152) );
  OAI21_X1 U22292 ( .B1(n20156), .B2(n20153), .A(n20152), .ZN(n20603) );
  OAI21_X1 U22293 ( .B1(n20154), .B2(n20601), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20155) );
  OAI21_X1 U22294 ( .B1(n20156), .B2(n20159), .A(n20155), .ZN(n20602) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20603), .B1(
        n20086), .B2(n20602), .ZN(n20157) );
  OAI211_X1 U22296 ( .C1(n20244), .C2(n20519), .A(n20158), .B(n20157), .ZN(
        P2_U3127) );
  NOR2_X1 U22297 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20159), .ZN(
        n20607) );
  AOI22_X1 U22298 ( .A1(n20608), .A2(n20265), .B1(n20263), .B2(n20607), .ZN(
        n20170) );
  NAND2_X1 U22299 ( .A1(n20519), .A2(n20619), .ZN(n20160) );
  AOI21_X1 U22300 ( .B1(n20160), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20254), 
        .ZN(n20165) );
  NOR2_X1 U22301 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20161), .ZN(
        n20204) );
  NAND2_X1 U22302 ( .A1(n20219), .A2(n20204), .ZN(n20174) );
  OAI21_X1 U22303 ( .B1(n20166), .B2(n20235), .A(n20162), .ZN(n20163) );
  AOI21_X1 U22304 ( .B1(n20165), .B2(n20174), .A(n20163), .ZN(n20164) );
  OAI21_X1 U22305 ( .B1(n20607), .B2(n20164), .A(n20257), .ZN(n20610) );
  INV_X1 U22306 ( .A(n20174), .ZN(n20613) );
  OAI21_X1 U22307 ( .B1(n20613), .B2(n20607), .A(n20165), .ZN(n20168) );
  OAI21_X1 U22308 ( .B1(n20166), .B2(n20607), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20167) );
  NAND2_X1 U22309 ( .A1(n20168), .A2(n20167), .ZN(n20609) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20610), .B1(
        n20609), .B2(n20086), .ZN(n20169) );
  OAI211_X1 U22311 ( .C1(n20244), .C2(n20619), .A(n20170), .B(n20169), .ZN(
        P2_U3119) );
  NAND2_X1 U22312 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20204), .ZN(
        n20179) );
  OAI21_X1 U22313 ( .B1(n20171), .B2(n20613), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20172) );
  OAI21_X1 U22314 ( .B1(n20179), .B2(n20254), .A(n20172), .ZN(n20614) );
  AOI22_X1 U22315 ( .A1(n20614), .A2(n20086), .B1(n20613), .B2(n20263), .ZN(
        n20178) );
  OAI21_X1 U22316 ( .B1(n20193), .B2(n20173), .A(n20179), .ZN(n20176) );
  OAI211_X1 U22317 ( .C1(n12577), .C2(n20209), .A(n20174), .B(n20254), .ZN(
        n20175) );
  NAND3_X1 U22318 ( .A1(n20176), .A2(n20257), .A3(n20175), .ZN(n20616) );
  INV_X1 U22319 ( .A(n20619), .ZN(n20289) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20616), .B1(
        n20289), .B2(n20265), .ZN(n20177) );
  OAI211_X1 U22321 ( .C1(n20244), .C2(n20625), .A(n20178), .B(n20177), .ZN(
        P2_U3111) );
  INV_X1 U22322 ( .A(n20204), .ZN(n20182) );
  INV_X1 U22323 ( .A(n12568), .ZN(n20180) );
  NOR2_X1 U22324 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20179), .ZN(
        n20620) );
  OAI21_X1 U22325 ( .B1(n20180), .B2(n20620), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20181) );
  OAI21_X1 U22326 ( .B1(n20182), .B2(n20233), .A(n20181), .ZN(n20621) );
  AOI22_X1 U22327 ( .A1(n20621), .A2(n20086), .B1(n20263), .B2(n20620), .ZN(
        n20190) );
  AOI21_X1 U22328 ( .B1(n20625), .B2(n20528), .A(n22410), .ZN(n20188) );
  NOR2_X1 U22329 ( .A1(n20183), .A2(n20182), .ZN(n20187) );
  NOR2_X1 U22330 ( .A1(n20184), .A2(n20620), .ZN(n20185) );
  OAI21_X1 U22331 ( .B1(n12568), .B2(n20209), .A(n20185), .ZN(n20186) );
  OAI211_X1 U22332 ( .C1(n20188), .C2(n20187), .A(n20257), .B(n20186), .ZN(
        n20622) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20622), .B1(
        n20615), .B2(n20265), .ZN(n20189) );
  OAI211_X1 U22334 ( .C1(n20244), .C2(n20528), .A(n20190), .B(n20189), .ZN(
        P2_U3103) );
  NAND2_X1 U22335 ( .A1(n20204), .A2(n20245), .ZN(n20199) );
  NOR2_X1 U22336 ( .A1(n20247), .A2(n20199), .ZN(n20626) );
  AOI22_X1 U22337 ( .A1(n20265), .A2(n20627), .B1(n20263), .B2(n20626), .ZN(
        n20202) );
  OAI21_X1 U22338 ( .B1(n20193), .B2(n20251), .A(n20222), .ZN(n20200) );
  INV_X1 U22339 ( .A(n20199), .ZN(n20196) );
  OAI21_X1 U22340 ( .B1(n20222), .B2(n20626), .A(n20257), .ZN(n20194) );
  OAI21_X1 U22341 ( .B1(n12576), .B2(n20209), .A(n20194), .ZN(n20195) );
  OAI21_X1 U22342 ( .B1(n20197), .B2(n20626), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20198) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20629), .B1(
        n20086), .B2(n20628), .ZN(n20201) );
  OAI211_X1 U22344 ( .C1(n20244), .C2(n20632), .A(n20202), .B(n20201), .ZN(
        P2_U3095) );
  NAND2_X1 U22345 ( .A1(n20205), .A2(n20204), .ZN(n20208) );
  INV_X1 U22346 ( .A(n20208), .ZN(n20633) );
  AOI22_X1 U22347 ( .A1(n20265), .A2(n20634), .B1(n20263), .B2(n20633), .ZN(
        n20217) );
  NOR2_X1 U22348 ( .A1(n20641), .A2(n20634), .ZN(n20206) );
  OAI21_X1 U22349 ( .B1(n20206), .B2(n22410), .A(n20222), .ZN(n20215) );
  NOR2_X1 U22350 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20207), .ZN(
        n20212) );
  OAI211_X1 U22351 ( .C1(n20210), .C2(n20209), .A(n20208), .B(n20254), .ZN(
        n20211) );
  OAI211_X1 U22352 ( .C1(n20215), .C2(n20212), .A(n20257), .B(n20211), .ZN(
        n20636) );
  INV_X1 U22353 ( .A(n20212), .ZN(n20214) );
  OAI21_X1 U22354 ( .B1(n11228), .B2(n20633), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20213) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20636), .B1(
        n20086), .B2(n20635), .ZN(n20216) );
  OAI211_X1 U22356 ( .C1(n20244), .C2(n20639), .A(n20217), .B(n20216), .ZN(
        P2_U3087) );
  AND2_X1 U22357 ( .A1(n20219), .A2(n20246), .ZN(n20640) );
  AOI22_X1 U22358 ( .A1(n20264), .A2(n20649), .B1(n20640), .B2(n20263), .ZN(
        n20231) );
  OAI21_X1 U22359 ( .B1(n20221), .B2(n20220), .A(n20222), .ZN(n20229) );
  NAND2_X1 U22360 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20246), .ZN(
        n20228) );
  INV_X1 U22361 ( .A(n20228), .ZN(n20225) );
  AOI211_X1 U22362 ( .C1(n20226), .C2(n20253), .A(n20222), .B(n20640), .ZN(
        n20223) );
  NOR2_X1 U22363 ( .A1(n20558), .A2(n20223), .ZN(n20224) );
  OAI21_X1 U22364 ( .B1(n20229), .B2(n20225), .A(n20224), .ZN(n20643) );
  OAI21_X1 U22365 ( .B1(n20226), .B2(n20640), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20227) );
  OAI21_X1 U22366 ( .B1(n20229), .B2(n20228), .A(n20227), .ZN(n20642) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20643), .B1(
        n20086), .B2(n20642), .ZN(n20230) );
  OAI211_X1 U22368 ( .C1(n20262), .C2(n20639), .A(n20231), .B(n20230), .ZN(
        P2_U3079) );
  NAND3_X1 U22369 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20246), .A3(
        n20247), .ZN(n20238) );
  AND2_X1 U22370 ( .A1(n12586), .A2(n20238), .ZN(n20236) );
  INV_X1 U22371 ( .A(n20233), .ZN(n20234) );
  NAND2_X1 U22372 ( .A1(n20234), .A2(n20246), .ZN(n20237) );
  INV_X1 U22373 ( .A(n20238), .ZN(n20647) );
  AOI22_X1 U22374 ( .A1(n20648), .A2(n20086), .B1(n20263), .B2(n20647), .ZN(
        n20243) );
  OAI221_X1 U22375 ( .B1(n22410), .B2(n20646), .C1(n22410), .C2(n20659), .A(
        n20237), .ZN(n20240) );
  OAI21_X1 U22376 ( .B1(n12586), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20238), 
        .ZN(n20239) );
  MUX2_X1 U22377 ( .A(n20240), .B(n20239), .S(n20254), .Z(n20241) );
  NAND2_X1 U22378 ( .A1(n20241), .A2(n20257), .ZN(n20650) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20650), .B1(
        n20649), .B2(n20265), .ZN(n20242) );
  OAI211_X1 U22380 ( .C1(n20244), .C2(n20659), .A(n20243), .B(n20242), .ZN(
        P2_U3071) );
  NAND2_X1 U22381 ( .A1(n20246), .A2(n20245), .ZN(n20250) );
  NOR2_X1 U22382 ( .A1(n20247), .A2(n20250), .ZN(n20654) );
  OAI21_X1 U22383 ( .B1(n12573), .B2(n20654), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20248) );
  OAI21_X1 U22384 ( .B1(n20250), .B2(n20254), .A(n20248), .ZN(n20655) );
  AOI22_X1 U22385 ( .A1(n20655), .A2(n20086), .B1(n20263), .B2(n20654), .ZN(
        n20261) );
  INV_X1 U22386 ( .A(n20249), .ZN(n20252) );
  OAI21_X1 U22387 ( .B1(n20252), .B2(n20251), .A(n20250), .ZN(n20259) );
  NAND2_X1 U22388 ( .A1(n12573), .A2(n20253), .ZN(n20256) );
  INV_X1 U22389 ( .A(n20654), .ZN(n20255) );
  NAND3_X1 U22390 ( .A1(n20256), .A2(n20255), .A3(n20254), .ZN(n20258) );
  NAND3_X1 U22391 ( .A1(n20259), .A2(n20258), .A3(n20257), .ZN(n20656) );
  AOI22_X1 U22392 ( .A1(n20668), .A2(n20264), .B1(n20656), .B2(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20260) );
  OAI211_X1 U22393 ( .C1(n20262), .C2(n20659), .A(n20261), .B(n20260), .ZN(
        P2_U3063) );
  AOI22_X1 U22394 ( .A1(n20264), .A2(n20663), .B1(n20662), .B2(n20263), .ZN(
        n20267) );
  AOI22_X1 U22395 ( .A1(n20086), .A2(n20666), .B1(n20668), .B2(n20265), .ZN(
        n20266) );
  OAI211_X1 U22396 ( .C1(n20672), .C2(n20268), .A(n20267), .B(n20266), .ZN(
        P2_U3055) );
  AOI22_X1 U22397 ( .A1(P2_EAX_REG_6__SCAN_IN), .A2(n20495), .B1(n20269), .B2(
        n20313), .ZN(n20270) );
  OAI21_X1 U22398 ( .B1(n20271), .B2(n20557), .A(n20270), .ZN(P2_U2913) );
  NOR2_X2 U22399 ( .A1(n13801), .A2(n20454), .ZN(n20306) );
  AOI22_X1 U22400 ( .A1(n20562), .A2(n20272), .B1(n20561), .B2(n20306), .ZN(
        n20274) );
  AOI22_X1 U22401 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20563), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20564), .ZN(n20305) );
  AOI22_X1 U22402 ( .A1(n20308), .A2(n20663), .B1(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n20565), .ZN(n20273) );
  OAI211_X1 U22403 ( .C1(n20302), .C2(n20568), .A(n20274), .B(n20273), .ZN(
        P2_U3174) );
  AOI22_X1 U22404 ( .A1(n20308), .A2(n20570), .B1(n20306), .B2(n20569), .ZN(
        n20276) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20572), .B1(
        n20272), .B2(n20571), .ZN(n20275) );
  OAI211_X1 U22406 ( .C1(n20302), .C2(n20580), .A(n20276), .B(n20275), .ZN(
        P2_U3166) );
  AOI22_X1 U22407 ( .A1(n20576), .A2(n20272), .B1(n20306), .B2(n20575), .ZN(
        n20278) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20577), .B1(
        n20507), .B2(n20308), .ZN(n20277) );
  OAI211_X1 U22409 ( .C1(n20302), .C2(n20510), .A(n20278), .B(n20277), .ZN(
        P2_U3158) );
  AOI22_X1 U22410 ( .A1(n20582), .A2(n20272), .B1(n20306), .B2(n20581), .ZN(
        n20280) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20308), .ZN(n20279) );
  OAI211_X1 U22412 ( .C1(n20302), .C2(n20593), .A(n20280), .B(n20279), .ZN(
        P2_U3150) );
  AOI22_X1 U22413 ( .A1(n20588), .A2(n20272), .B1(n20306), .B2(n20587), .ZN(
        n20282) );
  INV_X1 U22414 ( .A(n20302), .ZN(n20307) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20307), .ZN(n20281) );
  OAI211_X1 U22416 ( .C1(n20305), .C2(n20593), .A(n20282), .B(n20281), .ZN(
        P2_U3142) );
  AOI22_X1 U22417 ( .A1(n20307), .A2(n20595), .B1(n20306), .B2(n20594), .ZN(
        n20284) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20597), .B1(
        n20272), .B2(n20596), .ZN(n20283) );
  OAI211_X1 U22419 ( .C1(n20305), .C2(n20600), .A(n20284), .B(n20283), .ZN(
        P2_U3134) );
  AOI22_X1 U22420 ( .A1(n20308), .A2(n20595), .B1(n20306), .B2(n20601), .ZN(
        n20286) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20603), .B1(
        n20272), .B2(n20602), .ZN(n20285) );
  OAI211_X1 U22422 ( .C1(n20302), .C2(n20519), .A(n20286), .B(n20285), .ZN(
        P2_U3126) );
  AOI22_X1 U22423 ( .A1(n20308), .A2(n20608), .B1(n20306), .B2(n20607), .ZN(
        n20288) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20610), .B1(
        n20609), .B2(n20272), .ZN(n20287) );
  OAI211_X1 U22425 ( .C1(n20302), .C2(n20619), .A(n20288), .B(n20287), .ZN(
        P2_U3118) );
  AOI22_X1 U22426 ( .A1(n20614), .A2(n20272), .B1(n20613), .B2(n20306), .ZN(
        n20291) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20616), .B1(
        n20289), .B2(n20308), .ZN(n20290) );
  OAI211_X1 U22428 ( .C1(n20302), .C2(n20625), .A(n20291), .B(n20290), .ZN(
        P2_U3110) );
  AOI22_X1 U22429 ( .A1(n20621), .A2(n20272), .B1(n20306), .B2(n20620), .ZN(
        n20293) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20622), .B1(
        n20627), .B2(n20307), .ZN(n20292) );
  OAI211_X1 U22431 ( .C1(n20305), .C2(n20625), .A(n20293), .B(n20292), .ZN(
        P2_U3102) );
  AOI22_X1 U22432 ( .A1(n20308), .A2(n20627), .B1(n20306), .B2(n20626), .ZN(
        n20295) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20629), .B1(
        n20272), .B2(n20628), .ZN(n20294) );
  OAI211_X1 U22434 ( .C1(n20302), .C2(n20632), .A(n20295), .B(n20294), .ZN(
        P2_U3094) );
  AOI22_X1 U22435 ( .A1(n20308), .A2(n20634), .B1(n20633), .B2(n20306), .ZN(
        n20297) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20636), .B1(
        n20272), .B2(n20635), .ZN(n20296) );
  OAI211_X1 U22437 ( .C1(n20302), .C2(n20639), .A(n20297), .B(n20296), .ZN(
        P2_U3086) );
  AOI22_X1 U22438 ( .A1(n20307), .A2(n20649), .B1(n20640), .B2(n20306), .ZN(
        n20299) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20643), .B1(
        n20272), .B2(n20642), .ZN(n20298) );
  OAI211_X1 U22440 ( .C1(n20305), .C2(n20639), .A(n20299), .B(n20298), .ZN(
        P2_U3078) );
  AOI22_X1 U22441 ( .A1(n20648), .A2(n20272), .B1(n20306), .B2(n20647), .ZN(
        n20301) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20650), .B1(
        n20649), .B2(n20308), .ZN(n20300) );
  OAI211_X1 U22443 ( .C1(n20302), .C2(n20659), .A(n20301), .B(n20300), .ZN(
        P2_U3070) );
  AOI22_X1 U22444 ( .A1(n20655), .A2(n20272), .B1(n20306), .B2(n20654), .ZN(
        n20304) );
  AOI22_X1 U22445 ( .A1(n20668), .A2(n20307), .B1(n20656), .B2(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n20303) );
  OAI211_X1 U22446 ( .C1(n20305), .C2(n20659), .A(n20304), .B(n20303), .ZN(
        P2_U3062) );
  AOI22_X1 U22447 ( .A1(n20307), .A2(n20663), .B1(n20662), .B2(n20306), .ZN(
        n20310) );
  AOI22_X1 U22448 ( .A1(n20668), .A2(n20308), .B1(n20666), .B2(n20272), .ZN(
        n20309) );
  OAI211_X1 U22449 ( .C1(n20672), .C2(n20311), .A(n20310), .B(n20309), .ZN(
        P2_U3054) );
  INV_X1 U22450 ( .A(n20312), .ZN(n20314) );
  AOI22_X1 U22451 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n20495), .B1(n20314), .B2(
        n20313), .ZN(n20319) );
  INV_X1 U22452 ( .A(n20315), .ZN(n20316) );
  NAND3_X1 U22453 ( .A1(n20317), .A2(n20316), .A3(n20551), .ZN(n20318) );
  OAI211_X1 U22454 ( .C1(n20320), .C2(n20557), .A(n20319), .B(n20318), .ZN(
        P2_U2914) );
  AOI22_X1 U22455 ( .A1(n20562), .A2(n20321), .B1(n20561), .B2(n20355), .ZN(
        n20324) );
  AOI22_X1 U22456 ( .A1(n20663), .A2(n20357), .B1(n20565), .B2(
        P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20323) );
  OAI211_X1 U22457 ( .C1(n20351), .C2(n20568), .A(n20324), .B(n20323), .ZN(
        P2_U3173) );
  AOI22_X1 U22458 ( .A1(n20570), .A2(n20357), .B1(n20355), .B2(n20569), .ZN(
        n20326) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20572), .B1(
        n20321), .B2(n20571), .ZN(n20325) );
  OAI211_X1 U22460 ( .C1(n20351), .C2(n20580), .A(n20326), .B(n20325), .ZN(
        P2_U3165) );
  AOI22_X1 U22461 ( .A1(n20576), .A2(n20321), .B1(n20355), .B2(n20575), .ZN(
        n20328) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20577), .B1(
        n20583), .B2(n20356), .ZN(n20327) );
  OAI211_X1 U22463 ( .C1(n20354), .C2(n20580), .A(n20328), .B(n20327), .ZN(
        P2_U3157) );
  AOI22_X1 U22464 ( .A1(n20582), .A2(n20321), .B1(n20355), .B2(n20581), .ZN(
        n20330) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20357), .ZN(n20329) );
  OAI211_X1 U22466 ( .C1(n20351), .C2(n20593), .A(n20330), .B(n20329), .ZN(
        P2_U3149) );
  AOI22_X1 U22467 ( .A1(n20588), .A2(n20321), .B1(n20355), .B2(n20587), .ZN(
        n20332) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20356), .ZN(n20331) );
  OAI211_X1 U22469 ( .C1(n20354), .C2(n20593), .A(n20332), .B(n20331), .ZN(
        P2_U3141) );
  AOI22_X1 U22470 ( .A1(n20356), .A2(n20595), .B1(n20355), .B2(n20594), .ZN(
        n20334) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20597), .B1(
        n20321), .B2(n20596), .ZN(n20333) );
  OAI211_X1 U22472 ( .C1(n20354), .C2(n20600), .A(n20334), .B(n20333), .ZN(
        P2_U3133) );
  AOI22_X1 U22473 ( .A1(n20356), .A2(n20608), .B1(n20355), .B2(n20601), .ZN(
        n20336) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20603), .B1(
        n20321), .B2(n20602), .ZN(n20335) );
  OAI211_X1 U22475 ( .C1(n20354), .C2(n20606), .A(n20336), .B(n20335), .ZN(
        P2_U3125) );
  AOI22_X1 U22476 ( .A1(n20608), .A2(n20357), .B1(n20355), .B2(n20607), .ZN(
        n20338) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20610), .B1(
        n20609), .B2(n20321), .ZN(n20337) );
  OAI211_X1 U22478 ( .C1(n20351), .C2(n20619), .A(n20338), .B(n20337), .ZN(
        P2_U3117) );
  AOI22_X1 U22479 ( .A1(n20614), .A2(n20321), .B1(n20613), .B2(n20355), .ZN(
        n20340) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20616), .B1(
        n20615), .B2(n20356), .ZN(n20339) );
  OAI211_X1 U22481 ( .C1(n20354), .C2(n20619), .A(n20340), .B(n20339), .ZN(
        P2_U3109) );
  AOI22_X1 U22482 ( .A1(n20621), .A2(n20321), .B1(n20355), .B2(n20620), .ZN(
        n20342) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20622), .B1(
        n20615), .B2(n20357), .ZN(n20341) );
  OAI211_X1 U22484 ( .C1(n20351), .C2(n20528), .A(n20342), .B(n20341), .ZN(
        P2_U3101) );
  AOI22_X1 U22485 ( .A1(n20357), .A2(n20627), .B1(n20355), .B2(n20626), .ZN(
        n20344) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20629), .B1(
        n20321), .B2(n20628), .ZN(n20343) );
  OAI211_X1 U22487 ( .C1(n20351), .C2(n20632), .A(n20344), .B(n20343), .ZN(
        P2_U3093) );
  AOI22_X1 U22488 ( .A1(n20357), .A2(n20634), .B1(n20633), .B2(n20355), .ZN(
        n20346) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20636), .B1(
        n20321), .B2(n20635), .ZN(n20345) );
  OAI211_X1 U22490 ( .C1(n20351), .C2(n20639), .A(n20346), .B(n20345), .ZN(
        P2_U3085) );
  AOI22_X1 U22491 ( .A1(n20356), .A2(n20649), .B1(n20640), .B2(n20355), .ZN(
        n20348) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20643), .B1(
        n20321), .B2(n20642), .ZN(n20347) );
  OAI211_X1 U22493 ( .C1(n20354), .C2(n20639), .A(n20348), .B(n20347), .ZN(
        P2_U3077) );
  AOI22_X1 U22494 ( .A1(n20648), .A2(n20321), .B1(n20355), .B2(n20647), .ZN(
        n20350) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20650), .B1(
        n20649), .B2(n20357), .ZN(n20349) );
  OAI211_X1 U22496 ( .C1(n20351), .C2(n20659), .A(n20350), .B(n20349), .ZN(
        P2_U3069) );
  AOI22_X1 U22497 ( .A1(n20655), .A2(n20321), .B1(n20355), .B2(n20654), .ZN(
        n20353) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20656), .B1(
        n20356), .B2(n20668), .ZN(n20352) );
  OAI211_X1 U22499 ( .C1(n20354), .C2(n20659), .A(n20353), .B(n20352), .ZN(
        P2_U3061) );
  AOI22_X1 U22500 ( .A1(n20356), .A2(n20663), .B1(n20662), .B2(n20355), .ZN(
        n20359) );
  AOI22_X1 U22501 ( .A1(n20668), .A2(n20357), .B1(n20666), .B2(n20321), .ZN(
        n20358) );
  OAI211_X1 U22502 ( .C1(n20672), .C2(n20360), .A(n20359), .B(n20358), .ZN(
        P2_U3053) );
  NOR2_X2 U22503 ( .A1(n12014), .A2(n20454), .ZN(n20395) );
  AOI22_X1 U22504 ( .A1(n20562), .A2(n20362), .B1(n20561), .B2(n20395), .ZN(
        n20364) );
  AOI22_X1 U22505 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20563), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20564), .ZN(n20391) );
  AOI22_X1 U22506 ( .A1(n20396), .A2(n20570), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n20565), .ZN(n20363) );
  OAI211_X1 U22507 ( .C1(n20394), .C2(n20412), .A(n20364), .B(n20363), .ZN(
        P2_U3172) );
  AOI22_X1 U22508 ( .A1(n20396), .A2(n20507), .B1(n20395), .B2(n20569), .ZN(
        n20366) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20572), .B1(
        n20362), .B2(n20571), .ZN(n20365) );
  OAI211_X1 U22510 ( .C1(n20394), .C2(n20568), .A(n20366), .B(n20365), .ZN(
        P2_U3164) );
  AOI22_X1 U22511 ( .A1(n20576), .A2(n20362), .B1(n20395), .B2(n20575), .ZN(
        n20368) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20577), .B1(
        n20583), .B2(n20396), .ZN(n20367) );
  OAI211_X1 U22513 ( .C1(n20394), .C2(n20580), .A(n20368), .B(n20367), .ZN(
        P2_U3156) );
  AOI22_X1 U22514 ( .A1(n20582), .A2(n20362), .B1(n20395), .B2(n20581), .ZN(
        n20370) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20397), .ZN(n20369) );
  OAI211_X1 U22516 ( .C1(n20391), .C2(n20593), .A(n20370), .B(n20369), .ZN(
        P2_U3148) );
  AOI22_X1 U22517 ( .A1(n20588), .A2(n20362), .B1(n20395), .B2(n20587), .ZN(
        n20372) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20396), .ZN(n20371) );
  OAI211_X1 U22519 ( .C1(n20394), .C2(n20593), .A(n20372), .B(n20371), .ZN(
        P2_U3140) );
  AOI22_X1 U22520 ( .A1(n20396), .A2(n20595), .B1(n20395), .B2(n20594), .ZN(
        n20374) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20597), .B1(
        n20362), .B2(n20596), .ZN(n20373) );
  OAI211_X1 U22522 ( .C1(n20394), .C2(n20600), .A(n20374), .B(n20373), .ZN(
        P2_U3132) );
  AOI22_X1 U22523 ( .A1(n20396), .A2(n20608), .B1(n20395), .B2(n20601), .ZN(
        n20376) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20603), .B1(
        n20362), .B2(n20602), .ZN(n20375) );
  OAI211_X1 U22525 ( .C1(n20394), .C2(n20606), .A(n20376), .B(n20375), .ZN(
        P2_U3124) );
  AOI22_X1 U22526 ( .A1(n20608), .A2(n20397), .B1(n20395), .B2(n20607), .ZN(
        n20378) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20610), .B1(
        n20609), .B2(n20362), .ZN(n20377) );
  OAI211_X1 U22528 ( .C1(n20391), .C2(n20619), .A(n20378), .B(n20377), .ZN(
        P2_U3116) );
  AOI22_X1 U22529 ( .A1(n20614), .A2(n20362), .B1(n20613), .B2(n20395), .ZN(
        n20380) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20616), .B1(
        n20615), .B2(n20396), .ZN(n20379) );
  OAI211_X1 U22531 ( .C1(n20394), .C2(n20619), .A(n20380), .B(n20379), .ZN(
        P2_U3108) );
  AOI22_X1 U22532 ( .A1(n20621), .A2(n20362), .B1(n20395), .B2(n20620), .ZN(
        n20382) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20622), .B1(
        n20627), .B2(n20396), .ZN(n20381) );
  OAI211_X1 U22534 ( .C1(n20394), .C2(n20625), .A(n20382), .B(n20381), .ZN(
        P2_U3100) );
  AOI22_X1 U22535 ( .A1(n20396), .A2(n20634), .B1(n20395), .B2(n20626), .ZN(
        n20384) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20629), .B1(
        n20362), .B2(n20628), .ZN(n20383) );
  OAI211_X1 U22537 ( .C1(n20394), .C2(n20528), .A(n20384), .B(n20383), .ZN(
        P2_U3092) );
  AOI22_X1 U22538 ( .A1(n20397), .A2(n20634), .B1(n20395), .B2(n20633), .ZN(
        n20386) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20636), .B1(
        n20362), .B2(n20635), .ZN(n20385) );
  OAI211_X1 U22540 ( .C1(n20391), .C2(n20639), .A(n20386), .B(n20385), .ZN(
        P2_U3084) );
  AOI22_X1 U22541 ( .A1(n20397), .A2(n20641), .B1(n20640), .B2(n20395), .ZN(
        n20388) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20643), .B1(
        n20362), .B2(n20642), .ZN(n20387) );
  OAI211_X1 U22543 ( .C1(n20391), .C2(n20646), .A(n20388), .B(n20387), .ZN(
        P2_U3076) );
  AOI22_X1 U22544 ( .A1(n20648), .A2(n20362), .B1(n20395), .B2(n20647), .ZN(
        n20390) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20650), .B1(
        n20649), .B2(n20397), .ZN(n20389) );
  OAI211_X1 U22546 ( .C1(n20391), .C2(n20659), .A(n20390), .B(n20389), .ZN(
        P2_U3068) );
  AOI22_X1 U22547 ( .A1(n20655), .A2(n20362), .B1(n20395), .B2(n20654), .ZN(
        n20393) );
  AOI22_X1 U22548 ( .A1(n20656), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n20396), .B2(n20668), .ZN(n20392) );
  OAI211_X1 U22549 ( .C1(n20394), .C2(n20659), .A(n20393), .B(n20392), .ZN(
        P2_U3060) );
  AOI22_X1 U22550 ( .A1(n20396), .A2(n20663), .B1(n20662), .B2(n20395), .ZN(
        n20399) );
  AOI22_X1 U22551 ( .A1(n20668), .A2(n20397), .B1(n20666), .B2(n20362), .ZN(
        n20398) );
  OAI211_X1 U22552 ( .C1(n20672), .C2(n20400), .A(n20399), .B(n20398), .ZN(
        P2_U3052) );
  AOI22_X1 U22553 ( .A1(n20497), .A2(n20401), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20495), .ZN(n20408) );
  AOI21_X1 U22554 ( .B1(n20404), .B2(n20403), .A(n20402), .ZN(n20406) );
  OR2_X1 U22555 ( .A1(n20406), .A2(n20405), .ZN(n20407) );
  OAI211_X1 U22556 ( .C1(n20409), .C2(n20557), .A(n20408), .B(n20407), .ZN(
        P2_U2916) );
  AOI22_X1 U22557 ( .A1(n20562), .A2(n15775), .B1(n20561), .B2(n20441), .ZN(
        n20411) );
  AOI22_X1 U22558 ( .A1(n20442), .A2(n20570), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n20565), .ZN(n20410) );
  OAI211_X1 U22559 ( .C1(n20445), .C2(n20412), .A(n20411), .B(n20410), .ZN(
        P2_U3171) );
  AOI22_X1 U22560 ( .A1(n20437), .A2(n20570), .B1(n20441), .B2(n20569), .ZN(
        n20414) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20572), .B1(
        n15775), .B2(n20571), .ZN(n20413) );
  OAI211_X1 U22562 ( .C1(n20440), .C2(n20580), .A(n20414), .B(n20413), .ZN(
        P2_U3163) );
  AOI22_X1 U22563 ( .A1(n20576), .A2(n15775), .B1(n20441), .B2(n20575), .ZN(
        n20416) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20577), .B1(
        n20583), .B2(n20442), .ZN(n20415) );
  OAI211_X1 U22565 ( .C1(n20445), .C2(n20580), .A(n20416), .B(n20415), .ZN(
        P2_U3155) );
  AOI22_X1 U22566 ( .A1(n20582), .A2(n15775), .B1(n20441), .B2(n20581), .ZN(
        n20418) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20437), .ZN(n20417) );
  OAI211_X1 U22568 ( .C1(n20440), .C2(n20593), .A(n20418), .B(n20417), .ZN(
        P2_U3147) );
  AOI22_X1 U22569 ( .A1(n20588), .A2(n15775), .B1(n20441), .B2(n20587), .ZN(
        n20420) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20442), .ZN(n20419) );
  OAI211_X1 U22571 ( .C1(n20445), .C2(n20593), .A(n20420), .B(n20419), .ZN(
        P2_U3139) );
  AOI22_X1 U22572 ( .A1(n20437), .A2(n20589), .B1(n20441), .B2(n20594), .ZN(
        n20422) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20597), .B1(
        n15775), .B2(n20596), .ZN(n20421) );
  OAI211_X1 U22574 ( .C1(n20440), .C2(n20606), .A(n20422), .B(n20421), .ZN(
        P2_U3131) );
  AOI22_X1 U22575 ( .A1(n20437), .A2(n20595), .B1(n20441), .B2(n20601), .ZN(
        n20424) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20603), .B1(
        n15775), .B2(n20602), .ZN(n20423) );
  OAI211_X1 U22577 ( .C1(n20440), .C2(n20519), .A(n20424), .B(n20423), .ZN(
        P2_U3123) );
  AOI22_X1 U22578 ( .A1(n20437), .A2(n20608), .B1(n20441), .B2(n20607), .ZN(
        n20426) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20610), .B1(
        n20609), .B2(n15775), .ZN(n20425) );
  OAI211_X1 U22580 ( .C1(n20440), .C2(n20619), .A(n20426), .B(n20425), .ZN(
        P2_U3115) );
  AOI22_X1 U22581 ( .A1(n20614), .A2(n15775), .B1(n20441), .B2(n20613), .ZN(
        n20428) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20616), .B1(
        n20615), .B2(n20442), .ZN(n20427) );
  OAI211_X1 U22583 ( .C1(n20445), .C2(n20619), .A(n20428), .B(n20427), .ZN(
        P2_U3107) );
  AOI22_X1 U22584 ( .A1(n20621), .A2(n15775), .B1(n20441), .B2(n20620), .ZN(
        n20430) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20622), .B1(
        n20615), .B2(n20437), .ZN(n20429) );
  OAI211_X1 U22586 ( .C1(n20440), .C2(n20528), .A(n20430), .B(n20429), .ZN(
        P2_U3099) );
  AOI22_X1 U22587 ( .A1(n20442), .A2(n20634), .B1(n20441), .B2(n20626), .ZN(
        n20432) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20629), .B1(
        n15775), .B2(n20628), .ZN(n20431) );
  OAI211_X1 U22589 ( .C1(n20445), .C2(n20528), .A(n20432), .B(n20431), .ZN(
        P2_U3091) );
  AOI22_X1 U22590 ( .A1(n20437), .A2(n20634), .B1(n20441), .B2(n20633), .ZN(
        n20434) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20636), .B1(
        n15775), .B2(n20635), .ZN(n20433) );
  OAI211_X1 U22592 ( .C1(n20440), .C2(n20639), .A(n20434), .B(n20433), .ZN(
        P2_U3083) );
  AOI22_X1 U22593 ( .A1(n20442), .A2(n20649), .B1(n20441), .B2(n20640), .ZN(
        n20436) );
  AOI22_X1 U22594 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20643), .B1(
        n15775), .B2(n20642), .ZN(n20435) );
  OAI211_X1 U22595 ( .C1(n20445), .C2(n20639), .A(n20436), .B(n20435), .ZN(
        P2_U3075) );
  AOI22_X1 U22596 ( .A1(n20648), .A2(n15775), .B1(n20441), .B2(n20647), .ZN(
        n20439) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20650), .B1(
        n20649), .B2(n20437), .ZN(n20438) );
  OAI211_X1 U22598 ( .C1(n20440), .C2(n20659), .A(n20439), .B(n20438), .ZN(
        P2_U3067) );
  AOI22_X1 U22599 ( .A1(n20655), .A2(n15775), .B1(n20441), .B2(n20654), .ZN(
        n20444) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20656), .B1(
        n20442), .B2(n20668), .ZN(n20443) );
  OAI211_X1 U22601 ( .C1(n20445), .C2(n20659), .A(n20444), .B(n20443), .ZN(
        P2_U3059) );
  AOI22_X1 U22602 ( .A1(n20497), .A2(n20446), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n20495), .ZN(n20451) );
  XNOR2_X1 U22603 ( .A(n20448), .B(n20447), .ZN(n20449) );
  NAND2_X1 U22604 ( .A1(n20449), .A2(n20551), .ZN(n20450) );
  OAI211_X1 U22605 ( .C1(n20452), .C2(n20557), .A(n20451), .B(n20450), .ZN(
        P2_U2917) );
  NOR2_X2 U22606 ( .A1(n12046), .A2(n20454), .ZN(n20489) );
  AOI22_X1 U22607 ( .A1(n20562), .A2(n20453), .B1(n20561), .B2(n20489), .ZN(
        n20458) );
  AOI22_X1 U22608 ( .A1(n20663), .A2(n20491), .B1(n20565), .B2(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20457) );
  OAI211_X1 U22609 ( .C1(n20485), .C2(n20568), .A(n20458), .B(n20457), .ZN(
        P2_U3170) );
  INV_X1 U22610 ( .A(n20491), .ZN(n20488) );
  AOI22_X1 U22611 ( .A1(n20490), .A2(n20507), .B1(n20489), .B2(n20569), .ZN(
        n20460) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20572), .B1(
        n20453), .B2(n20571), .ZN(n20459) );
  OAI211_X1 U22613 ( .C1(n20488), .C2(n20568), .A(n20460), .B(n20459), .ZN(
        P2_U3162) );
  AOI22_X1 U22614 ( .A1(n20576), .A2(n20453), .B1(n20489), .B2(n20575), .ZN(
        n20462) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20577), .B1(
        n20507), .B2(n20491), .ZN(n20461) );
  OAI211_X1 U22616 ( .C1(n20485), .C2(n20510), .A(n20462), .B(n20461), .ZN(
        P2_U3154) );
  AOI22_X1 U22617 ( .A1(n20582), .A2(n20453), .B1(n20489), .B2(n20581), .ZN(
        n20464) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20491), .ZN(n20463) );
  OAI211_X1 U22619 ( .C1(n20485), .C2(n20593), .A(n20464), .B(n20463), .ZN(
        P2_U3146) );
  AOI22_X1 U22620 ( .A1(n20588), .A2(n20453), .B1(n20489), .B2(n20587), .ZN(
        n20466) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20490), .ZN(n20465) );
  OAI211_X1 U22622 ( .C1(n20488), .C2(n20593), .A(n20466), .B(n20465), .ZN(
        P2_U3138) );
  AOI22_X1 U22623 ( .A1(n20490), .A2(n20595), .B1(n20489), .B2(n20594), .ZN(
        n20468) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20597), .B1(
        n20453), .B2(n20596), .ZN(n20467) );
  OAI211_X1 U22625 ( .C1(n20488), .C2(n20600), .A(n20468), .B(n20467), .ZN(
        P2_U3130) );
  AOI22_X1 U22626 ( .A1(n20490), .A2(n20608), .B1(n20489), .B2(n20601), .ZN(
        n20470) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20603), .B1(
        n20453), .B2(n20602), .ZN(n20469) );
  OAI211_X1 U22628 ( .C1(n20488), .C2(n20606), .A(n20470), .B(n20469), .ZN(
        P2_U3122) );
  AOI22_X1 U22629 ( .A1(n20608), .A2(n20491), .B1(n20489), .B2(n20607), .ZN(
        n20472) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20610), .B1(
        n20609), .B2(n20453), .ZN(n20471) );
  OAI211_X1 U22631 ( .C1(n20485), .C2(n20619), .A(n20472), .B(n20471), .ZN(
        P2_U3114) );
  AOI22_X1 U22632 ( .A1(n20614), .A2(n20453), .B1(n20613), .B2(n20489), .ZN(
        n20474) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20616), .B1(
        n20615), .B2(n20490), .ZN(n20473) );
  OAI211_X1 U22634 ( .C1(n20488), .C2(n20619), .A(n20474), .B(n20473), .ZN(
        P2_U3106) );
  AOI22_X1 U22635 ( .A1(n20621), .A2(n20453), .B1(n20489), .B2(n20620), .ZN(
        n20476) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20622), .B1(
        n20627), .B2(n20490), .ZN(n20475) );
  OAI211_X1 U22637 ( .C1(n20488), .C2(n20625), .A(n20476), .B(n20475), .ZN(
        P2_U3098) );
  AOI22_X1 U22638 ( .A1(n20491), .A2(n20627), .B1(n20489), .B2(n20626), .ZN(
        n20478) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20629), .B1(
        n20453), .B2(n20628), .ZN(n20477) );
  OAI211_X1 U22640 ( .C1(n20485), .C2(n20632), .A(n20478), .B(n20477), .ZN(
        P2_U3090) );
  AOI22_X1 U22641 ( .A1(n20491), .A2(n20634), .B1(n20489), .B2(n20633), .ZN(
        n20480) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20636), .B1(
        n20453), .B2(n20635), .ZN(n20479) );
  OAI211_X1 U22643 ( .C1(n20485), .C2(n20639), .A(n20480), .B(n20479), .ZN(
        P2_U3082) );
  AOI22_X1 U22644 ( .A1(n20491), .A2(n20641), .B1(n20640), .B2(n20489), .ZN(
        n20482) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20643), .B1(
        n20453), .B2(n20642), .ZN(n20481) );
  OAI211_X1 U22646 ( .C1(n20485), .C2(n20646), .A(n20482), .B(n20481), .ZN(
        P2_U3074) );
  AOI22_X1 U22647 ( .A1(n20648), .A2(n20453), .B1(n20489), .B2(n20647), .ZN(
        n20484) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20650), .B1(
        n20649), .B2(n20491), .ZN(n20483) );
  OAI211_X1 U22649 ( .C1(n20485), .C2(n20659), .A(n20484), .B(n20483), .ZN(
        P2_U3066) );
  AOI22_X1 U22650 ( .A1(n20655), .A2(n20453), .B1(n20489), .B2(n20654), .ZN(
        n20487) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20656), .B1(
        n20490), .B2(n20668), .ZN(n20486) );
  OAI211_X1 U22652 ( .C1(n20488), .C2(n20659), .A(n20487), .B(n20486), .ZN(
        P2_U3058) );
  AOI22_X1 U22653 ( .A1(n20490), .A2(n20663), .B1(n20662), .B2(n20489), .ZN(
        n20493) );
  AOI22_X1 U22654 ( .A1(n20668), .A2(n20491), .B1(n20666), .B2(n20453), .ZN(
        n20492) );
  OAI211_X1 U22655 ( .C1(n20672), .C2(n20494), .A(n20493), .B(n20492), .ZN(
        P2_U3050) );
  AOI22_X1 U22656 ( .A1(n20497), .A2(n20496), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n20495), .ZN(n20501) );
  XOR2_X1 U22657 ( .A(n20550), .B(n20498), .Z(n20499) );
  NAND2_X1 U22658 ( .A1(n20499), .A2(n20551), .ZN(n20500) );
  OAI211_X1 U22659 ( .C1(n20502), .C2(n20557), .A(n20501), .B(n20500), .ZN(
        P2_U2918) );
  NOR2_X2 U22660 ( .A1(n20502), .A2(n20558), .ZN(n20541) );
  AOI22_X1 U22661 ( .A1(n20562), .A2(n20541), .B1(n20561), .B2(n20539), .ZN(
        n20504) );
  AOI22_X1 U22662 ( .A1(n20542), .A2(n20663), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n20565), .ZN(n20503) );
  OAI211_X1 U22663 ( .C1(n20535), .C2(n20568), .A(n20504), .B(n20503), .ZN(
        P2_U3169) );
  AOI22_X1 U22664 ( .A1(n20540), .A2(n20507), .B1(n20539), .B2(n20569), .ZN(
        n20506) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20572), .B1(
        n20541), .B2(n20571), .ZN(n20505) );
  OAI211_X1 U22666 ( .C1(n20538), .C2(n20568), .A(n20506), .B(n20505), .ZN(
        P2_U3161) );
  AOI22_X1 U22667 ( .A1(n20576), .A2(n20541), .B1(n20539), .B2(n20575), .ZN(
        n20509) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20577), .B1(
        n20507), .B2(n20542), .ZN(n20508) );
  OAI211_X1 U22669 ( .C1(n20535), .C2(n20510), .A(n20509), .B(n20508), .ZN(
        P2_U3153) );
  AOI22_X1 U22670 ( .A1(n20582), .A2(n20541), .B1(n20539), .B2(n20581), .ZN(
        n20512) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20542), .ZN(n20511) );
  OAI211_X1 U22672 ( .C1(n20535), .C2(n20593), .A(n20512), .B(n20511), .ZN(
        P2_U3145) );
  AOI22_X1 U22673 ( .A1(n20588), .A2(n20541), .B1(n20539), .B2(n20587), .ZN(
        n20514) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20540), .ZN(n20513) );
  OAI211_X1 U22675 ( .C1(n20538), .C2(n20593), .A(n20514), .B(n20513), .ZN(
        P2_U3137) );
  AOI22_X1 U22676 ( .A1(n20540), .A2(n20595), .B1(n20539), .B2(n20594), .ZN(
        n20516) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20597), .B1(
        n20541), .B2(n20596), .ZN(n20515) );
  OAI211_X1 U22678 ( .C1(n20538), .C2(n20600), .A(n20516), .B(n20515), .ZN(
        P2_U3129) );
  AOI22_X1 U22679 ( .A1(n20542), .A2(n20595), .B1(n20539), .B2(n20601), .ZN(
        n20518) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20603), .B1(
        n20541), .B2(n20602), .ZN(n20517) );
  OAI211_X1 U22681 ( .C1(n20535), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        P2_U3121) );
  AOI22_X1 U22682 ( .A1(n20542), .A2(n20608), .B1(n20539), .B2(n20607), .ZN(
        n20521) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20610), .B1(
        n20609), .B2(n20541), .ZN(n20520) );
  OAI211_X1 U22684 ( .C1(n20535), .C2(n20619), .A(n20521), .B(n20520), .ZN(
        P2_U3113) );
  AOI22_X1 U22685 ( .A1(n20614), .A2(n20541), .B1(n20613), .B2(n20539), .ZN(
        n20523) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20616), .B1(
        n20615), .B2(n20540), .ZN(n20522) );
  OAI211_X1 U22687 ( .C1(n20538), .C2(n20619), .A(n20523), .B(n20522), .ZN(
        P2_U3105) );
  AOI22_X1 U22688 ( .A1(n20621), .A2(n20541), .B1(n20539), .B2(n20620), .ZN(
        n20525) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20622), .B1(
        n20627), .B2(n20540), .ZN(n20524) );
  OAI211_X1 U22690 ( .C1(n20538), .C2(n20625), .A(n20525), .B(n20524), .ZN(
        P2_U3097) );
  AOI22_X1 U22691 ( .A1(n20540), .A2(n20634), .B1(n20539), .B2(n20626), .ZN(
        n20527) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20629), .B1(
        n20541), .B2(n20628), .ZN(n20526) );
  OAI211_X1 U22693 ( .C1(n20538), .C2(n20528), .A(n20527), .B(n20526), .ZN(
        P2_U3089) );
  AOI22_X1 U22694 ( .A1(n20542), .A2(n20634), .B1(n20539), .B2(n20633), .ZN(
        n20530) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20636), .B1(
        n20541), .B2(n20635), .ZN(n20529) );
  OAI211_X1 U22696 ( .C1(n20535), .C2(n20639), .A(n20530), .B(n20529), .ZN(
        P2_U3081) );
  AOI22_X1 U22697 ( .A1(n20542), .A2(n20641), .B1(n20640), .B2(n20539), .ZN(
        n20532) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20643), .B1(
        n20541), .B2(n20642), .ZN(n20531) );
  OAI211_X1 U22699 ( .C1(n20535), .C2(n20646), .A(n20532), .B(n20531), .ZN(
        P2_U3073) );
  AOI22_X1 U22700 ( .A1(n20648), .A2(n20541), .B1(n20539), .B2(n20647), .ZN(
        n20534) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20650), .B1(
        n20649), .B2(n20542), .ZN(n20533) );
  OAI211_X1 U22702 ( .C1(n20535), .C2(n20659), .A(n20534), .B(n20533), .ZN(
        P2_U3065) );
  AOI22_X1 U22703 ( .A1(n20655), .A2(n20541), .B1(n20539), .B2(n20654), .ZN(
        n20537) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20656), .B1(
        n20540), .B2(n20668), .ZN(n20536) );
  OAI211_X1 U22705 ( .C1(n20538), .C2(n20659), .A(n20537), .B(n20536), .ZN(
        P2_U3057) );
  AOI22_X1 U22706 ( .A1(n20540), .A2(n20663), .B1(n20662), .B2(n20539), .ZN(
        n20544) );
  AOI22_X1 U22707 ( .A1(n20668), .A2(n20542), .B1(n20666), .B2(n20541), .ZN(
        n20543) );
  OAI211_X1 U22708 ( .C1(n20672), .C2(n20545), .A(n20544), .B(n20543), .ZN(
        P2_U3049) );
  OAI22_X1 U22709 ( .A1(n20548), .A2(n20547), .B1(n20546), .B2(n18129), .ZN(
        n20549) );
  INV_X1 U22710 ( .A(n20549), .ZN(n20556) );
  INV_X1 U22711 ( .A(n20550), .ZN(n20552) );
  OAI211_X1 U22712 ( .C1(n20554), .C2(n20553), .A(n20552), .B(n20551), .ZN(
        n20555) );
  OAI211_X1 U22713 ( .C1(n20559), .C2(n20557), .A(n20556), .B(n20555), .ZN(
        P2_U2919) );
  NOR2_X2 U22714 ( .A1(n20559), .A2(n20558), .ZN(n20665) );
  AND2_X1 U22715 ( .A1(n12045), .A2(n20560), .ZN(n20661) );
  AOI22_X1 U22716 ( .A1(n20562), .A2(n20665), .B1(n20561), .B2(n20661), .ZN(
        n20567) );
  AOI22_X1 U22717 ( .A1(n20667), .A2(n20663), .B1(
        P2_INSTQUEUE_REG_15__0__SCAN_IN), .B2(n20565), .ZN(n20566) );
  OAI211_X1 U22718 ( .C1(n20653), .C2(n20568), .A(n20567), .B(n20566), .ZN(
        P2_U3168) );
  AOI22_X1 U22719 ( .A1(n20667), .A2(n20570), .B1(n20661), .B2(n20569), .ZN(
        n20574) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20572), .B1(
        n20665), .B2(n20571), .ZN(n20573) );
  OAI211_X1 U22721 ( .C1(n20653), .C2(n20580), .A(n20574), .B(n20573), .ZN(
        P2_U3160) );
  AOI22_X1 U22722 ( .A1(n20576), .A2(n20665), .B1(n20661), .B2(n20575), .ZN(
        n20579) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20577), .B1(
        n20583), .B2(n20664), .ZN(n20578) );
  OAI211_X1 U22724 ( .C1(n20660), .C2(n20580), .A(n20579), .B(n20578), .ZN(
        P2_U3152) );
  AOI22_X1 U22725 ( .A1(n20582), .A2(n20665), .B1(n20661), .B2(n20581), .ZN(
        n20586) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20584), .B1(
        n20583), .B2(n20667), .ZN(n20585) );
  OAI211_X1 U22727 ( .C1(n20653), .C2(n20593), .A(n20586), .B(n20585), .ZN(
        P2_U3144) );
  AOI22_X1 U22728 ( .A1(n20588), .A2(n20665), .B1(n20661), .B2(n20587), .ZN(
        n20592) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20664), .ZN(n20591) );
  OAI211_X1 U22730 ( .C1(n20660), .C2(n20593), .A(n20592), .B(n20591), .ZN(
        P2_U3136) );
  AOI22_X1 U22731 ( .A1(n20664), .A2(n20595), .B1(n20661), .B2(n20594), .ZN(
        n20599) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20597), .B1(
        n20665), .B2(n20596), .ZN(n20598) );
  OAI211_X1 U22733 ( .C1(n20660), .C2(n20600), .A(n20599), .B(n20598), .ZN(
        P2_U3128) );
  AOI22_X1 U22734 ( .A1(n20664), .A2(n20608), .B1(n20661), .B2(n20601), .ZN(
        n20605) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20603), .B1(
        n20665), .B2(n20602), .ZN(n20604) );
  OAI211_X1 U22736 ( .C1(n20660), .C2(n20606), .A(n20605), .B(n20604), .ZN(
        P2_U3120) );
  AOI22_X1 U22737 ( .A1(n20667), .A2(n20608), .B1(n20661), .B2(n20607), .ZN(
        n20612) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20610), .B1(
        n20609), .B2(n20665), .ZN(n20611) );
  OAI211_X1 U22739 ( .C1(n20653), .C2(n20619), .A(n20612), .B(n20611), .ZN(
        P2_U3112) );
  AOI22_X1 U22740 ( .A1(n20614), .A2(n20665), .B1(n20613), .B2(n20661), .ZN(
        n20618) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20616), .B1(
        n20615), .B2(n20664), .ZN(n20617) );
  OAI211_X1 U22742 ( .C1(n20660), .C2(n20619), .A(n20618), .B(n20617), .ZN(
        P2_U3104) );
  AOI22_X1 U22743 ( .A1(n20621), .A2(n20665), .B1(n20661), .B2(n20620), .ZN(
        n20624) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20622), .B1(
        n20627), .B2(n20664), .ZN(n20623) );
  OAI211_X1 U22745 ( .C1(n20660), .C2(n20625), .A(n20624), .B(n20623), .ZN(
        P2_U3096) );
  AOI22_X1 U22746 ( .A1(n20667), .A2(n20627), .B1(n20661), .B2(n20626), .ZN(
        n20631) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20629), .B1(
        n20665), .B2(n20628), .ZN(n20630) );
  OAI211_X1 U22748 ( .C1(n20653), .C2(n20632), .A(n20631), .B(n20630), .ZN(
        P2_U3088) );
  AOI22_X1 U22749 ( .A1(n20667), .A2(n20634), .B1(n20661), .B2(n20633), .ZN(
        n20638) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20636), .B1(
        n20665), .B2(n20635), .ZN(n20637) );
  OAI211_X1 U22751 ( .C1(n20653), .C2(n20639), .A(n20638), .B(n20637), .ZN(
        P2_U3080) );
  AOI22_X1 U22752 ( .A1(n20667), .A2(n20641), .B1(n20640), .B2(n20661), .ZN(
        n20645) );
  AOI22_X1 U22753 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20643), .B1(
        n20665), .B2(n20642), .ZN(n20644) );
  OAI211_X1 U22754 ( .C1(n20653), .C2(n20646), .A(n20645), .B(n20644), .ZN(
        P2_U3072) );
  AOI22_X1 U22755 ( .A1(n20648), .A2(n20665), .B1(n20661), .B2(n20647), .ZN(
        n20652) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20650), .B1(
        n20649), .B2(n20667), .ZN(n20651) );
  OAI211_X1 U22757 ( .C1(n20653), .C2(n20659), .A(n20652), .B(n20651), .ZN(
        P2_U3064) );
  AOI22_X1 U22758 ( .A1(n20655), .A2(n20665), .B1(n20661), .B2(n20654), .ZN(
        n20658) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20656), .B1(
        n20664), .B2(n20668), .ZN(n20657) );
  OAI211_X1 U22760 ( .C1(n20660), .C2(n20659), .A(n20658), .B(n20657), .ZN(
        P2_U3056) );
  AOI22_X1 U22761 ( .A1(n20664), .A2(n20663), .B1(n20662), .B2(n20661), .ZN(
        n20670) );
  AOI22_X1 U22762 ( .A1(n20668), .A2(n20667), .B1(n20666), .B2(n20665), .ZN(
        n20669) );
  OAI211_X1 U22763 ( .C1(n20672), .C2(n20671), .A(n20670), .B(n20669), .ZN(
        P2_U3048) );
  INV_X1 U22764 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20952) );
  INV_X1 U22765 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20673) );
  AOI222_X1 U22766 ( .A1(n20950), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n20952), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n20673), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20674) );
  INV_X1 U22767 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20676) );
  AOI22_X1 U22768 ( .A1(n20699), .A2(n20676), .B1(n20675), .B2(n20700), .ZN(
        U376) );
  OAI22_X1 U22769 ( .A1(n20700), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n20699), .ZN(n20677) );
  INV_X1 U22770 ( .A(n20677), .ZN(U365) );
  OAI22_X1 U22771 ( .A1(n20700), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n20699), .ZN(n20678) );
  INV_X1 U22772 ( .A(n20678), .ZN(U354) );
  OAI22_X1 U22773 ( .A1(n20700), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n20699), .ZN(n20679) );
  INV_X1 U22774 ( .A(n20679), .ZN(U353) );
  OAI22_X1 U22775 ( .A1(n20700), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n20699), .ZN(n20680) );
  INV_X1 U22776 ( .A(n20680), .ZN(U352) );
  OAI22_X1 U22777 ( .A1(n20700), .A2(P3_ADDRESS_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n20699), .ZN(n20681) );
  INV_X1 U22778 ( .A(n20681), .ZN(U351) );
  OAI22_X1 U22779 ( .A1(n20700), .A2(P3_ADDRESS_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n20699), .ZN(n20682) );
  INV_X1 U22780 ( .A(n20682), .ZN(U350) );
  OAI22_X1 U22781 ( .A1(n20700), .A2(P3_ADDRESS_REG_7__SCAN_IN), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(n20699), .ZN(n20683) );
  INV_X1 U22782 ( .A(n20683), .ZN(U349) );
  OAI22_X1 U22783 ( .A1(n20700), .A2(P3_ADDRESS_REG_8__SCAN_IN), .B1(
        P2_ADDRESS_REG_8__SCAN_IN), .B2(n20699), .ZN(n20684) );
  INV_X1 U22784 ( .A(n20684), .ZN(U348) );
  OAI22_X1 U22785 ( .A1(n20700), .A2(P3_ADDRESS_REG_9__SCAN_IN), .B1(
        P2_ADDRESS_REG_9__SCAN_IN), .B2(n20699), .ZN(n20685) );
  INV_X1 U22786 ( .A(n20685), .ZN(U347) );
  OAI22_X1 U22787 ( .A1(n20700), .A2(P3_ADDRESS_REG_10__SCAN_IN), .B1(
        P2_ADDRESS_REG_10__SCAN_IN), .B2(n20699), .ZN(n20686) );
  INV_X1 U22788 ( .A(n20686), .ZN(U375) );
  OAI22_X1 U22789 ( .A1(n20700), .A2(P3_ADDRESS_REG_11__SCAN_IN), .B1(
        P2_ADDRESS_REG_11__SCAN_IN), .B2(n20699), .ZN(n20687) );
  INV_X1 U22790 ( .A(n20687), .ZN(U374) );
  INV_X1 U22791 ( .A(n20700), .ZN(n20707) );
  OAI22_X1 U22792 ( .A1(n20700), .A2(P3_ADDRESS_REG_12__SCAN_IN), .B1(
        P2_ADDRESS_REG_12__SCAN_IN), .B2(n20707), .ZN(n20688) );
  INV_X1 U22793 ( .A(n20688), .ZN(U373) );
  OAI22_X1 U22794 ( .A1(n20700), .A2(P3_ADDRESS_REG_13__SCAN_IN), .B1(
        P2_ADDRESS_REG_13__SCAN_IN), .B2(n20699), .ZN(n20689) );
  INV_X1 U22795 ( .A(n20689), .ZN(U372) );
  OAI22_X1 U22796 ( .A1(n20700), .A2(P3_ADDRESS_REG_14__SCAN_IN), .B1(
        P2_ADDRESS_REG_14__SCAN_IN), .B2(n20699), .ZN(n20690) );
  INV_X1 U22797 ( .A(n20690), .ZN(U371) );
  OAI22_X1 U22798 ( .A1(n20700), .A2(P3_ADDRESS_REG_15__SCAN_IN), .B1(
        P2_ADDRESS_REG_15__SCAN_IN), .B2(n20699), .ZN(n20691) );
  INV_X1 U22799 ( .A(n20691), .ZN(U370) );
  OAI22_X1 U22800 ( .A1(n20700), .A2(P3_ADDRESS_REG_16__SCAN_IN), .B1(
        P2_ADDRESS_REG_16__SCAN_IN), .B2(n20707), .ZN(n20692) );
  INV_X1 U22801 ( .A(n20692), .ZN(U369) );
  OAI22_X1 U22802 ( .A1(n20700), .A2(P3_ADDRESS_REG_17__SCAN_IN), .B1(
        P2_ADDRESS_REG_17__SCAN_IN), .B2(n20699), .ZN(n20693) );
  INV_X1 U22803 ( .A(n20693), .ZN(U368) );
  OAI22_X1 U22804 ( .A1(n20700), .A2(P3_ADDRESS_REG_18__SCAN_IN), .B1(
        P2_ADDRESS_REG_18__SCAN_IN), .B2(n20699), .ZN(n20694) );
  INV_X1 U22805 ( .A(n20694), .ZN(U367) );
  OAI22_X1 U22806 ( .A1(n20700), .A2(P3_ADDRESS_REG_19__SCAN_IN), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(n20699), .ZN(n20695) );
  INV_X1 U22807 ( .A(n20695), .ZN(U366) );
  OAI22_X1 U22808 ( .A1(n20700), .A2(P3_ADDRESS_REG_20__SCAN_IN), .B1(
        P2_ADDRESS_REG_20__SCAN_IN), .B2(n20699), .ZN(n20696) );
  INV_X1 U22809 ( .A(n20696), .ZN(U364) );
  OAI22_X1 U22810 ( .A1(n20700), .A2(P3_ADDRESS_REG_21__SCAN_IN), .B1(
        P2_ADDRESS_REG_21__SCAN_IN), .B2(n20699), .ZN(n20697) );
  INV_X1 U22811 ( .A(n20697), .ZN(U363) );
  OAI22_X1 U22812 ( .A1(n20700), .A2(P3_ADDRESS_REG_22__SCAN_IN), .B1(
        P2_ADDRESS_REG_22__SCAN_IN), .B2(n20699), .ZN(n20698) );
  INV_X1 U22813 ( .A(n20698), .ZN(U362) );
  OAI22_X1 U22814 ( .A1(n20700), .A2(P3_ADDRESS_REG_23__SCAN_IN), .B1(
        P2_ADDRESS_REG_23__SCAN_IN), .B2(n20699), .ZN(n20701) );
  INV_X1 U22815 ( .A(n20701), .ZN(U361) );
  OAI22_X1 U22816 ( .A1(n20700), .A2(P3_ADDRESS_REG_24__SCAN_IN), .B1(
        P2_ADDRESS_REG_24__SCAN_IN), .B2(n20707), .ZN(n20702) );
  INV_X1 U22817 ( .A(n20702), .ZN(U360) );
  OAI22_X1 U22818 ( .A1(n20700), .A2(P3_ADDRESS_REG_25__SCAN_IN), .B1(
        P2_ADDRESS_REG_25__SCAN_IN), .B2(n20707), .ZN(n20703) );
  INV_X1 U22819 ( .A(n20703), .ZN(U359) );
  OAI22_X1 U22820 ( .A1(n20700), .A2(P3_ADDRESS_REG_26__SCAN_IN), .B1(
        P2_ADDRESS_REG_26__SCAN_IN), .B2(n20707), .ZN(n20704) );
  INV_X1 U22821 ( .A(n20704), .ZN(U358) );
  OAI22_X1 U22822 ( .A1(n20700), .A2(P3_ADDRESS_REG_27__SCAN_IN), .B1(
        P2_ADDRESS_REG_27__SCAN_IN), .B2(n20707), .ZN(n20705) );
  INV_X1 U22823 ( .A(n20705), .ZN(U357) );
  OAI22_X1 U22824 ( .A1(n20700), .A2(P3_ADDRESS_REG_28__SCAN_IN), .B1(
        P2_ADDRESS_REG_28__SCAN_IN), .B2(n20707), .ZN(n20706) );
  INV_X1 U22825 ( .A(n20706), .ZN(U356) );
  OAI22_X1 U22826 ( .A1(n20700), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n20707), .ZN(n20708) );
  INV_X1 U22827 ( .A(n20708), .ZN(U355) );
  AOI22_X1 U22828 ( .A1(n22106), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20710) );
  OAI21_X1 U22829 ( .B1(n20711), .B2(n20736), .A(n20710), .ZN(P1_U2936) );
  AOI22_X1 U22830 ( .A1(n20725), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20712) );
  OAI21_X1 U22831 ( .B1(n20713), .B2(n20736), .A(n20712), .ZN(P1_U2935) );
  AOI22_X1 U22832 ( .A1(n20725), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20714) );
  OAI21_X1 U22833 ( .B1(n20715), .B2(n20736), .A(n20714), .ZN(P1_U2934) );
  AOI22_X1 U22834 ( .A1(n20725), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20716) );
  OAI21_X1 U22835 ( .B1(n20717), .B2(n20736), .A(n20716), .ZN(P1_U2933) );
  AOI22_X1 U22836 ( .A1(n20725), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20718) );
  OAI21_X1 U22837 ( .B1(n20719), .B2(n20736), .A(n20718), .ZN(P1_U2932) );
  AOI22_X1 U22838 ( .A1(n20725), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20720) );
  OAI21_X1 U22839 ( .B1(n20721), .B2(n20736), .A(n20720), .ZN(P1_U2931) );
  AOI22_X1 U22840 ( .A1(n20725), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20722), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20723) );
  OAI21_X1 U22841 ( .B1(n13348), .B2(n20736), .A(n20723), .ZN(P1_U2930) );
  AOI22_X1 U22842 ( .A1(n22106), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20724) );
  OAI21_X1 U22843 ( .B1(n13357), .B2(n20736), .A(n20724), .ZN(P1_U2929) );
  AOI22_X1 U22844 ( .A1(n20725), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20726) );
  OAI21_X1 U22845 ( .B1(n15796), .B2(n20736), .A(n20726), .ZN(P1_U2928) );
  AOI22_X1 U22846 ( .A1(n22106), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20727) );
  OAI21_X1 U22847 ( .B1(n15694), .B2(n20736), .A(n20727), .ZN(P1_U2927) );
  AOI22_X1 U22848 ( .A1(n22106), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20728) );
  OAI21_X1 U22849 ( .B1(n15900), .B2(n20736), .A(n20728), .ZN(P1_U2926) );
  INV_X1 U22850 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20730) );
  AOI22_X1 U22851 ( .A1(n22106), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20729) );
  OAI21_X1 U22852 ( .B1(n20730), .B2(n20736), .A(n20729), .ZN(P1_U2925) );
  AOI22_X1 U22853 ( .A1(n22106), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20731) );
  OAI21_X1 U22854 ( .B1(n16835), .B2(n20736), .A(n20731), .ZN(P1_U2924) );
  AOI22_X1 U22855 ( .A1(n22106), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20732) );
  OAI21_X1 U22856 ( .B1(n16830), .B2(n20736), .A(n20732), .ZN(P1_U2923) );
  AOI22_X1 U22857 ( .A1(n22106), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20733) );
  OAI21_X1 U22858 ( .B1(n15954), .B2(n20736), .A(n20733), .ZN(P1_U2922) );
  AOI22_X1 U22859 ( .A1(n22106), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20734), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20735) );
  OAI21_X1 U22860 ( .B1(n20737), .B2(n20736), .A(n20735), .ZN(P1_U2921) );
  NAND2_X1 U22861 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22855), .ZN(n20794) );
  OAI222_X1 U22862 ( .A1(n20780), .A2(n22246), .B1(n20738), .B2(n22855), .C1(
        n22247), .C2(n22430), .ZN(P1_U3197) );
  INV_X1 U22863 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20739) );
  INV_X1 U22864 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20741) );
  OAI222_X1 U22865 ( .A1(n20794), .A2(n22246), .B1(n20739), .B2(n22855), .C1(
        n20741), .C2(n20780), .ZN(P1_U3198) );
  INV_X1 U22866 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20740) );
  OAI222_X1 U22867 ( .A1(n20794), .A2(n20741), .B1(n20740), .B2(n22855), .C1(
        n20743), .C2(n20780), .ZN(P1_U3199) );
  INV_X1 U22868 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20742) );
  INV_X1 U22869 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20745) );
  OAI222_X1 U22870 ( .A1(n22430), .A2(n20743), .B1(n20742), .B2(n22855), .C1(
        n20745), .C2(n20780), .ZN(P1_U3200) );
  INV_X1 U22871 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20744) );
  OAI222_X1 U22872 ( .A1(n22430), .A2(n20745), .B1(n20744), .B2(n22855), .C1(
        n22284), .C2(n20780), .ZN(P1_U3201) );
  INV_X1 U22873 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20746) );
  OAI222_X1 U22874 ( .A1(n20780), .A2(n22296), .B1(n20746), .B2(n22855), .C1(
        n22284), .C2(n22430), .ZN(P1_U3202) );
  INV_X1 U22875 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20747) );
  OAI222_X1 U22876 ( .A1(n20794), .A2(n22296), .B1(n20747), .B2(n22855), .C1(
        n20749), .C2(n20780), .ZN(P1_U3203) );
  INV_X1 U22877 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20748) );
  OAI222_X1 U22878 ( .A1(n20794), .A2(n20749), .B1(n20748), .B2(n22855), .C1(
        n20751), .C2(n20780), .ZN(P1_U3204) );
  INV_X1 U22879 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20750) );
  OAI222_X1 U22880 ( .A1(n20794), .A2(n20751), .B1(n20750), .B2(n22855), .C1(
        n20753), .C2(n20780), .ZN(P1_U3205) );
  INV_X1 U22881 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20752) );
  OAI222_X1 U22882 ( .A1(n22430), .A2(n20753), .B1(n20752), .B2(n22855), .C1(
        n20755), .C2(n20780), .ZN(P1_U3206) );
  INV_X1 U22883 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20754) );
  OAI222_X1 U22884 ( .A1(n20794), .A2(n20755), .B1(n20754), .B2(n22855), .C1(
        n20757), .C2(n20780), .ZN(P1_U3207) );
  INV_X1 U22885 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20756) );
  OAI222_X1 U22886 ( .A1(n22430), .A2(n20757), .B1(n20756), .B2(n22855), .C1(
        n22130), .C2(n20780), .ZN(P1_U3208) );
  INV_X1 U22887 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20758) );
  OAI222_X1 U22888 ( .A1(n20780), .A2(n20760), .B1(n20758), .B2(n22855), .C1(
        n22130), .C2(n22430), .ZN(P1_U3209) );
  INV_X1 U22889 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20759) );
  OAI222_X1 U22890 ( .A1(n20794), .A2(n20760), .B1(n20759), .B2(n22855), .C1(
        n20762), .C2(n20780), .ZN(P1_U3210) );
  INV_X1 U22891 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20761) );
  OAI222_X1 U22892 ( .A1(n20794), .A2(n20762), .B1(n20761), .B2(n22855), .C1(
        n20764), .C2(n20780), .ZN(P1_U3211) );
  INV_X1 U22893 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20763) );
  OAI222_X1 U22894 ( .A1(n20794), .A2(n20764), .B1(n20763), .B2(n22855), .C1(
        n20765), .C2(n20780), .ZN(P1_U3212) );
  INV_X1 U22895 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20766) );
  OAI222_X1 U22896 ( .A1(n20780), .A2(n20767), .B1(n20766), .B2(n22855), .C1(
        n20765), .C2(n22430), .ZN(P1_U3213) );
  INV_X1 U22897 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n22349) );
  INV_X1 U22898 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20768) );
  OAI222_X1 U22899 ( .A1(n20780), .A2(n22349), .B1(n20768), .B2(n22855), .C1(
        n20767), .C2(n22430), .ZN(P1_U3214) );
  INV_X1 U22900 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20769) );
  OAI222_X1 U22901 ( .A1(n20780), .A2(n20771), .B1(n20769), .B2(n22855), .C1(
        n22349), .C2(n22430), .ZN(P1_U3215) );
  INV_X1 U22902 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20770) );
  OAI222_X1 U22903 ( .A1(n22430), .A2(n20771), .B1(n20770), .B2(n22855), .C1(
        n20773), .C2(n20780), .ZN(P1_U3216) );
  INV_X1 U22904 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20772) );
  OAI222_X1 U22905 ( .A1(n22430), .A2(n20773), .B1(n20772), .B2(n22855), .C1(
        n20774), .C2(n20780), .ZN(P1_U3217) );
  INV_X1 U22906 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20775) );
  OAI222_X1 U22907 ( .A1(n20780), .A2(n20777), .B1(n20775), .B2(n22855), .C1(
        n20774), .C2(n22430), .ZN(P1_U3218) );
  INV_X1 U22908 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20776) );
  OAI222_X1 U22909 ( .A1(n22430), .A2(n20777), .B1(n20776), .B2(n22855), .C1(
        n20778), .C2(n20780), .ZN(P1_U3219) );
  INV_X1 U22910 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20779) );
  OAI222_X1 U22911 ( .A1(n20780), .A2(n20782), .B1(n20779), .B2(n22855), .C1(
        n20778), .C2(n22430), .ZN(P1_U3220) );
  INV_X1 U22912 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20781) );
  OAI222_X1 U22913 ( .A1(n20794), .A2(n20782), .B1(n20781), .B2(n22855), .C1(
        n20784), .C2(n20780), .ZN(P1_U3221) );
  INV_X1 U22914 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20783) );
  INV_X1 U22915 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20786) );
  OAI222_X1 U22916 ( .A1(n22430), .A2(n20784), .B1(n20783), .B2(n22855), .C1(
        n20786), .C2(n20780), .ZN(P1_U3222) );
  INV_X1 U22917 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20785) );
  OAI222_X1 U22918 ( .A1(n20794), .A2(n20786), .B1(n20785), .B2(n22855), .C1(
        n20787), .C2(n20780), .ZN(P1_U3223) );
  INV_X1 U22919 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20788) );
  OAI222_X1 U22920 ( .A1(n20780), .A2(n20790), .B1(n20788), .B2(n22855), .C1(
        n20787), .C2(n22430), .ZN(P1_U3224) );
  INV_X1 U22921 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20789) );
  OAI222_X1 U22922 ( .A1(n20794), .A2(n20790), .B1(n20789), .B2(n22855), .C1(
        n20793), .C2(n20780), .ZN(P1_U3225) );
  INV_X1 U22923 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20792) );
  OAI222_X1 U22924 ( .A1(n20794), .A2(n20793), .B1(n20792), .B2(n22855), .C1(
        n20791), .C2(n20780), .ZN(P1_U3226) );
  INV_X1 U22925 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20796) );
  INV_X1 U22926 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20795) );
  AOI22_X1 U22927 ( .A1(n22855), .A2(n20796), .B1(n20795), .B2(n22852), .ZN(
        P1_U3458) );
  INV_X1 U22928 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22407) );
  NOR3_X1 U22929 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20801) );
  AOI21_X1 U22930 ( .B1(n22247), .B2(n22407), .A(n20801), .ZN(n20797) );
  INV_X1 U22931 ( .A(n20804), .ZN(n20807) );
  AOI22_X1 U22932 ( .A1(n20804), .A2(n20797), .B1(n20796), .B2(n20807), .ZN(
        P1_U2808) );
  INV_X1 U22933 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20798) );
  AOI22_X1 U22934 ( .A1(n22855), .A2(n20799), .B1(n20798), .B2(n22852), .ZN(
        P1_U3459) );
  INV_X1 U22935 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20803) );
  INV_X1 U22936 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20800) );
  AOI22_X1 U22937 ( .A1(n22855), .A2(n20803), .B1(n20800), .B2(n22852), .ZN(
        P1_U3460) );
  OAI21_X1 U22938 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20801), .A(n20804), .ZN(
        n20802) );
  OAI21_X1 U22939 ( .B1(n20804), .B2(n20803), .A(n20802), .ZN(P1_U2807) );
  INV_X1 U22940 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20808) );
  INV_X1 U22941 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20805) );
  AOI22_X1 U22942 ( .A1(n22855), .A2(n20808), .B1(n20805), .B2(n22852), .ZN(
        P1_U3461) );
  NOR2_X1 U22943 ( .A1(n20807), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20806) );
  AOI22_X1 U22944 ( .A1(n20808), .A2(n20807), .B1(n22247), .B2(n20806), .ZN(
        P1_U3482) );
  OAI22_X1 U22945 ( .A1(n22232), .A2(n20812), .B1(n20828), .B2(n20809), .ZN(
        n20810) );
  INV_X1 U22946 ( .A(n20810), .ZN(n20811) );
  OAI21_X1 U22947 ( .B1(n20833), .B2(n22228), .A(n20811), .ZN(P1_U2870) );
  INV_X1 U22948 ( .A(n20812), .ZN(n20830) );
  INV_X1 U22949 ( .A(n20813), .ZN(n22326) );
  AOI22_X1 U22950 ( .A1(n22328), .A2(n20830), .B1(n20825), .B2(n22326), .ZN(
        n20814) );
  OAI21_X1 U22951 ( .B1(n20833), .B2(n20815), .A(n20814), .ZN(P1_U2860) );
  INV_X1 U22952 ( .A(n20816), .ZN(n20817) );
  AOI22_X1 U22953 ( .A1(n20844), .A2(n20830), .B1(n20825), .B2(n20817), .ZN(
        n20818) );
  OAI21_X1 U22954 ( .B1(n20833), .B2(n20819), .A(n20818), .ZN(P1_U2862) );
  INV_X1 U22955 ( .A(n20820), .ZN(n20863) );
  INV_X1 U22956 ( .A(n20821), .ZN(n20822) );
  AOI22_X1 U22957 ( .A1(n20863), .A2(n20830), .B1(n20825), .B2(n20822), .ZN(
        n20823) );
  OAI21_X1 U22958 ( .B1(n20833), .B2(n20824), .A(n20823), .ZN(P1_U2855) );
  INV_X1 U22959 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n20827) );
  AOI22_X1 U22960 ( .A1(n22305), .A2(n20830), .B1(n20825), .B2(n22302), .ZN(
        n20826) );
  OAI21_X1 U22961 ( .B1(n20833), .B2(n20827), .A(n20826), .ZN(P1_U2864) );
  INV_X1 U22962 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20832) );
  NOR2_X1 U22963 ( .A1(n20828), .A2(n22267), .ZN(n20829) );
  AOI21_X1 U22964 ( .B1(n22276), .B2(n20830), .A(n20829), .ZN(n20831) );
  OAI21_X1 U22965 ( .B1(n20833), .B2(n20832), .A(n20831), .ZN(P1_U2867) );
  INV_X1 U22966 ( .A(n22279), .ZN(n20834) );
  AOI222_X1 U22967 ( .A1(n20835), .A2(n20872), .B1(n20873), .B2(n22276), .C1(
        n20834), .C2(n20862), .ZN(n20837) );
  OAI211_X1 U22968 ( .C1(n20842), .C2(n22270), .A(n20837), .B(n20836), .ZN(
        P1_U2994) );
  INV_X1 U22969 ( .A(n22301), .ZN(n20838) );
  AOI222_X1 U22970 ( .A1(n20839), .A2(n20872), .B1(n20873), .B2(n22298), .C1(
        n20838), .C2(n20862), .ZN(n20841) );
  OAI211_X1 U22971 ( .C1(n20842), .C2(n22291), .A(n20841), .B(n20840), .ZN(
        P1_U2992) );
  AOI22_X1 U22972 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n22190), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20870), .ZN(n20846) );
  AOI22_X1 U22973 ( .A1(n20844), .A2(n20873), .B1(n20862), .B2(n20843), .ZN(
        n20845) );
  OAI211_X1 U22974 ( .C1(n22385), .C2(n20847), .A(n20846), .B(n20845), .ZN(
        P1_U2989) );
  AOI211_X1 U22975 ( .C1(n20870), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20850), .B(n20849), .ZN(n20851) );
  OAI21_X1 U22976 ( .B1(n20853), .B2(n20852), .A(n20851), .ZN(P1_U2988) );
  AOI22_X1 U22977 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n22202), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20870), .ZN(n20855) );
  AOI22_X1 U22978 ( .A1(n20862), .A2(n22329), .B1(n20873), .B2(n22328), .ZN(
        n20854) );
  OAI211_X1 U22979 ( .C1(n20856), .C2(n22385), .A(n20855), .B(n20854), .ZN(
        P1_U2987) );
  MUX2_X1 U22980 ( .A(n14256), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .S(
        n13229), .Z(n20857) );
  XNOR2_X1 U22981 ( .A(n20858), .B(n20857), .ZN(n22163) );
  AOI22_X1 U22982 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n22202), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20870), .ZN(n20860) );
  AOI22_X1 U22983 ( .A1(n22345), .A2(n20873), .B1(n20862), .B2(n22344), .ZN(
        n20859) );
  OAI211_X1 U22984 ( .C1(n22385), .C2(n22163), .A(n20860), .B(n20859), .ZN(
        P1_U2984) );
  AOI22_X1 U22985 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22202), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20870), .ZN(n20865) );
  AOI22_X1 U22986 ( .A1(n20863), .A2(n20873), .B1(n20862), .B2(n20861), .ZN(
        n20864) );
  OAI211_X1 U22987 ( .C1(n20866), .C2(n22385), .A(n20865), .B(n20864), .ZN(
        P1_U2982) );
  AOI22_X1 U22988 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n22202), .B1(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20870), .ZN(n20869) );
  AOI22_X1 U22989 ( .A1(n22363), .A2(n20873), .B1(n20872), .B2(n20867), .ZN(
        n20868) );
  OAI211_X1 U22990 ( .C1(n20877), .C2(n22351), .A(n20869), .B(n20868), .ZN(
        P1_U2980) );
  AOI22_X1 U22991 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22190), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20870), .ZN(n20876) );
  AOI22_X1 U22992 ( .A1(n20874), .A2(n20873), .B1(n20872), .B2(n20871), .ZN(
        n20875) );
  OAI211_X1 U22993 ( .C1(n20877), .C2(n22384), .A(n20876), .B(n20875), .ZN(
        P1_U2978) );
  INV_X1 U22994 ( .A(n20878), .ZN(n20879) );
  OAI21_X1 U22995 ( .B1(n20879), .B2(n22402), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20880) );
  OAI21_X1 U22996 ( .B1(n20881), .B2(n22392), .A(n20880), .ZN(P1_U2803) );
  INV_X1 U22997 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20882) );
  OAI222_X1 U22998 ( .A1(n22855), .A2(n20883), .B1(n22855), .B2(n20882), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(n22852), .ZN(P1_U2804) );
  INV_X1 U22999 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20886) );
  INV_X2 U23000 ( .A(U212), .ZN(n20931) );
  AOI22_X1 U23001 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n20947), .ZN(n20885) );
  OAI21_X1 U23002 ( .B1(n20886), .B2(n20933), .A(n20885), .ZN(U247) );
  AOI22_X1 U23003 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n20947), .ZN(n20887) );
  OAI21_X1 U23004 ( .B1(n20888), .B2(n20933), .A(n20887), .ZN(U246) );
  AOI22_X1 U23005 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n20947), .ZN(n20889) );
  OAI21_X1 U23006 ( .B1(n20890), .B2(n20933), .A(n20889), .ZN(U245) );
  AOI22_X1 U23007 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n20947), .ZN(n20891) );
  OAI21_X1 U23008 ( .B1(n20892), .B2(n20933), .A(n20891), .ZN(U244) );
  INV_X1 U23009 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20894) );
  AOI22_X1 U23010 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n20947), .ZN(n20893) );
  OAI21_X1 U23011 ( .B1(n20894), .B2(n20933), .A(n20893), .ZN(U243) );
  AOI22_X1 U23012 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n20947), .ZN(n20895) );
  OAI21_X1 U23013 ( .B1(n20896), .B2(n20933), .A(n20895), .ZN(U242) );
  AOI22_X1 U23014 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n20947), .ZN(n20897) );
  OAI21_X1 U23015 ( .B1(n20898), .B2(n20933), .A(n20897), .ZN(U241) );
  AOI22_X1 U23016 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n20947), .ZN(n20899) );
  OAI21_X1 U23017 ( .B1(n20900), .B2(n20933), .A(n20899), .ZN(U240) );
  AOI22_X1 U23018 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n20947), .ZN(n20901) );
  OAI21_X1 U23019 ( .B1(n20902), .B2(n20933), .A(n20901), .ZN(U239) );
  AOI22_X1 U23020 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n20947), .ZN(n20903) );
  OAI21_X1 U23021 ( .B1(n20904), .B2(n20933), .A(n20903), .ZN(U238) );
  AOI22_X1 U23022 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n20947), .ZN(n20905) );
  OAI21_X1 U23023 ( .B1(n20906), .B2(n20933), .A(n20905), .ZN(U237) );
  AOI22_X1 U23024 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n20947), .ZN(n20907) );
  OAI21_X1 U23025 ( .B1(n20908), .B2(n20933), .A(n20907), .ZN(U236) );
  AOI22_X1 U23026 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n20947), .ZN(n20909) );
  OAI21_X1 U23027 ( .B1(n20910), .B2(n20933), .A(n20909), .ZN(U235) );
  AOI22_X1 U23028 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n20947), .ZN(n20911) );
  OAI21_X1 U23029 ( .B1(n20912), .B2(n20933), .A(n20911), .ZN(U234) );
  AOI22_X1 U23030 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n20947), .ZN(n20913) );
  OAI21_X1 U23031 ( .B1(n20914), .B2(n20933), .A(n20913), .ZN(U233) );
  INV_X1 U23032 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20916) );
  AOI22_X1 U23033 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n20947), .ZN(n20915) );
  OAI21_X1 U23034 ( .B1(n20916), .B2(n20933), .A(n20915), .ZN(U232) );
  AOI22_X1 U23035 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20947), .ZN(n20917) );
  OAI21_X1 U23036 ( .B1(n20918), .B2(n20933), .A(n20917), .ZN(U231) );
  AOI22_X1 U23037 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n20947), .ZN(n20919) );
  OAI21_X1 U23038 ( .B1(n20920), .B2(n20933), .A(n20919), .ZN(U230) );
  AOI22_X1 U23039 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n20947), .ZN(n20921) );
  OAI21_X1 U23040 ( .B1(n20922), .B2(n20933), .A(n20921), .ZN(U229) );
  INV_X1 U23041 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U23042 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n20947), .ZN(n20923) );
  OAI21_X1 U23043 ( .B1(n20924), .B2(n20933), .A(n20923), .ZN(U228) );
  AOI22_X1 U23044 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n20947), .ZN(n20925) );
  OAI21_X1 U23045 ( .B1(n20926), .B2(n20933), .A(n20925), .ZN(U227) );
  AOI22_X1 U23046 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n20947), .ZN(n20927) );
  OAI21_X1 U23047 ( .B1(n20928), .B2(n20933), .A(n20927), .ZN(U226) );
  AOI22_X1 U23048 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n20947), .ZN(n20929) );
  OAI21_X1 U23049 ( .B1(n20930), .B2(n20933), .A(n20929), .ZN(U225) );
  AOI22_X1 U23050 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n20947), .ZN(n20932) );
  OAI21_X1 U23051 ( .B1(n20934), .B2(n20933), .A(n20932), .ZN(U224) );
  AOI22_X1 U23052 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n20947), .ZN(n20935) );
  OAI21_X1 U23053 ( .B1(n20936), .B2(n20933), .A(n20935), .ZN(U223) );
  AOI22_X1 U23054 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n20947), .ZN(n20937) );
  OAI21_X1 U23055 ( .B1(n20938), .B2(n20933), .A(n20937), .ZN(U222) );
  AOI22_X1 U23056 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n20947), .ZN(n20939) );
  OAI21_X1 U23057 ( .B1(n20940), .B2(n20933), .A(n20939), .ZN(U221) );
  AOI22_X1 U23058 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n20947), .ZN(n20941) );
  OAI21_X1 U23059 ( .B1(n20942), .B2(n20933), .A(n20941), .ZN(U220) );
  AOI22_X1 U23060 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n20947), .ZN(n20943) );
  OAI21_X1 U23061 ( .B1(n20944), .B2(n20933), .A(n20943), .ZN(U219) );
  AOI22_X1 U23062 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n20947), .ZN(n20945) );
  OAI21_X1 U23063 ( .B1(n20946), .B2(n20933), .A(n20945), .ZN(U218) );
  AOI22_X1 U23064 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n20931), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20947), .ZN(n20948) );
  OAI21_X1 U23065 ( .B1(n20949), .B2(n20933), .A(n20948), .ZN(U217) );
  OAI222_X1 U23066 ( .A1(U214), .A2(n20952), .B1(n20933), .B2(n20951), .C1(
        U212), .C2(n20950), .ZN(U216) );
  AOI22_X1 U23067 ( .A1(n22855), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20953), 
        .B2(n22852), .ZN(P1_U3483) );
  OAI21_X1 U23068 ( .B1(n22418), .B2(n20955), .A(n20954), .ZN(n20956) );
  AOI21_X1 U23069 ( .B1(n20957), .B2(n21653), .A(n20956), .ZN(n20965) );
  AOI21_X1 U23070 ( .B1(n20959), .B2(n22414), .A(n20958), .ZN(n20960) );
  OAI211_X1 U23071 ( .C1(n20961), .C2(n20960), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n22470), .ZN(n20962) );
  AOI21_X1 U23072 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20962), .A(n22088), 
        .ZN(n20964) );
  NAND2_X1 U23073 ( .A1(n20965), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20963) );
  OAI21_X1 U23074 ( .B1(n20965), .B2(n20964), .A(n20963), .ZN(P3_U3296) );
  NAND2_X2 U23075 ( .A1(n20967), .A2(n20966), .ZN(n21022) );
  INV_X1 U23076 ( .A(n21430), .ZN(n20968) );
  NOR2_X4 U23077 ( .A1(n20969), .A2(n20968), .ZN(n21008) );
  AOI22_X1 U23078 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20987), .ZN(n20970) );
  OAI21_X1 U23079 ( .B1(n20971), .B2(n21022), .A(n20970), .ZN(P3_U2768) );
  AOI22_X1 U23080 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20987), .ZN(n20972) );
  OAI21_X1 U23081 ( .B1(n20973), .B2(n21022), .A(n20972), .ZN(P3_U2769) );
  AOI22_X1 U23082 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20987), .ZN(n20974) );
  OAI21_X1 U23083 ( .B1(n20975), .B2(n21022), .A(n20974), .ZN(P3_U2770) );
  AOI22_X1 U23084 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20987), .ZN(n20977) );
  OAI21_X1 U23085 ( .B1(n21489), .B2(n21022), .A(n20977), .ZN(P3_U2771) );
  AOI22_X1 U23086 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20987), .ZN(n20978) );
  OAI21_X1 U23087 ( .B1(n21508), .B2(n21022), .A(n20978), .ZN(P3_U2772) );
  AOI22_X1 U23088 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20987), .ZN(n20979) );
  OAI21_X1 U23089 ( .B1(n21502), .B2(n21022), .A(n20979), .ZN(P3_U2773) );
  AOI22_X1 U23090 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20987), .ZN(n20980) );
  OAI21_X1 U23091 ( .B1(n21531), .B2(n21022), .A(n20980), .ZN(P3_U2774) );
  AOI22_X1 U23092 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20987), .ZN(n20981) );
  OAI21_X1 U23093 ( .B1(n20982), .B2(n21022), .A(n20981), .ZN(P3_U2775) );
  AOI22_X1 U23094 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20987), .ZN(n20983) );
  OAI21_X1 U23095 ( .B1(n20984), .B2(n21022), .A(n20983), .ZN(P3_U2776) );
  AOI22_X1 U23096 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20987), .ZN(n20985) );
  OAI21_X1 U23097 ( .B1(n20986), .B2(n21022), .A(n20985), .ZN(P3_U2777) );
  AOI22_X1 U23098 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n21020), .ZN(n20988) );
  OAI21_X1 U23099 ( .B1(n21540), .B2(n21022), .A(n20988), .ZN(P3_U2778) );
  AOI22_X1 U23100 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n21020), .ZN(n20989) );
  OAI21_X1 U23101 ( .B1(n20990), .B2(n21022), .A(n20989), .ZN(P3_U2779) );
  AOI22_X1 U23102 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n21020), .ZN(n20991) );
  OAI21_X1 U23103 ( .B1(n21558), .B2(n21022), .A(n20991), .ZN(P3_U2780) );
  AOI22_X1 U23104 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n21020), .ZN(n20992) );
  OAI21_X1 U23105 ( .B1(n20993), .B2(n21022), .A(n20992), .ZN(P3_U2781) );
  AOI22_X1 U23106 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21008), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n21020), .ZN(n20994) );
  OAI21_X1 U23107 ( .B1(n20995), .B2(n21022), .A(n20994), .ZN(P3_U2782) );
  AOI22_X1 U23108 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n21020), .ZN(n20996) );
  OAI21_X1 U23109 ( .B1(n21615), .B2(n21022), .A(n20996), .ZN(P3_U2783) );
  AOI22_X1 U23110 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n21020), .ZN(n20997) );
  OAI21_X1 U23111 ( .B1(n20998), .B2(n21022), .A(n20997), .ZN(P3_U2784) );
  AOI22_X1 U23112 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n21020), .ZN(n20999) );
  OAI21_X1 U23113 ( .B1(n21000), .B2(n21022), .A(n20999), .ZN(P3_U2785) );
  AOI22_X1 U23114 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n21020), .ZN(n21001) );
  OAI21_X1 U23115 ( .B1(n21002), .B2(n21022), .A(n21001), .ZN(P3_U2786) );
  AOI22_X1 U23116 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n21020), .ZN(n21003) );
  OAI21_X1 U23117 ( .B1(n21465), .B2(n21022), .A(n21003), .ZN(P3_U2787) );
  AOI22_X1 U23118 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n21020), .ZN(n21004) );
  OAI21_X1 U23119 ( .B1(n21005), .B2(n21022), .A(n21004), .ZN(P3_U2788) );
  AOI22_X1 U23120 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n21020), .ZN(n21006) );
  OAI21_X1 U23121 ( .B1(n21007), .B2(n21022), .A(n21006), .ZN(P3_U2789) );
  AOI22_X1 U23122 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n21020), .ZN(n21009) );
  OAI21_X1 U23123 ( .B1(n21010), .B2(n21022), .A(n21009), .ZN(P3_U2790) );
  AOI22_X1 U23124 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n21020), .ZN(n21011) );
  OAI21_X1 U23125 ( .B1(n21597), .B2(n21022), .A(n21011), .ZN(P3_U2791) );
  AOI22_X1 U23126 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n21020), .ZN(n21012) );
  OAI21_X1 U23127 ( .B1(n21457), .B2(n21022), .A(n21012), .ZN(P3_U2792) );
  AOI22_X1 U23128 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n21020), .ZN(n21013) );
  OAI21_X1 U23129 ( .B1(n21014), .B2(n21022), .A(n21013), .ZN(P3_U2793) );
  AOI22_X1 U23130 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n21020), .ZN(n21015) );
  OAI21_X1 U23131 ( .B1(n21450), .B2(n21022), .A(n21015), .ZN(P3_U2794) );
  AOI22_X1 U23132 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n21020), .ZN(n21016) );
  OAI21_X1 U23133 ( .B1(n21437), .B2(n21022), .A(n21016), .ZN(P3_U2795) );
  AOI22_X1 U23134 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n21020), .ZN(n21017) );
  OAI21_X1 U23135 ( .B1(n21018), .B2(n21022), .A(n21017), .ZN(P3_U2796) );
  AOI22_X1 U23136 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n21020), .ZN(n21019) );
  OAI21_X1 U23137 ( .B1(n21585), .B2(n21022), .A(n21019), .ZN(P3_U2797) );
  AOI22_X1 U23138 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n21008), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n21020), .ZN(n21021) );
  OAI21_X1 U23139 ( .B1(n21592), .B2(n21022), .A(n21021), .ZN(P3_U2798) );
  INV_X1 U23140 ( .A(n11262), .ZN(n21420) );
  INV_X1 U23141 ( .A(n21023), .ZN(n21621) );
  AOI22_X1 U23142 ( .A1(n21424), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n21621), .B2(
        n21421), .ZN(n21030) );
  INV_X1 U23143 ( .A(n21249), .ZN(n21400) );
  NOR2_X1 U23144 ( .A1(n21400), .A2(n21214), .ZN(n21410) );
  INV_X1 U23145 ( .A(n21410), .ZN(n21112) );
  OAI21_X1 U23146 ( .B1(n21113), .B2(n21112), .A(n21357), .ZN(n21028) );
  AOI21_X1 U23147 ( .B1(n21399), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21400), .ZN(n21026) );
  OAI22_X1 U23148 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n21419), .B1(n21397), 
        .B2(n21024), .ZN(n21025) );
  AOI221_X1 U23149 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21028), .C1(
        n21027), .C2(n21026), .A(n21025), .ZN(n21029) );
  OAI211_X1 U23150 ( .C1(n21420), .C2(n21687), .A(n21030), .B(n21029), .ZN(
        P3_U2670) );
  AOI22_X1 U23151 ( .A1(n21424), .A2(P3_EBX_REG_3__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n21404), .ZN(n21042) );
  NOR2_X1 U23152 ( .A1(n21064), .A2(n21419), .ZN(n21032) );
  OR2_X1 U23153 ( .A1(n18658), .A2(n21031), .ZN(n21635) );
  AOI22_X1 U23154 ( .A1(n21033), .A2(n21032), .B1(n21421), .B2(n21635), .ZN(
        n21041) );
  XNOR2_X1 U23155 ( .A(n21035), .B(n21034), .ZN(n21036) );
  OAI21_X1 U23156 ( .B1(n21064), .B2(n21327), .A(n21420), .ZN(n21053) );
  AOI22_X1 U23157 ( .A1(n11533), .A2(n21036), .B1(P3_REIP_REG_3__SCAN_IN), 
        .B2(n21053), .ZN(n21040) );
  NAND2_X1 U23158 ( .A1(n21038), .A2(n21037), .ZN(n21044) );
  OAI211_X1 U23159 ( .C1(n21038), .C2(n21037), .A(n21423), .B(n21044), .ZN(
        n21039) );
  NAND4_X1 U23160 ( .A1(n21042), .A2(n21041), .A3(n21040), .A4(n21039), .ZN(
        P3_U2668) );
  INV_X1 U23161 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n21057) );
  AOI221_X1 U23162 ( .B1(n21043), .B2(n21421), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n21421), .A(n22073), .ZN(
        n21050) );
  NAND2_X1 U23163 ( .A1(n21249), .A2(n21113), .ZN(n21172) );
  OAI21_X1 U23164 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n21172), .A(
        n21171), .ZN(n21047) );
  AOI211_X1 U23165 ( .C1(n21058), .C2(n21113), .A(n21048), .B(n21112), .ZN(
        n21046) );
  NOR2_X1 U23166 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n21044), .ZN(n21062) );
  AOI211_X1 U23167 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n21044), .A(n21062), .B(
        n21397), .ZN(n21045) );
  AOI211_X1 U23168 ( .C1(n21048), .C2(n21047), .A(n21046), .B(n21045), .ZN(
        n21049) );
  OAI211_X1 U23169 ( .C1(n21051), .C2(n21357), .A(n21050), .B(n21049), .ZN(
        n21052) );
  AOI21_X1 U23170 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n21053), .A(n21052), .ZN(
        n21056) );
  NAND3_X1 U23171 ( .A1(n21341), .A2(n21064), .A3(n21054), .ZN(n21055) );
  OAI211_X1 U23172 ( .C1(n21057), .C2(n21359), .A(n21056), .B(n21055), .ZN(
        P3_U2667) );
  AOI21_X1 U23173 ( .B1(n21058), .B2(n21113), .A(n21214), .ZN(n21060) );
  XOR2_X1 U23174 ( .A(n21060), .B(n21059), .Z(n21072) );
  INV_X1 U23175 ( .A(n21062), .ZN(n21061) );
  AOI21_X1 U23176 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n21061), .A(n21397), .ZN(
        n21063) );
  NAND2_X1 U23177 ( .A1(n21062), .A2(n21068), .ZN(n21079) );
  AOI22_X1 U23178 ( .A1(n21404), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n21063), .B2(n21079), .ZN(n21071) );
  NAND2_X1 U23179 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n21064), .ZN(n21067) );
  NOR2_X1 U23180 ( .A1(n21065), .A2(n21067), .ZN(n21087) );
  OAI21_X1 U23181 ( .B1(n21087), .B2(n21327), .A(n21420), .ZN(n21093) );
  INV_X1 U23182 ( .A(n21087), .ZN(n21073) );
  NAND2_X1 U23183 ( .A1(n21341), .A2(n21073), .ZN(n21066) );
  OAI22_X1 U23184 ( .A1(n21359), .A2(n21068), .B1(n21067), .B2(n21066), .ZN(
        n21069) );
  AOI211_X1 U23185 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n21093), .A(n22073), .B(
        n21069), .ZN(n21070) );
  OAI211_X1 U23186 ( .C1(n21400), .C2(n21072), .A(n21071), .B(n21070), .ZN(
        P3_U2666) );
  NOR3_X1 U23187 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n21419), .A3(n21073), .ZN(
        n21094) );
  AOI21_X1 U23188 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n21424), .A(n21094), .ZN(
        n21084) );
  OAI21_X1 U23189 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n21172), .A(
        n21171), .ZN(n21076) );
  AOI21_X1 U23190 ( .B1(n21074), .B2(n21113), .A(n21214), .ZN(n21086) );
  NOR2_X1 U23191 ( .A1(n21077), .A2(n21400), .ZN(n21075) );
  AOI22_X1 U23192 ( .A1(n21077), .A2(n21076), .B1(n21086), .B2(n21075), .ZN(
        n21083) );
  NOR2_X1 U23193 ( .A1(n21078), .A2(n21357), .ZN(n21081) );
  NOR2_X1 U23194 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n21079), .ZN(n21088) );
  AOI211_X1 U23195 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n21079), .A(n21088), .B(
        n21397), .ZN(n21080) );
  AOI211_X1 U23196 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n21093), .A(n21081), .B(
        n21080), .ZN(n21082) );
  NAND4_X1 U23197 ( .A1(n21084), .A2(n21083), .A3(n21082), .A4(n22049), .ZN(
        P3_U2665) );
  XOR2_X1 U23198 ( .A(n21086), .B(n21085), .Z(n21097) );
  NAND2_X1 U23199 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n21087), .ZN(n21098) );
  NOR3_X1 U23200 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n21419), .A3(n21098), .ZN(
        n21092) );
  NAND2_X1 U23201 ( .A1(n21088), .A2(n21090), .ZN(n21100) );
  OAI211_X1 U23202 ( .C1(n21088), .C2(n21090), .A(n21423), .B(n21100), .ZN(
        n21089) );
  OAI211_X1 U23203 ( .C1(n21359), .C2(n21090), .A(n22049), .B(n21089), .ZN(
        n21091) );
  AOI211_X1 U23204 ( .C1(n21404), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n21092), .B(n21091), .ZN(n21096) );
  OAI21_X1 U23205 ( .B1(n21094), .B2(n21093), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n21095) );
  OAI211_X1 U23206 ( .C1(n21097), .C2(n21400), .A(n21096), .B(n21095), .ZN(
        P3_U2664) );
  AOI22_X1 U23207 ( .A1(n21424), .A2(P3_EBX_REG_8__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n21404), .ZN(n21111) );
  NOR2_X1 U23208 ( .A1(n21099), .A2(n21098), .ZN(n21103) );
  NAND2_X1 U23209 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n21103), .ZN(n21126) );
  AND2_X1 U23210 ( .A1(n21126), .A2(n21341), .ZN(n21102) );
  AOI211_X1 U23211 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n21100), .A(n21118), .B(
        n21397), .ZN(n21101) );
  AOI211_X1 U23212 ( .C1(n21103), .C2(n21102), .A(n22073), .B(n21101), .ZN(
        n21110) );
  OAI21_X1 U23213 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21104), .A(
        n21399), .ZN(n21105) );
  XNOR2_X1 U23214 ( .A(n21106), .B(n21105), .ZN(n21108) );
  AOI21_X1 U23215 ( .B1(n21341), .B2(n21126), .A(n11262), .ZN(n21138) );
  INV_X1 U23216 ( .A(n21138), .ZN(n21107) );
  AOI22_X1 U23217 ( .A1(n11533), .A2(n21108), .B1(P3_REIP_REG_8__SCAN_IN), 
        .B2(n21107), .ZN(n21109) );
  NAND3_X1 U23218 ( .A1(n21111), .A2(n21110), .A3(n21109), .ZN(P3_U2663) );
  AOI211_X1 U23219 ( .C1(n21114), .C2(n21113), .A(n21116), .B(n21112), .ZN(
        n21124) );
  NAND2_X1 U23220 ( .A1(n21341), .A2(n21127), .ZN(n21137) );
  OAI21_X1 U23221 ( .B1(n21126), .B2(n21137), .A(n22049), .ZN(n21123) );
  OAI21_X1 U23222 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n21172), .A(
        n21171), .ZN(n21115) );
  AOI22_X1 U23223 ( .A1(n21424), .A2(P3_EBX_REG_9__SCAN_IN), .B1(n21116), .B2(
        n21115), .ZN(n21120) );
  NAND2_X1 U23224 ( .A1(n21118), .A2(n21117), .ZN(n21128) );
  OAI211_X1 U23225 ( .C1(n21118), .C2(n21117), .A(n21423), .B(n21128), .ZN(
        n21119) );
  OAI211_X1 U23226 ( .C1(n21357), .C2(n21121), .A(n21120), .B(n21119), .ZN(
        n21122) );
  NOR3_X1 U23227 ( .A1(n21124), .A2(n21123), .A3(n21122), .ZN(n21125) );
  OAI21_X1 U23228 ( .B1(n21138), .B2(n21127), .A(n21125), .ZN(P3_U2662) );
  NOR2_X1 U23229 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n21419), .ZN(n21135) );
  NOR2_X1 U23230 ( .A1(n21127), .A2(n21126), .ZN(n21140) );
  AOI211_X1 U23231 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n21128), .A(n21146), .B(
        n21397), .ZN(n21134) );
  OAI21_X1 U23232 ( .B1(n21129), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21399), .ZN(n21142) );
  XNOR2_X1 U23233 ( .A(n21142), .B(n21130), .ZN(n21132) );
  AOI22_X1 U23234 ( .A1(n21424), .A2(P3_EBX_REG_10__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n21404), .ZN(n21131) );
  OAI211_X1 U23235 ( .C1(n21400), .C2(n21132), .A(n21131), .B(n22049), .ZN(
        n21133) );
  AOI211_X1 U23236 ( .C1(n21135), .C2(n21140), .A(n21134), .B(n21133), .ZN(
        n21136) );
  OAI221_X1 U23237 ( .B1(n21139), .B2(n21138), .C1(n21139), .C2(n21137), .A(
        n21136), .ZN(P3_U2661) );
  NAND2_X1 U23238 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n21140), .ZN(n21141) );
  OAI21_X1 U23239 ( .B1(n21170), .B2(n21327), .A(n21420), .ZN(n21163) );
  OAI21_X1 U23240 ( .B1(n21327), .B2(n21141), .A(n21781), .ZN(n21151) );
  OAI21_X1 U23241 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n21214), .A(
        n21142), .ZN(n21144) );
  AOI21_X1 U23242 ( .B1(n21145), .B2(n21144), .A(n21400), .ZN(n21143) );
  OAI21_X1 U23243 ( .B1(n21145), .B2(n21144), .A(n21143), .ZN(n21148) );
  NAND2_X1 U23244 ( .A1(n21146), .A2(n21153), .ZN(n21158) );
  OAI211_X1 U23245 ( .C1(n21146), .C2(n21153), .A(n21423), .B(n21158), .ZN(
        n21147) );
  OAI211_X1 U23246 ( .C1(n21357), .C2(n21149), .A(n21148), .B(n21147), .ZN(
        n21150) );
  AOI21_X1 U23247 ( .B1(n21163), .B2(n21151), .A(n21150), .ZN(n21152) );
  OAI211_X1 U23248 ( .C1(n21359), .C2(n21153), .A(n21152), .B(n22049), .ZN(
        P3_U2660) );
  INV_X1 U23249 ( .A(n21154), .ZN(n21155) );
  AOI21_X1 U23250 ( .B1(n21155), .B2(n21195), .A(n21214), .ZN(n21157) );
  XOR2_X1 U23251 ( .A(n21157), .B(n21156), .Z(n21166) );
  AOI22_X1 U23252 ( .A1(n21424), .A2(P3_EBX_REG_12__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n21404), .ZN(n21165) );
  AOI211_X1 U23253 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n21158), .A(n21178), .B(
        n21397), .ZN(n21162) );
  INV_X1 U23254 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n21159) );
  NAND3_X1 U23255 ( .A1(n21341), .A2(n21170), .A3(n21159), .ZN(n21160) );
  NAND2_X1 U23256 ( .A1(n22049), .A2(n21160), .ZN(n21161) );
  AOI211_X1 U23257 ( .C1(n21163), .C2(P3_REIP_REG_12__SCAN_IN), .A(n21162), 
        .B(n21161), .ZN(n21164) );
  OAI211_X1 U23258 ( .C1(n21400), .C2(n21166), .A(n21165), .B(n21164), .ZN(
        P3_U2659) );
  AOI22_X1 U23259 ( .A1(n21424), .A2(P3_EBX_REG_13__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n21404), .ZN(n21182) );
  AOI21_X1 U23260 ( .B1(n21167), .B2(n21195), .A(n21214), .ZN(n21188) );
  NOR2_X1 U23261 ( .A1(n21175), .A2(n21400), .ZN(n21169) );
  NAND2_X1 U23262 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n21170), .ZN(n21184) );
  NOR3_X1 U23263 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n21419), .A3(n21184), 
        .ZN(n21168) );
  AOI211_X1 U23264 ( .C1(n21188), .C2(n21169), .A(n22073), .B(n21168), .ZN(
        n21181) );
  OAI221_X1 U23265 ( .B1(n21327), .B2(P3_REIP_REG_12__SCAN_IN), .C1(n21327), 
        .C2(n21170), .A(n21420), .ZN(n21176) );
  OAI21_X1 U23266 ( .B1(n21173), .B2(n21172), .A(n21171), .ZN(n21174) );
  AOI22_X1 U23267 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n21176), .B1(n21175), 
        .B2(n21174), .ZN(n21180) );
  NAND2_X1 U23268 ( .A1(n21178), .A2(n21177), .ZN(n21183) );
  OAI211_X1 U23269 ( .C1(n21178), .C2(n21177), .A(n21423), .B(n21183), .ZN(
        n21179) );
  NAND4_X1 U23270 ( .A1(n21182), .A2(n21181), .A3(n21180), .A4(n21179), .ZN(
        P3_U2658) );
  AOI211_X1 U23271 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n21183), .A(n21199), .B(
        n21397), .ZN(n21192) );
  NOR2_X1 U23272 ( .A1(n21185), .A2(n21184), .ZN(n21186) );
  AOI21_X1 U23273 ( .B1(n21341), .B2(n21186), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n21190) );
  NAND2_X1 U23274 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n21186), .ZN(n21206) );
  AOI21_X1 U23275 ( .B1(n21206), .B2(n21341), .A(n11262), .ZN(n21211) );
  XOR2_X1 U23276 ( .A(n21188), .B(n21187), .Z(n21189) );
  OAI22_X1 U23277 ( .A1(n21190), .A2(n21211), .B1(n21400), .B2(n21189), .ZN(
        n21191) );
  AOI211_X1 U23278 ( .C1(n21404), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n21192), .B(n21191), .ZN(n21193) );
  OAI211_X1 U23279 ( .C1(n21359), .C2(n21194), .A(n21193), .B(n22049), .ZN(
        P3_U2657) );
  NAND2_X1 U23280 ( .A1(n21196), .A2(n21195), .ZN(n21228) );
  INV_X1 U23281 ( .A(n21228), .ZN(n21215) );
  NOR2_X1 U23282 ( .A1(n21215), .A2(n21214), .ZN(n21198) );
  XOR2_X1 U23283 ( .A(n21198), .B(n21197), .Z(n21204) );
  INV_X1 U23284 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n21202) );
  NOR3_X1 U23285 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n21419), .A3(n21206), 
        .ZN(n21213) );
  AOI211_X1 U23286 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n21404), .A(
        n22073), .B(n21213), .ZN(n21201) );
  NAND2_X1 U23287 ( .A1(n21199), .A2(n21202), .ZN(n21209) );
  OAI211_X1 U23288 ( .C1(n21199), .C2(n21202), .A(n21423), .B(n21209), .ZN(
        n21200) );
  OAI211_X1 U23289 ( .C1(n21202), .C2(n21359), .A(n21201), .B(n21200), .ZN(
        n21203) );
  AOI21_X1 U23290 ( .B1(n21204), .B2(n11533), .A(n21203), .ZN(n21205) );
  OAI21_X1 U23291 ( .B1(n21207), .B2(n21211), .A(n21205), .ZN(P3_U2656) );
  NOR2_X1 U23292 ( .A1(n21207), .A2(n21206), .ZN(n21223) );
  NOR2_X1 U23293 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n21419), .ZN(n21208) );
  AOI22_X1 U23294 ( .A1(n21424), .A2(P3_EBX_REG_16__SCAN_IN), .B1(n21223), 
        .B2(n21208), .ZN(n21222) );
  AOI211_X1 U23295 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n21209), .A(n21233), .B(
        n21397), .ZN(n21210) );
  AOI211_X1 U23296 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n21404), .A(
        n22073), .B(n21210), .ZN(n21221) );
  INV_X1 U23297 ( .A(n21211), .ZN(n21212) );
  OAI21_X1 U23298 ( .B1(n21213), .B2(n21212), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n21220) );
  AOI21_X1 U23299 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n21215), .A(
        n21214), .ZN(n21217) );
  AOI21_X1 U23300 ( .B1(n21218), .B2(n21217), .A(n21400), .ZN(n21216) );
  OAI21_X1 U23301 ( .B1(n21218), .B2(n21217), .A(n21216), .ZN(n21219) );
  NAND4_X1 U23302 ( .A1(n21222), .A2(n21221), .A3(n21220), .A4(n21219), .ZN(
        P3_U2655) );
  NAND2_X1 U23303 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n21223), .ZN(n21226) );
  OAI21_X1 U23304 ( .B1(n21261), .B2(n21327), .A(n21420), .ZN(n21256) );
  OR2_X1 U23305 ( .A1(n21419), .A2(n21261), .ZN(n21225) );
  OAI22_X1 U23306 ( .A1(n21359), .A2(n21232), .B1(n21226), .B2(n21225), .ZN(
        n21227) );
  AOI211_X1 U23307 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n21256), .A(n22073), 
        .B(n21227), .ZN(n21237) );
  OAI211_X1 U23308 ( .C1(n21231), .C2(n21230), .A(n11533), .B(n21242), .ZN(
        n21236) );
  NAND2_X1 U23309 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n21404), .ZN(
        n21235) );
  NAND2_X1 U23310 ( .A1(n21233), .A2(n21232), .ZN(n21238) );
  OAI211_X1 U23311 ( .C1(n21233), .C2(n21232), .A(n21423), .B(n21238), .ZN(
        n21234) );
  NAND4_X1 U23312 ( .A1(n21237), .A2(n21236), .A3(n21235), .A4(n21234), .ZN(
        P3_U2654) );
  AOI211_X1 U23313 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n21238), .A(n21257), .B(
        n21397), .ZN(n21239) );
  AOI21_X1 U23314 ( .B1(n21404), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21239), .ZN(n21247) );
  NAND2_X1 U23315 ( .A1(n21341), .A2(n21261), .ZN(n21263) );
  OAI22_X1 U23316 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n21263), .B1(n21359), 
        .B2(n21240), .ZN(n21241) );
  AOI211_X1 U23317 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(n21256), .A(n22073), 
        .B(n21241), .ZN(n21246) );
  NAND2_X1 U23318 ( .A1(n21243), .A2(n21244), .ZN(n21248) );
  OAI211_X1 U23319 ( .C1(n21244), .C2(n21243), .A(n11533), .B(n21248), .ZN(
        n21245) );
  NAND3_X1 U23320 ( .A1(n21247), .A2(n21246), .A3(n21245), .ZN(P3_U2653) );
  INV_X1 U23321 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n21260) );
  NAND2_X1 U23322 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n21264) );
  OAI21_X1 U23323 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(P3_REIP_REG_19__SCAN_IN), 
        .A(n21264), .ZN(n21254) );
  AOI21_X1 U23324 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n21404), .A(
        n21869), .ZN(n21253) );
  NAND2_X1 U23325 ( .A1(n21399), .A2(n21248), .ZN(n21250) );
  NAND2_X1 U23326 ( .A1(n21250), .A2(n21251), .ZN(n21267) );
  OAI211_X1 U23327 ( .C1(n21251), .C2(n21250), .A(n21249), .B(n21267), .ZN(
        n21252) );
  OAI211_X1 U23328 ( .C1(n21263), .C2(n21254), .A(n21253), .B(n21252), .ZN(
        n21255) );
  AOI21_X1 U23329 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(n21256), .A(n21255), 
        .ZN(n21259) );
  NAND2_X1 U23330 ( .A1(n21257), .A2(n21260), .ZN(n21262) );
  OAI211_X1 U23331 ( .C1(n21257), .C2(n21260), .A(n21423), .B(n21262), .ZN(
        n21258) );
  OAI211_X1 U23332 ( .C1(n21260), .C2(n21359), .A(n21259), .B(n21258), .ZN(
        P3_U2652) );
  AOI22_X1 U23333 ( .A1(n21424), .A2(P3_EBX_REG_20__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21404), .ZN(n21272) );
  NAND4_X1 U23334 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n21261), .A3(
        P3_REIP_REG_18__SCAN_IN), .A4(P3_REIP_REG_19__SCAN_IN), .ZN(n21288) );
  AOI21_X1 U23335 ( .B1(n21341), .B2(n21288), .A(n11262), .ZN(n21297) );
  INV_X1 U23336 ( .A(n21297), .ZN(n21281) );
  AOI211_X1 U23337 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n21262), .A(n21276), .B(
        n21397), .ZN(n21266) );
  NOR3_X1 U23338 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n21264), .A3(n21263), 
        .ZN(n21265) );
  AOI211_X1 U23339 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n21281), .A(n21266), 
        .B(n21265), .ZN(n21271) );
  NAND2_X1 U23340 ( .A1(n21399), .A2(n21267), .ZN(n21268) );
  NAND2_X1 U23341 ( .A1(n21268), .A2(n21269), .ZN(n21273) );
  OAI211_X1 U23342 ( .C1(n21269), .C2(n21268), .A(n11533), .B(n21273), .ZN(
        n21270) );
  NAND3_X1 U23343 ( .A1(n21272), .A2(n21271), .A3(n21270), .ZN(P3_U2651) );
  NAND2_X1 U23344 ( .A1(n21399), .A2(n21273), .ZN(n21274) );
  NAND2_X1 U23345 ( .A1(n21274), .A2(n21275), .ZN(n21285) );
  OAI211_X1 U23346 ( .C1(n21275), .C2(n21274), .A(n11533), .B(n21285), .ZN(
        n21278) );
  NAND2_X1 U23347 ( .A1(n21276), .A2(n21283), .ZN(n21284) );
  OAI211_X1 U23348 ( .C1(n21276), .C2(n21283), .A(n21423), .B(n21284), .ZN(
        n21277) );
  OAI211_X1 U23349 ( .C1(n21357), .C2(n21279), .A(n21278), .B(n21277), .ZN(
        n21280) );
  AOI21_X1 U23350 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n21281), .A(n21280), 
        .ZN(n21282) );
  OR3_X1 U23351 ( .A1(n21327), .A2(n21288), .A3(P3_REIP_REG_21__SCAN_IN), .ZN(
        n21296) );
  OAI211_X1 U23352 ( .C1(n21283), .C2(n21359), .A(n21282), .B(n21296), .ZN(
        P3_U2650) );
  NOR2_X1 U23353 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n21284), .ZN(n21303) );
  AOI211_X1 U23354 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n21284), .A(n21303), .B(
        n21397), .ZN(n21294) );
  NAND2_X1 U23355 ( .A1(n21399), .A2(n21285), .ZN(n21286) );
  NAND2_X1 U23356 ( .A1(n21286), .A2(n21287), .ZN(n21307) );
  OAI211_X1 U23357 ( .C1(n21287), .C2(n21286), .A(n11533), .B(n21307), .ZN(
        n21291) );
  NOR2_X1 U23358 ( .A1(n21289), .A2(n21288), .ZN(n21299) );
  NAND3_X1 U23359 ( .A1(n21341), .A2(n21299), .A3(n21298), .ZN(n21290) );
  OAI211_X1 U23360 ( .C1(n21357), .C2(n21292), .A(n21291), .B(n21290), .ZN(
        n21293) );
  AOI211_X1 U23361 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n21424), .A(n21294), .B(
        n21293), .ZN(n21295) );
  OAI221_X1 U23362 ( .B1(n21298), .B2(n21297), .C1(n21298), .C2(n21296), .A(
        n21295), .ZN(P3_U2649) );
  NAND2_X1 U23363 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n21299), .ZN(n21301) );
  NOR2_X1 U23364 ( .A1(n21302), .A2(n21301), .ZN(n21325) );
  INV_X1 U23365 ( .A(n21325), .ZN(n21300) );
  AOI21_X1 U23366 ( .B1(n21341), .B2(n21300), .A(n11262), .ZN(n21326) );
  AOI221_X1 U23367 ( .B1(n21419), .B2(n21302), .C1(n21301), .C2(n21302), .A(
        n21326), .ZN(n21306) );
  INV_X1 U23368 ( .A(n21303), .ZN(n21304) );
  NOR2_X1 U23369 ( .A1(n21304), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n21313) );
  AOI211_X1 U23370 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n21304), .A(n21313), .B(
        n21397), .ZN(n21305) );
  AOI211_X1 U23371 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n21424), .A(n21306), .B(
        n21305), .ZN(n21311) );
  NAND2_X1 U23372 ( .A1(n21399), .A2(n21307), .ZN(n21308) );
  NAND2_X1 U23373 ( .A1(n21308), .A2(n21309), .ZN(n21319) );
  OAI211_X1 U23374 ( .C1(n21309), .C2(n21308), .A(n11533), .B(n21319), .ZN(
        n21310) );
  OAI211_X1 U23375 ( .C1(n21357), .C2(n21312), .A(n21311), .B(n21310), .ZN(
        P3_U2648) );
  NOR2_X1 U23376 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21419), .ZN(n21318) );
  INV_X1 U23377 ( .A(n21313), .ZN(n21314) );
  NOR2_X1 U23378 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n21314), .ZN(n21332) );
  AOI211_X1 U23379 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n21314), .A(n21332), .B(
        n21397), .ZN(n21317) );
  INV_X1 U23380 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21315) );
  OAI22_X1 U23381 ( .A1(n21359), .A2(n21315), .B1(n11527), .B2(n21357), .ZN(
        n21316) );
  AOI211_X1 U23382 ( .C1(n21318), .C2(n21325), .A(n21317), .B(n21316), .ZN(
        n21323) );
  NAND2_X1 U23383 ( .A1(n21399), .A2(n21319), .ZN(n21320) );
  NAND2_X1 U23384 ( .A1(n21320), .A2(n21321), .ZN(n21333) );
  OAI211_X1 U23385 ( .C1(n21321), .C2(n21320), .A(n11533), .B(n21333), .ZN(
        n21322) );
  OAI211_X1 U23386 ( .C1(n21326), .C2(n21324), .A(n21323), .B(n21322), .ZN(
        P3_U2647) );
  NAND2_X1 U23387 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21325), .ZN(n21339) );
  NOR2_X1 U23388 ( .A1(n21419), .A2(n21339), .ZN(n21330) );
  OAI21_X1 U23389 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n21327), .A(n21326), 
        .ZN(n21329) );
  OAI22_X1 U23390 ( .A1(n21359), .A2(n21331), .B1(n11526), .B2(n21357), .ZN(
        n21328) );
  AOI221_X1 U23391 ( .B1(n21330), .B2(n21340), .C1(n21329), .C2(
        P3_REIP_REG_25__SCAN_IN), .A(n21328), .ZN(n21338) );
  NAND2_X1 U23392 ( .A1(n21332), .A2(n21331), .ZN(n21343) );
  OAI211_X1 U23393 ( .C1(n21332), .C2(n21331), .A(n21423), .B(n21343), .ZN(
        n21337) );
  NAND2_X1 U23394 ( .A1(n21399), .A2(n21333), .ZN(n21334) );
  NAND2_X1 U23395 ( .A1(n21334), .A2(n21335), .ZN(n21350) );
  OAI211_X1 U23396 ( .C1(n21335), .C2(n21334), .A(n11533), .B(n21350), .ZN(
        n21336) );
  NAND3_X1 U23397 ( .A1(n21338), .A2(n21337), .A3(n21336), .ZN(P3_U2646) );
  NOR2_X1 U23398 ( .A1(n21340), .A2(n21339), .ZN(n21348) );
  NAND2_X1 U23399 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n21348), .ZN(n21356) );
  AND2_X1 U23400 ( .A1(n21356), .A2(n21341), .ZN(n21349) );
  NOR2_X1 U23401 ( .A1(n11262), .A2(n21349), .ZN(n21381) );
  NOR2_X1 U23402 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n21343), .ZN(n21362) );
  AOI211_X1 U23403 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n21343), .A(n21362), .B(
        n21397), .ZN(n21347) );
  INV_X1 U23404 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n21345) );
  OAI22_X1 U23405 ( .A1(n21359), .A2(n21345), .B1(n21344), .B2(n21357), .ZN(
        n21346) );
  AOI211_X1 U23406 ( .C1(n21349), .C2(n21348), .A(n21347), .B(n21346), .ZN(
        n21354) );
  NAND2_X1 U23407 ( .A1(n21399), .A2(n21350), .ZN(n21351) );
  NAND2_X1 U23408 ( .A1(n21352), .A2(n21351), .ZN(n21363) );
  OAI211_X1 U23409 ( .C1(n21352), .C2(n21351), .A(n11533), .B(n21363), .ZN(
        n21353) );
  OAI211_X1 U23410 ( .C1(n21381), .C2(n21355), .A(n21354), .B(n21353), .ZN(
        P3_U2645) );
  INV_X1 U23411 ( .A(n21381), .ZN(n21371) );
  AND2_X1 U23412 ( .A1(n21380), .A2(n21395), .ZN(n21372) );
  INV_X1 U23413 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21361) );
  OAI22_X1 U23414 ( .A1(n21359), .A2(n21361), .B1(n21358), .B2(n21357), .ZN(
        n21360) );
  AOI211_X1 U23415 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n21371), .A(n21372), 
        .B(n21360), .ZN(n21368) );
  NAND2_X1 U23416 ( .A1(n21362), .A2(n21361), .ZN(n21369) );
  OAI211_X1 U23417 ( .C1(n21362), .C2(n21361), .A(n21423), .B(n21369), .ZN(
        n21367) );
  NAND2_X1 U23418 ( .A1(n21399), .A2(n21363), .ZN(n21364) );
  NAND2_X1 U23419 ( .A1(n21364), .A2(n21365), .ZN(n21373) );
  OAI211_X1 U23420 ( .C1(n21365), .C2(n21364), .A(n11533), .B(n21373), .ZN(
        n21366) );
  NAND3_X1 U23421 ( .A1(n21368), .A2(n21367), .A3(n21366), .ZN(P3_U2644) );
  AOI22_X1 U23422 ( .A1(n21424), .A2(P3_EBX_REG_28__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21404), .ZN(n21379) );
  NOR2_X1 U23423 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21369), .ZN(n21384) );
  AOI211_X1 U23424 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n21369), .A(n21384), .B(
        n21397), .ZN(n21370) );
  AOI221_X1 U23425 ( .B1(n21372), .B2(P3_REIP_REG_28__SCAN_IN), .C1(n21371), 
        .C2(P3_REIP_REG_28__SCAN_IN), .A(n21370), .ZN(n21378) );
  NAND2_X1 U23426 ( .A1(n21399), .A2(n21373), .ZN(n21374) );
  NAND2_X1 U23427 ( .A1(n21375), .A2(n21374), .ZN(n21387) );
  OAI211_X1 U23428 ( .C1(n21375), .C2(n21374), .A(n11533), .B(n21387), .ZN(
        n21377) );
  NAND3_X1 U23429 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21395), .A3(n21954), 
        .ZN(n21376) );
  NAND4_X1 U23430 ( .A1(n21379), .A2(n21378), .A3(n21377), .A4(n21376), .ZN(
        P3_U2643) );
  AOI22_X1 U23431 ( .A1(n21424), .A2(P3_EBX_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21404), .ZN(n21394) );
  NOR3_X1 U23432 ( .A1(n21954), .A2(n21390), .A3(n21380), .ZN(n21382) );
  OAI21_X1 U23433 ( .B1(n21382), .B2(n21419), .A(n21381), .ZN(n21407) );
  INV_X1 U23434 ( .A(n21384), .ZN(n21385) );
  NAND2_X1 U23435 ( .A1(n21384), .A2(n21383), .ZN(n21396) );
  NAND2_X1 U23436 ( .A1(n21423), .A2(n21396), .ZN(n21401) );
  AOI21_X1 U23437 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n21385), .A(n21401), .ZN(
        n21386) );
  AOI21_X1 U23438 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(n21407), .A(n21386), 
        .ZN(n21393) );
  NAND2_X1 U23439 ( .A1(n21399), .A2(n21387), .ZN(n21388) );
  NAND2_X1 U23440 ( .A1(n21388), .A2(n21389), .ZN(n21398) );
  OAI211_X1 U23441 ( .C1(n21389), .C2(n21388), .A(n11533), .B(n21398), .ZN(
        n21392) );
  NAND4_X1 U23442 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n21395), .A4(n21390), .ZN(n21391) );
  NAND4_X1 U23443 ( .A1(n21394), .A2(n21393), .A3(n21392), .A4(n21391), .ZN(
        P3_U2642) );
  NAND4_X1 U23444 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n21395), .ZN(n21411) );
  AOI22_X1 U23445 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21404), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n21407), .ZN(n21403) );
  NOR2_X1 U23446 ( .A1(n21397), .A2(n21396), .ZN(n21406) );
  NAND2_X1 U23447 ( .A1(n21399), .A2(n21398), .ZN(n21408) );
  OAI211_X1 U23448 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n21411), .A(n21403), 
        .B(n21402), .ZN(P3_U2641) );
  AOI22_X1 U23449 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n21424), .B1(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21404), .ZN(n21418) );
  AOI22_X1 U23450 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n21407), .B1(n21406), 
        .B2(n21405), .ZN(n21417) );
  NAND3_X1 U23451 ( .A1(n21410), .A2(n21409), .A3(n21408), .ZN(n21416) );
  INV_X1 U23452 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21413) );
  AOI221_X1 U23453 ( .B1(n21413), .B2(n21412), .C1(P3_REIP_REG_30__SCAN_IN), 
        .C2(P3_REIP_REG_31__SCAN_IN), .A(n21411), .ZN(n21414) );
  INV_X1 U23454 ( .A(n21414), .ZN(n21415) );
  NAND4_X1 U23455 ( .A1(n21418), .A2(n21417), .A3(n21416), .A4(n21415), .ZN(
        P3_U2640) );
  NAND2_X1 U23456 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21420), .ZN(
        n21427) );
  NAND2_X1 U23457 ( .A1(n21420), .A2(n21419), .ZN(n21422) );
  AOI22_X1 U23458 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n21422), .B1(n21421), 
        .B2(n21618), .ZN(n21426) );
  OAI21_X1 U23459 ( .B1(n21424), .B2(n21423), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n21425) );
  OAI211_X1 U23460 ( .C1(n21634), .C2(n21427), .A(n21426), .B(n21425), .ZN(
        P3_U2671) );
  NOR2_X1 U23461 ( .A1(n21641), .A2(n21428), .ZN(n21432) );
  NOR2_X1 U23462 ( .A1(n21605), .A2(n21433), .ZN(n21612) );
  NAND2_X1 U23463 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n21434) );
  NAND2_X1 U23464 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n21493) );
  NAND3_X1 U23465 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .ZN(n21491) );
  NAND3_X1 U23466 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .ZN(n21490) );
  INV_X1 U23467 ( .A(n21605), .ZN(n21438) );
  NAND2_X1 U23468 ( .A1(n21435), .A2(n21438), .ZN(n21614) );
  NAND2_X1 U23469 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n21486), .ZN(n21474) );
  NAND2_X1 U23470 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21598), .ZN(n21456) );
  NOR2_X1 U23471 ( .A1(n21450), .A2(n21451), .ZN(n21443) );
  INV_X1 U23472 ( .A(n21443), .ZN(n21436) );
  NOR2_X1 U23473 ( .A1(n21434), .A2(n21436), .ZN(n21586) );
  NOR2_X1 U23474 ( .A1(n21437), .A2(n21436), .ZN(n21446) );
  AOI21_X1 U23475 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n21600), .A(n21446), .ZN(
        n21441) );
  AND2_X1 U23476 ( .A1(n21439), .A2(n21438), .ZN(n21611) );
  OAI222_X1 U23477 ( .A1(n21487), .A2(n21442), .B1(n21586), .B2(n21441), .C1(
        n21603), .C2(n21440), .ZN(P3_U2722) );
  AOI21_X1 U23478 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n21600), .A(n21443), .ZN(
        n21445) );
  OAI222_X1 U23479 ( .A1(n21487), .A2(n21447), .B1(n21446), .B2(n21445), .C1(
        n21603), .C2(n21444), .ZN(P3_U2723) );
  NAND2_X1 U23480 ( .A1(n21600), .A2(n21451), .ZN(n21454) );
  AOI22_X1 U23481 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21612), .B1(n21611), .B2(
        n21448), .ZN(n21449) );
  OAI221_X1 U23482 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n21451), .C1(n21450), 
        .C2(n21454), .A(n21449), .ZN(P3_U2724) );
  INV_X1 U23483 ( .A(n21456), .ZN(n21458) );
  AOI21_X1 U23484 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n21458), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n21453) );
  OAI222_X1 U23485 ( .A1(n21487), .A2(n21455), .B1(n21454), .B2(n21453), .C1(
        n21603), .C2(n21452), .ZN(P3_U2725) );
  NOR2_X1 U23486 ( .A1(n21457), .A2(n21456), .ZN(n21461) );
  AOI21_X1 U23487 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n21600), .A(n21458), .ZN(
        n21460) );
  OAI222_X1 U23488 ( .A1(n21487), .A2(n21462), .B1(n21461), .B2(n21460), .C1(
        n21603), .C2(n21459), .ZN(P3_U2726) );
  AOI21_X1 U23489 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n21600), .A(n21468), .ZN(
        n21463) );
  OAI222_X1 U23490 ( .A1(n21487), .A2(n21464), .B1(n21598), .B2(n21463), .C1(
        n21603), .C2(n21661), .ZN(P3_U2728) );
  NOR2_X1 U23491 ( .A1(n21465), .A2(n21474), .ZN(n21477) );
  AOI22_X1 U23492 ( .A1(n21477), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n21600), .ZN(n21467) );
  OAI222_X1 U23493 ( .A1(n21469), .A2(n21487), .B1(n21468), .B2(n21467), .C1(
        n21603), .C2(n21466), .ZN(P3_U2729) );
  AND2_X1 U23494 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n21477), .ZN(n21472) );
  AOI21_X1 U23495 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n21600), .A(n21477), .ZN(
        n21471) );
  OAI222_X1 U23496 ( .A1(n21473), .A2(n21487), .B1(n21472), .B2(n21471), .C1(
        n21603), .C2(n21470), .ZN(P3_U2730) );
  INV_X1 U23497 ( .A(n21474), .ZN(n21481) );
  AOI21_X1 U23498 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n21600), .A(n21481), .ZN(
        n21476) );
  OAI222_X1 U23499 ( .A1(n21478), .A2(n21487), .B1(n21477), .B2(n21476), .C1(
        n21603), .C2(n21475), .ZN(P3_U2731) );
  AOI21_X1 U23500 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21600), .A(n21486), .ZN(
        n21480) );
  OAI222_X1 U23501 ( .A1(n21482), .A2(n21487), .B1(n21481), .B2(n21480), .C1(
        n21603), .C2(n21479), .ZN(P3_U2732) );
  NAND2_X1 U23502 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n21483) );
  NOR2_X1 U23503 ( .A1(n21483), .A2(n21614), .ZN(n21609) );
  AOI21_X1 U23504 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n21600), .A(n21609), .ZN(
        n21485) );
  OAI222_X1 U23505 ( .A1(n21488), .A2(n21487), .B1(n21486), .B2(n21485), .C1(
        n21603), .C2(n21484), .ZN(P3_U2733) );
  NOR2_X1 U23506 ( .A1(n21508), .A2(n21489), .ZN(n21509) );
  NAND2_X1 U23507 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n21496) );
  NOR3_X1 U23508 ( .A1(n21605), .A2(n21491), .A3(n21490), .ZN(n21492) );
  NAND3_X1 U23509 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(n21492), .ZN(n21599) );
  NAND4_X1 U23510 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(n21494), .ZN(n21593) );
  INV_X1 U23511 ( .A(n21527), .ZN(n21495) );
  NAND2_X1 U23512 ( .A1(n21509), .A2(n21522), .ZN(n21503) );
  NAND2_X1 U23513 ( .A1(n21600), .A2(n21503), .ZN(n21511) );
  OAI22_X1 U23514 ( .A1(n21499), .A2(n21603), .B1(n21498), .B2(n21573), .ZN(
        n21500) );
  AOI21_X1 U23515 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21580), .A(n21500), .ZN(
        n21501) );
  OAI221_X1 U23516 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21503), .C1(n21502), 
        .C2(n21511), .A(n21501), .ZN(P3_U2714) );
  NAND2_X1 U23517 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n21522), .ZN(n21516) );
  OAI22_X1 U23518 ( .A1(n21505), .A2(n21603), .B1(n21504), .B2(n21573), .ZN(
        n21506) );
  AOI21_X1 U23519 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n21580), .A(n21506), .ZN(
        n21507) );
  OAI221_X1 U23520 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n21516), .C1(n21508), 
        .C2(n21511), .A(n21507), .ZN(P3_U2715) );
  NAND4_X1 U23521 ( .A1(n21509), .A2(P3_EAX_REG_17__SCAN_IN), .A3(
        P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_21__SCAN_IN), .ZN(n21532) );
  NAND2_X1 U23522 ( .A1(n21527), .A2(n21531), .ZN(n21515) );
  AOI22_X1 U23523 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n21579), .B1(n21611), .B2(
        n21510), .ZN(n21514) );
  OAI21_X1 U23524 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21614), .A(n21511), .ZN(
        n21512) );
  AOI22_X1 U23525 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n21580), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n21512), .ZN(n21513) );
  OAI211_X1 U23526 ( .C1(n21532), .C2(n21515), .A(n21514), .B(n21513), .ZN(
        P3_U2713) );
  AOI22_X1 U23527 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21580), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21579), .ZN(n21518) );
  OAI211_X1 U23528 ( .C1(n21522), .C2(P3_EAX_REG_19__SCAN_IN), .A(n21600), .B(
        n21516), .ZN(n21517) );
  OAI211_X1 U23529 ( .C1(n21519), .C2(n21603), .A(n21518), .B(n21517), .ZN(
        P3_U2716) );
  AOI22_X1 U23530 ( .A1(n21527), .A2(P3_EAX_REG_17__SCAN_IN), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n21600), .ZN(n21521) );
  OAI22_X1 U23531 ( .A1(n21522), .A2(n21521), .B1(n21520), .B2(n21573), .ZN(
        n21523) );
  AOI21_X1 U23532 ( .B1(BUF2_REG_2__SCAN_IN), .B2(n21580), .A(n21523), .ZN(
        n21524) );
  OAI21_X1 U23533 ( .B1(n21525), .B2(n21603), .A(n21524), .ZN(P3_U2717) );
  AOI22_X1 U23534 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21580), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21579), .ZN(n21529) );
  NAND2_X1 U23535 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n21527), .ZN(n21526) );
  OAI211_X1 U23536 ( .C1(n21527), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21600), .B(
        n21526), .ZN(n21528) );
  OAI211_X1 U23537 ( .C1(n21530), .C2(n21603), .A(n21529), .B(n21528), .ZN(
        P3_U2718) );
  AOI22_X1 U23538 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21580), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n21579), .ZN(n21536) );
  NAND2_X1 U23539 ( .A1(n21575), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21574) );
  NAND2_X1 U23540 ( .A1(n21570), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n21569) );
  OAI211_X1 U23541 ( .C1(n21534), .C2(P3_EAX_REG_25__SCAN_IN), .A(n21600), .B(
        n21539), .ZN(n21535) );
  OAI211_X1 U23542 ( .C1(n21537), .C2(n21603), .A(n21536), .B(n21535), .ZN(
        P3_U2710) );
  AOI22_X1 U23543 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21580), .B1(n21611), .B2(
        n21538), .ZN(n21543) );
  AOI211_X1 U23544 ( .C1(n21540), .C2(n21539), .A(n21564), .B(n21591), .ZN(
        n21541) );
  INV_X1 U23545 ( .A(n21541), .ZN(n21542) );
  OAI211_X1 U23546 ( .C1(n21573), .C2(n21544), .A(n21543), .B(n21542), .ZN(
        P3_U2709) );
  NAND2_X1 U23547 ( .A1(n21564), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n21563) );
  NAND2_X1 U23548 ( .A1(n21557), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n21552) );
  NAND2_X1 U23549 ( .A1(n21548), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n21547) );
  NAND2_X1 U23550 ( .A1(n21547), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n21546) );
  NAND2_X1 U23551 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n21579), .ZN(n21545) );
  OAI221_X1 U23552 ( .B1(n21547), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n21546), 
        .C2(n21591), .A(n21545), .ZN(P3_U2704) );
  AOI22_X1 U23553 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21580), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n21579), .ZN(n21550) );
  OAI211_X1 U23554 ( .C1(n21548), .C2(P3_EAX_REG_30__SCAN_IN), .A(n21600), .B(
        n21547), .ZN(n21549) );
  OAI211_X1 U23555 ( .C1(n21551), .C2(n21603), .A(n21550), .B(n21549), .ZN(
        P3_U2705) );
  AOI22_X1 U23556 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21580), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n21579), .ZN(n21554) );
  OAI211_X1 U23557 ( .C1(n21557), .C2(P3_EAX_REG_29__SCAN_IN), .A(n21600), .B(
        n21552), .ZN(n21553) );
  OAI211_X1 U23558 ( .C1(n21555), .C2(n21603), .A(n21554), .B(n21553), .ZN(
        P3_U2706) );
  AOI22_X1 U23559 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21580), .B1(n21611), .B2(
        n21556), .ZN(n21561) );
  AOI211_X1 U23560 ( .C1(n21558), .C2(n21563), .A(n21557), .B(n21591), .ZN(
        n21559) );
  INV_X1 U23561 ( .A(n21559), .ZN(n21560) );
  OAI211_X1 U23562 ( .C1(n21573), .C2(n21562), .A(n21561), .B(n21560), .ZN(
        P3_U2707) );
  AOI22_X1 U23563 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21580), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n21579), .ZN(n21566) );
  OAI211_X1 U23564 ( .C1(n21564), .C2(P3_EAX_REG_27__SCAN_IN), .A(n21600), .B(
        n21563), .ZN(n21565) );
  OAI211_X1 U23565 ( .C1(n21567), .C2(n21603), .A(n21566), .B(n21565), .ZN(
        P3_U2708) );
  AOI22_X1 U23566 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21580), .B1(n21611), .B2(
        n21568), .ZN(n21572) );
  OAI211_X1 U23567 ( .C1(n21570), .C2(P3_EAX_REG_24__SCAN_IN), .A(n21600), .B(
        n21569), .ZN(n21571) );
  OAI211_X1 U23568 ( .C1(n21573), .C2(n17354), .A(n21572), .B(n21571), .ZN(
        P3_U2711) );
  AOI22_X1 U23569 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21580), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n21579), .ZN(n21577) );
  OAI211_X1 U23570 ( .C1(n21575), .C2(P3_EAX_REG_23__SCAN_IN), .A(n21600), .B(
        n21574), .ZN(n21576) );
  OAI211_X1 U23571 ( .C1(n21578), .C2(n21603), .A(n21577), .B(n21576), .ZN(
        P3_U2712) );
  AOI22_X1 U23572 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21580), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n21579), .ZN(n21583) );
  OAI211_X1 U23573 ( .C1(n21590), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21600), .B(
        n21581), .ZN(n21582) );
  OAI211_X1 U23574 ( .C1(n21584), .C2(n21603), .A(n21583), .B(n21582), .ZN(
        P3_U2719) );
  AOI22_X1 U23575 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21612), .B1(n21586), .B2(
        n21585), .ZN(n21588) );
  NAND3_X1 U23576 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n21600), .A3(n21593), 
        .ZN(n21587) );
  OAI211_X1 U23577 ( .C1(n21589), .C2(n21603), .A(n21588), .B(n21587), .ZN(
        P3_U2721) );
  AOI211_X1 U23578 ( .C1(n21593), .C2(n21592), .A(n21591), .B(n21590), .ZN(
        n21594) );
  AOI21_X1 U23579 ( .B1(n21612), .B2(BUF2_REG_15__SCAN_IN), .A(n21594), .ZN(
        n21595) );
  OAI21_X1 U23580 ( .B1(n21596), .B2(n21603), .A(n21595), .ZN(P3_U2720) );
  AOI22_X1 U23581 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21612), .B1(n21598), .B2(
        n21597), .ZN(n21602) );
  NAND3_X1 U23582 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21600), .A3(n21599), .ZN(
        n21601) );
  OAI211_X1 U23583 ( .C1(n21604), .C2(n21603), .A(n21602), .B(n21601), .ZN(
        P3_U2727) );
  NOR2_X1 U23584 ( .A1(n21605), .A2(n21615), .ZN(n21616) );
  OAI21_X1 U23585 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n21616), .A(n21600), .ZN(
        n21608) );
  AOI22_X1 U23586 ( .A1(n21612), .A2(BUF2_REG_1__SCAN_IN), .B1(n21611), .B2(
        n21606), .ZN(n21607) );
  OAI21_X1 U23587 ( .B1(n21609), .B2(n21608), .A(n21607), .ZN(P3_U2734) );
  AOI22_X1 U23588 ( .A1(n21612), .A2(BUF2_REG_0__SCAN_IN), .B1(n21611), .B2(
        n21610), .ZN(n21613) );
  OAI221_X1 U23589 ( .B1(n21616), .B2(n21615), .C1(n21616), .C2(n21614), .A(
        n21613), .ZN(P3_U2735) );
  AOI22_X1 U23590 ( .A1(n21639), .A2(n21618), .B1(n21617), .B2(n21636), .ZN(
        P3_U3290) );
  AOI22_X1 U23591 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n18945), .B2(n21691), .ZN(
        n21627) );
  INV_X1 U23592 ( .A(n21627), .ZN(n21620) );
  NOR2_X1 U23593 ( .A1(n21619), .A2(n21834), .ZN(n21626) );
  AOI222_X1 U23594 ( .A1(n21622), .A2(n21634), .B1(n21621), .B2(n22087), .C1(
        n21620), .C2(n21626), .ZN(n21623) );
  AOI22_X1 U23595 ( .A1(n21639), .A2(n21624), .B1(n21623), .B2(n21636), .ZN(
        P3_U3289) );
  AOI222_X1 U23596 ( .A1(n21628), .A2(n21634), .B1(n21627), .B2(n21626), .C1(
        n21625), .C2(n22087), .ZN(n21632) );
  INV_X1 U23597 ( .A(n21629), .ZN(n21630) );
  AOI22_X1 U23598 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21639), .B1(
        n22087), .B2(n21630), .ZN(n21631) );
  OAI21_X1 U23599 ( .B1(n21639), .B2(n21632), .A(n21631), .ZN(P3_U3288) );
  AOI22_X1 U23600 ( .A1(n22087), .A2(n21635), .B1(n21634), .B2(n21633), .ZN(
        n21637) );
  AOI22_X1 U23601 ( .A1(n21639), .A2(n21638), .B1(n21637), .B2(n21636), .ZN(
        P3_U3285) );
  INV_X1 U23602 ( .A(n21640), .ZN(n21673) );
  NAND2_X1 U23603 ( .A1(n21642), .A2(n21641), .ZN(n21644) );
  OAI22_X1 U23604 ( .A1(n21645), .A2(n21644), .B1(n21654), .B2(n21643), .ZN(
        n21651) );
  NOR3_X1 U23605 ( .A1(n21648), .A2(n21647), .A3(n21646), .ZN(n21650) );
  AOI211_X1 U23606 ( .C1(n21652), .C2(n21651), .A(n21650), .B(n21649), .ZN(
        n21655) );
  AOI221_X4 U23607 ( .B1(n21656), .B2(n21655), .C1(n21654), .C2(n21655), .A(
        n21653), .ZN(n22048) );
  AOI22_X1 U23608 ( .A1(n22011), .A2(n21766), .B1(n21964), .B2(n21769), .ZN(
        n21776) );
  NAND2_X1 U23609 ( .A1(n22013), .A2(n21658), .ZN(n22015) );
  AOI21_X1 U23610 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21704) );
  AND3_X1 U23611 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21738) );
  NAND2_X1 U23612 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21738), .ZN(
        n21747) );
  NOR2_X1 U23613 ( .A1(n21704), .A2(n21747), .ZN(n21743) );
  NAND3_X1 U23614 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21743), .ZN(n21767) );
  NOR2_X1 U23615 ( .A1(n21660), .A2(n21767), .ZN(n21843) );
  NOR2_X1 U23616 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n22071), .ZN(
        n21680) );
  NOR2_X1 U23617 ( .A1(n11250), .A2(n21680), .ZN(n21702) );
  NAND2_X1 U23618 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21727) );
  NOR2_X1 U23619 ( .A1(n21747), .A2(n21727), .ZN(n21744) );
  NAND2_X1 U23620 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21744), .ZN(
        n22070) );
  NOR2_X1 U23621 ( .A1(n21756), .A2(n22070), .ZN(n22058) );
  INV_X1 U23622 ( .A(n22058), .ZN(n21815) );
  NOR2_X1 U23623 ( .A1(n21660), .A2(n21815), .ZN(n21832) );
  AOI22_X1 U23624 ( .A1(n22016), .A2(n21843), .B1(n21702), .B2(n21832), .ZN(
        n21883) );
  OAI21_X1 U23625 ( .B1(n21776), .B2(n21660), .A(n21883), .ZN(n21831) );
  NAND2_X1 U23626 ( .A1(n22048), .A2(n21831), .ZN(n21975) );
  NAND2_X1 U23627 ( .A1(n22048), .A2(n21932), .ZN(n21707) );
  AOI21_X1 U23628 ( .B1(n21832), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n22059), .ZN(n21662) );
  INV_X1 U23629 ( .A(n21662), .ZN(n21663) );
  OAI21_X1 U23630 ( .B1(n21843), .B2(n21894), .A(n21663), .ZN(n21983) );
  NOR2_X1 U23631 ( .A1(n22016), .A2(n22071), .ZN(n22060) );
  OAI22_X1 U23632 ( .A1(n21664), .A2(n22060), .B1(n21959), .B2(n21985), .ZN(
        n21665) );
  AOI211_X1 U23633 ( .C1(n22011), .C2(n21957), .A(n21983), .B(n21665), .ZN(
        n21835) );
  NAND2_X1 U23634 ( .A1(n21834), .A2(n21892), .ZN(n22012) );
  OAI211_X1 U23635 ( .C1(n21832), .C2(n22068), .A(n22048), .B(n22012), .ZN(
        n21984) );
  AOI21_X1 U23636 ( .B1(n21666), .B2(n21892), .A(n21984), .ZN(n21668) );
  AOI211_X1 U23637 ( .C1(n21835), .C2(n21668), .A(n22073), .B(n21667), .ZN(
        n21669) );
  AOI211_X1 U23638 ( .C1(n22079), .C2(n21671), .A(n21670), .B(n21669), .ZN(
        n21672) );
  OAI21_X1 U23639 ( .B1(n21673), .B2(n21975), .A(n21672), .ZN(P3_U2841) );
  NOR2_X1 U23640 ( .A1(n21947), .A2(n21985), .ZN(n21858) );
  INV_X1 U23641 ( .A(n21707), .ZN(n21751) );
  NAND2_X1 U23642 ( .A1(n22068), .A2(n21894), .ZN(n21897) );
  INV_X1 U23643 ( .A(n21897), .ZN(n22000) );
  AOI221_X1 U23644 ( .B1(n22059), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n22000), .C2(n21834), .A(n21947), .ZN(n21674) );
  AOI221_X1 U23645 ( .B1(n21858), .B2(n21676), .C1(n21751), .C2(n21675), .A(
        n21674), .ZN(n21678) );
  NAND2_X1 U23646 ( .A1(n21869), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n21677) );
  OAI211_X1 U23647 ( .C1(n21970), .C2(n21834), .A(n21678), .B(n21677), .ZN(
        P3_U2862) );
  AOI22_X1 U23648 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21962), .B1(
        n21751), .B2(n21679), .ZN(n21686) );
  INV_X1 U23649 ( .A(n21979), .ZN(n22038) );
  NOR3_X1 U23650 ( .A1(n22038), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n21680), .ZN(n21684) );
  NAND2_X1 U23651 ( .A1(n21834), .A2(n21897), .ZN(n21681) );
  OAI22_X1 U23652 ( .A1(n21682), .A2(n21985), .B1(n21691), .B2(n21681), .ZN(
        n21683) );
  OAI21_X1 U23653 ( .B1(n21684), .B2(n21683), .A(n22048), .ZN(n21685) );
  OAI211_X1 U23654 ( .C1(n21687), .C2(n22049), .A(n21686), .B(n21685), .ZN(
        P3_U2861) );
  AOI21_X1 U23655 ( .B1(n21751), .B2(n21689), .A(n21688), .ZN(n21698) );
  NAND2_X1 U23656 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21690) );
  INV_X1 U23657 ( .A(n21704), .ZN(n21700) );
  AOI221_X1 U23658 ( .B1(n21690), .B2(n21700), .C1(n21699), .C2(n21700), .A(
        n21894), .ZN(n21696) );
  INV_X1 U23659 ( .A(n22012), .ZN(n21746) );
  INV_X1 U23660 ( .A(n11250), .ZN(n22021) );
  OAI211_X1 U23661 ( .C1(n21746), .C2(n21691), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n22021), .ZN(n21693) );
  NAND3_X1 U23662 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21702), .A3(
        n21699), .ZN(n21692) );
  OAI211_X1 U23663 ( .C1(n21694), .C2(n21985), .A(n21693), .B(n21692), .ZN(
        n21695) );
  OAI21_X1 U23664 ( .B1(n21696), .B2(n21695), .A(n22048), .ZN(n21697) );
  OAI211_X1 U23665 ( .C1(n21970), .C2(n21699), .A(n21698), .B(n21697), .ZN(
        P3_U2860) );
  NOR2_X1 U23666 ( .A1(n21894), .A2(n21700), .ZN(n21726) );
  AOI211_X1 U23667 ( .C1(n22021), .C2(n21727), .A(n21746), .B(n21726), .ZN(
        n21701) );
  AOI21_X1 U23668 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21701), .A(
        n21947), .ZN(n21718) );
  INV_X1 U23669 ( .A(n21702), .ZN(n21703) );
  OAI22_X1 U23670 ( .A1(n21894), .A2(n21704), .B1(n21703), .B2(n21727), .ZN(
        n21711) );
  INV_X1 U23671 ( .A(n21858), .ZN(n21742) );
  OAI22_X1 U23672 ( .A1(n21707), .A2(n21706), .B1(n21742), .B2(n21705), .ZN(
        n21708) );
  AOI221_X1 U23673 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21718), .C1(
        n21711), .C2(n21718), .A(n21708), .ZN(n21710) );
  OAI211_X1 U23674 ( .C1(n21970), .C2(n21712), .A(n21710), .B(n21709), .ZN(
        P3_U2859) );
  INV_X1 U23675 ( .A(n21711), .ZN(n21748) );
  NOR4_X1 U23676 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21748), .A3(
        n21947), .A4(n21712), .ZN(n21716) );
  AOI22_X1 U23677 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21962), .B1(
        n21751), .B2(n21713), .ZN(n21714) );
  INV_X1 U23678 ( .A(n21714), .ZN(n21715) );
  NOR3_X1 U23679 ( .A1(n21717), .A2(n21716), .A3(n21715), .ZN(n21720) );
  NAND3_X1 U23680 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21718), .A3(
        n21979), .ZN(n21719) );
  OAI211_X1 U23681 ( .C1(n21721), .C2(n21742), .A(n21720), .B(n21719), .ZN(
        P3_U2858) );
  INV_X1 U23682 ( .A(n21722), .ZN(n21724) );
  AOI21_X1 U23683 ( .B1(n21724), .B2(n21858), .A(n21723), .ZN(n21734) );
  NAND2_X1 U23684 ( .A1(n22048), .A2(n22012), .ZN(n21725) );
  AOI211_X1 U23685 ( .C1(n22021), .C2(n21727), .A(n21726), .B(n21725), .ZN(
        n21728) );
  AOI221_X1 U23686 ( .B1(n22038), .B2(n21728), .C1(n21738), .C2(n21728), .A(
        n22073), .ZN(n21735) );
  AOI22_X1 U23687 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21735), .B1(
        n21751), .B2(n21729), .ZN(n21733) );
  NOR2_X1 U23688 ( .A1(n21748), .A2(n21947), .ZN(n21731) );
  NAND4_X1 U23689 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n21731), .A4(n21730), .ZN(
        n21732) );
  NAND3_X1 U23690 ( .A1(n21734), .A2(n21733), .A3(n21732), .ZN(P3_U2857) );
  AOI22_X1 U23691 ( .A1(n22057), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21735), .ZN(n21740) );
  NOR3_X1 U23692 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21748), .A3(
        n21947), .ZN(n21737) );
  AOI22_X1 U23693 ( .A1(n21738), .A2(n21737), .B1(n21751), .B2(n21736), .ZN(
        n21739) );
  OAI211_X1 U23694 ( .C1(n21742), .C2(n21741), .A(n21740), .B(n21739), .ZN(
        P3_U2856) );
  OAI22_X1 U23695 ( .A1(n11250), .A2(n21744), .B1(n21743), .B2(n21894), .ZN(
        n21745) );
  NOR3_X1 U23696 ( .A1(n21746), .A2(n21755), .A3(n21745), .ZN(n21757) );
  NOR2_X1 U23697 ( .A1(n21748), .A2(n21747), .ZN(n21775) );
  OAI21_X1 U23698 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21775), .A(
        n22048), .ZN(n21754) );
  AOI22_X1 U23699 ( .A1(n22073), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21962), .ZN(n21753) );
  AOI22_X1 U23700 ( .A1(n21751), .A2(n21750), .B1(n21858), .B2(n21749), .ZN(
        n21752) );
  OAI211_X1 U23701 ( .C1(n21757), .C2(n21754), .A(n21753), .B(n21752), .ZN(
        P3_U2855) );
  NOR2_X1 U23702 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21755), .ZN(
        n21761) );
  NOR3_X1 U23703 ( .A1(n22038), .A2(n21757), .A3(n21756), .ZN(n21760) );
  OAI22_X1 U23704 ( .A1(n21762), .A2(n21987), .B1(n21985), .B2(n21758), .ZN(
        n21759) );
  AOI211_X1 U23705 ( .C1(n21775), .C2(n21761), .A(n21760), .B(n21759), .ZN(
        n21765) );
  AOI22_X1 U23706 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21962), .B1(
        n22079), .B2(n21762), .ZN(n21764) );
  OAI211_X1 U23707 ( .C1(n21765), .C2(n21947), .A(n21764), .B(n21763), .ZN(
        P3_U2854) );
  NOR2_X1 U23708 ( .A1(n21964), .A2(n22011), .ZN(n22020) );
  INV_X1 U23709 ( .A(n21766), .ZN(n22010) );
  NAND2_X1 U23710 ( .A1(n22010), .A2(n22011), .ZN(n21768) );
  AND2_X1 U23711 ( .A1(n22016), .A2(n21767), .ZN(n21813) );
  NOR2_X1 U23712 ( .A1(n21813), .A2(n21947), .ZN(n22018) );
  OAI211_X1 U23713 ( .C1(n21769), .C2(n21985), .A(n21768), .B(n22018), .ZN(
        n21770) );
  INV_X1 U23714 ( .A(n21770), .ZN(n22075) );
  NOR2_X1 U23715 ( .A1(n21834), .A2(n21815), .ZN(n22066) );
  AOI21_X1 U23716 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n22066), .A(
        n22068), .ZN(n21771) );
  INV_X1 U23717 ( .A(n21771), .ZN(n21772) );
  OAI211_X1 U23718 ( .C1(n21779), .C2(n22020), .A(n22075), .B(n21772), .ZN(
        n22062) );
  NOR2_X1 U23719 ( .A1(n21790), .A2(n21894), .ZN(n21801) );
  NAND3_X1 U23720 ( .A1(n21779), .A2(n22058), .A3(n21894), .ZN(n21773) );
  OAI21_X1 U23721 ( .B1(n21801), .B2(n22071), .A(n21773), .ZN(n21786) );
  OAI21_X1 U23722 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n22068), .A(
        n21786), .ZN(n21774) );
  OAI21_X1 U23723 ( .B1(n22062), .B2(n21774), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21782) );
  NAND3_X1 U23724 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21775), .ZN(n21817) );
  NAND2_X1 U23725 ( .A1(n21776), .A2(n21817), .ZN(n21789) );
  NAND2_X1 U23726 ( .A1(n22048), .A2(n21789), .ZN(n22081) );
  NOR2_X1 U23727 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n22081), .ZN(
        n21778) );
  AOI22_X1 U23728 ( .A1(n21779), .A2(n21778), .B1(n22079), .B2(n21777), .ZN(
        n21780) );
  OAI221_X1 U23729 ( .B1(n22057), .B2(n21782), .C1(n22049), .C2(n21781), .A(
        n21780), .ZN(P3_U2851) );
  AOI21_X1 U23730 ( .B1(n21783), .B2(n22066), .A(n22068), .ZN(n21796) );
  AOI21_X1 U23731 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n22059), .ZN(n21784) );
  OAI211_X1 U23732 ( .C1(n21788), .C2(n21987), .A(n21787), .B(n21786), .ZN(
        n22051) );
  NOR3_X1 U23733 ( .A1(n21796), .A2(n22051), .A3(n21797), .ZN(n21795) );
  OAI221_X1 U23734 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21790), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n21789), .A(n22048), .ZN(
        n21794) );
  AOI22_X1 U23735 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21962), .B1(
        n22079), .B2(n21791), .ZN(n21793) );
  OAI211_X1 U23736 ( .C1(n21795), .C2(n21794), .A(n21793), .B(n21792), .ZN(
        P3_U2850) );
  OR2_X1 U23737 ( .A1(n21798), .A2(n21817), .ZN(n21806) );
  AOI21_X1 U23738 ( .B1(n22016), .B2(n21797), .A(n21796), .ZN(n22047) );
  OAI21_X1 U23739 ( .B1(n21798), .B2(n21815), .A(n22071), .ZN(n21799) );
  OAI211_X1 U23740 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n22000), .A(
        n22047), .B(n21799), .ZN(n21800) );
  NOR3_X1 U23741 ( .A1(n21813), .A2(n21801), .A3(n21800), .ZN(n21805) );
  AOI22_X1 U23742 ( .A1(n22011), .A2(n21803), .B1(n21964), .B2(n21802), .ZN(
        n21804) );
  OAI221_X1 U23743 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21806), 
        .C1(n21811), .C2(n21805), .A(n21804), .ZN(n21808) );
  AOI22_X1 U23744 ( .A1(n22048), .A2(n21808), .B1(n22079), .B2(n21807), .ZN(
        n21810) );
  OAI211_X1 U23745 ( .C1(n21970), .C2(n21811), .A(n21810), .B(n21809), .ZN(
        P3_U2848) );
  NOR2_X1 U23746 ( .A1(n21812), .A2(n21987), .ZN(n21819) );
  AOI22_X1 U23747 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n22068), .B1(
        n22013), .B2(n22066), .ZN(n21814) );
  AOI211_X1 U23748 ( .C1(n22071), .C2(n21815), .A(n21814), .B(n21813), .ZN(
        n21818) );
  OAI211_X1 U23749 ( .C1(n21822), .C2(n22060), .A(n22037), .B(n21818), .ZN(
        n21816) );
  NAND2_X1 U23750 ( .A1(n22049), .A2(n21816), .ZN(n22036) );
  NOR2_X1 U23751 ( .A1(n21818), .A2(n21817), .ZN(n21821) );
  AOI22_X1 U23752 ( .A1(n21822), .A2(n21821), .B1(n21820), .B2(n21819), .ZN(
        n21823) );
  OAI21_X1 U23753 ( .B1(n21985), .B2(n21824), .A(n21823), .ZN(n21826) );
  AOI22_X1 U23754 ( .A1(n22048), .A2(n21826), .B1(n22079), .B2(n21825), .ZN(
        n21828) );
  OAI211_X1 U23755 ( .C1(n22036), .C2(n21829), .A(n21828), .B(n21827), .ZN(
        P3_U2847) );
  AOI22_X1 U23756 ( .A1(n21869), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n22079), 
        .B2(n21830), .ZN(n21840) );
  NAND2_X1 U23757 ( .A1(n21842), .A2(n21831), .ZN(n21876) );
  INV_X1 U23758 ( .A(n21876), .ZN(n21838) );
  NAND2_X1 U23759 ( .A1(n21832), .A2(n21842), .ZN(n21890) );
  NOR2_X1 U23760 ( .A1(n21856), .A2(n21890), .ZN(n21845) );
  INV_X1 U23761 ( .A(n21845), .ZN(n21833) );
  OAI21_X1 U23762 ( .B1(n21834), .B2(n21833), .A(n21892), .ZN(n21836) );
  OAI211_X1 U23763 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n22060), .A(
        n21836), .B(n21835), .ZN(n21837) );
  OAI221_X1 U23764 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21838), 
        .C1(n21856), .C2(n21837), .A(n22048), .ZN(n21839) );
  OAI211_X1 U23765 ( .C1(n21970), .C2(n21856), .A(n21840), .B(n21839), .ZN(
        P3_U2840) );
  NOR2_X1 U23766 ( .A1(n21883), .A2(n21882), .ZN(n21850) );
  NOR2_X1 U23767 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21841), .ZN(
        n21849) );
  NAND2_X1 U23768 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21846) );
  NAND2_X1 U23769 ( .A1(n21843), .A2(n21842), .ZN(n21870) );
  INV_X1 U23770 ( .A(n21870), .ZN(n21844) );
  AOI21_X1 U23771 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21844), .A(
        n21894), .ZN(n21968) );
  OAI221_X1 U23772 ( .B1(n21845), .B2(n22068), .C1(n21845), .C2(n22059), .A(
        n22012), .ZN(n21961) );
  AOI211_X1 U23773 ( .C1(n21979), .C2(n21846), .A(n21968), .B(n21961), .ZN(
        n21863) );
  OAI22_X1 U23774 ( .A1(n21847), .A2(n21987), .B1(n21863), .B2(n21861), .ZN(
        n21848) );
  AOI21_X1 U23775 ( .B1(n21850), .B2(n21849), .A(n21848), .ZN(n21855) );
  AOI22_X1 U23776 ( .A1(n22057), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21962), .ZN(n21854) );
  AOI22_X1 U23777 ( .A1(n22079), .A2(n21852), .B1(n21858), .B2(n21851), .ZN(
        n21853) );
  OAI211_X1 U23778 ( .C1(n21855), .C2(n21947), .A(n21854), .B(n21853), .ZN(
        P3_U2837) );
  AND3_X1 U23779 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21871) );
  NOR2_X1 U23780 ( .A1(n21876), .A2(n21856), .ZN(n21971) );
  AOI21_X1 U23781 ( .B1(n21871), .B2(n21971), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21868) );
  AND2_X1 U23782 ( .A1(n21858), .A2(n21857), .ZN(n21878) );
  AND2_X1 U23783 ( .A1(n22011), .A2(n21873), .ZN(n21860) );
  AOI211_X1 U23784 ( .C1(n21979), .C2(n21861), .A(n21860), .B(n21859), .ZN(
        n21862) );
  AOI21_X1 U23785 ( .B1(n21863), .B2(n21862), .A(n21947), .ZN(n21864) );
  AOI211_X1 U23786 ( .C1(n21962), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n21878), .B(n21864), .ZN(n21867) );
  AOI22_X1 U23787 ( .A1(n22057), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n22079), 
        .B2(n21865), .ZN(n21866) );
  OAI21_X1 U23788 ( .B1(n21868), .B2(n21867), .A(n21866), .ZN(P3_U2836) );
  NAND2_X1 U23789 ( .A1(n21869), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21880) );
  OAI21_X1 U23790 ( .B1(n21891), .B2(n21870), .A(n22016), .ZN(n21906) );
  AND2_X1 U23791 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21906), .ZN(
        n21895) );
  OAI221_X1 U23792 ( .B1(n11250), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n11250), .C2(n21871), .A(n21895), .ZN(n21872) );
  AOI211_X1 U23793 ( .C1(n22011), .C2(n21873), .A(n21961), .B(n21872), .ZN(
        n21875) );
  OAI22_X1 U23794 ( .A1(n21875), .A2(n21947), .B1(n21874), .B2(n21970), .ZN(
        n21877) );
  NOR2_X1 U23795 ( .A1(n21876), .A2(n21891), .ZN(n21944) );
  OAI22_X1 U23796 ( .A1(n21878), .A2(n21877), .B1(n21944), .B2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21879) );
  OAI211_X1 U23797 ( .C1(n21881), .C2(n22044), .A(n21880), .B(n21879), .ZN(
        P3_U2835) );
  NOR3_X1 U23798 ( .A1(n21883), .A2(n21882), .A3(n21888), .ZN(n21919) );
  AOI21_X1 U23799 ( .B1(n21885), .B2(n22011), .A(n21919), .ZN(n21884) );
  OAI21_X1 U23800 ( .B1(n21985), .B2(n21940), .A(n21884), .ZN(n21910) );
  NAND3_X1 U23801 ( .A1(n21898), .A2(n22048), .A3(n21910), .ZN(n21904) );
  NAND2_X1 U23802 ( .A1(n21885), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21887) );
  AOI22_X1 U23803 ( .A1(n22011), .A2(n21887), .B1(n21964), .B2(n21886), .ZN(
        n21913) );
  OAI21_X1 U23804 ( .B1(n21888), .B2(n21890), .A(n22071), .ZN(n21889) );
  INV_X1 U23805 ( .A(n21889), .ZN(n21907) );
  NOR2_X1 U23806 ( .A1(n21891), .A2(n21890), .ZN(n21937) );
  NAND3_X1 U23807 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21937), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21893) );
  NAND2_X1 U23808 ( .A1(n21893), .A2(n21892), .ZN(n21905) );
  OAI211_X1 U23809 ( .C1(n21895), .C2(n21894), .A(n22048), .B(n21905), .ZN(
        n21896) );
  AOI211_X1 U23810 ( .C1(n21934), .C2(n21897), .A(n21907), .B(n21896), .ZN(
        n21899) );
  AOI211_X1 U23811 ( .C1(n21913), .C2(n21899), .A(n22073), .B(n21898), .ZN(
        n21900) );
  AOI211_X1 U23812 ( .C1(n22079), .C2(n21902), .A(n21901), .B(n21900), .ZN(
        n21903) );
  NAND2_X1 U23813 ( .A1(n21904), .A2(n21903), .ZN(P3_U2833) );
  NAND2_X1 U23814 ( .A1(n21906), .A2(n21905), .ZN(n21938) );
  AOI211_X1 U23815 ( .C1(n21979), .C2(n21908), .A(n21907), .B(n21938), .ZN(
        n21909) );
  NAND2_X1 U23816 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n21909), .ZN(
        n21922) );
  INV_X1 U23817 ( .A(n21922), .ZN(n21912) );
  AOI21_X1 U23818 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21910), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21911) );
  AOI211_X1 U23819 ( .C1(n21913), .C2(n21912), .A(n21947), .B(n21911), .ZN(
        n21914) );
  AOI21_X1 U23820 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n21962), .A(
        n21914), .ZN(n21916) );
  OAI211_X1 U23821 ( .C1(n21917), .C2(n22044), .A(n21916), .B(n21915), .ZN(
        P3_U2832) );
  NOR2_X1 U23822 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21918), .ZN(
        n21920) );
  AOI22_X1 U23823 ( .A1(n21964), .A2(n21921), .B1(n21920), .B2(n21919), .ZN(
        n21924) );
  NAND3_X1 U23824 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21979), .A3(
        n21922), .ZN(n21923) );
  OAI211_X1 U23825 ( .C1(n21925), .C2(n21987), .A(n21924), .B(n21923), .ZN(
        n21927) );
  AOI22_X1 U23826 ( .A1(n22048), .A2(n21927), .B1(n22079), .B2(n21926), .ZN(
        n21930) );
  INV_X1 U23827 ( .A(n21928), .ZN(n21929) );
  OAI211_X1 U23828 ( .C1(n18945), .C2(n21970), .A(n21930), .B(n21929), .ZN(
        P3_U2831) );
  OAI221_X1 U23829 ( .B1(n21935), .B2(n21934), .C1(n21945), .C2(n21934), .A(
        n21933), .ZN(n21936) );
  INV_X1 U23830 ( .A(n21936), .ZN(n21950) );
  INV_X1 U23831 ( .A(n21937), .ZN(n21939) );
  AOI211_X1 U23832 ( .C1(n22071), .C2(n21939), .A(n21962), .B(n21938), .ZN(
        n21943) );
  AOI22_X1 U23833 ( .A1(n22011), .A2(n21941), .B1(n21964), .B2(n21940), .ZN(
        n21942) );
  OAI211_X1 U23834 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n22060), .A(
        n21943), .B(n21942), .ZN(n21949) );
  OAI22_X1 U23835 ( .A1(n21950), .A2(n21949), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21948), .ZN(n21955) );
  OR3_X1 U23836 ( .A1(n21952), .A2(n22044), .A3(n21951), .ZN(n21953) );
  OAI221_X1 U23837 ( .B1(n22073), .B2(n21955), .C1(n22049), .C2(n21954), .A(
        n21953), .ZN(P3_U2834) );
  INV_X1 U23838 ( .A(n21956), .ZN(n21973) );
  NOR2_X1 U23839 ( .A1(n21958), .A2(n21957), .ZN(n21966) );
  NAND2_X1 U23840 ( .A1(n21960), .A2(n21959), .ZN(n21963) );
  OAI21_X1 U23841 ( .B1(n21966), .B2(n21987), .A(n21965), .ZN(n21978) );
  NOR3_X1 U23842 ( .A1(n21968), .A2(n21967), .A3(n21978), .ZN(n21969) );
  NOR2_X1 U23843 ( .A1(n21969), .A2(n22073), .ZN(n21977) );
  OAI221_X1 U23844 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21971), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n21970), .A(n21977), .ZN(
        n21972) );
  OAI211_X1 U23845 ( .C1(n21974), .C2(n22044), .A(n21973), .B(n21972), .ZN(
        P3_U2839) );
  INV_X1 U23846 ( .A(n21975), .ZN(n22004) );
  AOI22_X1 U23847 ( .A1(n22057), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n22004), 
        .B2(n21976), .ZN(n21981) );
  OAI211_X1 U23848 ( .C1(n21979), .C2(n21978), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21977), .ZN(n21980) );
  OAI211_X1 U23849 ( .C1(n21982), .C2(n22044), .A(n21981), .B(n21980), .ZN(
        P3_U2838) );
  INV_X1 U23850 ( .A(n21983), .ZN(n21992) );
  INV_X1 U23851 ( .A(n21984), .ZN(n21991) );
  OAI22_X1 U23852 ( .A1(n21988), .A2(n21987), .B1(n21986), .B2(n21985), .ZN(
        n21989) );
  INV_X1 U23853 ( .A(n21989), .ZN(n21990) );
  NAND3_X1 U23854 ( .A1(n21992), .A2(n21991), .A3(n21990), .ZN(n21993) );
  NAND2_X1 U23855 ( .A1(n22049), .A2(n21993), .ZN(n21999) );
  NAND2_X1 U23856 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21999), .ZN(
        n22001) );
  OAI21_X1 U23857 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n22004), .A(
        n22001), .ZN(n21995) );
  OAI211_X1 U23858 ( .C1(n21996), .C2(n22044), .A(n21995), .B(n21994), .ZN(
        P3_U2843) );
  INV_X1 U23859 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21997) );
  AOI221_X1 U23860 ( .B1(n22000), .B2(n21999), .C1(n21998), .C2(n21999), .A(
        n21997), .ZN(n22002) );
  AOI22_X1 U23861 ( .A1(n22004), .A2(n22003), .B1(n22002), .B2(n22001), .ZN(
        n22006) );
  OAI211_X1 U23862 ( .C1(n22044), .C2(n22007), .A(n22006), .B(n22005), .ZN(
        P3_U2842) );
  AOI211_X1 U23863 ( .C1(n22011), .C2(n22010), .A(n22009), .B(n22008), .ZN(
        n22019) );
  NAND4_X1 U23864 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n22013), .A3(
        n22058), .A4(n22012), .ZN(n22014) );
  AOI22_X1 U23865 ( .A1(n22016), .A2(n22015), .B1(n22021), .B2(n22014), .ZN(
        n22017) );
  OAI211_X1 U23866 ( .C1(n22020), .C2(n22019), .A(n22018), .B(n22017), .ZN(
        n22031) );
  OAI221_X1 U23867 ( .B1(n22031), .B2(n22021), .C1(n22031), .C2(n22028), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n22027) );
  NOR2_X1 U23868 ( .A1(n22022), .A2(n22081), .ZN(n22040) );
  AOI22_X1 U23869 ( .A1(n22079), .A2(n22024), .B1(n22040), .B2(n22023), .ZN(
        n22025) );
  OAI221_X1 U23870 ( .B1(n22057), .B2(n22027), .C1(n22049), .C2(n22026), .A(
        n22025), .ZN(P3_U2844) );
  NAND2_X1 U23871 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n22028), .ZN(
        n22035) );
  INV_X1 U23872 ( .A(n22040), .ZN(n22034) );
  AOI21_X1 U23873 ( .B1(n22079), .B2(n22030), .A(n22029), .ZN(n22033) );
  NAND3_X1 U23874 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n22049), .A3(
        n22031), .ZN(n22032) );
  OAI211_X1 U23875 ( .C1(n22035), .C2(n22034), .A(n22033), .B(n22032), .ZN(
        P3_U2845) );
  AOI21_X1 U23876 ( .B1(n22038), .B2(n22037), .A(n22036), .ZN(n22041) );
  AOI22_X1 U23877 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n22041), .B1(
        n22040), .B2(n22039), .ZN(n22043) );
  OAI211_X1 U23878 ( .C1(n22045), .C2(n22044), .A(n22043), .B(n22042), .ZN(
        P3_U2846) );
  AOI22_X1 U23879 ( .A1(n22057), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n22079), 
        .B2(n22046), .ZN(n22053) );
  NAND2_X1 U23880 ( .A1(n22048), .A2(n22047), .ZN(n22050) );
  OAI211_X1 U23881 ( .C1(n22051), .C2(n22050), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n22049), .ZN(n22052) );
  OAI211_X1 U23882 ( .C1(n22054), .C2(n22081), .A(n22053), .B(n22052), .ZN(
        P3_U2849) );
  NAND2_X1 U23883 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n22055), .ZN(
        n22065) );
  AOI22_X1 U23884 ( .A1(n22057), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n22079), 
        .B2(n22056), .ZN(n22064) );
  OAI22_X1 U23885 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n22060), .B1(
        n22059), .B2(n22058), .ZN(n22061) );
  OAI211_X1 U23886 ( .C1(n22062), .C2(n22061), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n22049), .ZN(n22063) );
  OAI211_X1 U23887 ( .C1(n22065), .C2(n22081), .A(n22064), .B(n22063), .ZN(
        P3_U2852) );
  AOI211_X1 U23888 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n22068), .A(
        n11250), .B(n22066), .ZN(n22069) );
  AOI21_X1 U23889 ( .B1(n22071), .B2(n22070), .A(n22069), .ZN(n22074) );
  AOI211_X1 U23890 ( .C1(n22075), .C2(n22074), .A(n22073), .B(n22072), .ZN(
        n22077) );
  AOI211_X1 U23891 ( .C1(n22079), .C2(n22078), .A(n22077), .B(n22076), .ZN(
        n22080) );
  OAI21_X1 U23892 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n22081), .A(
        n22080), .ZN(P3_U2853) );
  NOR2_X1 U23893 ( .A1(n22082), .A2(n22095), .ZN(n22085) );
  OAI21_X1 U23894 ( .B1(n22085), .B2(n22084), .A(n22083), .ZN(P3_U3282) );
  AOI211_X1 U23895 ( .C1(n22088), .C2(n22087), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n22086), .ZN(n22089) );
  AOI211_X1 U23896 ( .C1(n22097), .C2(n22091), .A(n22090), .B(n22089), .ZN(
        n22092) );
  OAI221_X1 U23897 ( .B1(n22095), .B2(n22094), .C1(n22095), .C2(n22093), .A(
        n22092), .ZN(P3_U2996) );
  NAND2_X1 U23898 ( .A1(n22097), .A2(n22096), .ZN(n22098) );
  INV_X1 U23899 ( .A(n22098), .ZN(n22103) );
  AOI22_X1 U23900 ( .A1(n22103), .A2(n22100), .B1(n22099), .B2(n22098), .ZN(
        P3_U3295) );
  OAI21_X1 U23901 ( .B1(n22103), .B2(n22102), .A(n22101), .ZN(P3_U2637) );
  AOI211_X1 U23902 ( .C1(n22106), .C2(n22424), .A(n22105), .B(n22104), .ZN(
        n22113) );
  INV_X1 U23903 ( .A(n22107), .ZN(n22108) );
  OAI211_X1 U23904 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n22109), .A(n22108), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n22110) );
  AOI21_X1 U23905 ( .B1(n22110), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n22397), 
        .ZN(n22112) );
  NAND2_X1 U23906 ( .A1(n22113), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n22111) );
  OAI21_X1 U23907 ( .B1(n22113), .B2(n22112), .A(n22111), .ZN(P1_U3485) );
  OAI22_X1 U23908 ( .A1(n22119), .A2(n22115), .B1(n22122), .B2(n22114), .ZN(
        n22187) );
  OAI221_X1 U23909 ( .B1(n22187), .B2(n22116), .C1(n22187), .C2(n22188), .A(
        n22138), .ZN(n22128) );
  OAI21_X1 U23910 ( .B1(n22138), .B2(n22122), .A(n22188), .ZN(n22117) );
  OAI211_X1 U23911 ( .C1(n22120), .C2(n22119), .A(n22118), .B(n22117), .ZN(
        n22121) );
  AOI21_X1 U23912 ( .B1(n22123), .B2(n22122), .A(n22121), .ZN(n22136) );
  OAI222_X1 U23913 ( .A1(n22125), .A2(n22214), .B1(n22138), .B2(n22136), .C1(
        n22218), .C2(n22124), .ZN(n22126) );
  INV_X1 U23914 ( .A(n22126), .ZN(n22127) );
  OAI211_X1 U23915 ( .C1(n22130), .C2(n22129), .A(n22128), .B(n22127), .ZN(
        P1_U3018) );
  INV_X1 U23916 ( .A(n22131), .ZN(n22133) );
  AOI22_X1 U23917 ( .A1(n22133), .A2(n22200), .B1(n22199), .B2(n22132), .ZN(
        n22143) );
  NAND2_X1 U23918 ( .A1(n22138), .A2(n22187), .ZN(n22135) );
  AOI21_X1 U23919 ( .B1(n22136), .B2(n22135), .A(n22134), .ZN(n22141) );
  NAND2_X1 U23920 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n22137) );
  NOR4_X1 U23921 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n22139), .A3(
        n22138), .A4(n22137), .ZN(n22140) );
  AOI211_X1 U23922 ( .C1(n22202), .C2(P1_REIP_REG_14__SCAN_IN), .A(n22141), 
        .B(n22140), .ZN(n22142) );
  NAND2_X1 U23923 ( .A1(n22143), .A2(n22142), .ZN(P1_U3017) );
  OAI21_X1 U23924 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n22144), .ZN(n22155) );
  AOI211_X1 U23925 ( .C1(n22148), .C2(n22147), .A(n22146), .B(n22145), .ZN(
        n22161) );
  INV_X1 U23926 ( .A(n22161), .ZN(n22149) );
  NAND2_X1 U23927 ( .A1(n22149), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n22151) );
  OAI211_X1 U23928 ( .C1(n22214), .C2(n22257), .A(n22151), .B(n22150), .ZN(
        n22152) );
  AOI21_X1 U23929 ( .B1(n22153), .B2(n22200), .A(n22152), .ZN(n22154) );
  OAI21_X1 U23930 ( .B1(n22162), .B2(n22155), .A(n22154), .ZN(P1_U3027) );
  INV_X1 U23931 ( .A(n22156), .ZN(n22159) );
  OAI21_X1 U23932 ( .B1(n22214), .B2(n22252), .A(n22157), .ZN(n22158) );
  AOI21_X1 U23933 ( .B1(n22159), .B2(n22200), .A(n22158), .ZN(n22160) );
  OAI221_X1 U23934 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n22162), .C1(
        n14216), .C2(n22161), .A(n22160), .ZN(P1_U3028) );
  INV_X1 U23935 ( .A(n22177), .ZN(n22165) );
  OAI22_X1 U23936 ( .A1(n22163), .A2(n22218), .B1(n22214), .B2(n22348), .ZN(
        n22164) );
  AOI21_X1 U23937 ( .B1(n14256), .B2(n22165), .A(n22164), .ZN(n22167) );
  NAND2_X1 U23938 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n22202), .ZN(n22166) );
  OAI211_X1 U23939 ( .C1(n22185), .C2(n14256), .A(n22167), .B(n22166), .ZN(
        P1_U3016) );
  NOR3_X1 U23940 ( .A1(n22177), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n22168), .ZN(n22171) );
  NOR2_X1 U23941 ( .A1(n22169), .A2(n22218), .ZN(n22170) );
  AOI211_X1 U23942 ( .C1(n22190), .C2(P1_REIP_REG_18__SCAN_IN), .A(n22171), 
        .B(n22170), .ZN(n22176) );
  INV_X1 U23943 ( .A(n22172), .ZN(n22174) );
  AOI22_X1 U23944 ( .A1(n22174), .A2(n22199), .B1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n22173), .ZN(n22175) );
  NAND2_X1 U23945 ( .A1(n22176), .A2(n22175), .ZN(P1_U3013) );
  AOI21_X1 U23946 ( .B1(n17098), .B2(n14256), .A(n22177), .ZN(n22179) );
  AOI22_X1 U23947 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n22190), .B1(n22179), 
        .B2(n22178), .ZN(n22184) );
  INV_X1 U23948 ( .A(n22180), .ZN(n22182) );
  AOI22_X1 U23949 ( .A1(n22182), .A2(n22200), .B1(n22199), .B2(n22181), .ZN(
        n22183) );
  OAI211_X1 U23950 ( .C1(n22185), .C2(n17098), .A(n22184), .B(n22183), .ZN(
        P1_U3015) );
  AOI221_X1 U23951 ( .B1(n22188), .B2(n17081), .C1(n22187), .C2(n17081), .A(
        n22186), .ZN(n22195) );
  NOR2_X1 U23952 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17081), .ZN(
        n22189) );
  AOI22_X1 U23953 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n22190), .B1(n22189), 
        .B2(n22206), .ZN(n22194) );
  AOI22_X1 U23954 ( .A1(n22192), .A2(n22200), .B1(n22199), .B2(n22191), .ZN(
        n22193) );
  OAI211_X1 U23955 ( .C1(n22196), .C2(n22195), .A(n22194), .B(n22193), .ZN(
        P1_U3011) );
  INV_X1 U23956 ( .A(n22197), .ZN(n22201) );
  AOI22_X1 U23957 ( .A1(n22201), .A2(n22200), .B1(n22199), .B2(n22198), .ZN(
        n22211) );
  NAND2_X1 U23958 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n22202), .ZN(n22210) );
  OAI21_X1 U23959 ( .B1(n22204), .B2(n22203), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n22209) );
  NAND3_X1 U23960 ( .A1(n22207), .A2(n22206), .A3(n22205), .ZN(n22208) );
  NAND4_X1 U23961 ( .A1(n22211), .A2(n22210), .A3(n22209), .A4(n22208), .ZN(
        P1_U3009) );
  OAI21_X1 U23962 ( .B1(n22214), .B2(n22213), .A(n22212), .ZN(n22215) );
  INV_X1 U23963 ( .A(n22215), .ZN(n22216) );
  OAI211_X1 U23964 ( .C1(n22219), .C2(n22218), .A(n22217), .B(n22216), .ZN(
        n22220) );
  INV_X1 U23965 ( .A(n22220), .ZN(n22221) );
  OAI221_X1 U23966 ( .B1(n11214), .B2(n22223), .C1(n11214), .C2(n22222), .A(
        n22221), .ZN(P1_U3031) );
  AOI21_X1 U23967 ( .B1(n22248), .B2(n22247), .A(n22238), .ZN(n22236) );
  INV_X1 U23968 ( .A(n22265), .ZN(n22225) );
  AOI22_X1 U23969 ( .A1(n22225), .A2(n22224), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n22371), .ZN(n22227) );
  NAND3_X1 U23970 ( .A1(n22248), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n22246), 
        .ZN(n22226) );
  OAI211_X1 U23971 ( .C1(n22374), .C2(n22228), .A(n22227), .B(n22226), .ZN(
        n22229) );
  AOI21_X1 U23972 ( .B1(n22327), .B2(n22230), .A(n22229), .ZN(n22235) );
  OAI22_X1 U23973 ( .A1(n22232), .A2(n22259), .B1(n22231), .B2(n22383), .ZN(
        n22233) );
  INV_X1 U23974 ( .A(n22233), .ZN(n22234) );
  OAI211_X1 U23975 ( .C1(n22236), .C2(n22246), .A(n22235), .B(n22234), .ZN(
        P1_U2838) );
  INV_X1 U23976 ( .A(n22237), .ZN(n22240) );
  AOI22_X1 U23977 ( .A1(n22371), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n22238), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n22239) );
  OAI21_X1 U23978 ( .B1(n22240), .B2(n22265), .A(n22239), .ZN(n22241) );
  AOI21_X1 U23979 ( .B1(n22358), .B2(P1_EBX_REG_3__SCAN_IN), .A(n22241), .ZN(
        n22242) );
  OAI21_X1 U23980 ( .B1(n22243), .B2(n22259), .A(n22242), .ZN(n22244) );
  AOI21_X1 U23981 ( .B1(n22245), .B2(n22353), .A(n22244), .ZN(n22251) );
  NOR2_X1 U23982 ( .A1(n22247), .A2(n22246), .ZN(n22249) );
  OAI211_X1 U23983 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(n22249), .A(n22248), .B(
        n22253), .ZN(n22250) );
  OAI211_X1 U23984 ( .C1(n22252), .C2(n22375), .A(n22251), .B(n22250), .ZN(
        P1_U2837) );
  NOR3_X1 U23985 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22323), .A3(n22253), .ZN(
        n22254) );
  AOI211_X1 U23986 ( .C1(n22371), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22325), .B(n22254), .ZN(n22264) );
  OAI21_X1 U23987 ( .B1(n22323), .B2(n22272), .A(n22255), .ZN(n22274) );
  OAI22_X1 U23988 ( .A1(n22375), .A2(n22257), .B1(n22374), .B2(n22256), .ZN(
        n22262) );
  OAI22_X1 U23989 ( .A1(n22260), .A2(n22259), .B1(n22258), .B2(n22383), .ZN(
        n22261) );
  AOI211_X1 U23990 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n22274), .A(n22262), .B(
        n22261), .ZN(n22263) );
  OAI211_X1 U23991 ( .C1(n22266), .C2(n22265), .A(n22264), .B(n22263), .ZN(
        P1_U2836) );
  NOR2_X1 U23992 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22323), .ZN(n22273) );
  INV_X1 U23993 ( .A(n22267), .ZN(n22268) );
  AOI22_X1 U23994 ( .A1(n22327), .A2(n22268), .B1(n22358), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n22269) );
  OAI211_X1 U23995 ( .C1(n22337), .C2(n22270), .A(n22269), .B(n22354), .ZN(
        n22271) );
  AOI21_X1 U23996 ( .B1(n22273), .B2(n22272), .A(n22271), .ZN(n22278) );
  AOI22_X1 U23997 ( .A1(n22276), .A2(n22275), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n22274), .ZN(n22277) );
  OAI211_X1 U23998 ( .C1(n22279), .C2(n22383), .A(n22278), .B(n22277), .ZN(
        P1_U2835) );
  OAI22_X1 U23999 ( .A1(n22375), .A2(n22281), .B1(n22374), .B2(n22280), .ZN(
        n22282) );
  AOI211_X1 U24000 ( .C1(n22371), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n22325), .B(n22282), .ZN(n22289) );
  NOR3_X1 U24001 ( .A1(n22284), .A2(n22323), .A3(n22285), .ZN(n22307) );
  INV_X1 U24002 ( .A(n22307), .ZN(n22283) );
  AND2_X1 U24003 ( .A1(n22339), .A2(n22283), .ZN(n22297) );
  OAI21_X1 U24004 ( .B1(n22323), .B2(n22285), .A(n22284), .ZN(n22286) );
  AOI22_X1 U24005 ( .A1(n22287), .A2(n22362), .B1(n22297), .B2(n22286), .ZN(
        n22288) );
  OAI211_X1 U24006 ( .C1(n22290), .C2(n22383), .A(n22289), .B(n22288), .ZN(
        P1_U2834) );
  OAI21_X1 U24007 ( .B1(n22337), .B2(n22291), .A(n22354), .ZN(n22295) );
  OAI22_X1 U24008 ( .A1(n22375), .A2(n22293), .B1(n22374), .B2(n22292), .ZN(
        n22294) );
  AOI211_X1 U24009 ( .C1(n22307), .C2(n22296), .A(n22295), .B(n22294), .ZN(
        n22300) );
  AOI22_X1 U24010 ( .A1(n22298), .A2(n22362), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n22297), .ZN(n22299) );
  OAI211_X1 U24011 ( .C1(n22301), .C2(n22383), .A(n22300), .B(n22299), .ZN(
        P1_U2833) );
  AOI22_X1 U24012 ( .A1(n22327), .A2(n22302), .B1(n22358), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n22311) );
  AOI21_X1 U24013 ( .B1(n22371), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n22325), .ZN(n22310) );
  INV_X1 U24014 ( .A(n22303), .ZN(n22304) );
  AOI22_X1 U24015 ( .A1(n22305), .A2(n22362), .B1(n22304), .B2(n22353), .ZN(
        n22309) );
  OAI221_X1 U24016 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(P1_REIP_REG_7__SCAN_IN), 
        .C1(P1_REIP_REG_8__SCAN_IN), .C2(n22307), .A(n22306), .ZN(n22308) );
  NAND4_X1 U24017 ( .A1(n22311), .A2(n22310), .A3(n22309), .A4(n22308), .ZN(
        P1_U2832) );
  NOR2_X1 U24018 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22323), .ZN(n22331) );
  AOI22_X1 U24019 ( .A1(n22327), .A2(n22313), .B1(n22312), .B2(n22331), .ZN(
        n22320) );
  INV_X1 U24020 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n22316) );
  NAND2_X1 U24021 ( .A1(n22330), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n22315) );
  AOI21_X1 U24022 ( .B1(n22371), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n22325), .ZN(n22314) );
  OAI211_X1 U24023 ( .C1(n22316), .C2(n22374), .A(n22315), .B(n22314), .ZN(
        n22317) );
  AOI21_X1 U24024 ( .B1(n22362), .B2(n22318), .A(n22317), .ZN(n22319) );
  OAI211_X1 U24025 ( .C1(n22321), .C2(n22383), .A(n22320), .B(n22319), .ZN(
        P1_U2829) );
  NOR3_X1 U24026 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n22323), .A3(n22322), 
        .ZN(n22324) );
  AOI211_X1 U24027 ( .C1(n22371), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n22325), .B(n22324), .ZN(n22335) );
  AOI22_X1 U24028 ( .A1(n22327), .A2(n22326), .B1(n22358), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n22334) );
  AOI22_X1 U24029 ( .A1(n22329), .A2(n22353), .B1(n22362), .B2(n22328), .ZN(
        n22333) );
  OAI21_X1 U24030 ( .B1(n22331), .B2(n22330), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n22332) );
  NAND4_X1 U24031 ( .A1(n22335), .A2(n22334), .A3(n22333), .A4(n22332), .ZN(
        P1_U2828) );
  OAI21_X1 U24032 ( .B1(n22337), .B2(n22336), .A(n22354), .ZN(n22343) );
  AOI21_X1 U24033 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n22339), .A(n22338), 
        .ZN(n22340) );
  NOR2_X1 U24034 ( .A1(n22341), .A2(n22340), .ZN(n22342) );
  AOI211_X1 U24035 ( .C1(P1_EBX_REG_15__SCAN_IN), .C2(n22358), .A(n22343), .B(
        n22342), .ZN(n22347) );
  AOI22_X1 U24036 ( .A1(n22345), .A2(n22362), .B1(n22353), .B2(n22344), .ZN(
        n22346) );
  OAI211_X1 U24037 ( .C1(n22375), .C2(n22348), .A(n22347), .B(n22346), .ZN(
        P1_U2825) );
  NAND3_X1 U24038 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n22350), .A3(n22349), 
        .ZN(n22360) );
  NAND2_X1 U24039 ( .A1(n22371), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n22356) );
  INV_X1 U24040 ( .A(n22351), .ZN(n22352) );
  NAND2_X1 U24041 ( .A1(n22353), .A2(n22352), .ZN(n22355) );
  NAND3_X1 U24042 ( .A1(n22356), .A2(n22355), .A3(n22354), .ZN(n22357) );
  AOI21_X1 U24043 ( .B1(n22358), .B2(P1_EBX_REG_19__SCAN_IN), .A(n22357), .ZN(
        n22359) );
  NAND2_X1 U24044 ( .A1(n22360), .A2(n22359), .ZN(n22361) );
  AOI21_X1 U24045 ( .B1(n22363), .B2(n22362), .A(n22361), .ZN(n22367) );
  OAI21_X1 U24046 ( .B1(n22365), .B2(n22364), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n22366) );
  OAI211_X1 U24047 ( .C1(n22368), .C2(n22375), .A(n22367), .B(n22366), .ZN(
        P1_U2821) );
  AOI22_X1 U24048 ( .A1(n22371), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n22370), .B2(n22369), .ZN(n22372) );
  OAI21_X1 U24049 ( .B1(n22374), .B2(n22373), .A(n22372), .ZN(n22380) );
  OAI22_X1 U24050 ( .A1(n22378), .A2(n22377), .B1(n22376), .B2(n22375), .ZN(
        n22379) );
  AOI211_X1 U24051 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n22381), .A(n22380), 
        .B(n22379), .ZN(n22382) );
  OAI21_X1 U24052 ( .B1(n22384), .B2(n22383), .A(n22382), .ZN(P1_U2819) );
  OAI21_X1 U24053 ( .B1(n22387), .B2(n22386), .A(n22385), .ZN(P1_U2806) );
  NOR2_X1 U24054 ( .A1(n22392), .A2(n22388), .ZN(n22390) );
  OAI21_X1 U24055 ( .B1(n22390), .B2(n22556), .A(n22389), .ZN(P1_U3163) );
  OAI22_X1 U24056 ( .A1(n22394), .A2(n22393), .B1(n22392), .B2(n22391), .ZN(
        P1_U3466) );
  AOI21_X1 U24057 ( .B1(n22397), .B2(n22396), .A(n22395), .ZN(n22398) );
  OAI22_X1 U24058 ( .A1(n22400), .A2(n22399), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22398), .ZN(n22401) );
  OAI21_X1 U24059 ( .B1(n22403), .B2(n22402), .A(n22401), .ZN(P1_U3161) );
  INV_X1 U24060 ( .A(n22404), .ZN(n22406) );
  OAI21_X1 U24061 ( .B1(n22408), .B2(n22405), .A(n22406), .ZN(P1_U2805) );
  OAI21_X1 U24062 ( .B1(n22408), .B2(n22407), .A(n22406), .ZN(P1_U3465) );
  INV_X1 U24063 ( .A(n22409), .ZN(n22411) );
  OAI21_X1 U24064 ( .B1(n22413), .B2(n22410), .A(n22411), .ZN(P2_U2818) );
  OAI21_X1 U24065 ( .B1(n22413), .B2(n22412), .A(n22411), .ZN(P2_U3592) );
  OAI21_X1 U24066 ( .B1(n22417), .B2(n22414), .A(n22415), .ZN(P3_U2636) );
  OAI21_X1 U24067 ( .B1(n22417), .B2(n22416), .A(n22415), .ZN(P3_U3281) );
  INV_X1 U24068 ( .A(HOLD), .ZN(n22462) );
  OAI21_X1 U24069 ( .B1(n22462), .B2(n22463), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22472) );
  AOI21_X1 U24070 ( .B1(HOLD), .B2(P3_STATE_REG_1__SCAN_IN), .A(n22472), .ZN(
        n22420) );
  NAND2_X1 U24071 ( .A1(n22418), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n22471) );
  AND2_X1 U24072 ( .A1(n22471), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n22478) );
  INV_X1 U24073 ( .A(NA), .ZN(n22456) );
  OAI21_X1 U24074 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n22456), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n22477) );
  INV_X1 U24075 ( .A(n22477), .ZN(n22419) );
  OAI22_X1 U24076 ( .A1(n22421), .A2(n22420), .B1(n22478), .B2(n22419), .ZN(
        P3_U3029) );
  NOR2_X1 U24077 ( .A1(NA), .A2(n22424), .ZN(n22423) );
  OAI21_X1 U24078 ( .B1(n22462), .B2(n22433), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22438) );
  OAI211_X1 U24079 ( .C1(n22423), .C2(n22422), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(n22438), .ZN(n22432) );
  NOR2_X1 U24080 ( .A1(n22437), .A2(n22424), .ZN(n22429) );
  INV_X1 U24081 ( .A(n22429), .ZN(n22425) );
  NOR2_X1 U24082 ( .A1(n22426), .A2(n22425), .ZN(n22427) );
  MUX2_X1 U24083 ( .A(P1_STATE_REG_2__SCAN_IN), .B(n22427), .S(
        P1_STATE_REG_0__SCAN_IN), .Z(n22428) );
  AOI22_X1 U24084 ( .A1(n22429), .A2(P1_STATE_REG_2__SCAN_IN), .B1(n22428), 
        .B2(n22456), .ZN(n22431) );
  OAI211_X1 U24085 ( .C1(n22432), .C2(n22462), .A(n22431), .B(n22430), .ZN(
        P1_U3196) );
  OAI221_X1 U24086 ( .B1(n22436), .B2(HOLD), .C1(n22436), .C2(n22433), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n22435) );
  OAI211_X1 U24087 ( .C1(n22440), .C2(n22438), .A(n22435), .B(n22434), .ZN(
        P1_U3195) );
  AOI21_X1 U24088 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n22436), .A(n22440), 
        .ZN(n22442) );
  NOR2_X1 U24089 ( .A1(n22462), .A2(n22437), .ZN(n22439) );
  AOI211_X1 U24090 ( .C1(NA), .C2(n22440), .A(n22439), .B(n22438), .ZN(n22441)
         );
  OAI22_X1 U24091 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22442), .B1(n22855), 
        .B2(n22441), .ZN(P1_U3194) );
  AOI22_X1 U24092 ( .A1(HOLD), .A2(n22443), .B1(NA), .B2(n22455), .ZN(n22448)
         );
  NOR2_X1 U24093 ( .A1(n22445), .A2(n22444), .ZN(n22454) );
  NOR2_X1 U24094 ( .A1(n22454), .A2(n22455), .ZN(n22447) );
  OAI222_X1 U24095 ( .A1(n22449), .A2(n22448), .B1(P2_STATE_REG_2__SCAN_IN), 
        .B2(n22447), .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n22446), .ZN(
        P2_U3209) );
  OAI211_X1 U24096 ( .C1(n22462), .C2(n22461), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22452) );
  INV_X1 U24097 ( .A(n22454), .ZN(n22457) );
  NAND2_X1 U24098 ( .A1(n22450), .A2(HOLD), .ZN(n22451) );
  NAND4_X1 U24099 ( .A1(n22453), .A2(n22452), .A3(n22457), .A4(n22451), .ZN(
        P2_U3210) );
  AOI221_X1 U24100 ( .B1(HOLD), .B2(P2_STATE_REG_0__SCAN_IN), .C1(n22456), 
        .C2(n22455), .A(n22454), .ZN(n22460) );
  OAI22_X1 U24101 ( .A1(NA), .A2(n22457), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22458) );
  OAI211_X1 U24102 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n22458), .ZN(n22459) );
  OAI221_X1 U24103 ( .B1(n22461), .B2(n22460), .C1(n22461), .C2(n18186), .A(
        n22459), .ZN(P2_U3211) );
  NOR2_X1 U24104 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22476)
         );
  OAI21_X1 U24105 ( .B1(n22462), .B2(n22463), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n22473) );
  OAI21_X1 U24106 ( .B1(n22476), .B2(n22473), .A(n22471), .ZN(n22467) );
  AOI221_X1 U24107 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n22472), .C1(n22464), 
        .C2(n22463), .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22466) );
  AOI211_X1 U24108 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(n22467), .A(n22466), 
        .B(n22465), .ZN(n22468) );
  OAI21_X1 U24109 ( .B1(n22470), .B2(n22469), .A(n22468), .ZN(P3_U3030) );
  NOR2_X1 U24110 ( .A1(NA), .A2(n22471), .ZN(n22474) );
  OAI221_X1 U24111 ( .B1(n22474), .B2(n22473), .C1(n22474), .C2(n22472), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n22475) );
  OAI22_X1 U24112 ( .A1(n22478), .A2(n22477), .B1(n22476), .B2(n22475), .ZN(
        P3_U3031) );
  NOR2_X1 U24113 ( .A1(n22480), .A2(n22479), .ZN(n22483) );
  AOI21_X1 U24114 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n22528), .A(n22483), 
        .ZN(n22481) );
  OAI21_X1 U24115 ( .B1(n22482), .B2(n22525), .A(n22481), .ZN(P1_U2945) );
  AOI21_X1 U24116 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n22528), .A(n22483), 
        .ZN(n22484) );
  OAI21_X1 U24117 ( .B1(n15796), .B2(n22525), .A(n22484), .ZN(P1_U2960) );
  INV_X1 U24118 ( .A(n22485), .ZN(n22486) );
  NAND2_X1 U24119 ( .A1(n22521), .A2(n22486), .ZN(n22490) );
  INV_X1 U24120 ( .A(n22490), .ZN(n22487) );
  AOI21_X1 U24121 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n22523), .A(n22487), 
        .ZN(n22488) );
  OAI21_X1 U24122 ( .B1(n22489), .B2(n22525), .A(n22488), .ZN(P1_U2946) );
  AOI22_X1 U24123 ( .A1(n22523), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(
        P1_EAX_REG_9__SCAN_IN), .B2(n22527), .ZN(n22491) );
  NAND2_X1 U24124 ( .A1(n22491), .A2(n22490), .ZN(P1_U2961) );
  INV_X1 U24125 ( .A(n22492), .ZN(n22493) );
  NAND2_X1 U24126 ( .A1(n22521), .A2(n22493), .ZN(n22497) );
  INV_X1 U24127 ( .A(n22497), .ZN(n22494) );
  AOI21_X1 U24128 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n22523), .A(n22494), 
        .ZN(n22495) );
  OAI21_X1 U24129 ( .B1(n22496), .B2(n22525), .A(n22495), .ZN(P1_U2947) );
  AOI22_X1 U24130 ( .A1(n22528), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(
        P1_EAX_REG_10__SCAN_IN), .B2(n22527), .ZN(n22498) );
  NAND2_X1 U24131 ( .A1(n22498), .A2(n22497), .ZN(P1_U2962) );
  NAND2_X1 U24132 ( .A1(n22521), .A2(n22499), .ZN(n22503) );
  INV_X1 U24133 ( .A(n22503), .ZN(n22500) );
  AOI21_X1 U24134 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n22523), .A(n22500), 
        .ZN(n22501) );
  OAI21_X1 U24135 ( .B1(n22502), .B2(n22525), .A(n22501), .ZN(P1_U2948) );
  AOI22_X1 U24136 ( .A1(n22528), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(
        P1_EAX_REG_11__SCAN_IN), .B2(n22527), .ZN(n22504) );
  NAND2_X1 U24137 ( .A1(n22504), .A2(n22503), .ZN(P1_U2963) );
  INV_X1 U24138 ( .A(n22505), .ZN(n22506) );
  NAND2_X1 U24139 ( .A1(n22521), .A2(n22506), .ZN(n22510) );
  INV_X1 U24140 ( .A(n22510), .ZN(n22507) );
  AOI21_X1 U24141 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n22523), .A(n22507), 
        .ZN(n22508) );
  OAI21_X1 U24142 ( .B1(n22509), .B2(n22525), .A(n22508), .ZN(P1_U2949) );
  AOI22_X1 U24143 ( .A1(n22528), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(
        P1_EAX_REG_12__SCAN_IN), .B2(n22527), .ZN(n22511) );
  NAND2_X1 U24144 ( .A1(n22511), .A2(n22510), .ZN(P1_U2964) );
  INV_X1 U24145 ( .A(n22512), .ZN(n22513) );
  NAND2_X1 U24146 ( .A1(n22521), .A2(n22513), .ZN(n22517) );
  INV_X1 U24147 ( .A(n22517), .ZN(n22514) );
  AOI21_X1 U24148 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n22523), .A(n22514), 
        .ZN(n22515) );
  OAI21_X1 U24149 ( .B1(n22516), .B2(n22525), .A(n22515), .ZN(P1_U2950) );
  AOI22_X1 U24150 ( .A1(n22528), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(
        P1_EAX_REG_13__SCAN_IN), .B2(n22527), .ZN(n22518) );
  NAND2_X1 U24151 ( .A1(n22518), .A2(n22517), .ZN(P1_U2965) );
  INV_X1 U24152 ( .A(n22519), .ZN(n22520) );
  NAND2_X1 U24153 ( .A1(n22521), .A2(n22520), .ZN(n22529) );
  INV_X1 U24154 ( .A(n22529), .ZN(n22522) );
  AOI21_X1 U24155 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n22523), .A(n22522), 
        .ZN(n22524) );
  OAI21_X1 U24156 ( .B1(n22526), .B2(n22525), .A(n22524), .ZN(P1_U2951) );
  AOI22_X1 U24157 ( .A1(n22528), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(
        P1_EAX_REG_14__SCAN_IN), .B2(n22527), .ZN(n22530) );
  NAND2_X1 U24158 ( .A1(n22530), .A2(n22529), .ZN(P1_U2966) );
  NOR3_X1 U24159 ( .A1(n22776), .A2(n22846), .A3(n22609), .ZN(n22531) );
  NOR2_X1 U24160 ( .A1(n22609), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22627) );
  NOR2_X1 U24161 ( .A1(n22531), .A2(n22627), .ZN(n22539) );
  INV_X1 U24162 ( .A(n22539), .ZN(n22533) );
  NOR2_X1 U24163 ( .A1(n22566), .A2(n22629), .ZN(n22538) );
  INV_X1 U24164 ( .A(n22536), .ZN(n22532) );
  NOR2_X1 U24165 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22534), .ZN(
        n22775) );
  AOI22_X1 U24166 ( .A1(n22846), .A2(n22655), .B1(n22775), .B2(n22652), .ZN(
        n22541) );
  INV_X1 U24167 ( .A(n22775), .ZN(n22535) );
  AOI22_X1 U24168 ( .A1(n22536), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22535), .ZN(n22537) );
  OAI211_X1 U24169 ( .C1(n22539), .C2(n22538), .A(n22622), .B(n22537), .ZN(
        n22777) );
  AOI22_X1 U24170 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22777), .B1(
        n22776), .B2(n22635), .ZN(n22540) );
  OAI211_X1 U24171 ( .C1(n22780), .C2(n22644), .A(n22541), .B(n22540), .ZN(
        P1_U3033) );
  INV_X1 U24172 ( .A(n22635), .ZN(n22660) );
  INV_X1 U24173 ( .A(n22542), .ZN(n22544) );
  AOI22_X1 U24174 ( .A1(n22544), .A2(n22654), .B1(n22652), .B2(n22543), .ZN(
        n22547) );
  AOI22_X1 U24175 ( .A1(n22545), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n22776), .B2(n22655), .ZN(n22546) );
  OAI211_X1 U24176 ( .C1(n22660), .C2(n22782), .A(n22547), .B(n22546), .ZN(
        P1_U3041) );
  NOR2_X1 U24177 ( .A1(n22789), .A2(n22609), .ZN(n22549) );
  AOI21_X1 U24178 ( .B1(n22549), .B2(n22782), .A(n22627), .ZN(n22559) );
  INV_X1 U24179 ( .A(n22559), .ZN(n22551) );
  NOR2_X1 U24180 ( .A1(n22566), .A2(n22611), .ZN(n22558) );
  NOR2_X1 U24181 ( .A1(n22550), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22586) );
  NAND3_X1 U24182 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n22553), .A3(
        n22552), .ZN(n22573) );
  NOR2_X1 U24183 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22573), .ZN(
        n22695) );
  INV_X1 U24184 ( .A(n22695), .ZN(n22781) );
  OAI22_X1 U24185 ( .A1(n22782), .A2(n22554), .B1(n22781), .B2(n22617), .ZN(
        n22555) );
  INV_X1 U24186 ( .A(n22555), .ZN(n22561) );
  NOR2_X1 U24187 ( .A1(n22586), .A2(n22556), .ZN(n22589) );
  AOI21_X1 U24188 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22781), .A(n22589), 
        .ZN(n22557) );
  OAI211_X1 U24189 ( .C1(n22559), .C2(n22558), .A(n22622), .B(n22557), .ZN(
        n22784) );
  AOI22_X1 U24190 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22784), .B1(
        n22789), .B2(n22635), .ZN(n22560) );
  OAI211_X1 U24191 ( .C1(n22787), .C2(n22644), .A(n22561), .B(n22560), .ZN(
        P1_U3049) );
  INV_X1 U24192 ( .A(n22573), .ZN(n22570) );
  INV_X1 U24193 ( .A(n22562), .ZN(n22564) );
  OAI21_X1 U24194 ( .B1(n22564), .B2(n22609), .A(n22563), .ZN(n22571) );
  NAND2_X1 U24195 ( .A1(n11162), .A2(n13313), .ZN(n22565) );
  OR2_X1 U24196 ( .A1(n22566), .A2(n22565), .ZN(n22569) );
  NOR2_X1 U24197 ( .A1(n22567), .A2(n22573), .ZN(n22788) );
  INV_X1 U24198 ( .A(n22788), .ZN(n22568) );
  NAND2_X1 U24199 ( .A1(n22569), .A2(n22568), .ZN(n22575) );
  AOI22_X1 U24200 ( .A1(n22789), .A2(n22655), .B1(n22788), .B2(n22652), .ZN(
        n22578) );
  INV_X1 U24201 ( .A(n22571), .ZN(n22576) );
  AOI21_X1 U24202 ( .B1(n22609), .B2(n22573), .A(n22572), .ZN(n22574) );
  AOI22_X1 U24203 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22791), .B1(
        n22790), .B2(n22635), .ZN(n22577) );
  OAI211_X1 U24204 ( .C1(n22794), .C2(n22644), .A(n22578), .B(n22577), .ZN(
        P1_U3057) );
  AOI22_X1 U24205 ( .A1(n22654), .A2(n22580), .B1(n22652), .B2(n22579), .ZN(
        n22583) );
  AOI22_X1 U24206 ( .A1(n22581), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n22790), .B2(n22655), .ZN(n22582) );
  OAI211_X1 U24207 ( .C1(n22660), .C2(n22800), .A(n22583), .B(n22582), .ZN(
        P1_U3065) );
  NOR3_X1 U24208 ( .A1(n22803), .A2(n22802), .A3(n22609), .ZN(n22584) );
  NOR2_X1 U24209 ( .A1(n22584), .A2(n22627), .ZN(n22593) );
  INV_X1 U24210 ( .A(n22593), .ZN(n22587) );
  AND2_X1 U24211 ( .A1(n22585), .A2(n22629), .ZN(n22592) );
  NOR2_X1 U24212 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22588), .ZN(
        n22801) );
  AOI22_X1 U24213 ( .A1(n22802), .A2(n22655), .B1(n22801), .B2(n22652), .ZN(
        n22595) );
  INV_X1 U24214 ( .A(n22801), .ZN(n22590) );
  AOI21_X1 U24215 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22590), .A(n22589), 
        .ZN(n22591) );
  OAI211_X1 U24216 ( .C1(n22593), .C2(n22592), .A(n22639), .B(n22591), .ZN(
        n22804) );
  AOI22_X1 U24217 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22804), .B1(
        n22803), .B2(n22635), .ZN(n22594) );
  OAI211_X1 U24218 ( .C1(n22807), .C2(n22644), .A(n22595), .B(n22594), .ZN(
        P1_U3081) );
  INV_X1 U24219 ( .A(n22596), .ZN(n22598) );
  AOI22_X1 U24220 ( .A1(n22598), .A2(n22654), .B1(n22597), .B2(n22652), .ZN(
        n22601) );
  AOI22_X1 U24221 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22599), .B1(
        n22803), .B2(n22655), .ZN(n22600) );
  OAI211_X1 U24222 ( .C1(n22660), .C2(n22602), .A(n22601), .B(n22600), .ZN(
        P1_U3089) );
  AOI22_X1 U24223 ( .A1(n22604), .A2(n22654), .B1(n22652), .B2(n22603), .ZN(
        n22608) );
  AOI22_X1 U24224 ( .A1(n22606), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n22605), .B2(n22655), .ZN(n22607) );
  OAI211_X1 U24225 ( .C1(n22660), .C2(n22814), .A(n22608), .B(n22607), .ZN(
        P1_U3097) );
  NOR3_X1 U24226 ( .A1(n22766), .A2(n22819), .A3(n22609), .ZN(n22610) );
  NOR2_X1 U24227 ( .A1(n22610), .A2(n22627), .ZN(n22624) );
  INV_X1 U24228 ( .A(n22624), .ZN(n22615) );
  NOR2_X1 U24229 ( .A1(n22612), .A2(n22611), .ZN(n22623) );
  NOR2_X1 U24230 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22616), .ZN(
        n22765) );
  INV_X1 U24231 ( .A(n22765), .ZN(n22816) );
  OAI22_X1 U24232 ( .A1(n22830), .A2(n22660), .B1(n22617), .B2(n22816), .ZN(
        n22618) );
  INV_X1 U24233 ( .A(n22618), .ZN(n22626) );
  INV_X1 U24234 ( .A(n22619), .ZN(n22620) );
  AOI21_X1 U24235 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22816), .A(n22620), 
        .ZN(n22621) );
  OAI211_X1 U24236 ( .C1(n22624), .C2(n22623), .A(n22622), .B(n22621), .ZN(
        n22820) );
  AOI22_X1 U24237 ( .A1(n22820), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22819), .B2(n22655), .ZN(n22625) );
  OAI211_X1 U24238 ( .C1(n22823), .C2(n22644), .A(n22626), .B(n22625), .ZN(
        P1_U3113) );
  NOR3_X1 U24239 ( .A1(n22834), .A2(n22832), .A3(n22609), .ZN(n22628) );
  NOR2_X1 U24240 ( .A1(n22628), .A2(n22627), .ZN(n22641) );
  INV_X1 U24241 ( .A(n22641), .ZN(n22633) );
  NOR2_X1 U24242 ( .A1(n22630), .A2(n22629), .ZN(n22640) );
  INV_X1 U24243 ( .A(n22637), .ZN(n22631) );
  NOR2_X1 U24244 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22634), .ZN(
        n22831) );
  AOI22_X1 U24245 ( .A1(n22832), .A2(n22635), .B1(n22652), .B2(n22831), .ZN(
        n22643) );
  INV_X1 U24246 ( .A(n22831), .ZN(n22636) );
  AOI22_X1 U24247 ( .A1(n22637), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22636), .ZN(n22638) );
  OAI211_X1 U24248 ( .C1(n22641), .C2(n22640), .A(n22639), .B(n22638), .ZN(
        n22835) );
  AOI22_X1 U24249 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n22834), .B2(n22655), .ZN(n22642) );
  OAI211_X1 U24250 ( .C1(n22839), .C2(n22644), .A(n22643), .B(n22642), .ZN(
        P1_U3129) );
  AOI22_X1 U24251 ( .A1(n22654), .A2(n22646), .B1(n22652), .B2(n22645), .ZN(
        n22649) );
  AOI22_X1 U24252 ( .A1(n22647), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n22832), .B2(n22655), .ZN(n22648) );
  OAI211_X1 U24253 ( .C1(n22660), .C2(n22650), .A(n22649), .B(n22648), .ZN(
        P1_U3137) );
  AOI22_X1 U24254 ( .A1(n22654), .A2(n22653), .B1(n22652), .B2(n22651), .ZN(
        n22659) );
  AOI22_X1 U24255 ( .A1(n22657), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n22656), .B2(n22655), .ZN(n22658) );
  OAI211_X1 U24256 ( .C1(n22660), .C2(n22850), .A(n22659), .B(n22658), .ZN(
        P1_U3145) );
  AOI22_X1 U24257 ( .A1(n22846), .A2(n11149), .B1(n22775), .B2(n22671), .ZN(
        n22662) );
  AOI22_X1 U24258 ( .A1(n22777), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n22776), .B2(n22672), .ZN(n22661) );
  OAI211_X1 U24259 ( .C1(n22780), .C2(n22676), .A(n22662), .B(n22661), .ZN(
        P1_U3034) );
  AOI22_X1 U24260 ( .A1(n22789), .A2(n22672), .B1(n22695), .B2(n22671), .ZN(
        n22664) );
  AOI22_X1 U24261 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n22696), .B2(n11149), .ZN(n22663) );
  OAI211_X1 U24262 ( .C1(n22787), .C2(n22676), .A(n22664), .B(n22663), .ZN(
        P1_U3050) );
  AOI22_X1 U24263 ( .A1(n22790), .A2(n22672), .B1(n22671), .B2(n22788), .ZN(
        n22666) );
  AOI22_X1 U24264 ( .A1(n22791), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n22789), .B2(n11149), .ZN(n22665) );
  OAI211_X1 U24265 ( .C1(n22794), .C2(n22676), .A(n22666), .B(n22665), .ZN(
        P1_U3058) );
  AOI22_X1 U24266 ( .A1(n22802), .A2(n11149), .B1(n22801), .B2(n22671), .ZN(
        n22668) );
  AOI22_X1 U24267 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n22803), .B2(n22672), .ZN(n22667) );
  OAI211_X1 U24268 ( .C1(n22807), .C2(n22676), .A(n22668), .B(n22667), .ZN(
        P1_U3082) );
  AOI22_X1 U24269 ( .A1(n11149), .A2(n22819), .B1(n22765), .B2(n22671), .ZN(
        n22670) );
  AOI22_X1 U24270 ( .A1(n22820), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n22766), .B2(n22672), .ZN(n22669) );
  OAI211_X1 U24271 ( .C1(n22823), .C2(n22676), .A(n22670), .B(n22669), .ZN(
        P1_U3114) );
  AOI22_X1 U24272 ( .A1(n22832), .A2(n22672), .B1(n22831), .B2(n22671), .ZN(
        n22675) );
  AOI22_X1 U24273 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n22834), .B2(n11149), .ZN(n22674) );
  OAI211_X1 U24274 ( .C1(n22839), .C2(n22676), .A(n22675), .B(n22674), .ZN(
        P1_U3130) );
  AOI22_X1 U24275 ( .A1(n22846), .A2(n22689), .B1(n22775), .B2(n22687), .ZN(
        n22678) );
  AOI22_X1 U24276 ( .A1(n22777), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n22776), .B2(n22688), .ZN(n22677) );
  OAI211_X1 U24277 ( .C1(n22780), .C2(n22692), .A(n22678), .B(n22677), .ZN(
        P1_U3035) );
  AOI22_X1 U24278 ( .A1(n22789), .A2(n22688), .B1(n22695), .B2(n22687), .ZN(
        n22680) );
  AOI22_X1 U24279 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n22696), .B2(n22689), .ZN(n22679) );
  OAI211_X1 U24280 ( .C1(n22787), .C2(n22692), .A(n22680), .B(n22679), .ZN(
        P1_U3051) );
  AOI22_X1 U24281 ( .A1(n22789), .A2(n22689), .B1(n22788), .B2(n22687), .ZN(
        n22682) );
  AOI22_X1 U24282 ( .A1(n22791), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n22790), .B2(n22688), .ZN(n22681) );
  OAI211_X1 U24283 ( .C1(n22794), .C2(n22692), .A(n22682), .B(n22681), .ZN(
        P1_U3059) );
  AOI22_X1 U24284 ( .A1(n22802), .A2(n22689), .B1(n22801), .B2(n22687), .ZN(
        n22684) );
  AOI22_X1 U24285 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22803), .B2(n22688), .ZN(n22683) );
  OAI211_X1 U24286 ( .C1(n22807), .C2(n22692), .A(n22684), .B(n22683), .ZN(
        P1_U3083) );
  AOI22_X1 U24287 ( .A1(n22819), .A2(n22689), .B1(n22765), .B2(n22687), .ZN(
        n22686) );
  AOI22_X1 U24288 ( .A1(n22820), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n22766), .B2(n22688), .ZN(n22685) );
  OAI211_X1 U24289 ( .C1(n22823), .C2(n22692), .A(n22686), .B(n22685), .ZN(
        P1_U3115) );
  AOI22_X1 U24290 ( .A1(n22832), .A2(n22688), .B1(n22831), .B2(n22687), .ZN(
        n22691) );
  AOI22_X1 U24291 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22834), .B2(n22689), .ZN(n22690) );
  OAI211_X1 U24292 ( .C1(n22839), .C2(n22692), .A(n22691), .B(n22690), .ZN(
        P1_U3131) );
  AOI22_X1 U24293 ( .A1(n22846), .A2(n22710), .B1(n22775), .B2(n22708), .ZN(
        n22694) );
  AOI22_X1 U24294 ( .A1(n22777), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n22776), .B2(n22709), .ZN(n22693) );
  OAI211_X1 U24295 ( .C1(n22780), .C2(n22713), .A(n22694), .B(n22693), .ZN(
        P1_U3036) );
  AOI22_X1 U24296 ( .A1(n22789), .A2(n22709), .B1(n22695), .B2(n22708), .ZN(
        n22698) );
  AOI22_X1 U24297 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n22696), .B2(n22710), .ZN(n22697) );
  OAI211_X1 U24298 ( .C1(n22787), .C2(n22713), .A(n22698), .B(n22697), .ZN(
        P1_U3052) );
  AOI22_X1 U24299 ( .A1(n22790), .A2(n22709), .B1(n22708), .B2(n22788), .ZN(
        n22700) );
  AOI22_X1 U24300 ( .A1(n22791), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22789), .B2(n22710), .ZN(n22699) );
  OAI211_X1 U24301 ( .C1(n22794), .C2(n22713), .A(n22700), .B(n22699), .ZN(
        P1_U3060) );
  AOI22_X1 U24302 ( .A1(n22803), .A2(n22709), .B1(n22801), .B2(n22708), .ZN(
        n22702) );
  AOI22_X1 U24303 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22802), .B2(n22710), .ZN(n22701) );
  OAI211_X1 U24304 ( .C1(n22807), .C2(n22713), .A(n22702), .B(n22701), .ZN(
        P1_U3084) );
  OAI22_X1 U24305 ( .A1(n22830), .A2(n22704), .B1(n22816), .B2(n22703), .ZN(
        n22705) );
  INV_X1 U24306 ( .A(n22705), .ZN(n22707) );
  AOI22_X1 U24307 ( .A1(n22820), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22819), .B2(n22710), .ZN(n22706) );
  OAI211_X1 U24308 ( .C1(n22823), .C2(n22713), .A(n22707), .B(n22706), .ZN(
        P1_U3116) );
  AOI22_X1 U24309 ( .A1(n22832), .A2(n22709), .B1(n22831), .B2(n22708), .ZN(
        n22712) );
  AOI22_X1 U24310 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22834), .B2(n22710), .ZN(n22711) );
  OAI211_X1 U24311 ( .C1(n22839), .C2(n22713), .A(n22712), .B(n22711), .ZN(
        P1_U3132) );
  AOI22_X1 U24312 ( .A1(n22846), .A2(n22729), .B1(n22775), .B2(n22727), .ZN(
        n22715) );
  AOI22_X1 U24313 ( .A1(n22777), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n22776), .B2(n22728), .ZN(n22714) );
  OAI211_X1 U24314 ( .C1(n22780), .C2(n22732), .A(n22715), .B(n22714), .ZN(
        P1_U3037) );
  OAI22_X1 U24315 ( .A1(n22782), .A2(n22717), .B1(n22781), .B2(n22716), .ZN(
        n22718) );
  INV_X1 U24316 ( .A(n22718), .ZN(n22720) );
  AOI22_X1 U24317 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n22789), .B2(n22728), .ZN(n22719) );
  OAI211_X1 U24318 ( .C1(n22787), .C2(n22732), .A(n22720), .B(n22719), .ZN(
        P1_U3053) );
  AOI22_X1 U24319 ( .A1(n22790), .A2(n22728), .B1(n22727), .B2(n22788), .ZN(
        n22722) );
  AOI22_X1 U24320 ( .A1(n22791), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22789), .B2(n22729), .ZN(n22721) );
  OAI211_X1 U24321 ( .C1(n22794), .C2(n22732), .A(n22722), .B(n22721), .ZN(
        P1_U3061) );
  AOI22_X1 U24322 ( .A1(n22802), .A2(n22729), .B1(n22801), .B2(n22727), .ZN(
        n22724) );
  AOI22_X1 U24323 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22803), .B2(n22728), .ZN(n22723) );
  OAI211_X1 U24324 ( .C1(n22807), .C2(n22732), .A(n22724), .B(n22723), .ZN(
        P1_U3085) );
  AOI22_X1 U24325 ( .A1(n22819), .A2(n22729), .B1(n22765), .B2(n22727), .ZN(
        n22726) );
  AOI22_X1 U24326 ( .A1(n22820), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n22766), .B2(n22728), .ZN(n22725) );
  OAI211_X1 U24327 ( .C1(n22823), .C2(n22732), .A(n22726), .B(n22725), .ZN(
        P1_U3117) );
  AOI22_X1 U24328 ( .A1(n22832), .A2(n22728), .B1(n22831), .B2(n22727), .ZN(
        n22731) );
  AOI22_X1 U24329 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22834), .B2(n22729), .ZN(n22730) );
  OAI211_X1 U24330 ( .C1(n22839), .C2(n22732), .A(n22731), .B(n22730), .ZN(
        P1_U3133) );
  AOI22_X1 U24331 ( .A1(n22846), .A2(n22750), .B1(n22775), .B2(n22748), .ZN(
        n22734) );
  AOI22_X1 U24332 ( .A1(n22777), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n22776), .B2(n22749), .ZN(n22733) );
  OAI211_X1 U24333 ( .C1(n22780), .C2(n22753), .A(n22734), .B(n22733), .ZN(
        P1_U3038) );
  OAI22_X1 U24334 ( .A1(n22782), .A2(n22735), .B1(n22781), .B2(n22743), .ZN(
        n22736) );
  INV_X1 U24335 ( .A(n22736), .ZN(n22738) );
  AOI22_X1 U24336 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n22789), .B2(n22749), .ZN(n22737) );
  OAI211_X1 U24337 ( .C1(n22787), .C2(n22753), .A(n22738), .B(n22737), .ZN(
        P1_U3054) );
  AOI22_X1 U24338 ( .A1(n22790), .A2(n22749), .B1(n22748), .B2(n22788), .ZN(
        n22740) );
  AOI22_X1 U24339 ( .A1(n22791), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22789), .B2(n22750), .ZN(n22739) );
  OAI211_X1 U24340 ( .C1(n22794), .C2(n22753), .A(n22740), .B(n22739), .ZN(
        P1_U3062) );
  AOI22_X1 U24341 ( .A1(n22802), .A2(n22750), .B1(n22801), .B2(n22748), .ZN(
        n22742) );
  AOI22_X1 U24342 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22803), .B2(n22749), .ZN(n22741) );
  OAI211_X1 U24343 ( .C1(n22807), .C2(n22753), .A(n22742), .B(n22741), .ZN(
        P1_U3086) );
  OAI22_X1 U24344 ( .A1(n22830), .A2(n22744), .B1(n22816), .B2(n22743), .ZN(
        n22745) );
  INV_X1 U24345 ( .A(n22745), .ZN(n22747) );
  AOI22_X1 U24346 ( .A1(n22820), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n22819), .B2(n22750), .ZN(n22746) );
  OAI211_X1 U24347 ( .C1(n22823), .C2(n22753), .A(n22747), .B(n22746), .ZN(
        P1_U3118) );
  AOI22_X1 U24348 ( .A1(n22832), .A2(n22749), .B1(n22831), .B2(n22748), .ZN(
        n22752) );
  AOI22_X1 U24349 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22834), .B2(n22750), .ZN(n22751) );
  OAI211_X1 U24350 ( .C1(n22839), .C2(n22753), .A(n22752), .B(n22751), .ZN(
        P1_U3134) );
  AOI22_X1 U24351 ( .A1(n22846), .A2(n22771), .B1(n22775), .B2(n22769), .ZN(
        n22755) );
  AOI22_X1 U24352 ( .A1(n22777), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n22776), .B2(n11150), .ZN(n22754) );
  OAI211_X1 U24353 ( .C1(n22780), .C2(n22774), .A(n22755), .B(n22754), .ZN(
        P1_U3039) );
  OAI22_X1 U24354 ( .A1(n22782), .A2(n22757), .B1(n22781), .B2(n22756), .ZN(
        n22758) );
  INV_X1 U24355 ( .A(n22758), .ZN(n22760) );
  AOI22_X1 U24356 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n22789), .B2(n11150), .ZN(n22759) );
  OAI211_X1 U24357 ( .C1(n22787), .C2(n22774), .A(n22760), .B(n22759), .ZN(
        P1_U3055) );
  AOI22_X1 U24358 ( .A1(n22790), .A2(n11150), .B1(n22769), .B2(n22788), .ZN(
        n22762) );
  AOI22_X1 U24359 ( .A1(n22791), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22789), .B2(n22771), .ZN(n22761) );
  OAI211_X1 U24360 ( .C1(n22794), .C2(n22774), .A(n22762), .B(n22761), .ZN(
        P1_U3063) );
  AOI22_X1 U24361 ( .A1(n11150), .A2(n22803), .B1(n22801), .B2(n22769), .ZN(
        n22764) );
  AOI22_X1 U24362 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22802), .B2(n22771), .ZN(n22763) );
  OAI211_X1 U24363 ( .C1(n22807), .C2(n22774), .A(n22764), .B(n22763), .ZN(
        P1_U3087) );
  AOI22_X1 U24364 ( .A1(n22819), .A2(n22771), .B1(n22765), .B2(n22769), .ZN(
        n22768) );
  AOI22_X1 U24365 ( .A1(n22820), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n22766), .B2(n11150), .ZN(n22767) );
  OAI211_X1 U24366 ( .C1(n22823), .C2(n22774), .A(n22768), .B(n22767), .ZN(
        P1_U3119) );
  AOI22_X1 U24367 ( .A1(n22832), .A2(n11150), .B1(n22831), .B2(n22769), .ZN(
        n22773) );
  AOI22_X1 U24368 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22834), .B2(n22771), .ZN(n22772) );
  OAI211_X1 U24369 ( .C1(n22839), .C2(n22774), .A(n22773), .B(n22772), .ZN(
        P1_U3135) );
  AOI22_X1 U24370 ( .A1(n22846), .A2(n22833), .B1(n22841), .B2(n22775), .ZN(
        n22779) );
  AOI22_X1 U24371 ( .A1(n22777), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n22776), .B2(n22845), .ZN(n22778) );
  OAI211_X1 U24372 ( .C1(n22780), .C2(n22838), .A(n22779), .B(n22778), .ZN(
        P1_U3040) );
  OAI22_X1 U24373 ( .A1(n22782), .A2(n22851), .B1(n22815), .B2(n22781), .ZN(
        n22783) );
  INV_X1 U24374 ( .A(n22783), .ZN(n22786) );
  AOI22_X1 U24375 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n22789), .B2(n22845), .ZN(n22785) );
  OAI211_X1 U24376 ( .C1(n22787), .C2(n22838), .A(n22786), .B(n22785), .ZN(
        P1_U3056) );
  AOI22_X1 U24377 ( .A1(n22789), .A2(n22833), .B1(n22841), .B2(n22788), .ZN(
        n22793) );
  AOI22_X1 U24378 ( .A1(n22791), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22790), .B2(n22845), .ZN(n22792) );
  OAI211_X1 U24379 ( .C1(n22794), .C2(n22838), .A(n22793), .B(n22792), .ZN(
        P1_U3064) );
  AOI22_X1 U24380 ( .A1(n22844), .A2(n22796), .B1(n22841), .B2(n22795), .ZN(
        n22799) );
  AOI22_X1 U24381 ( .A1(n22797), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n22802), .B2(n22845), .ZN(n22798) );
  OAI211_X1 U24382 ( .C1(n22851), .C2(n22800), .A(n22799), .B(n22798), .ZN(
        P1_U3080) );
  AOI22_X1 U24383 ( .A1(n22802), .A2(n22833), .B1(n22841), .B2(n22801), .ZN(
        n22806) );
  AOI22_X1 U24384 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22803), .B2(n22845), .ZN(n22805) );
  OAI211_X1 U24385 ( .C1(n22807), .C2(n22838), .A(n22806), .B(n22805), .ZN(
        P1_U3088) );
  INV_X1 U24386 ( .A(n22808), .ZN(n22810) );
  AOI22_X1 U24387 ( .A1(n22810), .A2(n22844), .B1(n22841), .B2(n22809), .ZN(
        n22813) );
  AOI22_X1 U24388 ( .A1(n22811), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n22819), .B2(n22845), .ZN(n22812) );
  OAI211_X1 U24389 ( .C1(n22851), .C2(n22814), .A(n22813), .B(n22812), .ZN(
        P1_U3112) );
  OAI22_X1 U24390 ( .A1(n22830), .A2(n22817), .B1(n22816), .B2(n22815), .ZN(
        n22818) );
  INV_X1 U24391 ( .A(n22818), .ZN(n22822) );
  AOI22_X1 U24392 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22820), .B1(
        n22819), .B2(n22833), .ZN(n22821) );
  OAI211_X1 U24393 ( .C1(n22823), .C2(n22838), .A(n22822), .B(n22821), .ZN(
        P1_U3120) );
  INV_X1 U24394 ( .A(n22824), .ZN(n22826) );
  AOI22_X1 U24395 ( .A1(n22826), .A2(n22844), .B1(n22841), .B2(n22825), .ZN(
        n22829) );
  AOI22_X1 U24396 ( .A1(n22827), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n22834), .B2(n22845), .ZN(n22828) );
  OAI211_X1 U24397 ( .C1(n22851), .C2(n22830), .A(n22829), .B(n22828), .ZN(
        P1_U3128) );
  AOI22_X1 U24398 ( .A1(n22832), .A2(n22845), .B1(n22831), .B2(n22841), .ZN(
        n22837) );
  AOI22_X1 U24399 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22835), .B1(
        n22834), .B2(n22833), .ZN(n22836) );
  OAI211_X1 U24400 ( .C1(n22839), .C2(n22838), .A(n22837), .B(n22836), .ZN(
        P1_U3136) );
  INV_X1 U24401 ( .A(n22840), .ZN(n22842) );
  AOI22_X1 U24402 ( .A1(n22844), .A2(n22843), .B1(n22842), .B2(n22841), .ZN(
        n22849) );
  AOI22_X1 U24403 ( .A1(n22847), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n22846), .B2(n22845), .ZN(n22848) );
  OAI211_X1 U24404 ( .C1(n22851), .C2(n22850), .A(n22849), .B(n22848), .ZN(
        P1_U3160) );
  INV_X1 U24405 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22854) );
  AOI22_X1 U24406 ( .A1(n22855), .A2(n22854), .B1(n22853), .B2(n22852), .ZN(
        P1_U3486) );
  AND2_X1 U14716 ( .A1(n12887), .A2(n14818), .ZN(n12900) );
  BUF_X1 U11650 ( .A(n12931), .Z(n13759) );
  NAND2_X2 U13825 ( .A1(n12044), .A2(n12079), .ZN(n12062) );
  NAND2_X1 U11346 ( .A1(n12093), .A2(n12092), .ZN(n12095) );
  OR2_X1 U15612 ( .A1(n19515), .A2(n15765), .ZN(n13819) );
  NAND2_X1 U15615 ( .A1(n13819), .A2(n13818), .ZN(n14658) );
  XNOR2_X1 U15616 ( .A(n14658), .B(n13825), .ZN(n14715) );
  AOI221_X1 U11256 ( .B1(n20162), .B2(n20146), .C1(n20162), .C2(n20601), .A(
        n20594), .ZN(n20141) );
  CLKBUF_X1 U11276 ( .A(n18617), .Z(n11157) );
  CLKBUF_X1 U11322 ( .A(n18927), .Z(n11152) );
  CLKBUF_X1 U11324 ( .A(n12460), .Z(n12476) );
  CLKBUF_X1 U11332 ( .A(n17451), .Z(n17452) );
  CLKBUF_X1 U11342 ( .A(n20722), .Z(n20734) );
  CLKBUF_X1 U11343 ( .A(n18146), .Z(n18154) );
  CLKBUF_X2 U11655 ( .A(n12041), .Z(n11259) );
  CLKBUF_X1 U11672 ( .A(n17571), .Z(n17581) );
  CLKBUF_X1 U11724 ( .A(n17633), .Z(n11230) );
  CLKBUF_X1 U11765 ( .A(n18184), .Z(n18192) );
  CLKBUF_X1 U12467 ( .A(n19208), .Z(n19215) );
  CLKBUF_X1 U12470 ( .A(n20987), .Z(n21020) );
  INV_X1 U12524 ( .A(n20709), .ZN(n20736) );
  CLKBUF_X1 U12597 ( .A(n22528), .Z(n22523) );
endmodule

