

module b22_C_gen_AntiSAT_k_256_8 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799;

  NAND2_X2 U7424 ( .A1(n9773), .A2(P3_U3151), .ZN(n13130) );
  AOI21_X1 U7425 ( .B1(n14124), .B2(n14121), .A(n14123), .ZN(n14346) );
  OR2_X1 U7426 ( .A1(n12804), .A2(n12802), .ZN(n12805) );
  AOI21_X1 U7427 ( .B1(n13816), .B2(n11804), .A(n11803), .ZN(n12194) );
  CLKBUF_X1 U7428 ( .A(n13987), .Z(n6884) );
  XNOR2_X1 U7429 ( .A(n7294), .B(n10631), .ZN(n10627) );
  AND2_X1 U7430 ( .A1(n9234), .A2(n9233), .ZN(n11120) );
  CLKBUF_X2 U7431 ( .A(n12358), .Z(n12378) );
  INV_X1 U7434 ( .A(n6690), .ZN(n7283) );
  AND2_X1 U7435 ( .A1(n7246), .A2(n11856), .ZN(n15299) );
  INV_X1 U7436 ( .A(n11858), .ZN(n6999) );
  CLKBUF_X1 U7437 ( .A(n15305), .Z(n6682) );
  INV_X1 U7439 ( .A(n12040), .ZN(n12026) );
  NAND2_X1 U7441 ( .A1(n11734), .A2(n7272), .ZN(n6676) );
  NAND2_X1 U7442 ( .A1(n11734), .A2(n7272), .ZN(n11723) );
  AND2_X2 U7443 ( .A1(n7349), .A2(n7348), .ZN(n10306) );
  INV_X1 U7444 ( .A(n9107), .ZN(n6677) );
  NOR2_X1 U7445 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9106) );
  BUF_X1 U7446 ( .A(n12026), .Z(n12177) );
  XNOR2_X1 U7447 ( .A(n11853), .B(n15305), .ZN(n11858) );
  INV_X1 U7448 ( .A(n11967), .ZN(n11959) );
  INV_X1 U7449 ( .A(n13226), .ZN(n13186) );
  CLKBUF_X2 U7450 ( .A(n10229), .Z(n13226) );
  OR2_X1 U7452 ( .A1(n11079), .A2(n11078), .ZN(n12625) );
  OAI21_X1 U7453 ( .B1(n12896), .B2(n12898), .A(n11924), .ZN(n12890) );
  INV_X1 U7454 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8681) );
  INV_X2 U7455 ( .A(n9571), .ZN(n9587) );
  OR2_X1 U7456 ( .A1(n10051), .A2(n9963), .ZN(n13651) );
  CLKBUF_X2 U7457 ( .A(n7885), .Z(n7922) );
  NOR2_X1 U7458 ( .A1(n14112), .A2(n12178), .ZN(n11808) );
  INV_X1 U7459 ( .A(n14071), .ZN(n14287) );
  AND2_X1 U7460 ( .A1(n7979), .A2(n7978), .ZN(n14846) );
  INV_X1 U7461 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8290) );
  XNOR2_X1 U7462 ( .A(n14502), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14539) );
  AND2_X1 U7463 ( .A1(n7045), .A2(n7282), .ZN(n10197) );
  NAND2_X1 U7464 ( .A1(n9468), .A2(n9467), .ZN(n13718) );
  XNOR2_X1 U7465 ( .A(n13491), .B(n13357), .ZN(n13485) );
  NAND2_X1 U7466 ( .A1(n9643), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9049) );
  BUF_X1 U7467 ( .A(n11814), .Z(n6899) );
  AND4_X1 U7468 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(n12059)
         );
  AOI211_X1 U7469 ( .C1(n12742), .C2(n15259), .A(n12741), .B(n12740), .ZN(
        n12748) );
  XNOR2_X1 U7470 ( .A(n8405), .B(n13117), .ZN(n8411) );
  AND2_X1 U7471 ( .A1(n9425), .A2(n9424), .ZN(n13799) );
  AND2_X1 U7472 ( .A1(n9338), .A2(n9337), .ZN(n13355) );
  XNOR2_X1 U7474 ( .A(n14573), .B(n14574), .ZN(n14709) );
  AND2_X1 U7475 ( .A1(n10259), .A2(n12016), .ZN(n11247) );
  AND2_X2 U7476 ( .A1(n10458), .A2(n15052), .ZN(n15067) );
  AND2_X2 U7477 ( .A1(n10847), .A2(n11120), .ZN(n11129) );
  INV_X1 U7478 ( .A(n10494), .ZN(n6678) );
  INV_X1 U7479 ( .A(n6678), .ZN(n6679) );
  INV_X1 U7480 ( .A(n6678), .ZN(n6680) );
  NAND2_X2 U7481 ( .A1(n7863), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7661) );
  AND3_X2 U7482 ( .A1(n9103), .A2(n9104), .A3(n9102), .ZN(n9118) );
  NAND2_X2 U7483 ( .A1(n8195), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7901) );
  AND2_X2 U7484 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  AND2_X2 U7485 ( .A1(n9393), .A2(n9394), .ZN(n9396) );
  NAND2_X2 U7486 ( .A1(n11041), .A2(n12205), .ZN(n11040) );
  NAND2_X2 U7487 ( .A1(n10546), .A2(n7945), .ZN(n11041) );
  XNOR2_X2 U7488 ( .A(n12021), .B(n7127), .ZN(n12201) );
  INV_X2 U7489 ( .A(n12022), .ZN(n7127) );
  XNOR2_X2 U7490 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14535) );
  NOR2_X2 U7491 ( .A1(n14614), .A2(n12672), .ZN(n12675) );
  NOR2_X2 U7492 ( .A1(n14615), .A2(n14616), .ZN(n14614) );
  OR2_X1 U7493 ( .A1(n7930), .A2(n9797), .ZN(n7919) );
  NOR2_X2 U7494 ( .A1(n11046), .A2(n12052), .ZN(n11094) );
  NAND2_X2 U7495 ( .A1(n7965), .A2(n7964), .ZN(n12052) );
  OR2_X2 U7496 ( .A1(n15240), .A2(n8695), .ZN(n6952) );
  XNOR2_X2 U7497 ( .A(n12702), .B(n12718), .ZN(n12695) );
  INV_X2 U7498 ( .A(n13692), .ZN(n13491) );
  OR2_X1 U7499 ( .A1(n8267), .A2(n11003), .ZN(n7890) );
  XNOR2_X2 U7500 ( .A(n8014), .B(n8013), .ZN(n9841) );
  XNOR2_X2 U7501 ( .A(n8181), .B(n8182), .ZN(n11256) );
  XNOR2_X2 U7502 ( .A(n8184), .B(n10454), .ZN(n8181) );
  NAND2_X1 U7503 ( .A1(n12023), .A2(n12025), .ZN(n12200) );
  INV_X1 U7505 ( .A(n8411), .ZN(n8410) );
  NAND2_X2 U7506 ( .A1(n15215), .A2(n12629), .ZN(n12631) );
  OAI21_X2 U7507 ( .B1(n8227), .B2(n7848), .A(n7847), .ZN(n8239) );
  NOR2_X2 U7508 ( .A1(n14629), .A2(n14628), .ZN(n14627) );
  NOR2_X2 U7509 ( .A1(n10232), .A2(n10231), .ZN(n10319) );
  OAI211_X1 U7510 ( .C1(n9719), .C2(n9692), .A(n8519), .B(n8518), .ZN(n15305)
         );
  OAI21_X2 U7511 ( .B1(n8146), .B2(n7075), .A(n7830), .ZN(n8160) );
  XNOR2_X2 U7512 ( .A(n7829), .B(SI_18_), .ZN(n8146) );
  INV_X1 U7513 ( .A(n12068), .ZN(n12070) );
  OAI22_X2 U7514 ( .A1(n11440), .A2(n11439), .B1(n11438), .B2(n11437), .ZN(
        n11618) );
  NAND2_X2 U7515 ( .A1(n8265), .A2(n8264), .ZN(n14133) );
  OAI21_X2 U7516 ( .B1(n8873), .B2(n8471), .A(n8472), .ZN(n8885) );
  OAI211_X2 U7517 ( .C1(n7891), .C2(n7355), .A(n7893), .B(n7354), .ZN(n10095)
         );
  AND2_X2 U7518 ( .A1(n6972), .A2(n6973), .ZN(n14573) );
  NAND2_X2 U7519 ( .A1(n12694), .A2(n12693), .ZN(n12702) );
  OR2_X2 U7520 ( .A1(n14471), .A2(n8290), .ZN(n7176) );
  XNOR2_X2 U7521 ( .A(n9049), .B(n9644), .ZN(n11827) );
  NOR2_X2 U7522 ( .A1(n10639), .A2(n9743), .ZN(n10638) );
  XNOR2_X2 U7523 ( .A(n9704), .B(n9745), .ZN(n10639) );
  OAI222_X1 U7524 ( .A1(P3_U3151), .A2(n9783), .B1(n13130), .B2(n9782), .C1(
        n11825), .C2(n9781), .ZN(P3_U3294) );
  NAND2_X2 U7525 ( .A1(n7806), .A2(n7805), .ZN(n8014) );
  BUF_X4 U7526 ( .A(n12331), .Z(n6683) );
  NAND2_X1 U7527 ( .A1(n10259), .A2(n10258), .ZN(n12331) );
  NAND2_X1 U7528 ( .A1(n8411), .A2(n13127), .ZN(n8494) );
  XNOR2_X2 U7529 ( .A(n6950), .B(n7217), .ZN(n15169) );
  XNOR2_X2 U7530 ( .A(n12668), .B(n12667), .ZN(n15224) );
  AND2_X2 U7531 ( .A1(n15203), .A2(n12666), .ZN(n12667) );
  AOI21_X2 U7532 ( .B1(n10595), .B2(n10533), .A(n10534), .ZN(n10536) );
  NAND2_X2 U7533 ( .A1(n8028), .A2(n8027), .ZN(n12080) );
  NAND2_X2 U7534 ( .A1(n14500), .A2(n6977), .ZN(n14502) );
  INV_X1 U7535 ( .A(n12651), .ZN(n6684) );
  INV_X1 U7536 ( .A(n8927), .ZN(n12651) );
  MUX2_X1 U7537 ( .A(n12964), .B(n12963), .S(n15396), .Z(n12968) );
  OAI21_X1 U7538 ( .B1(n14346), .B2(n14283), .A(n6891), .ZN(n7119) );
  OR2_X1 U7539 ( .A1(n12779), .A2(n12778), .ZN(n12973) );
  NAND2_X1 U7540 ( .A1(n13904), .A2(n13905), .ZN(n13903) );
  NAND2_X1 U7541 ( .A1(n14191), .A2(n7717), .ZN(n14173) );
  CLKBUF_X1 U7543 ( .A(n12531), .Z(n6912) );
  NAND2_X1 U7544 ( .A1(n14328), .A2(n14327), .ZN(n14326) );
  NAND2_X1 U7545 ( .A1(n12451), .A2(n7558), .ZN(n12611) );
  NAND2_X1 U7546 ( .A1(n12415), .A2(n7559), .ZN(n12451) );
  NAND2_X1 U7547 ( .A1(n8804), .A2(n8461), .ZN(n8812) );
  NAND2_X1 U7548 ( .A1(n9750), .A2(n9751), .ZN(n11057) );
  NOR2_X1 U7549 ( .A1(n10627), .A2(n9744), .ZN(n10626) );
  INV_X1 U7550 ( .A(n14037), .ZN(n11408) );
  INV_X4 U7551 ( .A(n9594), .ZN(n9435) );
  NAND2_X1 U7552 ( .A1(n15312), .A2(n15329), .ZN(n15301) );
  INV_X4 U7553 ( .A(n9593), .ZN(n6685) );
  AND4_X1 U7554 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n10664)
         );
  INV_X4 U7555 ( .A(n10749), .ZN(n13191) );
  NAND2_X1 U7556 ( .A1(n8345), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7899) );
  BUF_X2 U7557 ( .A(n11811), .Z(n6687) );
  INV_X4 U7558 ( .A(n13651), .ZN(n10749) );
  INV_X2 U7559 ( .A(n10950), .ZN(n8507) );
  CLKBUF_X2 U7560 ( .A(n10932), .Z(P3_U3897) );
  AND2_X1 U7561 ( .A1(n8376), .A2(n8383), .ZN(n8377) );
  INV_X1 U7562 ( .A(n7921), .ZN(n11811) );
  NAND2_X2 U7563 ( .A1(n9692), .A2(n9766), .ZN(n8815) );
  INV_X8 U7564 ( .A(n9766), .ZN(n9773) );
  OR2_X1 U7565 ( .A1(n9055), .A2(n9143), .ZN(n9030) );
  AND2_X1 U7566 ( .A1(n7750), .A2(n6944), .ZN(n8293) );
  CLKBUF_X1 U7567 ( .A(n9033), .Z(n9047) );
  INV_X4 U7568 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7569 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8289) );
  OR3_X1 U7570 ( .A1(n12235), .A2(n12199), .A3(n12227), .ZN(n7762) );
  AND2_X1 U7571 ( .A1(n6859), .A2(n6858), .ZN(n14438) );
  NAND2_X1 U7572 ( .A1(n13242), .A2(n7419), .ZN(n13327) );
  NAND2_X1 U7573 ( .A1(n13208), .A2(n13181), .ZN(n13283) );
  OAI21_X1 U7574 ( .B1(n6703), .B2(n6989), .A(n6778), .ZN(n7580) );
  NAND2_X1 U7575 ( .A1(n14173), .A2(n7715), .ZN(n14158) );
  NAND2_X1 U7576 ( .A1(n13443), .A2(n13442), .ZN(n13511) );
  AOI22_X1 U7577 ( .A1(n12520), .A2(n12521), .B1(n12605), .B2(n12444), .ZN(
        n12603) );
  AND2_X1 U7578 ( .A1(n6900), .A2(n13169), .ZN(n13310) );
  NAND2_X1 U7579 ( .A1(n6849), .A2(n13968), .ZN(n13971) );
  NAND2_X1 U7580 ( .A1(n13569), .A2(n13437), .ZN(n13555) );
  NAND2_X1 U7581 ( .A1(n14155), .A2(n8331), .ZN(n14139) );
  NOR2_X1 U7582 ( .A1(n13693), .A2(n7320), .ZN(n7058) );
  NAND2_X1 U7583 ( .A1(n8484), .A2(n8483), .ZN(n13035) );
  NAND2_X1 U7584 ( .A1(n12827), .A2(n12830), .ZN(n12829) );
  NAND2_X1 U7585 ( .A1(n8171), .A2(n8170), .ZN(n14246) );
  NAND2_X1 U7586 ( .A1(n8887), .A2(n8886), .ZN(n12787) );
  OAI211_X1 U7587 ( .C1(n13692), .C2(n13502), .A(n10749), .B(n13487), .ZN(
        n13691) );
  OR3_X1 U7588 ( .A1(n13517), .A2(n13491), .A3(n13503), .ZN(n13487) );
  NAND2_X1 U7589 ( .A1(n13320), .A2(n13152), .ZN(n13216) );
  NAND2_X1 U7590 ( .A1(n8476), .A2(n8475), .ZN(n8899) );
  AND2_X1 U7591 ( .A1(n14435), .A2(n14018), .ZN(n6932) );
  OAI21_X2 U7592 ( .B1(n8325), .B2(n7396), .A(n7394), .ZN(n14222) );
  NAND2_X1 U7593 ( .A1(n8253), .A2(n8252), .ZN(n13987) );
  XNOR2_X1 U7594 ( .A(n13718), .B(n13438), .ZN(n13560) );
  NAND2_X1 U7595 ( .A1(n8817), .A2(n8816), .ZN(n13070) );
  NAND2_X1 U7596 ( .A1(n8241), .A2(n8240), .ZN(n14167) );
  NAND2_X1 U7597 ( .A1(n8229), .A2(n8228), .ZN(n14185) );
  OAI21_X1 U7598 ( .B1(n8239), .B2(n7149), .A(n7147), .ZN(n8263) );
  NAND2_X1 U7599 ( .A1(n12882), .A2(n8800), .ZN(n12881) );
  NAND2_X1 U7600 ( .A1(n8806), .A2(n8805), .ZN(n12876) );
  OAI21_X1 U7601 ( .B1(n8812), .B2(n7586), .A(n7584), .ZN(n8838) );
  XNOR2_X1 U7602 ( .A(n7846), .B(SI_24_), .ZN(n8227) );
  NAND2_X1 U7603 ( .A1(n13893), .A2(n12255), .ZN(n13958) );
  INV_X1 U7604 ( .A(n14211), .ZN(n14454) );
  AOI21_X1 U7605 ( .B1(n9269), .B2(n6743), .A(n7505), .ZN(n9303) );
  XNOR2_X1 U7606 ( .A(n8189), .B(n8188), .ZN(n11341) );
  NAND2_X1 U7607 ( .A1(n6952), .A2(n6737), .ZN(n7224) );
  NAND2_X1 U7608 ( .A1(n8173), .A2(n8172), .ZN(n14251) );
  OAI21_X1 U7609 ( .B1(n12935), .B2(n8734), .A(n8735), .ZN(n12924) );
  NAND2_X1 U7610 ( .A1(n8460), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U7611 ( .A1(n7121), .A2(n6693), .ZN(n11463) );
  NAND2_X1 U7612 ( .A1(n15156), .A2(n12403), .ZN(n12404) );
  NAND2_X1 U7613 ( .A1(n8785), .A2(n8459), .ZN(n8460) );
  NAND2_X1 U7614 ( .A1(n8106), .A2(n8105), .ZN(n14421) );
  NAND2_X1 U7615 ( .A1(n8783), .A2(n8782), .ZN(n8785) );
  OAI21_X1 U7616 ( .B1(n7402), .B2(n7399), .A(n7397), .ZN(n11185) );
  NOR2_X1 U7617 ( .A1(n15189), .A2(n14650), .ZN(n15188) );
  NAND2_X1 U7618 ( .A1(n8769), .A2(n8768), .ZN(n8771) );
  INV_X1 U7619 ( .A(n11486), .ZN(n11489) );
  NOR2_X1 U7620 ( .A1(n8654), .A2(n15198), .ZN(n15197) );
  AND2_X1 U7621 ( .A1(n9273), .A2(n9272), .ZN(n11486) );
  NAND2_X1 U7622 ( .A1(n8045), .A2(n8044), .ZN(n12246) );
  NAND2_X1 U7623 ( .A1(n8076), .A2(n8075), .ZN(n14681) );
  XNOR2_X1 U7624 ( .A(n12661), .B(n12660), .ZN(n15189) );
  OR2_X1 U7625 ( .A1(n10853), .A2(n7303), .ZN(n7302) );
  NAND2_X1 U7626 ( .A1(n11057), .A2(n11056), .ZN(n15178) );
  AND2_X1 U7627 ( .A1(n6851), .A2(n6850), .ZN(n11440) );
  XNOR2_X1 U7628 ( .A(n8023), .B(n8022), .ZN(n9847) );
  NAND2_X1 U7629 ( .A1(n9257), .A2(n9256), .ZN(n11283) );
  NAND2_X1 U7630 ( .A1(n10871), .A2(n10870), .ZN(n10869) );
  NAND2_X1 U7631 ( .A1(n10819), .A2(n10818), .ZN(n10853) );
  NAND2_X1 U7632 ( .A1(n7064), .A2(n7062), .ZN(n8089) );
  OAI21_X1 U7633 ( .B1(n7065), .B2(n7066), .A(n7806), .ZN(n7064) );
  NOR2_X1 U7634 ( .A1(n14739), .A2(n14738), .ZN(n14737) );
  XNOR2_X1 U7635 ( .A(n8002), .B(n8001), .ZN(n9837) );
  NAND2_X1 U7636 ( .A1(n7992), .A2(n7991), .ZN(n12063) );
  NAND2_X1 U7637 ( .A1(n7293), .A2(n7292), .ZN(n11062) );
  OAI21_X2 U7638 ( .B1(n9966), .B2(n10645), .A(n15052), .ZN(n9967) );
  NAND2_X1 U7639 ( .A1(n8677), .A2(n8676), .ZN(n8679) );
  OAI22_X1 U7640 ( .A1(n7068), .A2(n6771), .B1(n7134), .B2(n6712), .ZN(n7063)
         );
  NOR2_X1 U7641 ( .A1(n15394), .A2(n15339), .ZN(n13016) );
  OAI211_X1 U7642 ( .C1(n12029), .C2(n7178), .A(n12202), .B(n12028), .ZN(n7177) );
  AND2_X1 U7643 ( .A1(n11865), .A2(n11862), .ZN(n11977) );
  AND2_X1 U7644 ( .A1(n9162), .A2(n9161), .ZN(n10661) );
  CLKBUF_X1 U7645 ( .A(n10381), .Z(n6878) );
  INV_X2 U7646 ( .A(n12484), .ZN(n12435) );
  NAND2_X1 U7647 ( .A1(n6874), .A2(n7789), .ZN(n7947) );
  CLKBUF_X1 U7648 ( .A(n14039), .Z(n6871) );
  INV_X1 U7649 ( .A(n14039), .ZN(n10788) );
  BUF_X1 U7650 ( .A(n7933), .Z(n12033) );
  INV_X1 U7651 ( .A(n10339), .ZN(n10963) );
  NAND4_X2 U7652 ( .A1(n8513), .A2(n8512), .A3(n8511), .A4(n8510), .ZN(n11853)
         );
  INV_X1 U7653 ( .A(n12059), .ZN(n14035) );
  NAND4_X1 U7654 ( .A1(n7927), .A2(n7926), .A3(n7925), .A4(n7924), .ZN(n14039)
         );
  NAND2_X1 U7655 ( .A1(n8615), .A2(n8614), .ZN(n8617) );
  AND2_X1 U7656 ( .A1(n7347), .A2(n7346), .ZN(n10131) );
  NAND2_X2 U7657 ( .A1(n8378), .A2(n8377), .ZN(n10259) );
  NAND2_X1 U7658 ( .A1(n6947), .A2(n14542), .ZN(n14546) );
  AND2_X1 U7659 ( .A1(n9562), .A2(n9661), .ZN(n10459) );
  AND3_X1 U7660 ( .A1(n8531), .A2(n8530), .A3(n8529), .ZN(n10764) );
  INV_X1 U7661 ( .A(n9428), .ZN(n9569) );
  NAND2_X2 U7662 ( .A1(n8410), .A2(n8409), .ZN(n8905) );
  NAND2_X1 U7663 ( .A1(n8411), .A2(n8409), .ZN(n8795) );
  INV_X2 U7664 ( .A(n8363), .ZN(n14423) );
  NAND2_X1 U7665 ( .A1(n9093), .A2(n9092), .ZN(n13375) );
  AND2_X1 U7666 ( .A1(n9562), .A2(n11827), .ZN(n9095) );
  OAI21_X1 U7667 ( .B1(n8580), .B2(n7592), .A(n7589), .ZN(n8615) );
  CLKBUF_X1 U7668 ( .A(n7923), .Z(n6943) );
  INV_X1 U7669 ( .A(n9111), .ZN(n9428) );
  NAND2_X1 U7670 ( .A1(n8429), .A2(n8428), .ZN(n8580) );
  INV_X1 U7671 ( .A(n9109), .ZN(n9567) );
  NOR2_X1 U7672 ( .A1(n8948), .A2(n11481), .ZN(n11798) );
  NAND2_X1 U7673 ( .A1(n8915), .A2(n8914), .ZN(n10677) );
  NOR2_X1 U7674 ( .A1(n8340), .A2(n12014), .ZN(n8363) );
  XNOR2_X1 U7675 ( .A(n8357), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8376) );
  INV_X2 U7676 ( .A(n13123), .ZN(n11825) );
  OR2_X1 U7677 ( .A1(n10593), .A2(n11018), .ZN(n10595) );
  NAND2_X1 U7678 ( .A1(n8919), .A2(n8918), .ZN(n10494) );
  INV_X1 U7679 ( .A(n12189), .ZN(n14496) );
  NAND2_X1 U7680 ( .A1(n9036), .A2(n9042), .ZN(n11268) );
  NAND2_X1 U7681 ( .A1(n12183), .A2(n12188), .ZN(n12016) );
  XNOR2_X1 U7682 ( .A(n8788), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12742) );
  AND2_X2 U7683 ( .A1(n9643), .A2(n9048), .ZN(n9661) );
  NAND2_X2 U7684 ( .A1(n9773), .A2(P2_U3088), .ZN(n13837) );
  NAND2_X1 U7685 ( .A1(n8352), .A2(n8294), .ZN(n12189) );
  XNOR2_X1 U7686 ( .A(n7792), .B(SI_5_), .ZN(n7946) );
  XNOR2_X1 U7687 ( .A(n7870), .B(n7869), .ZN(n14481) );
  XNOR2_X1 U7688 ( .A(n7788), .B(SI_4_), .ZN(n7939) );
  XNOR2_X1 U7689 ( .A(n8298), .B(n8297), .ZN(n12188) );
  MUX2_X1 U7690 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9043), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n9048) );
  NAND2_X1 U7691 ( .A1(n8293), .A2(n8292), .ZN(n8352) );
  NAND2_X1 U7692 ( .A1(n9047), .A2(n9046), .ZN(n9643) );
  NAND2_X1 U7693 ( .A1(n7159), .A2(SI_0_), .ZN(n7894) );
  NAND2_X1 U7694 ( .A1(n8946), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8482) );
  XNOR2_X1 U7695 ( .A(n6956), .B(n7862), .ZN(n14488) );
  OAI21_X1 U7696 ( .B1(n8161), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7688) );
  OR2_X1 U7697 ( .A1(n7867), .A2(n8290), .ZN(n7861) );
  NAND2_X1 U7698 ( .A1(n7915), .A2(n7914), .ZN(n10097) );
  OR2_X1 U7699 ( .A1(n10394), .A2(n9710), .ZN(n10395) );
  NOR2_X1 U7700 ( .A1(n10078), .A2(n10264), .ZN(n10086) );
  AND2_X1 U7701 ( .A1(n6984), .A2(n8740), .ZN(n7760) );
  OR2_X1 U7702 ( .A1(n10397), .A2(n9711), .ZN(n10399) );
  AND3_X2 U7703 ( .A1(n7310), .A2(n7311), .A3(n7309), .ZN(n9719) );
  AND2_X1 U7704 ( .A1(n8420), .A2(n8419), .ZN(n8515) );
  NOR2_X1 U7705 ( .A1(n7753), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n7752) );
  AND2_X1 U7706 ( .A1(n9029), .A2(n9028), .ZN(n7418) );
  AND2_X1 U7707 ( .A1(n9678), .A2(n8401), .ZN(n7277) );
  AND3_X1 U7708 ( .A1(n8400), .A2(n8560), .A3(n7535), .ZN(n7534) );
  NAND2_X1 U7709 ( .A1(n9771), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8420) );
  AND3_X1 U7710 ( .A1(n9021), .A2(n9020), .A3(n9654), .ZN(n9029) );
  AND2_X1 U7711 ( .A1(n6869), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14536) );
  AND2_X1 U7712 ( .A1(n9018), .A2(n9017), .ZN(n9039) );
  AND3_X1 U7713 ( .A1(n6983), .A2(n6982), .A3(n6981), .ZN(n8740) );
  AND3_X1 U7714 ( .A1(n9106), .A2(n9016), .A3(n9014), .ZN(n7479) );
  NOR2_X1 U7715 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n6986) );
  INV_X1 U7716 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7035) );
  NOR2_X1 U7717 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n6983) );
  INV_X4 U7718 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7719 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n6982) );
  INV_X1 U7720 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n12731) );
  NOR2_X1 U7721 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n6981) );
  INV_X1 U7722 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13405) );
  INV_X1 U7723 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14075) );
  NOR2_X1 U7724 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9011) );
  NOR2_X1 U7725 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n6988) );
  NOR2_X1 U7726 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n6987) );
  INV_X1 U7727 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7771) );
  NOR2_X2 U7728 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7892) );
  INV_X1 U7729 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9654) );
  INV_X1 U7730 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9649) );
  INV_X1 U7731 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n15553) );
  INV_X1 U7732 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n15698) );
  NOR2_X1 U7733 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n9021) );
  INV_X2 U7734 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8003) );
  INV_X4 U7735 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7736 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n9020) );
  INV_X1 U7737 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8560) );
  INV_X1 U7738 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8061) );
  NOR2_X2 U7739 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n9678) );
  NOR2_X1 U7740 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n9018) );
  NOR2_X2 U7741 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8058) );
  INV_X1 U7742 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U7743 ( .A1(n10459), .A2(n11827), .ZN(n9617) );
  AND4_X2 U7744 ( .A1(n7386), .A2(n7859), .A3(n7860), .A4(n7858), .ZN(n6724)
         );
  AND3_X1 U7745 ( .A1(n7760), .A2(n6934), .A3(n8612), .ZN(n8941) );
  AND3_X4 U7746 ( .A1(n7277), .A2(n7534), .A3(n7533), .ZN(n8612) );
  XNOR2_X2 U7747 ( .A(n13445), .B(n13485), .ZN(n13446) );
  NAND2_X1 U7748 ( .A1(n7868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7870) );
  NAND3_X2 U7749 ( .A1(n7897), .A2(n7896), .A3(n6793), .ZN(n6967) );
  XNOR2_X2 U7750 ( .A(n12717), .B(n12718), .ZN(n12684) );
  NAND2_X2 U7751 ( .A1(n12683), .A2(n12682), .ZN(n12717) );
  NAND2_X2 U7752 ( .A1(n10869), .A2(n8000), .ZN(n11025) );
  OAI21_X2 U7753 ( .B1(n10792), .B2(n7738), .A(n7736), .ZN(n11243) );
  OAI21_X2 U7754 ( .B1(n8184), .B2(n7141), .A(n7840), .ZN(n7841) );
  OAI21_X2 U7755 ( .B1(n8160), .B2(n8159), .A(n7834), .ZN(n8184) );
  NOR2_X2 U7756 ( .A1(n10224), .A2(n10963), .ZN(n10223) );
  AOI22_X2 U7757 ( .A1(n15191), .A2(n15190), .B1(n12660), .B2(n12645), .ZN(
        n15210) );
  NAND2_X4 U7758 ( .A1(n14488), .A2(n14483), .ZN(n8204) );
  AOI21_X2 U7759 ( .B1(n14970), .B2(n14567), .A(n14606), .ZN(n14706) );
  AND4_X2 U7760 ( .A1(n7890), .A2(n7889), .A3(n7888), .A4(n7887), .ZN(n7904)
         );
  OR2_X1 U7761 ( .A1(n7921), .A2(n7886), .ZN(n7887) );
  NOR2_X2 U7762 ( .A1(n7868), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n14471) );
  OAI211_X1 U7763 ( .C1(n9650), .C2(P2_IR_REG_27__SCAN_IN), .A(n9031), .B(
        n9662), .ZN(n6689) );
  OAI211_X2 U7764 ( .C1(n9650), .C2(P2_IR_REG_27__SCAN_IN), .A(n9031), .B(
        n9662), .ZN(n6690) );
  INV_X1 U7765 ( .A(n6689), .ZN(n9397) );
  NAND2_X1 U7766 ( .A1(n7872), .A2(n7871), .ZN(n8267) );
  NOR2_X4 U7767 ( .A1(n11463), .A2(n14681), .ZN(n11464) );
  NOR2_X1 U7769 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8401) );
  AOI21_X1 U7770 ( .B1(n7513), .B2(n7512), .A(n9283), .ZN(n7511) );
  OR2_X1 U7771 ( .A1(n11931), .A2(n11932), .ZN(n7018) );
  AOI21_X1 U7772 ( .B1(n7031), .B2(n7029), .A(n6775), .ZN(n7028) );
  INV_X1 U7773 ( .A(n11947), .ZN(n7029) );
  INV_X1 U7774 ( .A(n13127), .ZN(n8409) );
  OR2_X1 U7775 ( .A1(n13070), .A2(n8824), .ZN(n11942) );
  AND2_X1 U7776 ( .A1(n6691), .A2(n7054), .ZN(n7053) );
  INV_X1 U7777 ( .A(n10791), .ZN(n7741) );
  NOR2_X1 U7778 ( .A1(n14209), .A2(n7116), .ZN(n7115) );
  INV_X1 U7779 ( .A(n8327), .ZN(n7116) );
  OR2_X1 U7780 ( .A1(n14421), .A2(n14315), .ZN(n12100) );
  AOI21_X1 U7781 ( .B1(n6830), .B2(n7148), .A(n6719), .ZN(n7147) );
  NAND2_X1 U7782 ( .A1(n7150), .A2(n6830), .ZN(n7149) );
  NAND2_X1 U7783 ( .A1(n12484), .A2(n15329), .ZN(n10497) );
  INV_X1 U7784 ( .A(n8795), .ZN(n8832) );
  INV_X2 U7785 ( .A(n8832), .ZN(n10953) );
  AND2_X1 U7786 ( .A1(n8612), .A2(n8642), .ZN(n8741) );
  AND2_X1 U7787 ( .A1(n11985), .A2(n8668), .ZN(n7272) );
  OR2_X1 U7788 ( .A1(n12987), .A2(n12579), .ZN(n11950) );
  NAND2_X1 U7789 ( .A1(n13434), .A2(n7343), .ZN(n7342) );
  NOR2_X1 U7790 ( .A1(n13588), .A2(n7344), .ZN(n7343) );
  INV_X1 U7791 ( .A(n13433), .ZN(n7344) );
  OR2_X1 U7792 ( .A1(n13503), .A2(n13447), .ZN(n13444) );
  NAND2_X1 U7793 ( .A1(n14111), .A2(n8338), .ZN(n14112) );
  OR2_X1 U7794 ( .A1(n14596), .A2(n14595), .ZN(n6925) );
  NAND2_X1 U7795 ( .A1(n12027), .A2(n7681), .ZN(n12028) );
  NAND2_X1 U7796 ( .A1(n12024), .A2(n12026), .ZN(n12027) );
  NAND2_X1 U7797 ( .A1(n12048), .A2(n12051), .ZN(n7174) );
  NAND2_X1 U7798 ( .A1(n7490), .A2(n7486), .ZN(n7491) );
  AND2_X1 U7799 ( .A1(n7488), .A2(n7487), .ZN(n7486) );
  AOI22_X1 U7800 ( .A1(n9195), .A2(n9194), .B1(n9193), .B2(n9192), .ZN(n9211)
         );
  OR2_X1 U7801 ( .A1(n11864), .A2(n11967), .ZN(n6995) );
  AND2_X1 U7802 ( .A1(n9266), .A2(n9267), .ZN(n7513) );
  OAI22_X1 U7803 ( .A1(n11486), .A2(n9344), .B1(n11279), .B2(n6685), .ZN(n9282) );
  NAND2_X1 U7804 ( .A1(n9268), .A2(n7514), .ZN(n7512) );
  INV_X1 U7805 ( .A(n9333), .ZN(n7518) );
  NOR2_X1 U7806 ( .A1(n7495), .A2(n7496), .ZN(n7494) );
  NAND2_X1 U7807 ( .A1(n6713), .A2(n7018), .ZN(n7013) );
  NAND2_X1 U7808 ( .A1(n7016), .A2(n7019), .ZN(n7015) );
  AND2_X1 U7809 ( .A1(n7032), .A2(n7024), .ZN(n7023) );
  AND2_X1 U7810 ( .A1(n11955), .A2(n12802), .ZN(n7032) );
  NAND2_X1 U7811 ( .A1(n12176), .A2(n12174), .ZN(n7672) );
  AND2_X1 U7812 ( .A1(n7646), .A2(n6736), .ZN(n7645) );
  NAND2_X1 U7813 ( .A1(n11493), .A2(n8984), .ZN(n8988) );
  NAND2_X1 U7814 ( .A1(n7655), .A2(n7809), .ZN(n7654) );
  INV_X1 U7815 ( .A(n8022), .ZN(n7655) );
  INV_X1 U7816 ( .A(n7653), .ZN(n7652) );
  OAI21_X1 U7817 ( .B1(n7654), .B2(n7807), .A(n7813), .ZN(n7653) );
  NAND2_X1 U7818 ( .A1(n7810), .A2(n9800), .ZN(n7813) );
  NAND2_X1 U7819 ( .A1(n11062), .A2(n11061), .ZN(n6950) );
  NAND2_X1 U7820 ( .A1(n11073), .A2(n11072), .ZN(n7218) );
  NAND2_X1 U7821 ( .A1(n15309), .A2(n11858), .ZN(n7260) );
  NAND2_X1 U7822 ( .A1(n10280), .A2(n15340), .ZN(n7246) );
  NAND2_X1 U7823 ( .A1(n7259), .A2(n7257), .ZN(n12780) );
  INV_X1 U7824 ( .A(n8825), .ZN(n7251) );
  INV_X1 U7825 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U7826 ( .A1(n9770), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U7827 ( .A1(n10745), .A2(n10746), .ZN(n7457) );
  NOR2_X1 U7828 ( .A1(n11139), .A2(n10937), .ZN(n7468) );
  AND2_X1 U7829 ( .A1(n13140), .A2(n7448), .ZN(n7441) );
  AND2_X1 U7830 ( .A1(n11268), .A2(n9661), .ZN(n9922) );
  NOR2_X1 U7831 ( .A1(n13406), .A2(n13410), .ZN(n9614) );
  NAND2_X1 U7832 ( .A1(n13821), .A2(n9090), .ZN(n9111) );
  NOR2_X1 U7833 ( .A1(n13464), .A2(n7055), .ZN(n7054) );
  INV_X1 U7834 ( .A(n13463), .ZN(n7055) );
  AND2_X1 U7835 ( .A1(n7377), .A2(n13588), .ZN(n7376) );
  INV_X1 U7836 ( .A(n7768), .ZN(n7377) );
  OR2_X1 U7837 ( .A1(n13741), .A2(n13462), .ZN(n13430) );
  INV_X1 U7838 ( .A(n7368), .ZN(n7048) );
  AOI21_X1 U7839 ( .B1(n7370), .B2(n13662), .A(n6753), .ZN(n7368) );
  NAND2_X1 U7840 ( .A1(n7359), .A2(n7357), .ZN(n11285) );
  AOI21_X1 U7841 ( .B1(n7360), .B2(n10821), .A(n7358), .ZN(n7357) );
  OAI21_X1 U7842 ( .B1(n10799), .B2(n10812), .A(n10798), .ZN(n7367) );
  NAND2_X1 U7843 ( .A1(n13882), .A2(n13967), .ZN(n6849) );
  NAND2_X1 U7844 ( .A1(n7741), .A2(n6732), .ZN(n7738) );
  NOR2_X1 U7845 ( .A1(n14157), .A2(n7716), .ZN(n7715) );
  INV_X1 U7846 ( .A(n8237), .ZN(n7716) );
  AOI21_X1 U7847 ( .B1(n7093), .B2(n7097), .A(n7092), .ZN(n7091) );
  NAND2_X1 U7848 ( .A1(n11468), .A2(n7095), .ZN(n7094) );
  INV_X1 U7849 ( .A(n12100), .ZN(n7092) );
  AOI21_X1 U7850 ( .B1(n7853), .B2(n7671), .A(n7669), .ZN(n7668) );
  INV_X1 U7851 ( .A(n8277), .ZN(n7669) );
  INV_X1 U7852 ( .A(n6872), .ZN(n7975) );
  INV_X1 U7853 ( .A(n8117), .ZN(n7648) );
  INV_X1 U7854 ( .A(n7988), .ZN(n7800) );
  INV_X1 U7855 ( .A(n7958), .ZN(n7794) );
  NAND2_X1 U7856 ( .A1(n14513), .A2(n14512), .ZN(n14558) );
  OR2_X1 U7857 ( .A1(n14554), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14512) );
  INV_X1 U7858 ( .A(n7543), .ZN(n7542) );
  OAI21_X1 U7859 ( .B1(n11299), .B2(n7544), .A(n15136), .ZN(n7543) );
  OAI21_X1 U7860 ( .B1(n6817), .B2(n6695), .A(n7551), .ZN(n7550) );
  NAND2_X1 U7861 ( .A1(n6695), .A2(n7552), .ZN(n7551) );
  NAND2_X1 U7862 ( .A1(n7554), .A2(n6694), .ZN(n7552) );
  XNOR2_X1 U7863 ( .A(n15340), .B(n12484), .ZN(n10498) );
  NAND2_X1 U7864 ( .A1(n12611), .A2(n12421), .ZN(n12531) );
  AND4_X1 U7865 ( .A1(n8780), .A2(n8779), .A3(n8778), .A4(n8777), .ZN(n12543)
         );
  OR2_X1 U7866 ( .A1(n10953), .A2(n11058), .ZN(n8625) );
  AND4_X1 U7867 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(n15131)
         );
  OR2_X1 U7868 ( .A1(n8795), .A2(n15392), .ZN(n8606) );
  NAND2_X1 U7869 ( .A1(n9678), .A2(n8402), .ZN(n7311) );
  OR2_X1 U7870 ( .A1(n7311), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8543) );
  INV_X1 U7871 ( .A(n12522), .ZN(n12833) );
  INV_X1 U7872 ( .A(n12936), .ZN(n14640) );
  NAND2_X1 U7873 ( .A1(n11606), .A2(n6742), .ZN(n11734) );
  XNOR2_X1 U7874 ( .A(n12401), .B(n15153), .ZN(n11982) );
  NAND2_X1 U7875 ( .A1(n8930), .A2(n11959), .ZN(n15313) );
  NOR2_X1 U7876 ( .A1(n12820), .A2(n7623), .ZN(n7622) );
  INV_X1 U7877 ( .A(n11950), .ZN(n7623) );
  AOI21_X1 U7878 ( .B1(n7618), .B2(n7617), .A(n7616), .ZN(n7615) );
  INV_X1 U7879 ( .A(n11937), .ZN(n7617) );
  INV_X1 U7880 ( .A(n11942), .ZN(n7616) );
  OR2_X1 U7881 ( .A1(n12876), .A2(n12474), .ZN(n11937) );
  OAI21_X1 U7882 ( .B1(n12924), .B2(n12921), .A(n8753), .ZN(n12910) );
  INV_X1 U7883 ( .A(n8517), .ZN(n8790) );
  INV_X1 U7884 ( .A(n9692), .ZN(n8789) );
  INV_X1 U7885 ( .A(n8815), .ZN(n11840) );
  OAI22_X1 U7886 ( .A1(n11832), .A2(n11831), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n13824), .ZN(n11837) );
  NOR2_X1 U7887 ( .A1(n7263), .A2(n7262), .ZN(n7261) );
  AND2_X1 U7888 ( .A1(n6807), .A2(n7265), .ZN(n7264) );
  NAND2_X1 U7889 ( .A1(n8470), .A2(n8469), .ZN(n8873) );
  NAND2_X1 U7890 ( .A1(n8741), .A2(n6731), .ZN(n8757) );
  NAND2_X1 U7891 ( .A1(n8741), .A2(n7560), .ZN(n8786) );
  AND2_X1 U7892 ( .A1(n6731), .A2(n8758), .ZN(n7560) );
  NOR2_X1 U7893 ( .A1(n8543), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8561) );
  INV_X1 U7894 ( .A(n7425), .ZN(n7424) );
  OAI21_X1 U7895 ( .B1(n13200), .B2(n7428), .A(n7426), .ZN(n7425) );
  NAND2_X1 U7896 ( .A1(n7429), .A2(n7427), .ZN(n7426) );
  INV_X1 U7897 ( .A(n13224), .ZN(n7427) );
  OAI22_X1 U7898 ( .A1(n9818), .A2(n9766), .B1(n7662), .B2(n7845), .ZN(n7284)
         );
  NAND2_X1 U7899 ( .A1(n7469), .A2(n6832), .ZN(n7464) );
  NAND2_X1 U7900 ( .A1(n13444), .A2(n9624), .ZN(n13481) );
  XNOR2_X1 U7901 ( .A(n13522), .B(n13358), .ZN(n13514) );
  NAND2_X1 U7902 ( .A1(n7342), .A2(n7340), .ZN(n13569) );
  NOR2_X1 U7903 ( .A1(n13579), .A2(n7341), .ZN(n7340) );
  INV_X1 U7904 ( .A(n13436), .ZN(n7341) );
  NAND2_X1 U7905 ( .A1(n13599), .A2(n13431), .ZN(n13434) );
  OAI21_X1 U7906 ( .B1(n11325), .B2(n13364), .A(n11489), .ZN(n11287) );
  NAND2_X1 U7907 ( .A1(n7365), .A2(n10802), .ZN(n7038) );
  NOR2_X1 U7908 ( .A1(n7042), .A2(n7039), .ZN(n7037) );
  NAND2_X1 U7909 ( .A1(n7040), .A2(n7043), .ZN(n15059) );
  INV_X1 U7910 ( .A(n7365), .ZN(n7043) );
  NAND2_X1 U7911 ( .A1(n10799), .A2(n7041), .ZN(n7040) );
  NAND2_X1 U7912 ( .A1(n6689), .A2(n9773), .ZN(n9555) );
  INV_X1 U7914 ( .A(n9142), .ZN(n9255) );
  NAND2_X1 U7915 ( .A1(n6689), .A2(n9766), .ZN(n9142) );
  INV_X1 U7916 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9054) );
  NAND2_X1 U7917 ( .A1(n6848), .A2(n7743), .ZN(n7737) );
  AND2_X1 U7918 ( .A1(n13843), .A2(n7735), .ZN(n7734) );
  OR2_X1 U7919 ( .A1(n13990), .A2(n12366), .ZN(n7735) );
  AOI21_X1 U7920 ( .B1(n13865), .B2(n7730), .A(n7729), .ZN(n7728) );
  INV_X1 U7921 ( .A(n13866), .ZN(n7730) );
  INV_X1 U7922 ( .A(n12339), .ZN(n7729) );
  INV_X1 U7923 ( .A(n11808), .ZN(n14079) );
  NAND2_X1 U7924 ( .A1(n14145), .A2(n14142), .ZN(n7714) );
  AOI21_X1 U7925 ( .B1(n7115), .B2(n14225), .A(n6782), .ZN(n7113) );
  INV_X1 U7926 ( .A(n7115), .ZN(n7114) );
  AOI21_X1 U7927 ( .B1(n7395), .B2(n14262), .A(n6770), .ZN(n7394) );
  NAND2_X1 U7928 ( .A1(n9847), .A2(n11804), .ZN(n8028) );
  NAND2_X1 U7929 ( .A1(n13828), .A2(n7941), .ZN(n8265) );
  INV_X1 U7930 ( .A(n14202), .ZN(n14372) );
  OR2_X1 U7931 ( .A1(n9552), .A2(n9551), .ZN(n9554) );
  NAND2_X1 U7932 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6928), .ZN(n6927) );
  INV_X1 U7933 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6928) );
  AOI21_X1 U7934 ( .B1(n12773), .B2(n8894), .A(n8415), .ZN(n12782) );
  NAND2_X1 U7935 ( .A1(n13244), .A2(n13243), .ZN(n13242) );
  AND2_X1 U7936 ( .A1(n14130), .A2(n14131), .ZN(n6891) );
  NAND2_X1 U7937 ( .A1(n6946), .A2(n14538), .ZN(n14596) );
  NOR2_X1 U7938 ( .A1(n7181), .A2(n7180), .ZN(n7179) );
  INV_X1 U7939 ( .A(n12037), .ZN(n7180) );
  OR2_X1 U7940 ( .A1(n12051), .A2(n12048), .ZN(n7175) );
  OR2_X1 U7941 ( .A1(n9925), .A2(n9617), .ZN(n9115) );
  OR2_X1 U7942 ( .A1(n12055), .A2(n12056), .ZN(n12057) );
  NAND2_X1 U7943 ( .A1(n12071), .A2(n12072), .ZN(n7193) );
  INV_X1 U7944 ( .A(n9135), .ZN(n7478) );
  INV_X1 U7945 ( .A(n7191), .ZN(n7188) );
  AND2_X1 U7946 ( .A1(n9172), .A2(n9174), .ZN(n7485) );
  NAND2_X1 U7947 ( .A1(n9171), .A2(n7489), .ZN(n7488) );
  INV_X1 U7948 ( .A(n9174), .ZN(n7489) );
  AND2_X1 U7949 ( .A1(n6697), .A2(n7674), .ZN(n7196) );
  NAND2_X1 U7950 ( .A1(n12094), .A2(n6760), .ZN(n7674) );
  OAI21_X1 U7951 ( .B1(n6997), .B2(n11863), .A(n11862), .ZN(n6996) );
  NOR2_X1 U7952 ( .A1(n11857), .A2(n6998), .ZN(n6997) );
  INV_X1 U7953 ( .A(n9243), .ZN(n9246) );
  INV_X1 U7954 ( .A(n9284), .ZN(n7508) );
  INV_X1 U7955 ( .A(n7512), .ZN(n7509) );
  OAI21_X1 U7956 ( .B1(n11876), .B2(n11967), .A(n7005), .ZN(n7004) );
  AOI21_X1 U7957 ( .B1(n6758), .B2(n11967), .A(n7006), .ZN(n7005) );
  NAND2_X1 U7958 ( .A1(n12155), .A2(n7200), .ZN(n7199) );
  INV_X1 U7959 ( .A(n12154), .ZN(n7200) );
  NAND2_X1 U7960 ( .A1(n7518), .A2(n7517), .ZN(n7516) );
  MUX2_X1 U7961 ( .A(n11946), .B(n11945), .S(n11967), .Z(n11947) );
  NAND2_X1 U7962 ( .A1(n7013), .A2(n7014), .ZN(n7010) );
  NAND2_X1 U7963 ( .A1(n7018), .A2(n6708), .ZN(n7014) );
  AOI21_X1 U7964 ( .B1(n11947), .B2(n12845), .A(n11992), .ZN(n7031) );
  INV_X1 U7965 ( .A(n13588), .ZN(n7085) );
  NOR2_X1 U7966 ( .A1(n13620), .A2(n7082), .ZN(n7081) );
  NAND2_X1 U7967 ( .A1(n7084), .A2(n7083), .ZN(n7082) );
  NOR2_X1 U7968 ( .A1(n9637), .A2(n13646), .ZN(n7083) );
  NOR2_X1 U7969 ( .A1(n6716), .A2(n7642), .ZN(n7640) );
  AOI21_X1 U7970 ( .B1(n7023), .B2(n7026), .A(n6787), .ZN(n7021) );
  NAND2_X1 U7971 ( .A1(n7582), .A2(n11967), .ZN(n7581) );
  INV_X1 U7972 ( .A(n11965), .ZN(n7582) );
  INV_X1 U7973 ( .A(n7186), .ZN(n7162) );
  NOR3_X1 U7974 ( .A1(n7658), .A2(n12223), .A3(n8287), .ZN(n7657) );
  NAND2_X1 U7975 ( .A1(n6700), .A2(n14124), .ZN(n7658) );
  NAND2_X1 U7976 ( .A1(n11996), .A2(n11849), .ZN(n7626) );
  NOR2_X1 U7977 ( .A1(n11997), .A2(n11848), .ZN(n7628) );
  OR2_X1 U7978 ( .A1(n10562), .A2(n9701), .ZN(n7222) );
  OR2_X1 U7979 ( .A1(n15168), .A2(n11064), .ZN(n7337) );
  INV_X1 U7980 ( .A(n6950), .ZN(n11063) );
  OR2_X1 U7981 ( .A1(n8713), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U7982 ( .A1(n11882), .A2(n11979), .ZN(n8987) );
  NOR2_X1 U7983 ( .A1(n6698), .A2(n11870), .ZN(n7268) );
  INV_X1 U7984 ( .A(n8883), .ZN(n7256) );
  XNOR2_X1 U7985 ( .A(n12811), .B(n12821), .ZN(n12802) );
  OR2_X1 U7986 ( .A1(n13044), .A2(n12781), .ZN(n11961) );
  INV_X1 U7987 ( .A(n7250), .ZN(n7249) );
  OAI21_X1 U7988 ( .B1(n8823), .B2(n6721), .A(n8835), .ZN(n7250) );
  OR2_X1 U7989 ( .A1(n13054), .A2(n12833), .ZN(n11951) );
  OR2_X1 U7990 ( .A1(n13064), .A2(n12832), .ZN(n11945) );
  OR2_X1 U7991 ( .A1(n13080), .A2(n12868), .ZN(n11933) );
  OR2_X1 U7992 ( .A1(n13083), .A2(n12543), .ZN(n11924) );
  AND2_X1 U7993 ( .A1(n7267), .A2(n7265), .ZN(n6934) );
  INV_X1 U7994 ( .A(n8463), .ZN(n7588) );
  INV_X1 U7995 ( .A(n8811), .ZN(n7585) );
  INV_X1 U7996 ( .A(n7575), .ZN(n7574) );
  OAI21_X1 U7997 ( .B1(n8736), .B2(n7576), .A(n8454), .ZN(n7575) );
  INV_X1 U7998 ( .A(n8452), .ZN(n7576) );
  INV_X1 U7999 ( .A(n8433), .ZN(n7590) );
  NAND2_X1 U8000 ( .A1(n9829), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U8001 ( .A1(n9815), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8428) );
  INV_X1 U8002 ( .A(n11521), .ZN(n7432) );
  INV_X1 U8003 ( .A(n7435), .ZN(n7434) );
  CLKBUF_X1 U8004 ( .A(n9593), .Z(n9576) );
  NOR2_X1 U8005 ( .A1(n7504), .A2(n7502), .ZN(n7503) );
  NAND2_X1 U8006 ( .A1(n7504), .A2(n7502), .ZN(n7501) );
  INV_X1 U8007 ( .A(n6681), .ZN(n7383) );
  OR2_X1 U8008 ( .A1(n7329), .A2(n13545), .ZN(n6866) );
  AND2_X1 U8009 ( .A1(n13560), .A2(n13439), .ZN(n7329) );
  INV_X1 U8010 ( .A(n7370), .ZN(n7369) );
  INV_X1 U8011 ( .A(n13453), .ZN(n7051) );
  NAND2_X1 U8012 ( .A1(n7052), .A2(n6757), .ZN(n11546) );
  AOI21_X1 U8013 ( .B1(n10841), .B2(n7304), .A(n6774), .ZN(n7301) );
  NAND2_X1 U8014 ( .A1(n9923), .A2(n13400), .ZN(n11332) );
  AOI21_X1 U8015 ( .B1(n11113), .B2(n7361), .A(n6767), .ZN(n7360) );
  INV_X1 U8016 ( .A(n10804), .ZN(n7361) );
  AND2_X1 U8017 ( .A1(n15056), .A2(n10810), .ZN(n7285) );
  INV_X1 U8018 ( .A(n10813), .ZN(n7289) );
  NOR3_X1 U8019 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .A3(
        P2_IR_REG_18__SCAN_IN), .ZN(n9019) );
  NOR2_X1 U8020 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9012) );
  INV_X1 U8021 ( .A(n12269), .ZN(n7749) );
  AOI21_X1 U8022 ( .B1(n7722), .B2(n7720), .A(n11745), .ZN(n7719) );
  INV_X1 U8023 ( .A(n7722), .ZN(n7721) );
  INV_X1 U8024 ( .A(n11617), .ZN(n7720) );
  NAND2_X1 U8025 ( .A1(n11811), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7927) );
  NOR2_X1 U8026 ( .A1(n8202), .A2(n7713), .ZN(n7712) );
  INV_X1 U8027 ( .A(n8180), .ZN(n7713) );
  NOR2_X1 U8028 ( .A1(n12080), .A2(n7125), .ZN(n7124) );
  NAND2_X1 U8029 ( .A1(n14496), .A2(n14071), .ZN(n12012) );
  NOR2_X1 U8030 ( .A1(n14284), .A2(n14265), .ZN(n14264) );
  NAND3_X1 U8031 ( .A1(n11464), .A2(n14464), .A3(n6692), .ZN(n14284) );
  NOR2_X1 U8032 ( .A1(n7153), .A2(n7148), .ZN(n7146) );
  INV_X1 U8033 ( .A(n7151), .ZN(n7143) );
  AOI21_X1 U8034 ( .B1(n7154), .B2(n7152), .A(n6836), .ZN(n7151) );
  INV_X1 U8035 ( .A(n6830), .ZN(n7152) );
  NOR3_X1 U8036 ( .A1(n7153), .A2(n7148), .A3(n7150), .ZN(n7144) );
  AND3_X1 U8037 ( .A1(n8292), .A2(n7388), .A3(n7387), .ZN(n7386) );
  INV_X1 U8038 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7388) );
  OR2_X1 U8039 ( .A1(n7835), .A2(n7837), .ZN(n7141) );
  INV_X1 U8040 ( .A(n8145), .ZN(n7075) );
  INV_X1 U8041 ( .A(n7647), .ZN(n7646) );
  OAI21_X1 U8042 ( .B1(n7823), .B2(n7648), .A(n7827), .ZN(n7647) );
  NAND2_X1 U8043 ( .A1(n8089), .A2(n7819), .ZN(n7824) );
  INV_X1 U8044 ( .A(n7652), .ZN(n7140) );
  INV_X1 U8045 ( .A(n7137), .ZN(n7136) );
  NAND2_X1 U8046 ( .A1(n7652), .A2(n7139), .ZN(n7138) );
  AOI21_X1 U8047 ( .B1(n7652), .B2(n7654), .A(n7650), .ZN(n7649) );
  INV_X1 U8048 ( .A(n8001), .ZN(n7803) );
  NAND2_X1 U8049 ( .A1(n7808), .A2(SI_10_), .ZN(n7809) );
  NAND2_X1 U8050 ( .A1(n7813), .A2(n7812), .ZN(n8022) );
  XNOR2_X1 U8051 ( .A(n7808), .B(SI_10_), .ZN(n8013) );
  XNOR2_X1 U8052 ( .A(n7804), .B(SI_9_), .ZN(n8001) );
  XNOR2_X1 U8053 ( .A(n7785), .B(SI_3_), .ZN(n7929) );
  OAI21_X1 U8054 ( .B1(n7895), .B2(n7894), .A(n7780), .ZN(n7781) );
  INV_X1 U8055 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n15428) );
  AND2_X1 U8056 ( .A1(n7894), .A2(SI_2_), .ZN(n6868) );
  INV_X1 U8057 ( .A(n7226), .ZN(n7157) );
  OAI21_X1 U8058 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15187), .A(n14515), .ZN(
        n14517) );
  OAI21_X1 U8059 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14521), .A(n14520), .ZN(
        n14571) );
  NAND2_X1 U8060 ( .A1(n15135), .A2(n11582), .ZN(n12494) );
  NOR2_X1 U8061 ( .A1(n12529), .A2(n12937), .ZN(n7528) );
  NAND2_X1 U8062 ( .A1(n7530), .A2(n6816), .ZN(n7529) );
  INV_X1 U8063 ( .A(n6912), .ZN(n7530) );
  NAND2_X1 U8064 ( .A1(n10990), .A2(n6755), .ZN(n11106) );
  INV_X1 U8065 ( .A(n10994), .ZN(n10991) );
  NAND2_X1 U8066 ( .A1(n11587), .A2(n11586), .ZN(n12400) );
  AND2_X1 U8067 ( .A1(n12556), .A2(n7539), .ZN(n7538) );
  OR2_X1 U8068 ( .A1(n12472), .A2(n7540), .ZN(n7539) );
  INV_X1 U8069 ( .A(n12429), .ZN(n7540) );
  NAND2_X1 U8070 ( .A1(n12502), .A2(n12434), .ZN(n12462) );
  NAND2_X1 U8071 ( .A1(n7545), .A2(n11299), .ZN(n11580) );
  INV_X1 U8072 ( .A(n11301), .ZN(n7545) );
  INV_X1 U8073 ( .A(n12821), .ZN(n12605) );
  AND2_X1 U8074 ( .A1(n12453), .A2(n12414), .ZN(n7559) );
  OAI21_X1 U8075 ( .B1(n7580), .B2(n7579), .A(n11967), .ZN(n7578) );
  OR2_X1 U8076 ( .A1(n7580), .A2(n11967), .ZN(n7577) );
  AND3_X1 U8077 ( .A1(n8822), .A2(n8821), .A3(n8820), .ZN(n8824) );
  AND2_X1 U8078 ( .A1(n8810), .A2(n8809), .ZN(n12474) );
  AND4_X1 U8079 ( .A1(n8767), .A2(n8766), .A3(n8765), .A4(n8764), .ZN(n12596)
         );
  AND4_X1 U8080 ( .A1(n8752), .A2(n8751), .A3(n8750), .A4(n8749), .ZN(n12528)
         );
  AND4_X1 U8081 ( .A1(n8556), .A2(n8555), .A3(n8554), .A4(n8553), .ZN(n11303)
         );
  OR2_X1 U8082 ( .A1(n9698), .A2(n9778), .ZN(n9699) );
  OR2_X1 U8083 ( .A1(n9682), .A2(n9778), .ZN(n9683) );
  NAND2_X1 U8084 ( .A1(n9684), .A2(n10570), .ZN(n7312) );
  NOR2_X1 U8085 ( .A1(n10638), .A2(n9705), .ZN(n9707) );
  OR2_X1 U8086 ( .A1(n10626), .A2(n9689), .ZN(n7293) );
  NOR2_X1 U8087 ( .A1(n11075), .A2(n15171), .ZN(n11079) );
  INV_X1 U8088 ( .A(n7218), .ZN(n11074) );
  OR2_X1 U8089 ( .A1(n15217), .A2(n15218), .ZN(n15215) );
  XNOR2_X1 U8090 ( .A(n12631), .B(n15234), .ZN(n15240) );
  INV_X1 U8091 ( .A(n15260), .ZN(n7223) );
  INV_X1 U8092 ( .A(n12523), .ZN(n12781) );
  AND2_X1 U8093 ( .A1(n7259), .A2(n6730), .ZN(n7755) );
  OR2_X1 U8094 ( .A1(n8841), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8852) );
  OR2_X1 U8095 ( .A1(n8852), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8864) );
  INV_X1 U8096 ( .A(n12573), .ZN(n12832) );
  NAND2_X1 U8097 ( .A1(n12881), .A2(n8801), .ZN(n12867) );
  NAND2_X1 U8098 ( .A1(n8385), .A2(n15481), .ZN(n8696) );
  INV_X1 U8099 ( .A(n8669), .ZN(n8385) );
  AND4_X1 U8100 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n12583)
         );
  INV_X1 U8101 ( .A(n11368), .ZN(n7252) );
  NOR2_X1 U8102 ( .A1(n11980), .A2(n6727), .ZN(n7253) );
  NOR2_X1 U8103 ( .A1(n8584), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8604) );
  XNOR2_X1 U8104 ( .A(n12497), .B(n15276), .ZN(n15272) );
  AND4_X1 U8105 ( .A1(n8538), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n11317)
         );
  INV_X1 U8106 ( .A(n11977), .ZN(n8532) );
  AOI21_X1 U8107 ( .B1(n12788), .B2(n8894), .A(n8893), .ZN(n12766) );
  AND2_X1 U8108 ( .A1(n11961), .A2(n11960), .ZN(n12794) );
  NAND2_X1 U8109 ( .A1(n11951), .A2(n11952), .ZN(n12820) );
  NAND2_X1 U8110 ( .A1(n12856), .A2(n8823), .ZN(n12855) );
  INV_X1 U8111 ( .A(n7608), .ZN(n7607) );
  NAND2_X1 U8112 ( .A1(n7273), .A2(n8719), .ZN(n12935) );
  NAND2_X1 U8113 ( .A1(n12945), .A2(n12942), .ZN(n7273) );
  AOI21_X1 U8114 ( .B1(n7610), .B2(n11904), .A(n7609), .ZN(n7608) );
  INV_X1 U8115 ( .A(n11910), .ZN(n7609) );
  AND2_X1 U8116 ( .A1(n11918), .A2(n11912), .ZN(n12934) );
  INV_X1 U8117 ( .A(n15313), .ZN(n12946) );
  INV_X1 U8118 ( .A(n15315), .ZN(n12948) );
  INV_X1 U8119 ( .A(n15311), .ZN(n15322) );
  NAND2_X1 U8120 ( .A1(n8991), .A2(n8990), .ZN(n11598) );
  NAND2_X1 U8121 ( .A1(n11959), .A2(n8929), .ZN(n15315) );
  NAND2_X1 U8122 ( .A1(n8902), .A2(n8901), .ZN(n11832) );
  OR2_X1 U8123 ( .A1(n8899), .A2(n8898), .ZN(n8902) );
  NAND2_X1 U8124 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7602), .ZN(n7600) );
  NOR2_X1 U8125 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7602), .ZN(n7601) );
  AND2_X1 U8126 ( .A1(n7760), .A2(n7267), .ZN(n7266) );
  NAND2_X1 U8127 ( .A1(n8812), .A2(n8811), .ZN(n8814) );
  NAND2_X1 U8128 ( .A1(n8771), .A2(n8457), .ZN(n8783) );
  NAND2_X1 U8129 ( .A1(n8723), .A2(n8450), .ZN(n8737) );
  NAND2_X1 U8130 ( .A1(n8737), .A2(n8736), .ZN(n8739) );
  NAND2_X1 U8131 ( .A1(n8741), .A2(n8740), .ZN(n8743) );
  NAND2_X1 U8132 ( .A1(n8721), .A2(n8720), .ZN(n8723) );
  NAND2_X1 U8133 ( .A1(n7563), .A2(n10016), .ZN(n8446) );
  NAND2_X1 U8134 ( .A1(n8679), .A2(n8445), .ZN(n7563) );
  NAND2_X1 U8135 ( .A1(n8647), .A2(n8441), .ZN(n8663) );
  NAND2_X1 U8136 ( .A1(n8663), .A2(n8662), .ZN(n8665) );
  NAND2_X1 U8137 ( .A1(n8645), .A2(n8644), .ZN(n8647) );
  NOR2_X1 U8138 ( .A1(n8593), .A2(n7594), .ZN(n7593) );
  INV_X1 U8139 ( .A(n8431), .ZN(n7594) );
  NAND2_X1 U8140 ( .A1(n8580), .A2(n8430), .ZN(n7595) );
  NAND2_X1 U8141 ( .A1(n8423), .A2(n8422), .ZN(n8540) );
  AND2_X1 U8142 ( .A1(n8545), .A2(n8544), .ZN(n9728) );
  NAND2_X1 U8143 ( .A1(n8681), .A2(n8402), .ZN(n7309) );
  XNOR2_X1 U8144 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8491) );
  NAND2_X1 U8145 ( .A1(n7158), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U8146 ( .A1(n11529), .A2(n11526), .ZN(n7435) );
  INV_X1 U8147 ( .A(n13216), .ZN(n13154) );
  NAND2_X1 U8148 ( .A1(n13229), .A2(n13224), .ZN(n7428) );
  NAND2_X1 U8149 ( .A1(n13327), .A2(n13195), .ZN(n13198) );
  NOR2_X1 U8150 ( .A1(n10488), .A2(n10326), .ZN(n7456) );
  INV_X1 U8151 ( .A(n7457), .ZN(n7454) );
  OAI21_X1 U8152 ( .B1(n13154), .B2(n7437), .A(n7436), .ZN(n13236) );
  NAND2_X1 U8153 ( .A1(n13170), .A2(n13300), .ZN(n7437) );
  OR2_X1 U8154 ( .A1(n7438), .A2(n13162), .ZN(n7436) );
  OR2_X1 U8155 ( .A1(n13138), .A2(n13139), .ZN(n13140) );
  CLKBUF_X1 U8156 ( .A(n10939), .Z(n6898) );
  NAND2_X1 U8157 ( .A1(n7462), .A2(n7466), .ZN(n7460) );
  AND2_X1 U8158 ( .A1(n7464), .A2(n6723), .ZN(n7462) );
  NAND2_X1 U8159 ( .A1(n13216), .A2(n13300), .ZN(n6929) );
  NAND2_X1 U8160 ( .A1(n6898), .A2(n7468), .ZN(n7467) );
  INV_X1 U8161 ( .A(n13374), .ZN(n10196) );
  OAI21_X1 U8162 ( .B1(n7447), .B2(n7445), .A(n7444), .ZN(n13319) );
  AOI21_X1 U8163 ( .B1(n13272), .B2(n13271), .A(n6705), .ZN(n7444) );
  INV_X1 U8164 ( .A(n13271), .ZN(n7445) );
  NAND2_X1 U8165 ( .A1(n7069), .A2(n6747), .ZN(n6961) );
  AND2_X1 U8166 ( .A1(n9433), .A2(n9432), .ZN(n13465) );
  AND2_X1 U8167 ( .A1(n9392), .A2(n9391), .ZN(n13457) );
  AND2_X1 U8168 ( .A1(n9373), .A2(n9372), .ZN(n13455) );
  AND3_X1 U8169 ( .A1(n9332), .A2(n9331), .A3(n9330), .ZN(n11560) );
  AND4_X1 U8170 ( .A1(n9228), .A2(n9227), .A3(n9226), .A4(n9225), .ZN(n10823)
         );
  NAND2_X1 U8171 ( .A1(n9587), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9126) );
  NOR2_X1 U8172 ( .A1(n9111), .A2(n13376), .ZN(n7414) );
  INV_X1 U8173 ( .A(n13540), .ZN(n7330) );
  AND2_X1 U8174 ( .A1(n13545), .A2(n13474), .ZN(n7385) );
  NAND2_X1 U8175 ( .A1(n13555), .A2(n13439), .ZN(n7326) );
  AOI21_X1 U8176 ( .B1(n7374), .B2(n6691), .A(n6710), .ZN(n7373) );
  NAND2_X1 U8177 ( .A1(n6696), .A2(n6681), .ZN(n13559) );
  NAND2_X1 U8178 ( .A1(n7057), .A2(n7376), .ZN(n13587) );
  NAND2_X1 U8179 ( .A1(n7297), .A2(n7295), .ZN(n13599) );
  AOI21_X1 U8180 ( .B1(n6704), .B2(n7300), .A(n7296), .ZN(n7295) );
  INV_X1 U8181 ( .A(n13430), .ZN(n7296) );
  NAND2_X1 U8182 ( .A1(n13430), .A2(n13429), .ZN(n13620) );
  NAND2_X1 U8183 ( .A1(n13460), .A2(n13459), .ZN(n13612) );
  NAND2_X1 U8184 ( .A1(n13629), .A2(n13427), .ZN(n13631) );
  AND2_X1 U8185 ( .A1(n13646), .A2(n13456), .ZN(n7370) );
  NAND2_X1 U8186 ( .A1(n13663), .A2(n13665), .ZN(n7371) );
  NAND2_X1 U8187 ( .A1(n13454), .A2(n13453), .ZN(n13663) );
  NAND2_X1 U8188 ( .A1(n11540), .A2(n11539), .ZN(n11563) );
  NAND2_X1 U8189 ( .A1(n11285), .A2(n11284), .ZN(n11325) );
  NAND2_X1 U8190 ( .A1(n11277), .A2(n11276), .ZN(n11328) );
  XNOR2_X1 U8191 ( .A(n15054), .B(n7290), .ZN(n15056) );
  NAND2_X1 U8192 ( .A1(n10654), .A2(n10653), .ZN(n10799) );
  NAND2_X1 U8193 ( .A1(n9547), .A2(n9546), .ZN(n13406) );
  NAND2_X1 U8194 ( .A1(n9445), .A2(n9444), .ZN(n13730) );
  AND2_X1 U8195 ( .A1(n9180), .A2(n9179), .ZN(n15089) );
  INV_X1 U8196 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9016) );
  INV_X1 U8197 ( .A(n9286), .ZN(n7480) );
  INV_X1 U8198 ( .A(n9026), .ZN(n7417) );
  NAND2_X1 U8199 ( .A1(n9056), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U8200 ( .A1(n9663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9650) );
  OR2_X1 U8201 ( .A1(n9651), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9656) );
  NAND2_X1 U8202 ( .A1(n9040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9041) );
  INV_X1 U8203 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7158) );
  INV_X1 U8204 ( .A(n7863), .ZN(n7790) );
  NAND2_X1 U8205 ( .A1(n12262), .A2(n6845), .ZN(n13850) );
  NOR2_X1 U8206 ( .A1(n13853), .A2(n6846), .ZN(n6845) );
  INV_X1 U8207 ( .A(n12261), .ZN(n6846) );
  NAND2_X1 U8208 ( .A1(n7742), .A2(n7741), .ZN(n7740) );
  INV_X1 U8209 ( .A(n11239), .ZN(n6847) );
  INV_X1 U8210 ( .A(n12322), .ZN(n12375) );
  AND2_X1 U8211 ( .A1(n11626), .A2(n6729), .ZN(n7722) );
  AND2_X1 U8212 ( .A1(n13940), .A2(n7725), .ZN(n7724) );
  NAND2_X1 U8213 ( .A1(n7728), .A2(n7731), .ZN(n7725) );
  INV_X1 U8214 ( .A(n6939), .ZN(n6938) );
  OAI21_X1 U8215 ( .B1(n10381), .B2(n12017), .A(n10262), .ZN(n6939) );
  AOI21_X1 U8216 ( .B1(n12358), .B2(n10446), .A(n6783), .ZN(n10260) );
  NAND2_X1 U8217 ( .A1(n11790), .A2(n11789), .ZN(n7744) );
  INV_X1 U8218 ( .A(n11398), .ZN(n6870) );
  AND4_X1 U8219 ( .A1(n8083), .A2(n8082), .A3(n8081), .A4(n8080), .ZN(n13959)
         );
  OAI21_X1 U8220 ( .B1(n10095), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6975), .ZN(
        n10072) );
  MUX2_X1 U8221 ( .A(n10088), .B(P1_REG2_REG_2__SCAN_IN), .S(n10097), .Z(
        n10089) );
  MUX2_X1 U8222 ( .A(n10096), .B(P1_REG1_REG_2__SCAN_IN), .S(n10097), .Z(
        n10253) );
  OR2_X1 U8223 ( .A1(n10306), .A2(n10305), .ZN(n7347) );
  NOR2_X1 U8224 ( .A1(n10138), .A2(n7350), .ZN(n10121) );
  AND2_X1 U8225 ( .A1(n10144), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7350) );
  NAND2_X1 U8226 ( .A1(n8281), .A2(n8280), .ZN(n12178) );
  AOI21_X1 U8227 ( .B1(n6720), .B2(n7393), .A(n7391), .ZN(n7390) );
  INV_X1 U8228 ( .A(n8333), .ZN(n7391) );
  NAND2_X1 U8229 ( .A1(n7714), .A2(n6756), .ZN(n14122) );
  NOR2_X1 U8230 ( .A1(n14177), .A2(n7718), .ZN(n7717) );
  INV_X1 U8231 ( .A(n8225), .ZN(n7718) );
  AOI21_X1 U8232 ( .B1(n7113), .B2(n7114), .A(n14192), .ZN(n7112) );
  OR2_X1 U8233 ( .A1(n14246), .A2(n14247), .ZN(n14244) );
  AOI21_X1 U8234 ( .B1(n7108), .B2(n7106), .A(n6759), .ZN(n7105) );
  INV_X1 U8235 ( .A(n7108), .ZN(n7107) );
  INV_X1 U8236 ( .A(n8323), .ZN(n7106) );
  NAND2_X1 U8237 ( .A1(n8325), .A2(n8324), .ZN(n14259) );
  INV_X1 U8238 ( .A(n14025), .ZN(n14304) );
  NAND2_X1 U8239 ( .A1(n8116), .A2(n8115), .ZN(n14328) );
  INV_X1 U8240 ( .A(n8084), .ZN(n12094) );
  NAND2_X1 U8241 ( .A1(n12100), .A2(n12101), .ZN(n12218) );
  NAND2_X1 U8242 ( .A1(n12096), .A2(n12095), .ZN(n8084) );
  AOI21_X1 U8243 ( .B1(n7102), .B2(n7104), .A(n6766), .ZN(n7100) );
  NAND2_X1 U8244 ( .A1(n12215), .A2(n11185), .ZN(n7101) );
  OR2_X1 U8245 ( .A1(n12080), .A2(n12073), .ZN(n7123) );
  NOR2_X1 U8246 ( .A1(n12213), .A2(n7401), .ZN(n7400) );
  INV_X1 U8247 ( .A(n8315), .ZN(n7401) );
  NAND2_X1 U8248 ( .A1(n7402), .A2(n7698), .ZN(n11026) );
  INV_X1 U8249 ( .A(n8012), .ZN(n7699) );
  NAND2_X1 U8250 ( .A1(n11025), .A2(n7398), .ZN(n11024) );
  INV_X1 U8251 ( .A(n7698), .ZN(n7398) );
  AND4_X1 U8252 ( .A1(n8011), .A2(n8010), .A3(n8009), .A4(n8008), .ZN(n12069)
         );
  AOI21_X1 U8253 ( .B1(n10681), .B2(n7692), .A(n6763), .ZN(n7691) );
  INV_X1 U8254 ( .A(n10681), .ZN(n7693) );
  NAND2_X1 U8255 ( .A1(n7951), .A2(n7950), .ZN(n12047) );
  INV_X1 U8256 ( .A(n14038), .ZN(n12039) );
  NAND2_X1 U8257 ( .A1(n12201), .A2(n7920), .ZN(n7700) );
  NAND2_X1 U8258 ( .A1(n10614), .A2(n10615), .ZN(n10613) );
  CLKBUF_X1 U8259 ( .A(n8363), .Z(n14248) );
  AND2_X2 U8260 ( .A1(n14495), .A2(n8204), .ZN(n14211) );
  OAI21_X1 U8261 ( .B1(n8263), .B2(n7667), .A(n7665), .ZN(n9540) );
  NAND2_X1 U8262 ( .A1(n7164), .A2(n7975), .ZN(n8133) );
  NAND2_X1 U8263 ( .A1(n7841), .A2(SI_22_), .ZN(n7842) );
  XNOR2_X1 U8264 ( .A(n8296), .B(P1_IR_REG_21__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U8265 ( .A1(n6944), .A2(n7752), .ZN(n8295) );
  NAND2_X1 U8266 ( .A1(n14509), .A2(n14508), .ZN(n14551) );
  NAND2_X1 U8267 ( .A1(n14543), .A2(n14544), .ZN(n14508) );
  NAND2_X1 U8268 ( .A1(n6919), .A2(n6918), .ZN(n14592) );
  NAND2_X1 U8269 ( .A1(n14585), .A2(n15045), .ZN(n6918) );
  AND4_X1 U8270 ( .A1(n8701), .A2(n8700), .A3(n8699), .A4(n8698), .ZN(n12562)
         );
  NAND2_X1 U8271 ( .A1(n8840), .A2(n8839), .ZN(n12987) );
  NAND2_X1 U8272 ( .A1(n12592), .A2(n12427), .ZN(n12473) );
  NAND2_X1 U8273 ( .A1(n12504), .A2(n12503), .ZN(n12502) );
  NOR2_X1 U8274 ( .A1(n6706), .A2(n15146), .ZN(n7547) );
  NAND2_X1 U8275 ( .A1(n7550), .A2(n7553), .ZN(n7549) );
  NAND2_X1 U8276 ( .A1(n6695), .A2(n7554), .ZN(n7553) );
  XNOR2_X1 U8277 ( .A(n12462), .B(n12460), .ZN(n12574) );
  AND4_X2 U8278 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(n15312)
         );
  OAI21_X2 U8279 ( .B1(n12531), .B2(n7522), .A(n7520), .ZN(n12592) );
  INV_X1 U8280 ( .A(n7523), .ZN(n7522) );
  AOI21_X1 U8281 ( .B1(n7523), .B2(n7525), .A(n7521), .ZN(n7520) );
  INV_X1 U8282 ( .A(n12593), .ZN(n7521) );
  INV_X1 U8283 ( .A(n15159), .ZN(n12619) );
  INV_X1 U8284 ( .A(n10772), .ZN(n12004) );
  INV_X1 U8285 ( .A(n8824), .ZN(n12869) );
  INV_X1 U8286 ( .A(n12543), .ZN(n12912) );
  INV_X1 U8287 ( .A(n12528), .ZN(n12937) );
  NAND4_X1 U8288 ( .A1(n8641), .A2(n8640), .A3(n8639), .A4(n8638), .ZN(n12401)
         );
  OR2_X1 U8289 ( .A1(n8795), .A2(n11076), .ZN(n8638) );
  OR2_X1 U8290 ( .A1(n8494), .A2(n8509), .ZN(n8510) );
  NAND2_X1 U8291 ( .A1(n15162), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15161) );
  INV_X1 U8292 ( .A(n9774), .ZN(n10570) );
  OR2_X1 U8293 ( .A1(n12636), .A2(n12637), .ZN(n12683) );
  NOR2_X1 U8294 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  NAND2_X1 U8295 ( .A1(n7621), .A2(n11990), .ZN(n13000) );
  INV_X1 U8296 ( .A(n12878), .ZN(n7621) );
  OR2_X1 U8297 ( .A1(n10453), .A2(n8815), .ZN(n8806) );
  NAND2_X1 U8298 ( .A1(n8762), .A2(n8761), .ZN(n13089) );
  NAND2_X1 U8299 ( .A1(n7636), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8480) );
  NAND2_X1 U8300 ( .A1(n7459), .A2(n10486), .ZN(n7458) );
  INV_X1 U8301 ( .A(n10487), .ZN(n7459) );
  INV_X1 U8302 ( .A(n13804), .ZN(n13637) );
  NOR2_X1 U8303 ( .A1(n6709), .A2(n13339), .ZN(n7421) );
  NAND2_X1 U8304 ( .A1(n7424), .A2(n7428), .ZN(n7423) );
  INV_X1 U8305 ( .A(n13198), .ZN(n13201) );
  AND2_X1 U8306 ( .A1(n9219), .A2(n9218), .ZN(n15103) );
  NAND2_X1 U8307 ( .A1(n13281), .A2(n13185), .ZN(n13244) );
  NAND2_X1 U8308 ( .A1(n9070), .A2(n9069), .ZN(n15078) );
  INV_X1 U8309 ( .A(n13230), .ZN(n13357) );
  NAND2_X1 U8310 ( .A1(n9506), .A2(n9505), .ZN(n13522) );
  NAND2_X1 U8311 ( .A1(n13828), .A2(n9579), .ZN(n9506) );
  NAND2_X1 U8312 ( .A1(n15127), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7322) );
  NAND2_X1 U8313 ( .A1(n13694), .A2(n7317), .ZN(n7316) );
  NOR2_X1 U8314 ( .A1(n7320), .A2(n7318), .ZN(n7317) );
  INV_X1 U8315 ( .A(n7322), .ZN(n7318) );
  AND2_X1 U8316 ( .A1(n9557), .A2(n9556), .ZN(n13775) );
  OR2_X1 U8317 ( .A1(n14479), .A2(n9555), .ZN(n9557) );
  NAND2_X1 U8318 ( .A1(n9581), .A2(n9580), .ZN(n13503) );
  CLKBUF_X1 U8319 ( .A(n11618), .Z(n11444) );
  OAI21_X1 U8320 ( .B1(n13989), .B2(n12366), .A(n7734), .ZN(n13842) );
  INV_X1 U8321 ( .A(n14014), .ZN(n13991) );
  AND2_X1 U8322 ( .A1(n9987), .A2(n10268), .ZN(n14238) );
  NOR2_X1 U8323 ( .A1(n10141), .A2(n6913), .ZN(n10110) );
  AND2_X1 U8324 ( .A1(n10144), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6913) );
  OR2_X1 U8325 ( .A1(n14731), .A2(n10077), .ZN(n14789) );
  NAND2_X1 U8326 ( .A1(n8216), .A2(n8215), .ZN(n14202) );
  AND2_X1 U8327 ( .A1(n10888), .A2(n14071), .ZN(n14333) );
  INV_X1 U8328 ( .A(n14309), .ZN(n14319) );
  OR2_X1 U8329 ( .A1(n9796), .A2(n11805), .ZN(n7918) );
  AND2_X1 U8330 ( .A1(n14343), .A2(n14342), .ZN(n6976) );
  NAND2_X1 U8331 ( .A1(n11807), .A2(n11806), .ZN(n14431) );
  OR2_X1 U8332 ( .A1(n14479), .A2(n11805), .ZN(n11807) );
  NAND2_X1 U8333 ( .A1(n6862), .A2(n6754), .ZN(n9672) );
  NAND2_X1 U8334 ( .A1(n7865), .A2(n7864), .ZN(n14435) );
  NAND2_X1 U8335 ( .A1(n13825), .A2(n11804), .ZN(n7865) );
  NAND2_X1 U8336 ( .A1(n14348), .A2(n14842), .ZN(n6858) );
  OAI21_X1 U8337 ( .B1(n6926), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n6925), .ZN(
        n6924) );
  AND2_X1 U8338 ( .A1(n14596), .A2(n14595), .ZN(n6926) );
  INV_X1 U8339 ( .A(n14560), .ZN(n7241) );
  NOR2_X1 U8340 ( .A1(n14715), .A2(n14716), .ZN(n14714) );
  NOR2_X1 U8341 ( .A1(n14720), .A2(n14719), .ZN(n14718) );
  NAND2_X1 U8342 ( .A1(n14592), .A2(n14591), .ZN(n7245) );
  OR2_X1 U8343 ( .A1(n14043), .A2(n12016), .ZN(n12018) );
  NOR2_X1 U8344 ( .A1(n12032), .A2(n7182), .ZN(n7181) );
  NAND2_X1 U8345 ( .A1(n7172), .A2(n7174), .ZN(n12055) );
  NAND2_X1 U8346 ( .A1(n12049), .A2(n7174), .ZN(n7170) );
  NAND2_X1 U8347 ( .A1(n7171), .A2(n7174), .ZN(n6949) );
  NOR2_X1 U8348 ( .A1(n12071), .A2(n12072), .ZN(n7191) );
  AND2_X1 U8349 ( .A1(n7193), .A2(n12066), .ZN(n7192) );
  NAND2_X1 U8350 ( .A1(n6921), .A2(n6920), .ZN(n12086) );
  NAND2_X1 U8351 ( .A1(n12081), .A2(n12083), .ZN(n6920) );
  INV_X1 U8352 ( .A(n12093), .ZN(n7676) );
  NAND2_X1 U8353 ( .A1(n7491), .A2(n9175), .ZN(n9177) );
  NAND2_X1 U8354 ( .A1(n7490), .A2(n7488), .ZN(n6942) );
  NAND2_X1 U8355 ( .A1(n7000), .A2(n15308), .ZN(n6998) );
  NAND2_X1 U8356 ( .A1(n11859), .A2(n11860), .ZN(n7000) );
  AOI21_X1 U8357 ( .B1(n7197), .B2(n6697), .A(n6786), .ZN(n7195) );
  INV_X1 U8358 ( .A(n12102), .ZN(n7197) );
  NAND2_X1 U8359 ( .A1(n6994), .A2(n6993), .ZN(n11871) );
  AND2_X1 U8360 ( .A1(n11976), .A2(n6828), .ZN(n6993) );
  NAND2_X1 U8361 ( .A1(n6996), .A2(n6995), .ZN(n6994) );
  INV_X1 U8362 ( .A(n9231), .ZN(n7493) );
  NAND2_X1 U8363 ( .A1(n15268), .A2(n7007), .ZN(n7006) );
  NAND2_X1 U8364 ( .A1(n11967), .A2(n7008), .ZN(n7007) );
  INV_X1 U8365 ( .A(n11877), .ZN(n7008) );
  INV_X1 U8366 ( .A(n7511), .ZN(n7510) );
  NAND2_X1 U8367 ( .A1(n12145), .A2(n12147), .ZN(n6907) );
  NAND2_X1 U8368 ( .A1(n7003), .A2(n7001), .ZN(n11889) );
  NOR2_X1 U8369 ( .A1(n7002), .A2(n8635), .ZN(n7001) );
  INV_X1 U8370 ( .A(n11884), .ZN(n7002) );
  NAND2_X1 U8371 ( .A1(n7202), .A2(n12154), .ZN(n7201) );
  INV_X1 U8372 ( .A(n12155), .ZN(n7202) );
  INV_X1 U8373 ( .A(n11922), .ZN(n7020) );
  NAND2_X1 U8374 ( .A1(n11928), .A2(n11926), .ZN(n7019) );
  NAND2_X1 U8375 ( .A1(n12164), .A2(n7683), .ZN(n7682) );
  OR2_X1 U8376 ( .A1(n12164), .A2(n7683), .ZN(n6806) );
  NAND2_X1 U8377 ( .A1(n7012), .A2(n7009), .ZN(n11936) );
  AND2_X1 U8378 ( .A1(n7011), .A2(n7010), .ZN(n7009) );
  INV_X1 U8379 ( .A(n7028), .ZN(n7025) );
  INV_X1 U8380 ( .A(n12820), .ZN(n7033) );
  NAND2_X1 U8381 ( .A1(n7028), .A2(n7030), .ZN(n7027) );
  INV_X1 U8382 ( .A(n7031), .ZN(n7030) );
  NAND2_X1 U8383 ( .A1(n12175), .A2(n7673), .ZN(n7163) );
  INV_X1 U8384 ( .A(n12174), .ZN(n7673) );
  INV_X1 U8385 ( .A(n6734), .ZN(n7026) );
  INV_X1 U8386 ( .A(n12096), .ZN(n7098) );
  NAND2_X1 U8387 ( .A1(n7345), .A2(n7079), .ZN(n7078) );
  NOR2_X1 U8388 ( .A1(n13602), .A2(n7080), .ZN(n7079) );
  NAND2_X1 U8389 ( .A1(n7085), .A2(n7081), .ZN(n7080) );
  NOR2_X1 U8390 ( .A1(n11118), .A2(n7305), .ZN(n7304) );
  INV_X1 U8391 ( .A(n10820), .ZN(n7305) );
  OR2_X1 U8392 ( .A1(n12094), .A2(n7098), .ZN(n7097) );
  AND2_X1 U8393 ( .A1(n8319), .A2(n7098), .ZN(n7093) );
  NOR2_X1 U8394 ( .A1(n7853), .A2(n6719), .ZN(n7154) );
  INV_X1 U8395 ( .A(n7154), .ZN(n7153) );
  NAND2_X1 U8396 ( .A1(n7639), .A2(n7637), .ZN(n7846) );
  INV_X1 U8397 ( .A(n7638), .ZN(n7637) );
  OAI21_X1 U8398 ( .B1(n7842), .B2(n6716), .A(n7844), .ZN(n7638) );
  NAND2_X1 U8399 ( .A1(n7643), .A2(n7644), .ZN(n7829) );
  AOI21_X1 U8400 ( .B1(n7646), .B2(n6707), .A(n6825), .ZN(n7644) );
  NAND2_X1 U8401 ( .A1(n7824), .A2(n7645), .ZN(n7643) );
  NOR2_X1 U8402 ( .A1(n7136), .A2(n15723), .ZN(n7068) );
  NOR2_X1 U8403 ( .A1(n7068), .A2(n8055), .ZN(n7065) );
  NOR2_X1 U8404 ( .A1(n7137), .A2(SI_13_), .ZN(n7066) );
  INV_X1 U8405 ( .A(n8038), .ZN(n7650) );
  INV_X1 U8406 ( .A(n7805), .ZN(n7139) );
  OAI21_X1 U8407 ( .B1(n7845), .B2(P2_DATAO_REG_11__SCAN_IN), .A(n6906), .ZN(
        n7810) );
  NAND2_X1 U8408 ( .A1(n7845), .A2(n9850), .ZN(n6906) );
  INV_X1 U8409 ( .A(n6679), .ZN(n9002) );
  NAND2_X1 U8410 ( .A1(n6990), .A2(n12776), .ZN(n6989) );
  NOR2_X1 U8411 ( .A1(n12762), .A2(n11966), .ZN(n7579) );
  NAND2_X1 U8412 ( .A1(n6784), .A2(n8490), .ZN(n7216) );
  INV_X1 U8413 ( .A(n10582), .ZN(n7221) );
  NAND2_X1 U8414 ( .A1(n7337), .A2(n7336), .ZN(n12659) );
  INV_X1 U8415 ( .A(n11067), .ZN(n7336) );
  OR2_X1 U8416 ( .A1(n12787), .A2(n12766), .ZN(n11966) );
  NAND2_X1 U8417 ( .A1(n8391), .A2(n8390), .ZN(n8793) );
  INV_X1 U8418 ( .A(n8775), .ZN(n8391) );
  NAND2_X1 U8419 ( .A1(n8568), .A2(n8567), .ZN(n11315) );
  INV_X1 U8420 ( .A(n10677), .ZN(n11855) );
  NAND2_X1 U8421 ( .A1(n12877), .A2(n11937), .ZN(n7620) );
  NAND2_X1 U8422 ( .A1(n7608), .A2(n7611), .ZN(n7606) );
  NOR2_X1 U8423 ( .A1(n11984), .A2(n7634), .ZN(n7633) );
  INV_X1 U8424 ( .A(n8988), .ZN(n8985) );
  INV_X1 U8425 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7265) );
  INV_X1 U8426 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8404) );
  AND2_X1 U8427 ( .A1(n7631), .A2(n8403), .ZN(n7267) );
  INV_X1 U8428 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8403) );
  NAND4_X1 U8429 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(n7262)
         );
  AND2_X1 U8430 ( .A1(n8417), .A2(n8420), .ZN(n7568) );
  NAND2_X1 U8431 ( .A1(n9795), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8425) );
  AND2_X1 U8432 ( .A1(n13301), .A2(n7439), .ZN(n7438) );
  NAND2_X1 U8433 ( .A1(n13217), .A2(n13300), .ZN(n7439) );
  NOR2_X1 U8434 ( .A1(n9367), .A2(n13277), .ZN(n9366) );
  AND2_X1 U8435 ( .A1(n9366), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9383) );
  AOI21_X1 U8436 ( .B1(n13406), .B2(n13410), .A(n9614), .ZN(n9641) );
  NAND2_X1 U8437 ( .A1(n7086), .A2(n7076), .ZN(n9638) );
  NOR2_X1 U8438 ( .A1(n7330), .A2(n7077), .ZN(n7076) );
  INV_X1 U8439 ( .A(n13535), .ZN(n7086) );
  OR2_X1 U8440 ( .A1(n6681), .A2(n7078), .ZN(n7077) );
  AND2_X1 U8441 ( .A1(n9640), .A2(n7073), .ZN(n7072) );
  AND2_X1 U8442 ( .A1(n13485), .A2(n13514), .ZN(n7073) );
  NOR2_X1 U8443 ( .A1(n13590), .A2(n13471), .ZN(n7236) );
  NOR2_X1 U8444 ( .A1(n13561), .A2(n13788), .ZN(n7234) );
  INV_X1 U8445 ( .A(n7376), .ZN(n7374) );
  INV_X1 U8446 ( .A(n13468), .ZN(n7375) );
  NOR2_X1 U8447 ( .A1(n9446), .A2(n13313), .ZN(n9462) );
  NAND2_X1 U8448 ( .A1(n7299), .A2(n13627), .ZN(n7298) );
  INV_X1 U8449 ( .A(n13427), .ZN(n7299) );
  OR2_X1 U8450 ( .A1(n13637), .A2(n13428), .ZN(n13459) );
  AND2_X1 U8451 ( .A1(n9235), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9258) );
  NOR2_X1 U8452 ( .A1(n11489), .A2(n11283), .ZN(n7229) );
  NOR2_X1 U8453 ( .A1(n9237), .A2(n9236), .ZN(n9235) );
  INV_X1 U8454 ( .A(n10802), .ZN(n7039) );
  NAND2_X1 U8455 ( .A1(n10801), .A2(n7366), .ZN(n7365) );
  NAND2_X1 U8456 ( .A1(n10798), .A2(n10812), .ZN(n7366) );
  NOR2_X1 U8457 ( .A1(n9183), .A2(n9182), .ZN(n9181) );
  AND2_X1 U8458 ( .A1(n10223), .A2(n10661), .ZN(n10655) );
  INV_X1 U8459 ( .A(n7236), .ZN(n13574) );
  OR2_X1 U8460 ( .A1(n13604), .A2(n13730), .ZN(n13590) );
  NAND2_X1 U8461 ( .A1(n15061), .A2(n15089), .ZN(n15060) );
  INV_X1 U8462 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9017) );
  AND2_X1 U8463 ( .A1(n12333), .A2(n12332), .ZN(n12335) );
  OR2_X1 U8464 ( .A1(n14372), .A2(n6683), .ZN(n12333) );
  AND2_X1 U8465 ( .A1(n12285), .A2(n12284), .ZN(n12287) );
  INV_X1 U8466 ( .A(n6683), .ZN(n12358) );
  NAND2_X1 U8467 ( .A1(n7162), .A2(n7161), .ZN(n7160) );
  INV_X1 U8468 ( .A(n12179), .ZN(n7161) );
  XNOR2_X1 U8469 ( .A(n7656), .B(n14071), .ZN(n12226) );
  XNOR2_X1 U8470 ( .A(n14431), .B(n14017), .ZN(n7659) );
  OR2_X1 U8471 ( .A1(n14762), .A2(n7351), .ZN(n14049) );
  AND2_X1 U8472 ( .A1(n14060), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7351) );
  AOI21_X1 U8473 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14063), .A(n14804), .ZN(
        n14053) );
  OR2_X1 U8474 ( .A1(n14144), .A2(n7393), .ZN(n7392) );
  INV_X1 U8475 ( .A(n14126), .ZN(n7393) );
  OR2_X1 U8476 ( .A1(n14133), .A2(n8272), .ZN(n8273) );
  AND2_X1 U8477 ( .A1(n7109), .A2(n14278), .ZN(n7108) );
  NAND2_X1 U8478 ( .A1(n14302), .A2(n8323), .ZN(n7109) );
  INV_X1 U8479 ( .A(n7103), .ZN(n7102) );
  OAI21_X1 U8480 ( .B1(n12215), .B2(n7104), .A(n11420), .ZN(n7103) );
  INV_X1 U8481 ( .A(n8316), .ZN(n7104) );
  NOR2_X1 U8482 ( .A1(n7993), .A2(n7873), .ZN(n8006) );
  INV_X1 U8483 ( .A(n8310), .ZN(n7404) );
  NAND2_X1 U8484 ( .A1(n10679), .A2(n7693), .ZN(n7405) );
  NAND2_X1 U8485 ( .A1(n10519), .A2(n7905), .ZN(n10614) );
  NAND2_X1 U8486 ( .A1(n7898), .A2(n11001), .ZN(n12023) );
  NAND2_X1 U8487 ( .A1(n12189), .A2(n12013), .ZN(n8340) );
  AOI21_X1 U8488 ( .B1(n7668), .B2(n7670), .A(n7666), .ZN(n7665) );
  INV_X1 U8489 ( .A(n9535), .ZN(n7666) );
  INV_X1 U8490 ( .A(n7668), .ZN(n7667) );
  NOR2_X1 U8491 ( .A1(n7751), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n7750) );
  INV_X2 U8492 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n15539) );
  AOI21_X1 U8493 ( .B1(n7136), .B2(n7140), .A(n7135), .ZN(n7134) );
  INV_X1 U8494 ( .A(n7817), .ZN(n7135) );
  OR2_X1 U8495 ( .A1(n8024), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8025) );
  CLKBUF_X1 U8496 ( .A(n7975), .Z(n7976) );
  XNOR2_X1 U8497 ( .A(n7801), .B(SI_8_), .ZN(n7988) );
  NAND2_X1 U8498 ( .A1(n7060), .A2(n7799), .ZN(n7989) );
  INV_X1 U8499 ( .A(n7971), .ZN(n7797) );
  XNOR2_X1 U8500 ( .A(n7798), .B(SI_7_), .ZN(n7971) );
  XNOR2_X1 U8501 ( .A(n7795), .B(SI_6_), .ZN(n7958) );
  NAND2_X1 U8502 ( .A1(n7061), .A2(n7793), .ZN(n7959) );
  INV_X1 U8503 ( .A(n7946), .ZN(n7791) );
  OR2_X1 U8504 ( .A1(n7948), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7960) );
  INV_X1 U8505 ( .A(n7929), .ZN(n7784) );
  OAI21_X1 U8506 ( .B1(n7863), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7660), .ZN(
        n7772) );
  NAND2_X1 U8507 ( .A1(n7863), .A2(n7662), .ZN(n7660) );
  NAND2_X1 U8508 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6978), .ZN(n6977) );
  INV_X1 U8509 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6978) );
  NAND2_X1 U8510 ( .A1(n14505), .A2(n14506), .ZN(n14507) );
  XNOR2_X1 U8511 ( .A(n14507), .B(n6979), .ZN(n14543) );
  OAI21_X1 U8512 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n15500), .A(n14510), .ZN(
        n14511) );
  NAND2_X1 U8513 ( .A1(n8389), .A2(n8388), .ZN(n8747) );
  INV_X1 U8514 ( .A(n8728), .ZN(n8389) );
  INV_X1 U8515 ( .A(n6817), .ZN(n7554) );
  OR2_X1 U8516 ( .A1(n8793), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8807) );
  AOI21_X1 U8517 ( .B1(n7527), .B2(n7524), .A(n6824), .ZN(n7523) );
  INV_X1 U8518 ( .A(n6816), .ZN(n7524) );
  AND2_X1 U8519 ( .A1(n10957), .A2(n10956), .ZN(n11844) );
  NOR2_X1 U8520 ( .A1(n9716), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9679) );
  INV_X1 U8521 ( .A(n7337), .ZN(n11068) );
  NAND2_X1 U8522 ( .A1(n7339), .A2(n7338), .ZN(n15203) );
  INV_X1 U8523 ( .A(n15205), .ZN(n7338) );
  NAND2_X1 U8524 ( .A1(n15246), .A2(n12650), .ZN(n7307) );
  OR2_X1 U8525 ( .A1(n12669), .A2(n12670), .ZN(n7308) );
  AND2_X1 U8526 ( .A1(n15262), .A2(n7209), .ZN(n6980) );
  NOR2_X1 U8527 ( .A1(n12746), .A2(n12744), .ZN(n7209) );
  INV_X1 U8528 ( .A(n12720), .ZN(n7215) );
  NOR2_X1 U8529 ( .A1(n8786), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8912) );
  OR2_X1 U8530 ( .A1(n8888), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U8531 ( .A1(n8397), .A2(n15555), .ZN(n8888) );
  INV_X1 U8532 ( .A(n8876), .ZN(n8397) );
  OAI21_X1 U8533 ( .B1(n12856), .B2(n6721), .A(n7249), .ZN(n12831) );
  NAND2_X1 U8534 ( .A1(n8394), .A2(n8393), .ZN(n8841) );
  NAND2_X1 U8535 ( .A1(n8392), .A2(n15658), .ZN(n8818) );
  INV_X1 U8536 ( .A(n8807), .ZN(n8392) );
  NAND2_X1 U8537 ( .A1(n8387), .A2(n8386), .ZN(n8713) );
  AND4_X1 U8538 ( .A1(n8675), .A2(n8674), .A3(n8673), .A4(n8672), .ZN(n14639)
         );
  OR2_X1 U8539 ( .A1(n8983), .A2(n8982), .ZN(n11493) );
  OR2_X1 U8540 ( .A1(n7270), .A2(n6698), .ZN(n7269) );
  AND2_X1 U8541 ( .A1(n6794), .A2(n8570), .ZN(n7270) );
  NAND2_X1 U8542 ( .A1(n11883), .A2(n11882), .ZN(n11979) );
  INV_X1 U8543 ( .A(n15272), .ZN(n15268) );
  OR2_X1 U8544 ( .A1(n8571), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8584) );
  AND2_X1 U8545 ( .A1(n11877), .A2(n11874), .ZN(n15283) );
  NAND2_X1 U8546 ( .A1(n11315), .A2(n8570), .ZN(n15284) );
  NOR2_X1 U8547 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8551) );
  INV_X1 U8548 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8550) );
  AND3_X1 U8549 ( .A1(n8566), .A2(n8565), .A3(n8564), .ZN(n11311) );
  AND3_X1 U8550 ( .A1(n8548), .A2(n8547), .A3(n8546), .ZN(n11158) );
  INV_X1 U8551 ( .A(n11152), .ZN(n11976) );
  NAND2_X1 U8552 ( .A1(n7260), .A2(n8520), .ZN(n11015) );
  OR2_X1 U8553 ( .A1(n8815), .A2(n9787), .ZN(n8519) );
  CLKBUF_X1 U8554 ( .A(n6999), .Z(n15308) );
  AND2_X1 U8555 ( .A1(n10415), .A2(n10414), .ZN(n10475) );
  NAND2_X1 U8556 ( .A1(n11842), .A2(n11841), .ZN(n11849) );
  AND2_X1 U8557 ( .A1(n8896), .A2(n7255), .ZN(n7254) );
  NAND2_X1 U8558 ( .A1(n7257), .A2(n7256), .ZN(n7255) );
  AOI21_X1 U8559 ( .B1(n7249), .B2(n6721), .A(n12830), .ZN(n7247) );
  AND2_X1 U8560 ( .A1(n11851), .A2(n8935), .ZN(n15311) );
  INV_X1 U8561 ( .A(n11982), .ZN(n11597) );
  OR2_X1 U8562 ( .A1(n10473), .A2(n8970), .ZN(n10291) );
  INV_X1 U8563 ( .A(n10476), .ZN(n10413) );
  INV_X1 U8564 ( .A(n15328), .ZN(n15339) );
  INV_X1 U8565 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8479) );
  OR2_X1 U8566 ( .A1(n8885), .A2(n8474), .ZN(n8476) );
  NOR2_X1 U8567 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7631) );
  INV_X1 U8568 ( .A(n7587), .ZN(n7586) );
  AOI21_X1 U8569 ( .B1(n7585), .B2(n7587), .A(n6837), .ZN(n7584) );
  NOR2_X1 U8570 ( .A1(n8826), .A2(n7588), .ZN(n7587) );
  OR2_X1 U8571 ( .A1(n8916), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8918) );
  OAI21_X1 U8572 ( .B1(n8460), .B2(P1_DATAO_REG_20__SCAN_IN), .A(n8461), .ZN(
        n8802) );
  AOI21_X1 U8573 ( .B1(n7574), .B2(n7576), .A(n7573), .ZN(n7572) );
  INV_X1 U8574 ( .A(n8455), .ZN(n7573) );
  NAND2_X1 U8575 ( .A1(n8679), .A2(n6821), .ZN(n7566) );
  NAND2_X1 U8576 ( .A1(n7565), .A2(n10016), .ZN(n7564) );
  INV_X1 U8577 ( .A(n8445), .ZN(n7565) );
  NAND2_X1 U8578 ( .A1(n8665), .A2(n8443), .ZN(n8677) );
  AND2_X1 U8579 ( .A1(n8445), .A2(n8444), .ZN(n8676) );
  NAND2_X1 U8580 ( .A1(n8439), .A2(n8438), .ZN(n8645) );
  AND2_X1 U8581 ( .A1(n8441), .A2(n8440), .ZN(n8644) );
  AOI21_X1 U8582 ( .B1(n7593), .B2(n7591), .A(n7590), .ZN(n7589) );
  INV_X1 U8583 ( .A(n7593), .ZN(n7592) );
  INV_X1 U8584 ( .A(n8430), .ZN(n7591) );
  AND2_X1 U8585 ( .A1(n8435), .A2(n8434), .ZN(n8614) );
  AND2_X1 U8586 ( .A1(n8541), .A2(n8402), .ZN(n7533) );
  INV_X1 U8587 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7535) );
  AND2_X1 U8588 ( .A1(n8541), .A2(n8560), .ZN(n7532) );
  AND2_X1 U8589 ( .A1(n8400), .A2(n8402), .ZN(n7531) );
  AND2_X1 U8590 ( .A1(n8428), .A2(n8427), .ZN(n8557) );
  AND2_X1 U8591 ( .A1(n8422), .A2(n8421), .ZN(n8525) );
  NAND2_X1 U8592 ( .A1(n8418), .A2(n8417), .ZN(n8516) );
  NAND2_X1 U8593 ( .A1(n9426), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U8594 ( .A1(n13308), .A2(n13177), .ZN(n13180) );
  AND2_X1 U8595 ( .A1(n13174), .A2(n13166), .ZN(n6901) );
  NAND2_X1 U8596 ( .A1(n11137), .A2(n7471), .ZN(n7470) );
  INV_X1 U8597 ( .A(n11138), .ZN(n7471) );
  NOR2_X1 U8598 ( .A1(n13330), .A2(n13189), .ZN(n7419) );
  AND2_X1 U8599 ( .A1(n9667), .A2(n9661), .ZN(n9958) );
  NAND2_X1 U8600 ( .A1(n7433), .A2(n7430), .ZN(n13138) );
  OAI21_X1 U8601 ( .B1(n7435), .B2(n7432), .A(n13134), .ZN(n7431) );
  OAI211_X1 U8602 ( .C1(n13771), .C2(n9617), .A(n9616), .B(n9615), .ZN(n9618)
         );
  NOR2_X1 U8603 ( .A1(n9533), .A2(n7503), .ZN(n7500) );
  AND2_X1 U8604 ( .A1(n7763), .A2(n7499), .ZN(n7498) );
  NAND2_X1 U8605 ( .A1(n9534), .A2(n6761), .ZN(n7499) );
  INV_X1 U8606 ( .A(n9623), .ZN(n7483) );
  AND4_X1 U8607 ( .A1(n9575), .A2(n9574), .A3(n9573), .A4(n9572), .ZN(n13230)
         );
  AND2_X1 U8608 ( .A1(n9409), .A2(n9408), .ZN(n9626) );
  AND3_X1 U8609 ( .A1(n9343), .A2(n9342), .A3(n9341), .ZN(n13137) );
  AND4_X1 U8610 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), .ZN(n11531)
         );
  AND4_X1 U8611 ( .A1(n9281), .A2(n9280), .A3(n9279), .A4(n9278), .ZN(n11279)
         );
  AND4_X1 U8612 ( .A1(n9242), .A2(n9241), .A3(n9240), .A4(n9239), .ZN(n11115)
         );
  OR2_X1 U8613 ( .A1(n10172), .A2(n10171), .ZN(n11667) );
  OR2_X1 U8614 ( .A1(n14972), .A2(n14971), .ZN(n14974) );
  AND2_X1 U8615 ( .A1(n15034), .A2(n15033), .ZN(n15037) );
  AOI21_X1 U8616 ( .B1(n13511), .B2(n13514), .A(n6864), .ZN(n13496) );
  AND2_X1 U8617 ( .A1(n13522), .A2(n13480), .ZN(n6864) );
  INV_X1 U8618 ( .A(n13481), .ZN(n13500) );
  NOR2_X1 U8619 ( .A1(n13517), .A2(n13503), .ZN(n13502) );
  OAI21_X1 U8620 ( .B1(n6696), .B2(n7384), .A(n7382), .ZN(n13534) );
  AOI21_X1 U8621 ( .B1(n7385), .B2(n7383), .A(n6764), .ZN(n7382) );
  INV_X1 U8622 ( .A(n7385), .ZN(n7384) );
  INV_X1 U8623 ( .A(n6865), .ZN(n7327) );
  NAND2_X1 U8624 ( .A1(n7236), .A2(n7235), .ZN(n13561) );
  INV_X1 U8625 ( .A(n7234), .ZN(n13547) );
  AND2_X1 U8626 ( .A1(n13617), .A2(n13635), .ZN(n13614) );
  NAND2_X1 U8627 ( .A1(n7049), .A2(n7047), .ZN(n13626) );
  AOI21_X1 U8628 ( .B1(n7050), .B2(n11698), .A(n7048), .ZN(n7047) );
  NOR2_X1 U8629 ( .A1(n7369), .A2(n7051), .ZN(n7050) );
  AND3_X1 U8630 ( .A1(n11568), .A2(n6702), .A3(n7232), .ZN(n13652) );
  NOR2_X1 U8631 ( .A1(n13749), .A2(n13672), .ZN(n7232) );
  OR2_X1 U8632 ( .A1(n13813), .A2(n13451), .ZN(n13664) );
  OR2_X1 U8633 ( .A1(n11692), .A2(n11698), .ZN(n13454) );
  NAND2_X1 U8634 ( .A1(n11568), .A2(n13355), .ZN(n11694) );
  NAND2_X1 U8635 ( .A1(n11568), .A2(n6702), .ZN(n13671) );
  INV_X1 U8636 ( .A(n11699), .ZN(n7334) );
  NOR2_X1 U8637 ( .A1(n11566), .A2(n7332), .ZN(n7331) );
  NAND2_X1 U8638 ( .A1(n11564), .A2(n11698), .ZN(n7332) );
  NOR2_X1 U8639 ( .A1(n11566), .A2(n7333), .ZN(n7335) );
  AND4_X1 U8640 ( .A1(n7229), .A2(n14668), .A3(n7228), .A4(n11129), .ZN(n11548) );
  AND2_X1 U8641 ( .A1(n11648), .A2(n11548), .ZN(n11568) );
  INV_X1 U8642 ( .A(n7279), .ZN(n7278) );
  OAI21_X1 U8643 ( .B1(n6735), .B2(n11278), .A(n11380), .ZN(n7279) );
  OR2_X1 U8644 ( .A1(n9294), .A2(n9293), .ZN(n9310) );
  NAND2_X1 U8645 ( .A1(n11129), .A2(n15112), .ZN(n11333) );
  NAND2_X1 U8646 ( .A1(n6909), .A2(n7358), .ZN(n11277) );
  CLKBUF_X1 U8647 ( .A(n11332), .Z(n6873) );
  OAI21_X1 U8648 ( .B1(n10844), .B2(n10821), .A(n7360), .ZN(n11116) );
  OR2_X1 U8649 ( .A1(n9222), .A2(n9221), .ZN(n9237) );
  OR2_X1 U8650 ( .A1(n15060), .A2(n10817), .ZN(n10845) );
  NOR2_X1 U8651 ( .A1(n10845), .A2(n10850), .ZN(n10847) );
  AND2_X1 U8652 ( .A1(n7287), .A2(n6810), .ZN(n7286) );
  AND2_X1 U8653 ( .A1(n10655), .A2(n10798), .ZN(n15061) );
  NAND2_X1 U8654 ( .A1(n10211), .A2(n10210), .ZN(n7356) );
  NAND2_X1 U8655 ( .A1(n7044), .A2(n10178), .ZN(n10190) );
  INV_X1 U8656 ( .A(n10182), .ZN(n7044) );
  CLKBUF_X1 U8657 ( .A(n9562), .Z(n10460) );
  NAND2_X1 U8658 ( .A1(n7056), .A2(n13463), .ZN(n13603) );
  NAND2_X1 U8659 ( .A1(n7087), .A2(n9032), .ZN(n13741) );
  NAND2_X1 U8660 ( .A1(n11256), .A2(n9579), .ZN(n7087) );
  NAND2_X1 U8661 ( .A1(n9323), .A2(n9322), .ZN(n11553) );
  NAND2_X1 U8662 ( .A1(n7367), .A2(n10800), .ZN(n15057) );
  NAND2_X1 U8663 ( .A1(n10799), .A2(n10812), .ZN(n10800) );
  OAI21_X1 U8664 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n15068) );
  NOR2_X1 U8665 ( .A1(n7281), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7280) );
  INV_X1 U8666 ( .A(n9029), .ZN(n7281) );
  INV_X1 U8667 ( .A(n9656), .ZN(n9653) );
  CLKBUF_X1 U8668 ( .A(n9286), .Z(n9287) );
  OR2_X1 U8669 ( .A1(n9214), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9216) );
  OR2_X1 U8670 ( .A1(n9216), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9251) );
  OR2_X1 U8671 ( .A1(n9158), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9288) );
  AND2_X1 U8672 ( .A1(n6677), .A2(n9014), .ZN(n9144) );
  INV_X1 U8673 ( .A(n8205), .ZN(n8218) );
  NAND2_X1 U8674 ( .A1(n7747), .A2(n7745), .ZN(n13882) );
  NOR2_X1 U8675 ( .A1(n13883), .A2(n7746), .ZN(n7745) );
  INV_X1 U8676 ( .A(n12311), .ZN(n7746) );
  NAND2_X1 U8677 ( .A1(n13949), .A2(n13948), .ZN(n7747) );
  NAND2_X1 U8678 ( .A1(n13938), .A2(n12348), .ZN(n13904) );
  NAND2_X1 U8679 ( .A1(n13850), .A2(n7748), .ZN(n12282) );
  NOR2_X1 U8680 ( .A1(n6746), .A2(n7749), .ZN(n7748) );
  AND3_X1 U8681 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7966) );
  AND2_X1 U8682 ( .A1(n8123), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8137) );
  XNOR2_X1 U8683 ( .A(n11243), .B(n11241), .ZN(n11259) );
  NOR2_X1 U8684 ( .A1(n8175), .A2(n8174), .ZN(n8192) );
  OR3_X1 U8685 ( .A1(n8031), .A2(n8029), .A3(n8030), .ZN(n8047) );
  OAI21_X1 U8686 ( .B1(n7904), .B2(n6683), .A(n6966), .ZN(n10372) );
  NAND2_X1 U8687 ( .A1(n11247), .A2(n6967), .ZN(n6966) );
  OR2_X1 U8688 ( .A1(n8267), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U8689 ( .A1(n10072), .A2(n6744), .ZN(n10093) );
  OR2_X1 U8690 ( .A1(n10246), .A2(n6964), .ZN(n6963) );
  AND2_X1 U8691 ( .A1(n10250), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U8692 ( .A1(n6963), .A2(n6962), .ZN(n7349) );
  INV_X1 U8693 ( .A(n10091), .ZN(n6962) );
  NAND2_X1 U8694 ( .A1(n10116), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7346) );
  OR2_X1 U8695 ( .A1(n10154), .A2(n10155), .ZN(n6911) );
  NOR2_X1 U8696 ( .A1(n11168), .A2(n7352), .ZN(n14739) );
  AND2_X1 U8697 ( .A1(n11174), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7352) );
  NOR2_X1 U8698 ( .A1(n11173), .A2(n6914), .ZN(n14735) );
  AND2_X1 U8699 ( .A1(n11174), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6914) );
  NAND2_X1 U8700 ( .A1(n14735), .A2(n14734), .ZN(n14733) );
  NAND2_X1 U8701 ( .A1(n11177), .A2(n11178), .ZN(n14057) );
  XNOR2_X1 U8702 ( .A(n14061), .B(n8104), .ZN(n14773) );
  NAND2_X1 U8703 ( .A1(n14758), .A2(n6915), .ZN(n14061) );
  OR2_X1 U8704 ( .A1(n14060), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6915) );
  AOI21_X1 U8705 ( .B1(n14795), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14790), .ZN(
        n14806) );
  NOR2_X1 U8706 ( .A1(n14816), .A2(n14817), .ZN(n14815) );
  NOR2_X1 U8707 ( .A1(n14821), .A2(n14822), .ZN(n14820) );
  OAI21_X1 U8708 ( .B1(n14139), .B2(n7393), .A(n6720), .ZN(n14125) );
  AND2_X1 U8709 ( .A1(n14140), .A2(n7118), .ZN(n14128) );
  AND2_X1 U8710 ( .A1(n14127), .A2(n14126), .ZN(n7118) );
  NAND2_X1 U8711 ( .A1(n14139), .A2(n14144), .ZN(n14140) );
  NAND2_X1 U8712 ( .A1(n14158), .A2(n8248), .ZN(n14145) );
  NAND2_X1 U8713 ( .A1(n7132), .A2(n7131), .ZN(n14160) );
  NAND2_X1 U8714 ( .A1(n14213), .A2(n14372), .ZN(n14196) );
  AOI21_X1 U8715 ( .B1(n14247), .B2(n7712), .A(n6765), .ZN(n7711) );
  NAND2_X1 U8716 ( .A1(n8164), .A2(n8163), .ZN(n14265) );
  NOR2_X1 U8717 ( .A1(n7704), .A2(n7703), .ZN(n7702) );
  INV_X1 U8718 ( .A(n8129), .ZN(n7703) );
  OAI21_X1 U8719 ( .B1(n14314), .B2(n14327), .A(n8320), .ZN(n14303) );
  NAND2_X1 U8720 ( .A1(n7110), .A2(n14294), .ZN(n14307) );
  INV_X1 U8721 ( .A(n14303), .ZN(n7110) );
  NAND2_X1 U8722 ( .A1(n11464), .A2(n6701), .ZN(n14332) );
  NAND2_X1 U8723 ( .A1(n11464), .A2(n8337), .ZN(n14330) );
  INV_X1 U8724 ( .A(n12216), .ZN(n11456) );
  AOI21_X1 U8725 ( .B1(n7400), .B2(n7398), .A(n6768), .ZN(n7397) );
  INV_X1 U8726 ( .A(n7400), .ZN(n7399) );
  NAND2_X1 U8727 ( .A1(n8006), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U8728 ( .A1(n7405), .A2(n8310), .ZN(n11086) );
  NAND2_X1 U8729 ( .A1(n10548), .A2(n12038), .ZN(n11045) );
  NOR2_X1 U8730 ( .A1(n10622), .A2(n12033), .ZN(n10548) );
  INV_X1 U8731 ( .A(n10888), .ZN(n14091) );
  INV_X1 U8732 ( .A(n12201), .ZN(n10615) );
  NAND2_X1 U8733 ( .A1(n7128), .A2(n7127), .ZN(n10622) );
  INV_X1 U8734 ( .A(n8217), .ZN(n11810) );
  OR2_X1 U8735 ( .A1(n14043), .A2(n12017), .ZN(n12019) );
  AND2_X1 U8736 ( .A1(n8339), .A2(n14079), .ZN(n14088) );
  INV_X1 U8737 ( .A(n14251), .ZN(n14459) );
  INV_X1 U8738 ( .A(n14855), .ZN(n14684) );
  INV_X1 U8739 ( .A(n14239), .ZN(n14395) );
  NAND2_X1 U8740 ( .A1(n9554), .A2(n9542), .ZN(n9545) );
  NAND2_X1 U8741 ( .A1(n7664), .A2(n7668), .ZN(n9536) );
  NAND2_X1 U8742 ( .A1(n8263), .A2(n7671), .ZN(n7664) );
  AND2_X1 U8743 ( .A1(n7709), .A2(n7862), .ZN(n7707) );
  INV_X1 U8744 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7866) );
  XNOR2_X1 U8745 ( .A(n8279), .B(n8278), .ZN(n13825) );
  NAND2_X1 U8746 ( .A1(n7145), .A2(n7142), .ZN(n8279) );
  NOR2_X1 U8747 ( .A1(n7144), .A2(n7143), .ZN(n7142) );
  INV_X1 U8748 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7862) );
  INV_X1 U8749 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7709) );
  XNOR2_X1 U8750 ( .A(n8360), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U8751 ( .A1(n6724), .A2(n7708), .ZN(n8359) );
  INV_X1 U8752 ( .A(n8133), .ZN(n7708) );
  OAI21_X1 U8753 ( .B1(n8239), .B2(n8238), .A(n7852), .ZN(n8251) );
  XNOR2_X1 U8754 ( .A(n8227), .B(n8226), .ZN(n11635) );
  NAND2_X1 U8755 ( .A1(n8186), .A2(n8185), .ZN(n8189) );
  NAND2_X1 U8756 ( .A1(n8289), .A2(n7754), .ZN(n7753) );
  OAI21_X1 U8757 ( .B1(n7824), .B2(n7648), .A(n7646), .ZN(n8132) );
  NAND2_X1 U8758 ( .A1(n7824), .A2(n7823), .ZN(n8118) );
  XNOR2_X1 U8759 ( .A(n8094), .B(n8093), .ZN(n10334) );
  NAND2_X1 U8760 ( .A1(n7133), .A2(n7136), .ZN(n8041) );
  OR2_X1 U8761 ( .A1(n7806), .A2(n7140), .ZN(n7133) );
  NAND2_X1 U8762 ( .A1(n7651), .A2(n7809), .ZN(n8023) );
  NAND2_X1 U8763 ( .A1(n8014), .A2(n7807), .ZN(n7651) );
  XNOR2_X1 U8764 ( .A(n7959), .B(n7958), .ZN(n9820) );
  INV_X1 U8765 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n15757) );
  XNOR2_X1 U8766 ( .A(n7779), .B(SI_1_), .ZN(n7895) );
  OAI211_X1 U8767 ( .C1(n7227), .C2(n7158), .A(n7156), .B(n7155), .ZN(n7159)
         );
  NAND2_X1 U8768 ( .A1(n7157), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7156) );
  XNOR2_X1 U8769 ( .A(n14532), .B(n7242), .ZN(n14541) );
  XNOR2_X1 U8770 ( .A(n14543), .B(n14544), .ZN(n14545) );
  NAND2_X1 U8771 ( .A1(n7238), .A2(n14552), .ZN(n14553) );
  OAI21_X1 U8772 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15687), .A(n14514), .ZN(
        n14562) );
  NAND2_X1 U8773 ( .A1(n14519), .A2(n14518), .ZN(n14568) );
  OAI21_X1 U8774 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15208), .A(n14522), .ZN(
        n14530) );
  NAND2_X1 U8775 ( .A1(n11580), .A2(n11579), .ZN(n15137) );
  AND2_X1 U8776 ( .A1(n12415), .A2(n12414), .ZN(n12452) );
  NAND2_X1 U8777 ( .A1(n12400), .A2(n12399), .ZN(n15148) );
  NAND2_X1 U8778 ( .A1(n12400), .A2(n7556), .ZN(n15156) );
  NOR2_X1 U8779 ( .A1(n15147), .A2(n7557), .ZN(n7556) );
  INV_X1 U8780 ( .A(n12399), .ZN(n7557) );
  NAND2_X1 U8781 ( .A1(n12473), .A2(n12472), .ZN(n12471) );
  NAND2_X1 U8782 ( .A1(n7537), .A2(n7536), .ZN(n12504) );
  AOI21_X1 U8783 ( .B1(n7538), .B2(n7540), .A(n6776), .ZN(n7536) );
  NAND2_X1 U8784 ( .A1(n8863), .A2(n8862), .ZN(n12811) );
  NAND2_X1 U8785 ( .A1(n7529), .A2(n7526), .ZN(n12538) );
  INV_X1 U8786 ( .A(n7528), .ZN(n7526) );
  NAND2_X1 U8787 ( .A1(n7529), .A2(n7527), .ZN(n12539) );
  AND3_X1 U8788 ( .A1(n8634), .A2(n8633), .A3(n8632), .ZN(n11885) );
  NAND2_X1 U8789 ( .A1(n12471), .A2(n12429), .ZN(n12557) );
  OAI21_X1 U8790 ( .B1(n12473), .B2(n7540), .A(n7538), .ZN(n12555) );
  AND2_X1 U8791 ( .A1(n8667), .A2(n8666), .ZN(n12587) );
  NAND2_X1 U8792 ( .A1(n7519), .A2(n7523), .ZN(n12594) );
  NAND2_X1 U8793 ( .A1(n6912), .A2(n7527), .ZN(n7519) );
  AND2_X1 U8794 ( .A1(n12612), .A2(n12418), .ZN(n7558) );
  AND2_X1 U8795 ( .A1(n12451), .A2(n12418), .ZN(n12613) );
  INV_X1 U8796 ( .A(n11844), .ZN(n12752) );
  AND2_X1 U8797 ( .A1(n10957), .A2(n8925), .ZN(n11845) );
  AND2_X1 U8798 ( .A1(n10957), .A2(n8909), .ZN(n12767) );
  NAND2_X1 U8799 ( .A1(n8870), .A2(n8869), .ZN(n12821) );
  NAND2_X1 U8800 ( .A1(n8858), .A2(n8857), .ZN(n12522) );
  INV_X1 U8801 ( .A(n14639), .ZN(n12566) );
  NAND4_X1 U8802 ( .A1(n8627), .A2(n8626), .A3(n8625), .A4(n8624), .ZN(n12496)
         );
  NAND4_X1 U8803 ( .A1(n8589), .A2(n8588), .A3(n8587), .A4(n8586), .ZN(n12497)
         );
  NAND2_X1 U8804 ( .A1(n15161), .A2(n6844), .ZN(n15163) );
  XNOR2_X1 U8805 ( .A(n9719), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10692) );
  AND2_X1 U8806 ( .A1(n8528), .A2(n8543), .ZN(n10611) );
  NAND2_X1 U8807 ( .A1(n9727), .A2(n10604), .ZN(n10608) );
  NAND2_X1 U8808 ( .A1(n9738), .A2(n10555), .ZN(n10575) );
  NAND2_X1 U8809 ( .A1(n9749), .A2(n10632), .ZN(n10637) );
  INV_X1 U8810 ( .A(n9706), .ZN(n7219) );
  INV_X1 U8811 ( .A(n9690), .ZN(n7292) );
  INV_X1 U8812 ( .A(n7293), .ZN(n9691) );
  INV_X1 U8813 ( .A(n7339), .ZN(n15206) );
  AND2_X1 U8814 ( .A1(n8685), .A2(n8708), .ZN(n15214) );
  INV_X1 U8815 ( .A(n6952), .ZN(n15239) );
  INV_X1 U8816 ( .A(n7224), .ZN(n15261) );
  NOR2_X1 U8817 ( .A1(n15223), .A2(n12669), .ZN(n15247) );
  NOR2_X1 U8818 ( .A1(n14627), .A2(n12634), .ZN(n12636) );
  AND2_X1 U8819 ( .A1(n12721), .A2(n12720), .ZN(n12722) );
  AND2_X1 U8820 ( .A1(n12702), .A2(n12718), .ZN(n6965) );
  OAI21_X1 U8821 ( .B1(n15289), .B2(n12786), .A(n12785), .ZN(n12972) );
  AND2_X1 U8822 ( .A1(n12871), .A2(n12870), .ZN(n13002) );
  AND2_X1 U8823 ( .A1(n11734), .A2(n8668), .ZN(n11724) );
  AND2_X1 U8824 ( .A1(n11606), .A2(n8651), .ZN(n11735) );
  INV_X1 U8825 ( .A(n14652), .ZN(n12953) );
  NOR2_X1 U8826 ( .A1(n7252), .A2(n6727), .ZN(n11496) );
  INV_X1 U8827 ( .A(n6992), .ZN(n6991) );
  OAI22_X1 U8828 ( .A1(n8815), .A2(n9781), .B1(n9692), .B2(n9783), .ZN(n6992)
         );
  AND2_X1 U8829 ( .A1(n10480), .A2(n15307), .ZN(n15337) );
  INV_X1 U8830 ( .A(n15307), .ZN(n15332) );
  NAND2_X1 U8831 ( .A1(n8904), .A2(n8903), .ZN(n12965) );
  INV_X2 U8832 ( .A(n15394), .ZN(n15396) );
  INV_X1 U8833 ( .A(n11849), .ZN(n13027) );
  NAND2_X1 U8834 ( .A1(n11835), .A2(n11834), .ZN(n13028) );
  NAND2_X1 U8835 ( .A1(n8875), .A2(n8874), .ZN(n13044) );
  AOI21_X1 U8836 ( .B1(n12797), .B2(n15322), .A(n12796), .ZN(n13042) );
  XOR2_X1 U8837 ( .A(n12794), .B(n12793), .Z(n13047) );
  NAND2_X1 U8838 ( .A1(n12829), .A2(n11950), .ZN(n12818) );
  NAND2_X1 U8839 ( .A1(n12855), .A2(n8825), .ZN(n12844) );
  OR2_X1 U8840 ( .A1(n10675), .A2(n8815), .ZN(n8817) );
  AND2_X1 U8841 ( .A1(n12862), .A2(n12861), .ZN(n13068) );
  NAND2_X1 U8842 ( .A1(n13000), .A2(n11937), .ZN(n12854) );
  NAND2_X1 U8843 ( .A1(n8792), .A2(n8791), .ZN(n13080) );
  NAND2_X1 U8844 ( .A1(n8774), .A2(n8773), .ZN(n13083) );
  AND2_X1 U8845 ( .A1(n12914), .A2(n12913), .ZN(n13088) );
  NAND2_X1 U8846 ( .A1(n8746), .A2(n8745), .ZN(n13095) );
  NAND2_X1 U8847 ( .A1(n8727), .A2(n8726), .ZN(n13102) );
  INV_X1 U8848 ( .A(n13114), .ZN(n13101) );
  NAND2_X1 U8849 ( .A1(n7605), .A2(n7608), .ZN(n12933) );
  NAND2_X1 U8850 ( .A1(n14634), .A2(n7610), .ZN(n7605) );
  NAND2_X1 U8851 ( .A1(n8712), .A2(n8711), .ZN(n13113) );
  NAND2_X1 U8852 ( .A1(n7612), .A2(n11905), .ZN(n12943) );
  NAND2_X1 U8853 ( .A1(n7614), .A2(n7613), .ZN(n7612) );
  INV_X1 U8854 ( .A(n14634), .ZN(n7614) );
  AND2_X1 U8855 ( .A1(n15382), .A2(n15368), .ZN(n13109) );
  INV_X1 U8856 ( .A(n12587), .ZN(n14651) );
  OAI211_X1 U8857 ( .C1(n11083), .C2(n9692), .A(n8649), .B(n8648), .ZN(n15153)
         );
  CLKBUF_X1 U8858 ( .A(n10481), .Z(n6935) );
  AND2_X1 U8859 ( .A1(n8953), .A2(n8952), .ZN(n13116) );
  AND2_X1 U8860 ( .A1(n10283), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13115) );
  NAND2_X1 U8861 ( .A1(n13121), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U8862 ( .A1(n8467), .A2(n11637), .ZN(n7603) );
  NAND2_X1 U8863 ( .A1(n7599), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U8864 ( .A1(n8814), .A2(n8463), .ZN(n8827) );
  NAND2_X1 U8865 ( .A1(n8739), .A2(n8452), .ZN(n8755) );
  INV_X1 U8866 ( .A(SI_16_), .ZN(n15453) );
  INV_X1 U8867 ( .A(SI_12_), .ZN(n15480) );
  INV_X1 U8868 ( .A(SI_11_), .ZN(n9800) );
  AND2_X1 U8869 ( .A1(n8596), .A2(n8595), .ZN(n9789) );
  NAND2_X1 U8870 ( .A1(n7595), .A2(n7593), .ZN(n8596) );
  NAND2_X1 U8871 ( .A1(n7595), .A2(n8431), .ZN(n8594) );
  OR2_X1 U8872 ( .A1(n8563), .A2(n8562), .ZN(n9774) );
  INV_X1 U8873 ( .A(n9728), .ZN(n10539) );
  INV_X1 U8874 ( .A(n10611), .ZN(n9778) );
  INV_X1 U8875 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9810) );
  OR2_X1 U8876 ( .A1(n11528), .A2(n7435), .ZN(n13135) );
  NOR2_X1 U8877 ( .A1(n11528), .A2(n11527), .ZN(n11530) );
  XNOR2_X1 U8878 ( .A(n13180), .B(n13178), .ZN(n13210) );
  NAND2_X1 U8879 ( .A1(n13210), .A2(n13209), .ZN(n13208) );
  NAND2_X1 U8880 ( .A1(n6898), .A2(n10938), .ZN(n11140) );
  INV_X1 U8881 ( .A(n7453), .ZN(n7452) );
  AND2_X1 U8882 ( .A1(n7451), .A2(n10752), .ZN(n7450) );
  NAND2_X1 U8883 ( .A1(n7453), .A2(n6726), .ZN(n7451) );
  OAI21_X1 U8884 ( .B1(n7449), .B2(n6726), .A(n7453), .ZN(n10753) );
  INV_X1 U8885 ( .A(n7455), .ZN(n7449) );
  NAND2_X1 U8886 ( .A1(n9397), .A2(n13377), .ZN(n7282) );
  NOR2_X1 U8887 ( .A1(n9928), .A2(n9927), .ZN(n9971) );
  NAND2_X1 U8888 ( .A1(n7463), .A2(n7464), .ZN(n11353) );
  NAND2_X1 U8889 ( .A1(n7467), .A2(n7465), .ZN(n7463) );
  NAND2_X1 U8890 ( .A1(n7442), .A2(n7446), .ZN(n7443) );
  NAND2_X1 U8891 ( .A1(n13283), .A2(n13282), .ZN(n13281) );
  NOR2_X1 U8892 ( .A1(n11522), .A2(n11521), .ZN(n11528) );
  NAND2_X1 U8893 ( .A1(n7467), .A2(n7470), .ZN(n11347) );
  NAND2_X1 U8894 ( .A1(n13151), .A2(n13150), .ZN(n13320) );
  NAND2_X1 U8895 ( .A1(n13242), .A2(n13190), .ZN(n13329) );
  CLKBUF_X1 U8896 ( .A(n13341), .Z(n13342) );
  NAND2_X1 U8897 ( .A1(n6788), .A2(n7482), .ZN(n7481) );
  INV_X1 U8898 ( .A(n6961), .ZN(n7482) );
  INV_X1 U8899 ( .A(n11560), .ZN(n13361) );
  OR2_X1 U8900 ( .A1(n9558), .A2(n9124), .ZN(n9125) );
  NOR2_X1 U8901 ( .A1(n7414), .A2(n7381), .ZN(n7413) );
  INV_X1 U8902 ( .A(n13775), .ZN(n13418) );
  INV_X1 U8903 ( .A(n13487), .ZN(n13414) );
  AOI21_X1 U8904 ( .B1(n13482), .B2(n13331), .A(n7324), .ZN(n7323) );
  NOR2_X1 U8905 ( .A1(n13450), .A2(n13449), .ZN(n7324) );
  NAND2_X1 U8906 ( .A1(n13503), .A2(n13482), .ZN(n13483) );
  NAND2_X1 U8907 ( .A1(n13559), .A2(n7385), .ZN(n13544) );
  AND2_X1 U8908 ( .A1(n13559), .A2(n13474), .ZN(n13546) );
  NAND2_X1 U8909 ( .A1(n7326), .A2(n7328), .ZN(n13539) );
  NAND2_X1 U8910 ( .A1(n7342), .A2(n13436), .ZN(n13571) );
  NAND2_X1 U8911 ( .A1(n13587), .A2(n13468), .ZN(n13580) );
  NOR2_X1 U8912 ( .A1(n13466), .A2(n7768), .ZN(n13589) );
  NAND2_X1 U8913 ( .A1(n13434), .A2(n13433), .ZN(n13584) );
  INV_X1 U8914 ( .A(n13741), .ZN(n13617) );
  NAND2_X1 U8915 ( .A1(n13631), .A2(n13627), .ZN(n13619) );
  NAND2_X1 U8916 ( .A1(n7371), .A2(n13456), .ZN(n13657) );
  NAND2_X1 U8917 ( .A1(n7364), .A2(n11561), .ZN(n11689) );
  NAND2_X1 U8918 ( .A1(n11326), .A2(n11278), .ZN(n11379) );
  NAND2_X1 U8919 ( .A1(n11287), .A2(n11286), .ZN(n11383) );
  NAND2_X1 U8920 ( .A1(n7306), .A2(n10820), .ZN(n11119) );
  NAND2_X1 U8921 ( .A1(n10853), .A2(n10852), .ZN(n7306) );
  NAND2_X1 U8922 ( .A1(n15059), .A2(n10802), .ZN(n10828) );
  NAND2_X1 U8923 ( .A1(n7291), .A2(n10813), .ZN(n15046) );
  INV_X1 U8924 ( .A(n15062), .ZN(n13673) );
  NAND2_X1 U8925 ( .A1(n11340), .A2(n10644), .ZN(n13609) );
  OR2_X1 U8926 ( .A1(n9796), .A2(n9555), .ZN(n9134) );
  INV_X1 U8927 ( .A(n13406), .ZN(n13771) );
  INV_X1 U8928 ( .A(n7323), .ZN(n7320) );
  NAND2_X1 U8929 ( .A1(n7319), .A2(n7325), .ZN(n7321) );
  INV_X1 U8930 ( .A(n13522), .ZN(n13784) );
  AND2_X1 U8931 ( .A1(n9400), .A2(n9399), .ZN(n13804) );
  INV_X1 U8932 ( .A(n11553), .ZN(n11648) );
  AND3_X1 U8933 ( .A1(n9150), .A2(n9149), .A3(n9148), .ZN(n10339) );
  AND4_X1 U8934 ( .A1(n7480), .A2(n9015), .A3(n7479), .A4(n7758), .ZN(n7415)
         );
  MUX2_X1 U8935 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9035), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n9036) );
  INV_X1 U8936 ( .A(n9094), .ZN(n13400) );
  INV_X1 U8937 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9850) );
  INV_X1 U8938 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9840) );
  INV_X1 U8939 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9833) );
  INV_X1 U8940 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9831) );
  INV_X1 U8941 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9821) );
  INV_X1 U8942 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9815) );
  INV_X1 U8943 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9795) );
  INV_X1 U8944 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U8945 ( .A1(n12262), .A2(n12261), .ZN(n13852) );
  NAND2_X1 U8946 ( .A1(n7727), .A2(n13865), .ZN(n13868) );
  NAND2_X1 U8947 ( .A1(n6940), .A2(n13866), .ZN(n7727) );
  INV_X1 U8948 ( .A(n7737), .ZN(n7739) );
  NAND2_X1 U8949 ( .A1(n7740), .A2(n7743), .ZN(n10793) );
  INV_X1 U8950 ( .A(n6848), .ZN(n10794) );
  AOI21_X1 U8951 ( .B1(n7734), .B2(n12366), .A(n12374), .ZN(n7733) );
  NAND2_X1 U8952 ( .A1(n7723), .A2(n7722), .ZN(n11746) );
  NAND2_X1 U8953 ( .A1(n11444), .A2(n11617), .ZN(n7723) );
  NAND2_X1 U8954 ( .A1(n10374), .A2(n6876), .ZN(n10376) );
  NAND2_X1 U8955 ( .A1(n6877), .A2(n12329), .ZN(n6876) );
  INV_X1 U8956 ( .A(n10375), .ZN(n6877) );
  NAND2_X1 U8957 ( .A1(n7747), .A2(n12311), .ZN(n13884) );
  NAND2_X1 U8958 ( .A1(n7744), .A2(n6750), .ZN(n13893) );
  AND3_X1 U8959 ( .A1(n8158), .A2(n8157), .A3(n8156), .ZN(n14305) );
  OAI21_X1 U8960 ( .B1(n6940), .B2(n7731), .A(n7728), .ZN(n13939) );
  OR2_X1 U8961 ( .A1(n10352), .A2(n10351), .ZN(n13996) );
  INV_X1 U8962 ( .A(n7744), .ZN(n13892) );
  NAND2_X1 U8963 ( .A1(n6853), .A2(n6852), .ZN(n6850) );
  OAI21_X1 U8964 ( .B1(n6853), .B2(n6852), .A(n6870), .ZN(n6851) );
  AND2_X1 U8965 ( .A1(n10784), .A2(n12240), .ZN(n14010) );
  OR2_X1 U8966 ( .A1(n10352), .A2(n10350), .ZN(n14014) );
  AND2_X1 U8967 ( .A1(n12198), .A2(n6745), .ZN(n12234) );
  INV_X1 U8968 ( .A(n12240), .ZN(n6895) );
  NAND2_X1 U8969 ( .A1(n8195), .A2(n7408), .ZN(n7407) );
  INV_X1 U8970 ( .A(n7349), .ZN(n10113) );
  INV_X1 U8971 ( .A(n6963), .ZN(n10092) );
  AND2_X1 U8972 ( .A1(n10101), .A2(n10100), .ZN(n10106) );
  NAND2_X1 U8973 ( .A1(n10114), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7348) );
  INV_X1 U8974 ( .A(n7347), .ZN(n10304) );
  AOI21_X1 U8975 ( .B1(n10114), .B2(P1_REG1_REG_3__SCAN_IN), .A(n10106), .ZN(
        n10303) );
  INV_X1 U8976 ( .A(n6911), .ZN(n10153) );
  AND2_X1 U8977 ( .A1(n6911), .A2(n6910), .ZN(n10143) );
  NAND2_X1 U8978 ( .A1(n10156), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8979 ( .A1(n10110), .A2(n10109), .ZN(n10430) );
  AND2_X1 U8980 ( .A1(n10732), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7353) );
  NAND2_X1 U8981 ( .A1(n14057), .A2(n6974), .ZN(n14747) );
  OR2_X1 U8982 ( .A1(n14058), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6974) );
  AOI21_X1 U8983 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n14754), .A(n14746), .ZN(
        n14760) );
  OAI211_X1 U8984 ( .C1(n14070), .C2(n14789), .A(n14828), .B(n14068), .ZN(
        n6890) );
  INV_X1 U8985 ( .A(n14072), .ZN(n6887) );
  OAI21_X1 U8986 ( .B1(n14075), .B2(n14832), .A(n14074), .ZN(n6886) );
  INV_X1 U8987 ( .A(n14106), .ZN(n6959) );
  NAND2_X1 U8988 ( .A1(n14191), .A2(n8225), .ZN(n14175) );
  OAI21_X1 U8989 ( .B1(n14222), .B2(n7114), .A(n7113), .ZN(n14195) );
  NAND2_X1 U8990 ( .A1(n14222), .A2(n8202), .ZN(n7117) );
  NAND2_X1 U8991 ( .A1(n14244), .A2(n8180), .ZN(n14226) );
  NAND2_X1 U8992 ( .A1(n14259), .A2(n7395), .ZN(n14236) );
  NAND2_X1 U8993 ( .A1(n14326), .A2(n8129), .ZN(n14295) );
  NAND2_X1 U8994 ( .A1(n11468), .A2(n12094), .ZN(n7096) );
  NOR2_X1 U8995 ( .A1(n11213), .A2(n12073), .ZN(n11192) );
  NAND2_X1 U8996 ( .A1(n11026), .A2(n7400), .ZN(n11209) );
  NAND2_X1 U8997 ( .A1(n11026), .A2(n8315), .ZN(n11208) );
  OAI21_X1 U8998 ( .B1(n11025), .B2(n7699), .A(n7696), .ZN(n11211) );
  NAND2_X1 U8999 ( .A1(n11024), .A2(n8012), .ZN(n11212) );
  OAI21_X1 U9000 ( .B1(n11040), .B2(n7693), .A(n7691), .ZN(n11088) );
  NAND2_X1 U9001 ( .A1(n10682), .A2(n10681), .ZN(n10680) );
  NAND2_X1 U9002 ( .A1(n11040), .A2(n7957), .ZN(n10682) );
  NAND2_X1 U9003 ( .A1(n10613), .A2(n7920), .ZN(n10512) );
  AND2_X1 U9004 ( .A1(n14319), .A2(n10886), .ZN(n14329) );
  INV_X1 U9005 ( .A(n14333), .ZN(n14253) );
  INV_X1 U9006 ( .A(n14300), .ZN(n14325) );
  INV_X1 U9007 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7411) );
  AND2_X1 U9008 ( .A1(n14863), .A2(n14680), .ZN(n14345) );
  INV_X1 U9009 ( .A(n8004), .ZN(n6875) );
  NAND2_X1 U9010 ( .A1(n9554), .A2(n9553), .ZN(n14479) );
  NAND2_X1 U9011 ( .A1(n8356), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8357) );
  NAND2_X1 U9012 ( .A1(n9443), .A2(n9442), .ZN(n7641) );
  XNOR2_X1 U9013 ( .A(n8203), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14495) );
  INV_X1 U9014 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10300) );
  INV_X1 U9015 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9842) );
  INV_X1 U9016 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9838) );
  INV_X1 U9017 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9835) );
  INV_X1 U9018 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9829) );
  AND2_X1 U9019 ( .A1(n7977), .A2(n6872), .ZN(n10144) );
  INV_X1 U9020 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9824) );
  INV_X1 U9021 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9817) );
  INV_X1 U9022 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9793) );
  INV_X1 U9023 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9768) );
  INV_X1 U9024 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9797) );
  MUX2_X1 U9025 ( .A(n8290), .B(n7911), .S(P1_IR_REG_2__SCAN_IN), .Z(n7912) );
  NAND2_X1 U9026 ( .A1(n7355), .A2(n8290), .ZN(n7354) );
  CLKBUF_X1 U9027 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n6889) );
  INV_X1 U9028 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6923) );
  AOI21_X1 U9029 ( .B1(n15796), .B2(n14540), .A(n15793), .ZN(n15787) );
  XNOR2_X1 U9030 ( .A(n14553), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15792) );
  NAND2_X1 U9031 ( .A1(n7240), .A2(n14561), .ZN(n14604) );
  NOR2_X1 U9032 ( .A1(n14706), .A2(n14705), .ZN(n14704) );
  AND2_X1 U9033 ( .A1(n6917), .A2(n6916), .ZN(n14720) );
  AOI21_X1 U9034 ( .B1(n15027), .B2(n14580), .A(n14722), .ZN(n14612) );
  NAND2_X1 U9035 ( .A1(n7549), .A2(n15134), .ZN(n7548) );
  NAND2_X1 U9036 ( .A1(n10990), .A2(n10989), .ZN(n10993) );
  OR2_X1 U9037 ( .A1(n12006), .A2(n12005), .ZN(n6905) );
  AOI21_X1 U9038 ( .B1(n15259), .B2(P3_IR_REG_0__SCAN_IN), .A(n7225), .ZN(
        n15166) );
  AND2_X1 U9039 ( .A1(P3_U3151), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7225) );
  OAI211_X1 U9040 ( .C1(n12700), .C2(n15241), .A(n6951), .B(n6728), .ZN(
        P3_U3199) );
  AOI21_X1 U9041 ( .B1(n12699), .B2(n12698), .A(n12697), .ZN(n6951) );
  AOI21_X1 U9042 ( .B1(n12966), .B2(n12893), .A(n7275), .ZN(n7274) );
  OR2_X1 U9043 ( .A1(n12393), .A2(n6839), .ZN(n7275) );
  INV_X1 U9044 ( .A(n13206), .ZN(n6930) );
  NAND2_X1 U9045 ( .A1(n7423), .A2(n13343), .ZN(n7422) );
  NAND2_X1 U9046 ( .A1(n13261), .A2(n10327), .ZN(n10489) );
  OAI21_X1 U9047 ( .B1(n13446), .B2(n6838), .A(n7314), .ZN(P2_U3528) );
  OAI21_X1 U9048 ( .B1(n13693), .B2(n7316), .A(n7315), .ZN(n7314) );
  NAND2_X1 U9049 ( .A1(n7322), .A2(n15127), .ZN(n7315) );
  NAND2_X1 U9050 ( .A1(n13503), .A2(n13766), .ZN(n6867) );
  NAND2_X1 U9051 ( .A1(n13503), .A2(n13814), .ZN(n6863) );
  INV_X1 U9052 ( .A(n6903), .ZN(n6902) );
  OAI21_X1 U9053 ( .B1(n14440), .B2(n14002), .A(n13849), .ZN(n6903) );
  NAND2_X1 U9054 ( .A1(n6888), .A2(n6885), .ZN(P1_U3262) );
  OR2_X1 U9055 ( .A1(n14073), .A2(n14071), .ZN(n6888) );
  AOI21_X1 U9056 ( .B1(n6887), .B2(n14071), .A(n6886), .ZN(n6885) );
  INV_X1 U9057 ( .A(n6890), .ZN(n14073) );
  NAND2_X1 U9058 ( .A1(n7119), .A2(n14319), .ZN(n14138) );
  NAND2_X1 U9059 ( .A1(n14861), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U9060 ( .A1(n7412), .A2(n7409), .ZN(P1_U3556) );
  AOI21_X1 U9061 ( .B1(n14435), .B2(n14345), .A(n7410), .ZN(n7409) );
  NAND2_X1 U9062 ( .A1(n14433), .A2(n14863), .ZN(n7412) );
  NOR2_X1 U9063 ( .A1(n14863), .A2(n7411), .ZN(n7410) );
  OAI21_X1 U9064 ( .B1(n14438), .B2(n14861), .A(n6855), .ZN(P1_U3555) );
  NOR2_X1 U9065 ( .A1(n6857), .A2(n6856), .ZN(n6855) );
  NOR2_X1 U9066 ( .A1(n14863), .A2(n14349), .ZN(n6856) );
  NOR2_X1 U9067 ( .A1(n14440), .A2(n14419), .ZN(n6857) );
  NAND2_X1 U9068 ( .A1(n6937), .A2(n6936), .ZN(n14434) );
  NAND2_X1 U9069 ( .A1(n9673), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6936) );
  INV_X1 U9070 ( .A(n6954), .ZN(n6953) );
  OAI22_X1 U9071 ( .A1(n14440), .A2(n14469), .B1(n14857), .B2(n14439), .ZN(
        n6954) );
  INV_X1 U9072 ( .A(n6925), .ZN(n14594) );
  NAND2_X1 U9073 ( .A1(n6971), .A2(n7245), .ZN(n6970) );
  XNOR2_X1 U9074 ( .A(n15785), .B(n15784), .ZN(n7243) );
  NOR2_X1 U9075 ( .A1(n13472), .A2(n7375), .ZN(n6691) );
  INV_X2 U9076 ( .A(n12177), .ZN(n12195) );
  AND2_X1 U9077 ( .A1(n6701), .A2(n14301), .ZN(n6692) );
  AND2_X1 U9078 ( .A1(n7124), .A2(n7122), .ZN(n6693) );
  AND2_X1 U9079 ( .A1(n12464), .A2(n12579), .ZN(n6694) );
  NAND2_X2 U9080 ( .A1(n9292), .A2(n9291), .ZN(n11384) );
  INV_X1 U9081 ( .A(n11384), .ZN(n7228) );
  XOR2_X1 U9082 ( .A(n12550), .B(n12833), .Z(n6695) );
  AND2_X1 U9083 ( .A1(n7372), .A2(n7373), .ZN(n6696) );
  OR3_X1 U9084 ( .A1(n12109), .A2(n12108), .A3(n12114), .ZN(n6697) );
  OAI21_X2 U9085 ( .B1(n6690), .B2(P2_IR_REG_0__SCAN_IN), .A(n9098), .ZN(n9926) );
  NOR2_X1 U9086 ( .A1(n8602), .A2(n8601), .ZN(n6698) );
  INV_X1 U9087 ( .A(n11121), .ZN(n7358) );
  OR3_X1 U9088 ( .A1(n13517), .A2(n13503), .A3(n6777), .ZN(n6699) );
  AND4_X1 U9089 ( .A1(n14144), .A2(n12222), .A3(n14157), .A4(n14177), .ZN(
        n6700) );
  NAND2_X1 U9090 ( .A1(n7266), .A2(n8612), .ZN(n8938) );
  OR2_X1 U9091 ( .A1(n10747), .A2(n7454), .ZN(n7453) );
  AND2_X1 U9092 ( .A1(n8337), .A2(n7129), .ZN(n6701) );
  AND2_X1 U9093 ( .A1(n13355), .A2(n13452), .ZN(n6702) );
  AND2_X1 U9094 ( .A1(n11963), .A2(n11962), .ZN(n6703) );
  INV_X1 U9095 ( .A(n13794), .ZN(n13471) );
  AND2_X1 U9096 ( .A1(n9461), .A2(n9460), .ZN(n13794) );
  AND2_X1 U9097 ( .A1(n13429), .A2(n7298), .ZN(n6704) );
  NAND2_X1 U9098 ( .A1(n11965), .A2(n9001), .ZN(n12762) );
  INV_X1 U9099 ( .A(n12762), .ZN(n6990) );
  AND2_X1 U9100 ( .A1(n13147), .A2(n13146), .ZN(n6705) );
  AND2_X1 U9101 ( .A1(n7550), .A2(n6749), .ZN(n6706) );
  AND2_X1 U9102 ( .A1(n6736), .A2(n7648), .ZN(n6707) );
  AND2_X1 U9103 ( .A1(n7019), .A2(n11921), .ZN(n6708) );
  AND2_X1 U9104 ( .A1(n7424), .A2(n6773), .ZN(n6709) );
  AND2_X1 U9105 ( .A1(n9565), .A2(n9564), .ZN(n13692) );
  AND2_X1 U9106 ( .A1(n13794), .A2(n13469), .ZN(n6710) );
  AND2_X1 U9107 ( .A1(n10386), .A2(n10387), .ZN(n6711) );
  AND2_X1 U9108 ( .A1(n8055), .A2(SI_13_), .ZN(n6712) );
  INV_X1 U9109 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7632) );
  AND2_X1 U9110 ( .A1(n8150), .A2(n8149), .ZN(n14464) );
  INV_X1 U9111 ( .A(n14464), .ZN(n14290) );
  AND2_X1 U9112 ( .A1(n9382), .A2(n9381), .ZN(n13656) );
  NAND2_X1 U9113 ( .A1(n7015), .A2(n8996), .ZN(n6713) );
  AND2_X1 U9114 ( .A1(n9618), .A2(n9621), .ZN(n6714) );
  NAND2_X1 U9115 ( .A1(n9618), .A2(n10460), .ZN(n6715) );
  AND2_X1 U9116 ( .A1(n7843), .A2(n15478), .ZN(n6716) );
  INV_X1 U9117 ( .A(n12579), .ZN(n12846) );
  NAND2_X1 U9118 ( .A1(n8063), .A2(n8062), .ZN(n13964) );
  INV_X1 U9119 ( .A(n13964), .ZN(n7122) );
  OR2_X1 U9120 ( .A1(n7123), .A2(n11213), .ZN(n6717) );
  AND2_X1 U9121 ( .A1(n11129), .A2(n7229), .ZN(n6718) );
  INV_X1 U9122 ( .A(n8238), .ZN(n7150) );
  AND2_X1 U9123 ( .A1(n8249), .A2(n15673), .ZN(n6719) );
  AND2_X1 U9124 ( .A1(n14124), .A2(n7392), .ZN(n6720) );
  INV_X2 U9125 ( .A(n11805), .ZN(n7941) );
  OR2_X1 U9126 ( .A1(n13612), .A2(n13461), .ZN(n7056) );
  NAND2_X1 U9127 ( .A1(n7630), .A2(n7760), .ZN(n8914) );
  INV_X1 U9128 ( .A(n12376), .ZN(n12329) );
  OR2_X1 U9129 ( .A1(n7251), .A2(n8836), .ZN(n6721) );
  AND2_X1 U9130 ( .A1(n14208), .A2(n8211), .ZN(n6722) );
  INV_X1 U9131 ( .A(n11399), .ZN(n6852) );
  INV_X1 U9132 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15514) );
  NAND2_X1 U9133 ( .A1(n11348), .A2(n11349), .ZN(n6723) );
  NAND2_X1 U9134 ( .A1(n8492), .A2(n6991), .ZN(n15329) );
  INV_X1 U9135 ( .A(n15329), .ZN(n15340) );
  OR2_X1 U9136 ( .A1(n9701), .A2(n6933), .ZN(n6725) );
  NAND2_X1 U9137 ( .A1(n9033), .A2(n9045), .ZN(n9042) );
  XNOR2_X1 U9138 ( .A(n9057), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9090) );
  OR2_X1 U9139 ( .A1(n8993), .A2(n11898), .ZN(n7611) );
  NAND2_X1 U9140 ( .A1(n7457), .A2(n7458), .ZN(n6726) );
  AND2_X1 U9141 ( .A1(n15131), .A2(n8620), .ZN(n6727) );
  INV_X1 U9142 ( .A(n9334), .ZN(n7517) );
  INV_X1 U9143 ( .A(n7396), .ZN(n7395) );
  NAND2_X1 U9144 ( .A1(n14247), .A2(n12133), .ZN(n7396) );
  INV_X1 U9145 ( .A(n12202), .ZN(n7182) );
  XNOR2_X1 U9146 ( .A(n9545), .B(n9544), .ZN(n13816) );
  OR2_X1 U9147 ( .A1(n12696), .A2(n15266), .ZN(n6728) );
  NAND2_X1 U9148 ( .A1(n11616), .A2(n11615), .ZN(n6729) );
  NAND2_X1 U9149 ( .A1(n13044), .A2(n12523), .ZN(n6730) );
  XNOR2_X1 U9150 ( .A(n11571), .B(n13360), .ZN(n11688) );
  AND2_X1 U9151 ( .A1(n8740), .A2(n6985), .ZN(n6731) );
  NAND2_X1 U9152 ( .A1(n11240), .A2(n11239), .ZN(n6732) );
  NAND2_X1 U9153 ( .A1(n14307), .A2(n8323), .ZN(n14277) );
  AND2_X1 U9154 ( .A1(n9365), .A2(n9364), .ZN(n13810) );
  NAND2_X1 U9155 ( .A1(n7117), .A2(n8327), .ZN(n14207) );
  AND2_X1 U9156 ( .A1(n9283), .A2(n7512), .ZN(n6733) );
  AND2_X1 U9157 ( .A1(n7033), .A2(n7027), .ZN(n6734) );
  NOR2_X1 U9158 ( .A1(n11384), .A2(n11381), .ZN(n6735) );
  OR2_X1 U9159 ( .A1(n7828), .A2(SI_17_), .ZN(n6736) );
  OR2_X1 U9160 ( .A1(n12668), .A2(n12630), .ZN(n6737) );
  AND4_X1 U9161 ( .A1(n9189), .A2(n9188), .A3(n9187), .A4(n9186), .ZN(n10814)
         );
  AND2_X1 U9162 ( .A1(n10156), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6738) );
  XNOR2_X1 U9163 ( .A(n12178), .B(n14105), .ZN(n12224) );
  INV_X1 U9164 ( .A(n12224), .ZN(n8287) );
  INV_X1 U9165 ( .A(n13579), .ZN(n7345) );
  AND2_X1 U9166 ( .A1(n10117), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6739) );
  AND2_X1 U9167 ( .A1(n12717), .A2(n12718), .ZN(n6740) );
  OR2_X1 U9168 ( .A1(n13027), .A2(n12752), .ZN(n6741) );
  AND3_X1 U9169 ( .A1(n15428), .A2(n7355), .A3(n7684), .ZN(n7913) );
  AND2_X1 U9170 ( .A1(n11872), .A2(n11867), .ZN(n11870) );
  INV_X1 U9171 ( .A(n12165), .ZN(n7683) );
  AND2_X1 U9172 ( .A1(n11984), .A2(n8651), .ZN(n6742) );
  OR2_X1 U9173 ( .A1(n7507), .A2(n6733), .ZN(n6743) );
  AND2_X2 U9174 ( .A1(n9090), .A2(n9058), .ZN(n9109) );
  AND2_X1 U9175 ( .A1(n6889), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U9176 ( .A1(n8333), .A2(n8273), .ZN(n14127) );
  NAND2_X1 U9177 ( .A1(n12197), .A2(n12196), .ZN(n6745) );
  NOR2_X1 U9178 ( .A1(n13916), .A2(n13915), .ZN(n6746) );
  INV_X1 U9179 ( .A(n14301), .ZN(n14409) );
  AND2_X1 U9180 ( .A1(n8136), .A2(n8135), .ZN(n14301) );
  OR2_X1 U9181 ( .A1(n9618), .A2(n7483), .ZN(n6747) );
  AND2_X1 U9182 ( .A1(n9612), .A2(n9611), .ZN(n6748) );
  OR2_X1 U9183 ( .A1(n6695), .A2(n6694), .ZN(n6749) );
  NOR2_X1 U9184 ( .A1(n13890), .A2(n13891), .ZN(n6750) );
  AND2_X1 U9185 ( .A1(n7905), .A2(n7920), .ZN(n6751) );
  INV_X1 U9186 ( .A(n13452), .ZN(n13813) );
  AND2_X1 U9187 ( .A1(n9355), .A2(n9354), .ZN(n13452) );
  INV_X1 U9188 ( .A(n7132), .ZN(n14184) );
  NOR2_X1 U9189 ( .A1(n14196), .A2(n14185), .ZN(n7132) );
  AND2_X1 U9190 ( .A1(n7321), .A2(n7323), .ZN(n6752) );
  AND2_X1 U9191 ( .A1(n13656), .A2(n13457), .ZN(n6753) );
  AND2_X1 U9192 ( .A1(n12339), .A2(n12338), .ZN(n13865) );
  INV_X1 U9193 ( .A(n13865), .ZN(n7731) );
  AND2_X1 U9194 ( .A1(n8351), .A2(n8350), .ZN(n6754) );
  INV_X1 U9195 ( .A(n14192), .ZN(n14194) );
  AND2_X1 U9196 ( .A1(n10991), .A2(n10989), .ZN(n6755) );
  AND2_X1 U9197 ( .A1(n14127), .A2(n8260), .ZN(n6756) );
  AND2_X1 U9198 ( .A1(n11966), .A2(n12758), .ZN(n12776) );
  INV_X1 U9199 ( .A(n9361), .ZN(n7495) );
  AND2_X1 U9200 ( .A1(n11385), .A2(n7230), .ZN(n6757) );
  AND3_X1 U9201 ( .A1(n11868), .A2(n11874), .A3(n11867), .ZN(n6758) );
  INV_X1 U9202 ( .A(n11992), .ZN(n12830) );
  XNOR2_X1 U9203 ( .A(n12987), .B(n12579), .ZN(n11992) );
  AND2_X1 U9204 ( .A1(n14464), .A2(n14023), .ZN(n6759) );
  INV_X1 U9205 ( .A(n7042), .ZN(n7041) );
  NOR2_X1 U9206 ( .A1(n10798), .A2(n10812), .ZN(n7042) );
  AND2_X1 U9207 ( .A1(n12092), .A2(n7676), .ZN(n6760) );
  INV_X1 U9208 ( .A(n13272), .ZN(n7446) );
  INV_X1 U9209 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8402) );
  INV_X1 U9210 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U9211 ( .A1(n9502), .A2(n7501), .ZN(n6761) );
  INV_X1 U9212 ( .A(n11921), .ZN(n7017) );
  AND2_X1 U9213 ( .A1(n7371), .A2(n7370), .ZN(n6762) );
  NOR2_X1 U9214 ( .A1(n12052), .A2(n14036), .ZN(n6763) );
  NOR2_X1 U9215 ( .A1(n13788), .A2(n13475), .ZN(n6764) );
  NOR2_X1 U9216 ( .A1(n14240), .A2(n14386), .ZN(n6765) );
  NOR2_X1 U9217 ( .A1(n12246), .A2(n12244), .ZN(n6766) );
  NOR2_X1 U9218 ( .A1(n11120), .A2(n11115), .ZN(n6767) );
  NOR2_X1 U9219 ( .A1(n12073), .A2(n11765), .ZN(n6768) );
  OR2_X1 U9220 ( .A1(n12092), .A2(n7676), .ZN(n6769) );
  INV_X1 U9221 ( .A(n7466), .ZN(n7465) );
  NAND2_X1 U9222 ( .A1(n7469), .A2(n7470), .ZN(n7466) );
  AND2_X1 U9223 ( .A1(n6897), .A2(n14269), .ZN(n6770) );
  OR2_X1 U9224 ( .A1(n8055), .A2(SI_13_), .ZN(n6771) );
  OR2_X1 U9225 ( .A1(n8161), .A2(n7753), .ZN(n6772) );
  NAND2_X1 U9226 ( .A1(n13200), .A2(n7429), .ZN(n6773) );
  AND2_X1 U9227 ( .A1(n11120), .A2(n13366), .ZN(n6774) );
  AND2_X1 U9228 ( .A1(n11949), .A2(n12987), .ZN(n6775) );
  AND2_X1 U9229 ( .A1(n12431), .A2(n12505), .ZN(n6776) );
  INV_X1 U9230 ( .A(n13810), .ZN(n13672) );
  NAND2_X1 U9231 ( .A1(n13692), .A2(n13775), .ZN(n6777) );
  AND2_X1 U9232 ( .A1(n7583), .A2(n7581), .ZN(n6778) );
  NAND3_X1 U9233 ( .A1(n8612), .A2(n7760), .A3(n7631), .ZN(n6779) );
  AND2_X1 U9234 ( .A1(n7606), .A2(n12934), .ZN(n6780) );
  AND2_X1 U9235 ( .A1(n14173), .A2(n8237), .ZN(n6781) );
  AND2_X1 U9236 ( .A1(n14211), .A2(n12321), .ZN(n6782) );
  AND2_X1 U9237 ( .A1(n10782), .A2(n6889), .ZN(n6783) );
  INV_X1 U9238 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8975) );
  AND2_X1 U9239 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9810), .ZN(n6784) );
  INV_X1 U9240 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8297) );
  INV_X1 U9241 ( .A(n7258), .ZN(n7257) );
  NAND2_X1 U9242 ( .A1(n8895), .A2(n6730), .ZN(n7258) );
  AND2_X1 U9243 ( .A1(n7169), .A2(n7168), .ZN(n6785) );
  NAND2_X1 U9244 ( .A1(n12125), .A2(n12124), .ZN(n6786) );
  INV_X1 U9245 ( .A(n7619), .ZN(n7618) );
  NAND2_X1 U9246 ( .A1(n11941), .A2(n7620), .ZN(n7619) );
  INV_X1 U9247 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9848) );
  INV_X1 U9248 ( .A(n11564), .ZN(n7333) );
  OAI21_X1 U9249 ( .B1(n7017), .B2(n7020), .A(n12907), .ZN(n7016) );
  NAND2_X1 U9250 ( .A1(n7056), .A2(n7054), .ZN(n7057) );
  NAND2_X1 U9251 ( .A1(n12794), .A2(n11958), .ZN(n6787) );
  AND2_X1 U9252 ( .A1(n9642), .A2(n7483), .ZN(n6788) );
  INV_X1 U9253 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15475) );
  OR2_X1 U9254 ( .A1(n9231), .A2(n9230), .ZN(n6789) );
  INV_X1 U9255 ( .A(n12076), .ZN(n7189) );
  INV_X1 U9256 ( .A(n12136), .ZN(n7168) );
  NAND2_X1 U9257 ( .A1(n11924), .A2(n11929), .ZN(n12898) );
  OR2_X1 U9258 ( .A1(n7493), .A2(n9229), .ZN(n6790) );
  INV_X1 U9259 ( .A(n9176), .ZN(n7487) );
  OR2_X1 U9260 ( .A1(n12226), .A2(n12225), .ZN(n6791) );
  OR2_X1 U9261 ( .A1(n14573), .A2(n14574), .ZN(n6792) );
  OR2_X1 U9262 ( .A1(n8204), .A2(n10095), .ZN(n6793) );
  NOR2_X1 U9263 ( .A1(n15283), .A2(n8602), .ZN(n6794) );
  NOR2_X1 U9264 ( .A1(n12073), .A2(n14032), .ZN(n6795) );
  OR2_X1 U9265 ( .A1(n12965), .A2(n12767), .ZN(n11968) );
  INV_X1 U9266 ( .A(n11968), .ZN(n7629) );
  NOR2_X1 U9267 ( .A1(n7189), .A2(n7191), .ZN(n6796) );
  AND2_X1 U9268 ( .A1(n8084), .A2(n8070), .ZN(n6797) );
  AND2_X1 U9269 ( .A1(n7659), .A2(n7657), .ZN(n6798) );
  AND2_X1 U9270 ( .A1(n9308), .A2(n9307), .ZN(n14668) );
  INV_X1 U9271 ( .A(n14668), .ZN(n7230) );
  AND2_X1 U9272 ( .A1(n14259), .A2(n12133), .ZN(n6799) );
  AND2_X1 U9273 ( .A1(n12094), .A2(n6769), .ZN(n6800) );
  INV_X1 U9274 ( .A(n11579), .ZN(n7544) );
  AND2_X1 U9275 ( .A1(n10539), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6801) );
  AND2_X1 U9276 ( .A1(n8532), .A2(n8520), .ZN(n6802) );
  OR2_X1 U9277 ( .A1(n12083), .A2(n12081), .ZN(n6803) );
  OR2_X1 U9278 ( .A1(n12147), .A2(n12145), .ZN(n6804) );
  AND2_X1 U9279 ( .A1(n11566), .A2(n11561), .ZN(n6805) );
  AND2_X1 U9280 ( .A1(n8404), .A2(n8481), .ZN(n6807) );
  AND2_X1 U9281 ( .A1(n8479), .A2(n8407), .ZN(n6808) );
  OR2_X1 U9282 ( .A1(n7518), .A2(n7517), .ZN(n6809) );
  OR2_X1 U9283 ( .A1(n15089), .A2(n7290), .ZN(n6810) );
  NAND2_X1 U9284 ( .A1(n13788), .A2(n13440), .ZN(n6811) );
  INV_X1 U9285 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U9286 ( .A1(n11384), .A2(n13363), .ZN(n6812) );
  INV_X1 U9287 ( .A(n15180), .ZN(n7217) );
  INV_X1 U9288 ( .A(n9428), .ZN(n9586) );
  NAND2_X1 U9289 ( .A1(n13850), .A2(n12269), .ZN(n13914) );
  NAND2_X1 U9290 ( .A1(n12909), .A2(n8781), .ZN(n12882) );
  INV_X1 U9291 ( .A(n13718), .ZN(n7235) );
  NAND2_X1 U9292 ( .A1(n11768), .A2(n7769), .ZN(n11790) );
  INV_X1 U9293 ( .A(n14167), .ZN(n7131) );
  AND2_X1 U9294 ( .A1(n13154), .A2(n13153), .ZN(n6813) );
  AND3_X1 U9295 ( .A1(n11568), .A2(n6702), .A3(n13810), .ZN(n6814) );
  INV_X1 U9296 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7684) );
  NOR3_X1 U9297 ( .A1(n13614), .A2(n13613), .A3(n13651), .ZN(n6815) );
  NAND2_X1 U9298 ( .A1(n12529), .A2(n12937), .ZN(n6816) );
  INV_X1 U9299 ( .A(n9504), .ZN(n7502) );
  AND2_X1 U9300 ( .A1(n12465), .A2(n12846), .ZN(n6817) );
  NOR2_X1 U9301 ( .A1(n9037), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n9335) );
  INV_X1 U9302 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7663) );
  NAND2_X1 U9303 ( .A1(n7096), .A2(n12096), .ZN(n11505) );
  NAND2_X1 U9304 ( .A1(n7101), .A2(n8316), .ZN(n11419) );
  INV_X1 U9305 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7387) );
  INV_X1 U9306 ( .A(n13627), .ZN(n7300) );
  AND2_X1 U9307 ( .A1(n14754), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U9308 ( .A1(n9480), .A2(n9479), .ZN(n13707) );
  INV_X1 U9309 ( .A(n13707), .ZN(n7233) );
  INV_X1 U9310 ( .A(n11890), .ZN(n7634) );
  NAND2_X1 U9311 ( .A1(n11937), .A2(n11938), .ZN(n12877) );
  AND2_X1 U9312 ( .A1(n10437), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6819) );
  AND2_X1 U9313 ( .A1(n7443), .A2(n13271), .ZN(n6820) );
  AND2_X1 U9314 ( .A1(n8445), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6821) );
  INV_X1 U9315 ( .A(n12464), .ZN(n12465) );
  NAND2_X1 U9316 ( .A1(n11464), .A2(n6692), .ZN(n7130) );
  INV_X1 U9317 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7242) );
  NOR2_X1 U9318 ( .A1(n15247), .A2(n15246), .ZN(n6822) );
  AND2_X1 U9319 ( .A1(n11565), .A2(n11564), .ZN(n6823) );
  AND2_X1 U9320 ( .A1(n12424), .A2(n12423), .ZN(n6824) );
  AND2_X1 U9321 ( .A1(n7828), .A2(SI_17_), .ZN(n6825) );
  INV_X1 U9322 ( .A(n7183), .ZN(n7178) );
  INV_X1 U9323 ( .A(n12200), .ZN(n7183) );
  AND2_X1 U9324 ( .A1(n11176), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6826) );
  AND2_X1 U9325 ( .A1(n9144), .A2(n9015), .ZN(n6827) );
  OR2_X1 U9326 ( .A1(n11865), .A2(n11967), .ZN(n6828) );
  AND2_X1 U9327 ( .A1(n13459), .A2(n13458), .ZN(n13628) );
  INV_X1 U9328 ( .A(n13628), .ZN(n7084) );
  AND2_X1 U9329 ( .A1(n12570), .A2(n12562), .ZN(n11904) );
  INV_X1 U9330 ( .A(n11904), .ZN(n7613) );
  AND2_X1 U9331 ( .A1(n8071), .A2(n8070), .ZN(n6829) );
  INV_X1 U9332 ( .A(n15129), .ZN(n15127) );
  INV_X1 U9333 ( .A(n13339), .ZN(n13343) );
  INV_X1 U9334 ( .A(n12073), .ZN(n7126) );
  OR2_X1 U9335 ( .A1(n8249), .A2(n15673), .ZN(n6830) );
  INV_X1 U9336 ( .A(n14413), .ZN(n7129) );
  AND2_X1 U9337 ( .A1(n7121), .A2(n7124), .ZN(n6831) );
  INV_X1 U9338 ( .A(n9442), .ZN(n7642) );
  NAND2_X1 U9339 ( .A1(n10844), .A2(n10804), .ZN(n11114) );
  INV_X1 U9340 ( .A(n6853), .ZN(n11400) );
  INV_X1 U9341 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7754) );
  INV_X1 U9342 ( .A(n7852), .ZN(n7148) );
  INV_X1 U9343 ( .A(n13300), .ZN(n7440) );
  AND2_X1 U9344 ( .A1(n11142), .A2(n11141), .ZN(n6832) );
  AND2_X1 U9345 ( .A1(n10677), .A2(n9002), .ZN(n6833) );
  OR2_X1 U9346 ( .A1(n11032), .A2(n12070), .ZN(n11213) );
  INV_X1 U9347 ( .A(n11213), .ZN(n7121) );
  INV_X1 U9348 ( .A(n7527), .ZN(n7525) );
  NOR2_X1 U9349 ( .A1(n12537), .A2(n7528), .ZN(n7527) );
  INV_X1 U9350 ( .A(n7671), .ZN(n7670) );
  NOR2_X1 U9351 ( .A1(n8278), .A2(n6836), .ZN(n7671) );
  AND2_X1 U9352 ( .A1(n7635), .A2(n11890), .ZN(n6834) );
  AND2_X1 U9353 ( .A1(n7740), .A2(n7739), .ZN(n6835) );
  AND2_X1 U9354 ( .A1(n7854), .A2(SI_27_), .ZN(n6836) );
  INV_X1 U9355 ( .A(n7611), .ZN(n7610) );
  AND2_X1 U9356 ( .A1(n11829), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U9357 ( .A1(n15129), .A2(n7325), .ZN(n6838) );
  NOR2_X1 U9358 ( .A1(n15335), .A2(n12392), .ZN(n6839) );
  NAND3_X1 U9359 ( .A1(n7630), .A2(n7760), .A3(n7632), .ZN(n6840) );
  AND2_X1 U9360 ( .A1(n7723), .A2(n6729), .ZN(n6841) );
  XNOR2_X1 U9361 ( .A(n8480), .B(n8479), .ZN(n8926) );
  INV_X1 U9362 ( .A(n14863), .ZN(n14861) );
  INV_X1 U9363 ( .A(n15146), .ZN(n15134) );
  INV_X1 U9364 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7602) );
  INV_X1 U9365 ( .A(n13331), .ZN(n13448) );
  AND2_X1 U9366 ( .A1(n9958), .A2(n9873), .ZN(n13331) );
  INV_X1 U9367 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6854) );
  NAND2_X2 U9368 ( .A1(n11855), .A2(n12004), .ZN(n11967) );
  NAND2_X1 U9369 ( .A1(n12017), .A2(n11001), .ZN(n10621) );
  INV_X1 U9370 ( .A(n10621), .ZN(n7128) );
  AND2_X1 U9371 ( .A1(n12720), .A2(n12743), .ZN(n6842) );
  AND2_X1 U9372 ( .A1(n12746), .A2(n7215), .ZN(n6843) );
  INV_X1 U9373 ( .A(n12742), .ZN(n7624) );
  INV_X1 U9374 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6979) );
  OR2_X1 U9375 ( .A1(n15162), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n6844) );
  INV_X1 U9376 ( .A(n11267), .ZN(n7408) );
  INV_X1 U9377 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7239) );
  INV_X1 U9378 ( .A(n13622), .ZN(n7325) );
  AND2_X1 U9379 ( .A1(n10259), .A2(n9909), .ZN(n12237) );
  NAND2_X1 U9380 ( .A1(n8361), .A2(n8383), .ZN(n9904) );
  XNOR2_X1 U9381 ( .A(n11240), .B(n6847), .ZN(n6848) );
  XNOR2_X1 U9382 ( .A(n10787), .B(n12376), .ZN(n11240) );
  NAND2_X2 U9383 ( .A1(n13903), .A2(n12357), .ZN(n13989) );
  NAND2_X1 U9384 ( .A1(n7726), .A2(n7724), .ZN(n13938) );
  OR2_X2 U9385 ( .A1(n11258), .A2(n11246), .ZN(n6853) );
  NOR2_X1 U9386 ( .A1(n11259), .A2(n11260), .ZN(n11258) );
  AND3_X2 U9387 ( .A1(n7164), .A2(n7975), .A3(n6854), .ZN(n6944) );
  NAND2_X1 U9388 ( .A1(n13872), .A2(n12302), .ZN(n13876) );
  NAND2_X1 U9389 ( .A1(n13980), .A2(n13981), .ZN(n13872) );
  INV_X1 U9390 ( .A(n11247), .ZN(n10381) );
  NAND2_X1 U9391 ( .A1(n8144), .A2(n8321), .ZN(n14276) );
  OAI21_X1 U9392 ( .B1(n8133), .B2(n7705), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6956) );
  INV_X1 U9393 ( .A(n7957), .ZN(n7692) );
  NAND2_X1 U9394 ( .A1(n11417), .A2(n8054), .ZN(n11457) );
  NOR2_X1 U9395 ( .A1(n7119), .A2(n14347), .ZN(n6859) );
  NAND2_X1 U9396 ( .A1(n7710), .A2(n7711), .ZN(n14210) );
  NAND2_X1 U9397 ( .A1(n7695), .A2(n7694), .ZN(n11191) );
  NAND2_X1 U9398 ( .A1(n14433), .A2(n14857), .ZN(n6937) );
  NOR2_X1 U9399 ( .A1(n14108), .A2(n14107), .ZN(n14110) );
  NAND2_X1 U9400 ( .A1(n6861), .A2(n6860), .ZN(P1_U3557) );
  NAND2_X1 U9401 ( .A1(n9672), .A2(n14863), .ZN(n6861) );
  NAND2_X1 U9402 ( .A1(n14087), .A2(n14855), .ZN(n6862) );
  NAND2_X1 U9403 ( .A1(n13779), .A2(n6863), .ZN(P2_U3495) );
  INV_X1 U9404 ( .A(n6866), .ZN(n7328) );
  OAI21_X1 U9405 ( .B1(n6866), .B2(n13439), .A(n6811), .ZN(n6865) );
  NAND2_X1 U9406 ( .A1(n13699), .A2(n6867), .ZN(P2_U3527) );
  NAND2_X1 U9407 ( .A1(n7780), .A2(n6868), .ZN(n7778) );
  NAND2_X1 U9408 ( .A1(n7070), .A2(n11342), .ZN(n9642) );
  NAND2_X1 U9409 ( .A1(n7059), .A2(n7784), .ZN(n7089) );
  NAND2_X1 U9410 ( .A1(n7783), .A2(n7782), .ZN(n7059) );
  NAND2_X1 U9411 ( .A1(n11189), .A2(n8037), .ZN(n11418) );
  NAND2_X1 U9412 ( .A1(n11191), .A2(n11190), .ZN(n11189) );
  NAND2_X1 U9413 ( .A1(n7698), .A2(n8012), .ZN(n7697) );
  NAND2_X1 U9414 ( .A1(n14576), .A2(n14998), .ZN(n6916) );
  NOR2_X1 U9415 ( .A1(n14723), .A2(n14724), .ZN(n14722) );
  NOR2_X1 U9416 ( .A1(n14711), .A2(n14712), .ZN(n14710) );
  INV_X1 U9417 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6869) );
  INV_X1 U9418 ( .A(n14610), .ZN(n6919) );
  NAND2_X1 U9419 ( .A1(n14499), .A2(n6927), .ZN(n14533) );
  NAND4_X1 U9420 ( .A1(n7892), .A2(n7687), .A3(n7685), .A4(n7686), .ZN(n6872)
         );
  NAND2_X1 U9421 ( .A1(n12291), .A2(n13928), .ZN(n13931) );
  NAND2_X1 U9422 ( .A1(n11090), .A2(n7987), .ZN(n10871) );
  INV_X1 U9423 ( .A(n7885), .ZN(n11814) );
  NAND2_X1 U9424 ( .A1(n13262), .A2(n13263), .ZN(n13261) );
  NAND2_X1 U9425 ( .A1(n6929), .A2(n7438), .ZN(n13171) );
  NAND2_X1 U9426 ( .A1(n10915), .A2(n10916), .ZN(n10939) );
  NAND2_X1 U9427 ( .A1(n13302), .A2(n6901), .ZN(n6900) );
  OAI21_X1 U9428 ( .B1(n7455), .B2(n7452), .A(n7450), .ZN(n10914) );
  NAND2_X1 U9429 ( .A1(n7787), .A2(n7940), .ZN(n6874) );
  NAND2_X1 U9430 ( .A1(n9841), .A2(n11804), .ZN(n7120) );
  AOI21_X2 U9431 ( .B1(n9837), .B2(n11804), .A(n6875), .ZN(n12068) );
  INV_X1 U9432 ( .A(n12212), .ZN(n7698) );
  NOR2_X1 U9433 ( .A1(n9773), .A2(n9808), .ZN(n7903) );
  INV_X2 U9434 ( .A(n7845), .ZN(n9766) );
  OAI21_X1 U9435 ( .B1(n12322), .B2(n10261), .A(n10260), .ZN(n10373) );
  NOR2_X1 U9436 ( .A1(n10526), .A2(n6801), .ZN(n9700) );
  AOI21_X2 U9437 ( .B1(n10598), .B2(n10527), .A(n10528), .ZN(n10526) );
  OAI21_X2 U9438 ( .B1(n11618), .B2(n7721), .A(n7719), .ZN(n11761) );
  OAI21_X1 U9439 ( .B1(n14634), .B2(n7607), .A(n6780), .ZN(n8994) );
  NAND2_X1 U9440 ( .A1(n11010), .A2(n11865), .ZN(n11149) );
  NAND2_X1 U9441 ( .A1(n12920), .A2(n11920), .ZN(n12908) );
  NAND2_X1 U9442 ( .A1(n11732), .A2(n11895), .ZN(n11722) );
  NAND2_X1 U9443 ( .A1(n8981), .A2(n11872), .ZN(n15282) );
  NAND2_X1 U9444 ( .A1(n6879), .A2(n11960), .ZN(n12777) );
  OAI21_X2 U9445 ( .B1(n12878), .B2(n7619), .A(n7615), .ZN(n12843) );
  OAI21_X1 U9446 ( .B1(n11850), .B2(n11851), .A(n12002), .ZN(n6922) );
  NAND2_X1 U9447 ( .A1(n12793), .A2(n11961), .ZN(n6879) );
  NAND2_X1 U9448 ( .A1(n8941), .A2(n8404), .ZN(n8946) );
  INV_X1 U9449 ( .A(n6922), .ZN(n7598) );
  NAND2_X2 U9450 ( .A1(n6880), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7227) );
  NAND3_X1 U9451 ( .A1(n14075), .A2(n13405), .A3(n7771), .ZN(n6880) );
  NAND2_X1 U9452 ( .A1(n7641), .A2(n7842), .ZN(n8214) );
  NAND2_X1 U9453 ( .A1(n14156), .A2(n14157), .ZN(n14155) );
  NAND2_X1 U9454 ( .A1(n7112), .A2(n7111), .ZN(n14193) );
  NOR2_X2 U9455 ( .A1(n9684), .A2(n10570), .ZN(n9685) );
  NOR2_X1 U9456 ( .A1(n10561), .A2(n9734), .ZN(n10560) );
  INV_X1 U9457 ( .A(n9688), .ZN(n7294) );
  NOR2_X2 U9458 ( .A1(n15172), .A2(n11058), .ZN(n15171) );
  OAI21_X2 U9459 ( .B1(n15223), .B2(n7308), .A(n7307), .ZN(n12671) );
  NOR2_X2 U9460 ( .A1(n15224), .A2(n8694), .ZN(n15223) );
  OAI21_X1 U9461 ( .B1(n11843), .B2(n7629), .A(n7628), .ZN(n7627) );
  NOR2_X2 U9462 ( .A1(n9037), .A2(n7416), .ZN(n9055) );
  NAND3_X2 U9463 ( .A1(n7480), .A2(n7479), .A3(n9015), .ZN(n9037) );
  NAND2_X1 U9464 ( .A1(n9118), .A2(n9119), .ZN(n9117) );
  OAI21_X2 U9465 ( .B1(n9320), .B2(n7515), .A(n7516), .ZN(n9347) );
  AOI22_X1 U9466 ( .A1(n9423), .A2(n9422), .B1(n9421), .B2(n9420), .ZN(n9438)
         );
  NAND2_X1 U9467 ( .A1(n9123), .A2(n9122), .ZN(n7477) );
  NAND2_X1 U9468 ( .A1(n9177), .A2(n6941), .ZN(n9190) );
  OAI22_X2 U9469 ( .A1(n6881), .A2(n9349), .B1(n9362), .B2(n9361), .ZN(n9377)
         );
  NAND2_X1 U9470 ( .A1(n6942), .A2(n9176), .ZN(n6941) );
  NAND2_X1 U9471 ( .A1(n9613), .A2(n6748), .ZN(n9619) );
  INV_X1 U9472 ( .A(n7284), .ZN(n7046) );
  NAND2_X1 U9473 ( .A1(n7046), .A2(n6690), .ZN(n7045) );
  NOR2_X1 U9474 ( .A1(n9348), .A2(n7494), .ZN(n6882) );
  AOI21_X1 U9475 ( .B1(n6948), .B2(n7166), .A(n6785), .ZN(n12139) );
  NAND2_X2 U9476 ( .A1(n7090), .A2(n7802), .ZN(n8002) );
  MUX2_X1 U9477 ( .A(n14025), .B(n14413), .S(n12177), .Z(n12120) );
  NAND2_X1 U9478 ( .A1(n7186), .A2(n12179), .ZN(n7185) );
  AOI21_X1 U9479 ( .B1(n7206), .B2(n12186), .A(n12185), .ZN(n12187) );
  NAND2_X1 U9480 ( .A1(n7089), .A2(n7786), .ZN(n7940) );
  INV_X1 U9481 ( .A(n6882), .ZN(n6881) );
  NAND2_X1 U9482 ( .A1(n7088), .A2(n7796), .ZN(n7972) );
  OAI21_X1 U9483 ( .B1(n9319), .B2(n9318), .A(n6809), .ZN(n7515) );
  NAND2_X2 U9484 ( .A1(n7872), .A2(n14481), .ZN(n8217) );
  OAI211_X1 U9485 ( .C1(n9619), .C2(n7481), .A(n6883), .B(n11395), .ZN(n9669)
         );
  NAND2_X1 U9486 ( .A1(n9619), .A2(n6960), .ZN(n6883) );
  AOI22_X1 U9487 ( .A1(n7507), .A2(n7510), .B1(n6733), .B2(n7513), .ZN(n7506)
         );
  XNOR2_X1 U9488 ( .A(n12080), .B(n14031), .ZN(n12215) );
  NAND2_X1 U9489 ( .A1(n11418), .A2(n12214), .ZN(n11417) );
  XNOR2_X2 U9490 ( .A(n12073), .B(n11765), .ZN(n12213) );
  NAND2_X2 U9491 ( .A1(n7120), .A2(n8017), .ZN(n12073) );
  NAND2_X1 U9492 ( .A1(n12229), .A2(n6798), .ZN(n7656) );
  NAND2_X1 U9493 ( .A1(n6791), .A2(n12233), .ZN(n7204) );
  NOR2_X1 U9494 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  NOR2_X1 U9495 ( .A1(n10121), .A2(n10120), .ZN(n10436) );
  NOR2_X1 U9496 ( .A1(n10248), .A2(n10247), .ZN(n10246) );
  NAND2_X1 U9497 ( .A1(n11169), .A2(n11170), .ZN(n14045) );
  NOR2_X1 U9498 ( .A1(n10140), .A2(n10139), .ZN(n10138) );
  NOR2_X1 U9499 ( .A1(n10729), .A2(n10728), .ZN(n11168) );
  NOR2_X1 U9500 ( .A1(n14764), .A2(n14763), .ZN(n14762) );
  NAND2_X2 U9501 ( .A1(n7227), .A2(n7226), .ZN(n7863) );
  NOR2_X1 U9502 ( .A1(n10436), .A2(n6819), .ZN(n10439) );
  NAND2_X1 U9503 ( .A1(n14775), .A2(n14050), .ZN(n14792) );
  AOI21_X1 U9504 ( .B1(n7691), .B2(n7693), .A(n12208), .ZN(n7689) );
  NOR2_X1 U9505 ( .A1(n10129), .A2(n6739), .ZN(n10152) );
  NOR2_X1 U9506 ( .A1(n10726), .A2(n7353), .ZN(n10729) );
  NOR2_X1 U9507 ( .A1(n14749), .A2(n6818), .ZN(n14764) );
  NOR2_X1 U9508 ( .A1(n10150), .A2(n6738), .ZN(n10140) );
  NAND3_X1 U9509 ( .A1(n6893), .A2(n6892), .A3(n7199), .ZN(n7198) );
  NAND2_X1 U9510 ( .A1(n12153), .A2(n12152), .ZN(n6892) );
  NAND2_X1 U9511 ( .A1(n12149), .A2(n12148), .ZN(n6893) );
  NAND2_X1 U9512 ( .A1(n7185), .A2(n12180), .ZN(n7184) );
  NOR2_X2 U9513 ( .A1(n12686), .A2(n12685), .ZN(n12689) );
  NOR3_X2 U9514 ( .A1(n12689), .A2(n12688), .A3(n12687), .ZN(n12707) );
  NAND2_X1 U9515 ( .A1(n6894), .A2(n12239), .ZN(P1_U3242) );
  NAND2_X1 U9516 ( .A1(n6896), .A2(n6895), .ZN(n6894) );
  NAND2_X1 U9517 ( .A1(n7203), .A2(n7762), .ZN(n6896) );
  NAND2_X1 U9518 ( .A1(n7187), .A2(n7672), .ZN(n7186) );
  OR2_X1 U9519 ( .A1(n10393), .A2(n15161), .ZN(n10392) );
  NAND2_X1 U9520 ( .A1(n6908), .A2(n6907), .ZN(n12150) );
  NOR2_X2 U9521 ( .A1(n15254), .A2(n15255), .ZN(n15252) );
  AOI21_X2 U9522 ( .B1(n15178), .B2(n15174), .A(n15175), .ZN(n12643) );
  NOR2_X2 U9523 ( .A1(n10376), .A2(n10377), .ZN(n10385) );
  NAND2_X1 U9524 ( .A1(n10395), .A2(n7216), .ZN(n10694) );
  AND2_X1 U9525 ( .A1(n9700), .A2(n10570), .ZN(n6933) );
  NAND2_X1 U9526 ( .A1(n6904), .A2(n6902), .ZN(P1_U3214) );
  OR2_X1 U9527 ( .A1(n10790), .A2(n10789), .ZN(n7743) );
  NAND2_X1 U9528 ( .A1(n6958), .A2(n13991), .ZN(n6904) );
  NAND2_X1 U9529 ( .A1(n11457), .A2(n11456), .ZN(n8071) );
  OAI21_X1 U9530 ( .B1(n12008), .B2(n12007), .A(n6905), .ZN(P3_U3296) );
  OAI211_X1 U9531 ( .C1(n8515), .C2(n7570), .A(n7567), .B(n8525), .ZN(n8423)
         );
  NAND2_X1 U9532 ( .A1(n6734), .A2(n7025), .ZN(n7024) );
  NAND2_X1 U9533 ( .A1(n13341), .A2(n7441), .ZN(n7447) );
  NAND2_X1 U9534 ( .A1(n11972), .A2(n11973), .ZN(n7597) );
  INV_X1 U9535 ( .A(n11346), .ZN(n7469) );
  NAND2_X1 U9536 ( .A1(n7578), .A2(n7577), .ZN(n11970) );
  NAND2_X1 U9537 ( .A1(n7022), .A2(n7021), .ZN(n11963) );
  NAND3_X1 U9538 ( .A1(n10939), .A2(n7468), .A3(n7462), .ZN(n7461) );
  INV_X1 U9539 ( .A(n7063), .ZN(n7062) );
  NAND2_X1 U9540 ( .A1(n7649), .A2(n7138), .ZN(n7137) );
  AOI211_X2 U9541 ( .C1(n13697), .C2(n15099), .A(n13696), .B(n13695), .ZN(
        n13777) );
  OAI21_X1 U9542 ( .B1(n11326), .B2(n6735), .A(n7278), .ZN(n11538) );
  INV_X1 U9543 ( .A(n11122), .ZN(n6909) );
  INV_X1 U9544 ( .A(n7304), .ZN(n7303) );
  NAND3_X1 U9545 ( .A1(n12144), .A2(n12143), .A3(n6804), .ZN(n6908) );
  NAND2_X1 U9546 ( .A1(n7234), .A2(n7233), .ZN(n13529) );
  NAND2_X1 U9547 ( .A1(n12200), .A2(n10520), .ZN(n10519) );
  OAI22_X1 U9548 ( .A1(n10788), .A2(n6683), .B1(n10381), .B2(n12034), .ZN(
        n10787) );
  OAI21_X2 U9549 ( .B1(n13555), .B2(n6866), .A(n7327), .ZN(n13526) );
  NAND2_X1 U9550 ( .A1(n8912), .A2(n8911), .ZN(n8916) );
  AOI21_X1 U9551 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14063), .A(n14800), .ZN(
        n14064) );
  AOI21_X1 U9552 ( .B1(n14795), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14786), .ZN(
        n14802) );
  NAND2_X1 U9553 ( .A1(n14533), .A2(n14534), .ZN(n14500) );
  INV_X1 U9554 ( .A(n14714), .ZN(n6917) );
  OAI21_X1 U9555 ( .B1(n7680), .B2(n12062), .A(n12061), .ZN(n7679) );
  NAND3_X1 U9556 ( .A1(n12078), .A2(n12079), .A3(n6803), .ZN(n6921) );
  MUX2_X2 U9557 ( .A(n12020), .B(n12019), .S(n12040), .Z(n12029) );
  INV_X1 U9558 ( .A(n12049), .ZN(n7173) );
  NAND2_X1 U9559 ( .A1(n7604), .A2(n7603), .ZN(n8849) );
  INV_X1 U9560 ( .A(n8467), .ZN(n7599) );
  NAND2_X1 U9561 ( .A1(n7190), .A2(n7188), .ZN(n12077) );
  NOR2_X2 U9562 ( .A1(n10385), .A2(n6711), .ZN(n10792) );
  INV_X2 U9563 ( .A(n6967), .ZN(n11001) );
  NAND2_X2 U9564 ( .A1(n8204), .A2(n9766), .ZN(n11805) );
  OAI21_X1 U9565 ( .B1(n14709), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6792), .ZN(
        n7237) );
  OAI21_X1 U9566 ( .B1(n15783), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n7245), .ZN(
        n7244) );
  XNOR2_X1 U9567 ( .A(n14537), .B(n6923), .ZN(n15798) );
  XNOR2_X1 U9568 ( .A(n14536), .B(n14535), .ZN(n14537) );
  INV_X1 U9569 ( .A(n6924), .ZN(n15795) );
  NOR2_X1 U9570 ( .A1(n13843), .A2(n12366), .ZN(n6969) );
  NAND2_X1 U9571 ( .A1(n7959), .A2(n7794), .ZN(n7088) );
  NAND2_X1 U9572 ( .A1(n6931), .A2(n6930), .ZN(P2_U3186) );
  NAND2_X1 U9573 ( .A1(n13225), .A2(n13207), .ZN(n6931) );
  NAND2_X1 U9574 ( .A1(n10373), .A2(n10375), .ZN(n10374) );
  INV_X1 U9575 ( .A(n7431), .ZN(n7430) );
  NOR2_X1 U9576 ( .A1(n14110), .A2(n6932), .ZN(n8288) );
  AOI21_X2 U9577 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9457) );
  OAI21_X1 U9578 ( .B1(n9417), .B2(n9416), .A(n9415), .ZN(n9419) );
  NOR2_X1 U9579 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  XNOR2_X1 U9580 ( .A(n12633), .B(n14626), .ZN(n14629) );
  NOR2_X2 U9581 ( .A1(n10581), .A2(n9703), .ZN(n9704) );
  NOR2_X1 U9582 ( .A1(n9733), .A2(n6725), .ZN(n10562) );
  NAND3_X1 U9583 ( .A1(n7321), .A2(n7058), .A3(n13694), .ZN(n13776) );
  NAND2_X1 U9584 ( .A1(n11598), .A2(n11597), .ZN(n7635) );
  NAND2_X1 U9585 ( .A1(n12816), .A2(n11952), .ZN(n12803) );
  NAND2_X2 U9586 ( .A1(n8992), .A2(n11899), .ZN(n14634) );
  NAND2_X1 U9587 ( .A1(n11460), .A2(n8085), .ZN(n11504) );
  NAND2_X1 U9588 ( .A1(n14122), .A2(n8274), .ZN(n14108) );
  NAND2_X1 U9589 ( .A1(n10263), .A2(n6938), .ZN(n10375) );
  NAND2_X1 U9590 ( .A1(n7477), .A2(n7478), .ZN(n7476) );
  NAND2_X1 U9591 ( .A1(n7737), .A2(n6732), .ZN(n7736) );
  NAND2_X1 U9592 ( .A1(n7492), .A2(n6790), .ZN(n9243) );
  AOI22_X1 U9593 ( .A1(n9157), .A2(n9156), .B1(n9155), .B2(n9154), .ZN(n9173)
         );
  NAND2_X1 U9594 ( .A1(n7484), .A2(n6715), .ZN(n7069) );
  XNOR2_X1 U9595 ( .A(n7071), .B(n9094), .ZN(n7070) );
  INV_X1 U9596 ( .A(n9641), .ZN(n7074) );
  NOR2_X1 U9597 ( .A1(n6714), .A2(n6961), .ZN(n6960) );
  NAND2_X1 U9598 ( .A1(n9540), .A2(n9539), .ZN(n9552) );
  INV_X1 U9599 ( .A(n6944), .ZN(n8161) );
  INV_X1 U9600 ( .A(n7752), .ZN(n7751) );
  NAND2_X1 U9601 ( .A1(n13876), .A2(n12307), .ZN(n13949) );
  NAND2_X1 U9602 ( .A1(n6945), .A2(n7682), .ZN(n12168) );
  NAND3_X1 U9603 ( .A1(n12163), .A2(n12162), .A3(n6806), .ZN(n6945) );
  NAND2_X1 U9604 ( .A1(n15798), .A2(n15799), .ZN(n6946) );
  NAND2_X1 U9605 ( .A1(n15787), .A2(n15786), .ZN(n6947) );
  OAI21_X1 U9606 ( .B1(n7168), .B2(n7169), .A(n12134), .ZN(n7167) );
  NOR2_X1 U9607 ( .A1(n12187), .A2(n7205), .ZN(n12235) );
  NAND2_X1 U9608 ( .A1(n12131), .A2(n12130), .ZN(n6948) );
  NOR2_X1 U9609 ( .A1(n7206), .A2(n12186), .ZN(n7205) );
  NAND2_X1 U9610 ( .A1(n12139), .A2(n12140), .ZN(n12138) );
  NAND2_X1 U9611 ( .A1(n12086), .A2(n12087), .ZN(n12085) );
  NAND2_X1 U9612 ( .A1(n12058), .A2(n12057), .ZN(n7680) );
  AOI21_X1 U9613 ( .B1(n12235), .B2(n12234), .A(n7204), .ZN(n7203) );
  NAND3_X1 U9614 ( .A1(n7170), .A2(n6949), .A3(n12056), .ZN(n12054) );
  NAND2_X1 U9615 ( .A1(n13931), .A2(n12292), .ZN(n13980) );
  AOI21_X2 U9616 ( .B1(n7224), .B2(n7223), .A(n12652), .ZN(n12633) );
  AND2_X2 U9617 ( .A1(n12659), .A2(n12658), .ZN(n12661) );
  NAND2_X1 U9618 ( .A1(n10691), .A2(n10692), .ZN(n10690) );
  NOR2_X1 U9619 ( .A1(n10578), .A2(n10579), .ZN(n10577) );
  NAND2_X1 U9620 ( .A1(n6955), .A2(n6953), .ZN(P1_U3523) );
  OR2_X1 U9621 ( .A1(n14438), .A2(n9673), .ZN(n6955) );
  NOR2_X1 U9622 ( .A1(n15169), .A2(n11500), .ZN(n15168) );
  NAND2_X1 U9623 ( .A1(n7690), .A2(n7689), .ZN(n11090) );
  NAND2_X1 U9624 ( .A1(n7313), .A2(n7312), .ZN(n10561) );
  NOR2_X1 U9625 ( .A1(n12695), .A2(n12915), .ZN(n12701) );
  XNOR2_X1 U9626 ( .A(n12671), .B(n14626), .ZN(n14615) );
  NAND2_X1 U9627 ( .A1(n8514), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7310) );
  NOR2_X2 U9628 ( .A1(n7165), .A2(n6957), .ZN(n7164) );
  NAND4_X1 U9629 ( .A1(n15553), .A2(n15539), .A3(n8095), .A4(n15698), .ZN(
        n6957) );
  NAND2_X1 U9630 ( .A1(n6968), .A2(n13842), .ZN(n6958) );
  NAND2_X1 U9631 ( .A1(n13261), .A2(n7456), .ZN(n7455) );
  OR2_X1 U9632 ( .A1(n11538), .A2(n11537), .ZN(n11540) );
  NAND2_X1 U9633 ( .A1(n7417), .A2(n7418), .ZN(n7416) );
  NAND2_X1 U9634 ( .A1(n7302), .A2(n7301), .ZN(n11122) );
  INV_X1 U9635 ( .A(n13446), .ZN(n7319) );
  NAND2_X1 U9636 ( .A1(n14532), .A2(n7242), .ZN(n14505) );
  NAND2_X1 U9637 ( .A1(n14600), .A2(n14599), .ZN(n7238) );
  NAND2_X1 U9638 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8489) );
  NOR2_X2 U9639 ( .A1(n12716), .A2(n6740), .ZN(n12721) );
  OAI21_X1 U9640 ( .B1(n6784), .B2(n9783), .A(n7216), .ZN(n10394) );
  XNOR2_X1 U9641 ( .A(n14559), .B(n7241), .ZN(n14601) );
  OAI21_X2 U9642 ( .B1(n14539), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14503), .ZN(
        n14504) );
  NAND2_X1 U9643 ( .A1(n14222), .A2(n7113), .ZN(n7111) );
  AOI21_X2 U9644 ( .B1(n14103), .B2(n14688), .A(n6959), .ZN(n14343) );
  XNOR2_X2 U9645 ( .A(n14454), .B(n14224), .ZN(n14209) );
  NAND2_X1 U9646 ( .A1(n13988), .A2(n6969), .ZN(n6968) );
  AOI21_X1 U9647 ( .B1(n7511), .B2(n7509), .A(n7508), .ZN(n7507) );
  NAND2_X1 U9648 ( .A1(n14776), .A2(n11510), .ZN(n14775) );
  NOR2_X1 U9649 ( .A1(n14737), .A2(n6826), .ZN(n11169) );
  INV_X1 U9650 ( .A(n14049), .ZN(n14048) );
  NAND2_X1 U9651 ( .A1(n7461), .A2(n7460), .ZN(n11355) );
  OAI21_X1 U9652 ( .B1(n8014), .B2(n7654), .A(n7652), .ZN(n8039) );
  INV_X1 U9653 ( .A(n9685), .ZN(n7313) );
  NOR2_X2 U9654 ( .A1(n12704), .A2(n12703), .ZN(n12728) );
  NOR2_X2 U9655 ( .A1(n12701), .A2(n6965), .ZN(n12704) );
  XNOR2_X1 U9656 ( .A(n10384), .B(n10383), .ZN(n10377) );
  XNOR2_X1 U9657 ( .A(n14549), .B(n7239), .ZN(n14600) );
  NAND2_X1 U9658 ( .A1(n14601), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7240) );
  XNOR2_X1 U9659 ( .A(n6970), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  INV_X1 U9660 ( .A(n15783), .ZN(n6971) );
  NAND2_X1 U9661 ( .A1(n14570), .A2(n14707), .ZN(n6972) );
  INV_X1 U9662 ( .A(n14704), .ZN(n6973) );
  INV_X4 U9663 ( .A(n7790), .ZN(n7845) );
  INV_X1 U9664 ( .A(n7506), .ZN(n7505) );
  NAND2_X1 U9665 ( .A1(n10095), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6975) );
  XNOR2_X1 U9666 ( .A(n11761), .B(n11759), .ZN(n11749) );
  INV_X1 U9667 ( .A(n7262), .ZN(n6984) );
  NAND2_X1 U9668 ( .A1(n8995), .A2(n11923), .ZN(n12896) );
  XNOR2_X1 U9669 ( .A(n7625), .B(n7624), .ZN(n11850) );
  OAI211_X1 U9670 ( .C1(n11972), .C2(n10421), .A(n7598), .B(n7597), .ZN(n7596)
         );
  INV_X1 U9671 ( .A(n7596), .ZN(n12008) );
  AOI21_X1 U9672 ( .B1(n7696), .B2(n7699), .A(n6795), .ZN(n7694) );
  OAI21_X2 U9673 ( .B1(n14344), .B2(n14684), .A(n6976), .ZN(n14433) );
  INV_X1 U9674 ( .A(n7237), .ZN(n14712) );
  XNOR2_X1 U9675 ( .A(n7244), .B(n7243), .ZN(SUB_1596_U4) );
  NAND2_X1 U9676 ( .A1(n8071), .A2(n6797), .ZN(n11460) );
  NAND2_X1 U9677 ( .A1(n12721), .A2(n6980), .ZN(n7208) );
  INV_X1 U9678 ( .A(n9707), .ZN(n7220) );
  INV_X2 U9679 ( .A(n8217), .ZN(n7923) );
  NOR2_X2 U9680 ( .A1(n8133), .A2(n7706), .ZN(n7867) );
  NAND3_X1 U9681 ( .A1(n7004), .A2(n11880), .A3(n11881), .ZN(n7003) );
  NAND3_X1 U9682 ( .A1(n11917), .A2(n7013), .A3(n11967), .ZN(n7011) );
  NAND2_X1 U9683 ( .A1(n11916), .A2(n7013), .ZN(n7012) );
  NAND2_X1 U9684 ( .A1(n11948), .A2(n7023), .ZN(n7022) );
  NAND2_X2 U9685 ( .A1(n7034), .A2(n12731), .ZN(n7226) );
  NAND3_X1 U9686 ( .A1(n7035), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7034) );
  NAND2_X1 U9687 ( .A1(n10799), .A2(n7037), .ZN(n7036) );
  NAND3_X1 U9688 ( .A1(n7038), .A2(n10833), .A3(n7036), .ZN(n10827) );
  INV_X2 U9689 ( .A(n10197), .ZN(n9925) );
  XNOR2_X2 U9690 ( .A(n13374), .B(n10197), .ZN(n10182) );
  NAND2_X1 U9691 ( .A1(n11692), .A2(n7050), .ZN(n7049) );
  NAND3_X1 U9692 ( .A1(n11287), .A2(n6812), .A3(n11286), .ZN(n7052) );
  NAND2_X1 U9693 ( .A1(n7052), .A2(n11385), .ZN(n11545) );
  NAND2_X1 U9694 ( .A1(n7056), .A2(n7053), .ZN(n7372) );
  INV_X1 U9695 ( .A(n7057), .ZN(n13466) );
  XNOR2_X1 U9696 ( .A(n7059), .B(n7929), .ZN(n9767) );
  NAND2_X1 U9697 ( .A1(n7989), .A2(n7800), .ZN(n7090) );
  NAND2_X1 U9698 ( .A1(n7972), .A2(n7797), .ZN(n7060) );
  NAND2_X1 U9699 ( .A1(n7947), .A2(n7791), .ZN(n7061) );
  NAND2_X1 U9700 ( .A1(n7067), .A2(n7134), .ZN(n8057) );
  NAND2_X1 U9701 ( .A1(n7806), .A2(n7136), .ZN(n7067) );
  NAND3_X1 U9702 ( .A1(n9639), .A2(n7074), .A3(n7072), .ZN(n7071) );
  NAND2_X2 U9703 ( .A1(n8002), .A2(n7803), .ZN(n7806) );
  NAND2_X1 U9704 ( .A1(n7094), .A2(n7091), .ZN(n14314) );
  AND2_X1 U9705 ( .A1(n7097), .A2(n8319), .ZN(n7095) );
  NAND2_X1 U9706 ( .A1(n11185), .A2(n7102), .ZN(n7099) );
  NAND2_X1 U9707 ( .A1(n7099), .A2(n7100), .ZN(n11451) );
  OAI21_X1 U9708 ( .B1(n14303), .B2(n7107), .A(n7105), .ZN(n14261) );
  AND2_X2 U9709 ( .A1(n11094), .A2(n14846), .ZN(n11095) );
  OR2_X1 U9710 ( .A1(n11045), .A2(n12047), .ZN(n11046) );
  NAND2_X1 U9711 ( .A1(n7126), .A2(n13902), .ZN(n7125) );
  INV_X1 U9712 ( .A(n7130), .ZN(n14296) );
  NOR2_X2 U9713 ( .A1(n14227), .A2(n14211), .ZN(n14213) );
  NOR2_X2 U9714 ( .A1(n14146), .A2(n14133), .ZN(n14111) );
  NAND2_X1 U9715 ( .A1(n8239), .A2(n7146), .ZN(n7145) );
  NAND3_X1 U9716 ( .A1(n7227), .A2(n7226), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n7155) );
  INV_X1 U9717 ( .A(n7894), .ZN(n7775) );
  AND2_X2 U9718 ( .A1(n7184), .A2(n7160), .ZN(n7206) );
  NAND3_X1 U9719 ( .A1(n12173), .A2(n12172), .A3(n7163), .ZN(n7187) );
  NAND4_X1 U9720 ( .A1(n8058), .A2(n8061), .A3(n8003), .A4(n8101), .ZN(n7165)
         );
  INV_X1 U9721 ( .A(n7167), .ZN(n7166) );
  INV_X1 U9722 ( .A(n12135), .ZN(n7169) );
  NAND2_X1 U9723 ( .A1(n7173), .A2(n7175), .ZN(n7172) );
  INV_X1 U9724 ( .A(n7175), .ZN(n7171) );
  XNOR2_X2 U9725 ( .A(n7176), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U9726 ( .A1(n7179), .A2(n7177), .ZN(n12044) );
  NAND2_X1 U9727 ( .A1(n7677), .A2(n7192), .ZN(n7190) );
  NAND2_X1 U9728 ( .A1(n7190), .A2(n6796), .ZN(n12075) );
  NAND3_X1 U9729 ( .A1(n7675), .A2(n12099), .A3(n7196), .ZN(n7194) );
  NAND2_X1 U9730 ( .A1(n7194), .A2(n7195), .ZN(n12129) );
  NAND2_X1 U9731 ( .A1(n7198), .A2(n7201), .ZN(n12156) );
  INV_X1 U9732 ( .A(n7207), .ZN(n12747) );
  OAI211_X1 U9733 ( .C1(n12721), .C2(n7212), .A(n7210), .B(n7208), .ZN(n7207)
         );
  NAND2_X1 U9734 ( .A1(n15262), .A2(n7211), .ZN(n7210) );
  INV_X1 U9735 ( .A(n7213), .ZN(n7211) );
  NAND2_X1 U9736 ( .A1(n15262), .A2(n6843), .ZN(n7212) );
  NOR2_X1 U9737 ( .A1(n12721), .A2(n12720), .ZN(n12745) );
  OAI21_X1 U9738 ( .B1(n12746), .B2(n6842), .A(n7214), .ZN(n7213) );
  NAND2_X1 U9739 ( .A1(n12746), .A2(n12743), .ZN(n7214) );
  XNOR2_X2 U9740 ( .A(n7218), .B(n7217), .ZN(n15172) );
  INV_X1 U9741 ( .A(n7222), .ZN(n10583) );
  AND2_X2 U9742 ( .A1(n7222), .A2(n7221), .ZN(n10581) );
  NOR2_X2 U9743 ( .A1(n12684), .A2(n13010), .ZN(n12716) );
  NAND3_X1 U9744 ( .A1(n7229), .A2(n11129), .A3(n7228), .ZN(n7231) );
  INV_X1 U9745 ( .A(n7231), .ZN(n11390) );
  NOR2_X2 U9746 ( .A1(n14547), .A2(n14548), .ZN(n14549) );
  NOR2_X2 U9747 ( .A1(n14555), .A2(n14556), .ZN(n14559) );
  XNOR2_X2 U9748 ( .A(n14504), .B(n15701), .ZN(n14532) );
  NAND2_X1 U9749 ( .A1(n7246), .A2(n15301), .ZN(n15324) );
  AND2_X1 U9750 ( .A1(n7246), .A2(n11854), .ZN(n11860) );
  NAND2_X1 U9751 ( .A1(n12856), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U9752 ( .A1(n7248), .A2(n7247), .ZN(n8848) );
  NAND2_X1 U9753 ( .A1(n11368), .A2(n7253), .ZN(n11602) );
  NAND2_X1 U9754 ( .A1(n11602), .A2(n11599), .ZN(n8650) );
  NAND2_X1 U9755 ( .A1(n12795), .A2(n8883), .ZN(n7259) );
  OAI21_X2 U9756 ( .B1(n12795), .B2(n7258), .A(n7254), .ZN(n12764) );
  NAND2_X1 U9757 ( .A1(n7260), .A2(n6802), .ZN(n11013) );
  NAND2_X1 U9758 ( .A1(n7264), .A2(n8740), .ZN(n7263) );
  NAND3_X1 U9759 ( .A1(n8612), .A2(n7267), .A3(n7261), .ZN(n7636) );
  NAND2_X1 U9760 ( .A1(n8568), .A2(n7268), .ZN(n7271) );
  NAND2_X1 U9761 ( .A1(n7271), .A2(n7269), .ZN(n11369) );
  NAND2_X1 U9762 ( .A1(n8478), .A2(n8479), .ZN(n8406) );
  NAND2_X1 U9763 ( .A1(n8478), .A2(n6808), .ZN(n13121) );
  NAND2_X1 U9764 ( .A1(n7276), .A2(n7274), .ZN(P3_U3204) );
  NAND2_X1 U9765 ( .A1(n12391), .A2(n15335), .ZN(n7276) );
  NAND3_X1 U9766 ( .A1(n7277), .A2(n7531), .A3(n7532), .ZN(n8610) );
  NAND2_X1 U9767 ( .A1(n9033), .A2(n7280), .ZN(n9663) );
  INV_X1 U9768 ( .A(n9663), .ZN(n9025) );
  NAND2_X1 U9769 ( .A1(n10811), .A2(n7285), .ZN(n7288) );
  NAND2_X1 U9770 ( .A1(n15056), .A2(n7289), .ZN(n7287) );
  NAND2_X1 U9771 ( .A1(n7288), .A2(n7286), .ZN(n10834) );
  NAND2_X1 U9772 ( .A1(n10811), .A2(n10810), .ZN(n7291) );
  INV_X1 U9773 ( .A(n15056), .ZN(n10801) );
  INV_X1 U9774 ( .A(n10814), .ZN(n7290) );
  NAND2_X1 U9775 ( .A1(n13629), .A2(n6704), .ZN(n7297) );
  OAI21_X1 U9776 ( .B1(n13555), .B2(n6681), .A(n13439), .ZN(n13541) );
  AOI22_X2 U9777 ( .A1(n11565), .A2(n7331), .B1(n11698), .B2(n7334), .ZN(
        n13666) );
  NAND2_X1 U9778 ( .A1(n11565), .A2(n7335), .ZN(n11701) );
  OR2_X2 U9779 ( .A1(n15188), .A2(n12662), .ZN(n7339) );
  MUX2_X1 U9780 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10076), .S(n10095), .Z(
        n10078) );
  NAND2_X1 U9781 ( .A1(n7356), .A2(n10191), .ZN(n10222) );
  OAI21_X1 U9782 ( .B1(n10211), .B2(n10210), .A(n7356), .ZN(n10864) );
  NAND2_X1 U9783 ( .A1(n10844), .A2(n7360), .ZN(n7359) );
  NAND2_X1 U9784 ( .A1(n11559), .A2(n11558), .ZN(n7364) );
  NAND2_X1 U9785 ( .A1(n11547), .A2(n11546), .ZN(n11559) );
  OAI211_X1 U9786 ( .C1(n11547), .C2(n11541), .A(n7362), .B(n6805), .ZN(n11691) );
  NAND2_X1 U9787 ( .A1(n7363), .A2(n11558), .ZN(n7362) );
  INV_X1 U9788 ( .A(n11546), .ZN(n7363) );
  INV_X1 U9789 ( .A(n9090), .ZN(n7378) );
  INV_X1 U9790 ( .A(n9058), .ZN(n13821) );
  NAND2_X2 U9791 ( .A1(n7378), .A2(n9058), .ZN(n9571) );
  OR2_X1 U9792 ( .A1(n9090), .A2(n9058), .ZN(n9558) );
  AOI21_X1 U9793 ( .B1(n7380), .B2(n7379), .A(n9090), .ZN(n7381) );
  NAND2_X1 U9794 ( .A1(n9058), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7379) );
  OR2_X1 U9795 ( .A1(n9058), .A2(n10925), .ZN(n7380) );
  OAI21_X1 U9796 ( .B1(n13534), .B2(n13478), .A(n13477), .ZN(n13479) );
  OAI22_X1 U9797 ( .A1(n13516), .A2(n13514), .B1(n13784), .B2(n13480), .ZN(
        n13501) );
  NAND2_X1 U9798 ( .A1(n10190), .A2(n10189), .ZN(n10211) );
  NAND2_X1 U9799 ( .A1(n11691), .A2(n11690), .ZN(n11692) );
  NAND2_X1 U9800 ( .A1(n10221), .A2(n10192), .ZN(n10194) );
  XNOR2_X2 U9801 ( .A(n9030), .B(n9054), .ZN(n9662) );
  NAND2_X1 U9802 ( .A1(n10222), .A2(n10225), .ZN(n10221) );
  XNOR2_X2 U9803 ( .A(n13372), .B(n9974), .ZN(n10214) );
  XNOR2_X2 U9804 ( .A(n8489), .B(n8490), .ZN(n9783) );
  AOI21_X1 U9805 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10539), .A(n10536), .ZN(
        n9684) );
  NOR2_X2 U9806 ( .A1(n14592), .A2(n14591), .ZN(n15783) );
  NAND2_X1 U9807 ( .A1(n14139), .A2(n6720), .ZN(n7389) );
  NAND2_X1 U9808 ( .A1(n7389), .A2(n7390), .ZN(n14102) );
  INV_X1 U9809 ( .A(n11028), .ZN(n7402) );
  NAND2_X1 U9810 ( .A1(n7405), .A2(n7403), .ZN(n7406) );
  NOR2_X1 U9811 ( .A1(n8311), .A2(n7404), .ZN(n7403) );
  NAND2_X1 U9812 ( .A1(n7406), .A2(n8312), .ZN(n10873) );
  INV_X2 U9813 ( .A(n8195), .ZN(n8282) );
  NAND4_X1 U9814 ( .A1(n7938), .A2(n7936), .A3(n7937), .A4(n7407), .ZN(n14038)
         );
  NAND2_X2 U9815 ( .A1(n9112), .A2(n7413), .ZN(n13374) );
  NAND3_X1 U9816 ( .A1(n7415), .A2(n7417), .A3(n7418), .ZN(n13818) );
  NAND2_X1 U9817 ( .A1(n13201), .A2(n7421), .ZN(n7420) );
  OAI211_X1 U9818 ( .C1(n13201), .C2(n7422), .A(n13233), .B(n7420), .ZN(
        P2_U3192) );
  NAND2_X1 U9819 ( .A1(n13201), .A2(n13200), .ZN(n13225) );
  INV_X1 U9820 ( .A(n13229), .ZN(n7429) );
  NAND2_X1 U9821 ( .A1(n11522), .A2(n7434), .ZN(n7433) );
  CLKBUF_X1 U9822 ( .A(n7447), .Z(n7442) );
  NAND2_X1 U9823 ( .A1(n13342), .A2(n13140), .ZN(n13251) );
  INV_X1 U9824 ( .A(n7442), .ZN(n13273) );
  INV_X1 U9825 ( .A(n13252), .ZN(n7448) );
  NAND2_X1 U9826 ( .A1(n7455), .A2(n7458), .ZN(n10748) );
  INV_X1 U9827 ( .A(n9152), .ZN(n9155) );
  NAND2_X1 U9828 ( .A1(n7474), .A2(n7472), .ZN(n9152) );
  NAND2_X1 U9829 ( .A1(n7473), .A2(n9135), .ZN(n7472) );
  INV_X1 U9830 ( .A(n7477), .ZN(n7473) );
  NAND2_X1 U9831 ( .A1(n7476), .A2(n7475), .ZN(n7474) );
  INV_X1 U9832 ( .A(n9136), .ZN(n7475) );
  NAND2_X1 U9833 ( .A1(n6827), .A2(n7480), .ZN(n9285) );
  INV_X1 U9834 ( .A(n9642), .ZN(n7484) );
  OR2_X2 U9835 ( .A1(n9173), .A2(n7485), .ZN(n7490) );
  NAND3_X1 U9836 ( .A1(n9213), .A2(n9212), .A3(n6789), .ZN(n7492) );
  AOI21_X1 U9837 ( .B1(n9377), .B2(n9376), .A(n9374), .ZN(n9375) );
  INV_X1 U9838 ( .A(n9362), .ZN(n7496) );
  NAND2_X1 U9839 ( .A1(n7497), .A2(n7498), .ZN(n9613) );
  NAND3_X1 U9840 ( .A1(n9459), .A2(n9458), .A3(n7500), .ZN(n7497) );
  INV_X1 U9841 ( .A(n9503), .ZN(n7504) );
  INV_X1 U9842 ( .A(n9266), .ZN(n7514) );
  NAND2_X1 U9843 ( .A1(n12473), .A2(n7538), .ZN(n7537) );
  NAND2_X1 U9844 ( .A1(n11301), .A2(n11579), .ZN(n7541) );
  NAND2_X1 U9845 ( .A1(n7541), .A2(n7542), .ZN(n15135) );
  NAND2_X1 U9846 ( .A1(n12548), .A2(n7547), .ZN(n7546) );
  OAI211_X1 U9847 ( .C1(n12548), .C2(n7548), .A(n7546), .B(n12554), .ZN(
        P3_U3169) );
  XNOR2_X1 U9848 ( .A(n12548), .B(n12465), .ZN(n12549) );
  AND2_X4 U9849 ( .A1(n10496), .A2(n7555), .ZN(n12484) );
  NAND3_X1 U9850 ( .A1(n10677), .A2(n9002), .A3(n13116), .ZN(n7555) );
  NAND2_X1 U9851 ( .A1(n11106), .A2(n11105), .ZN(n11294) );
  XNOR2_X1 U9852 ( .A(n12404), .B(n12405), .ZN(n12584) );
  INV_X1 U9853 ( .A(n8679), .ZN(n7561) );
  NAND2_X1 U9854 ( .A1(n7561), .A2(n10016), .ZN(n7562) );
  NAND3_X1 U9855 ( .A1(n7566), .A2(n7564), .A3(n7562), .ZN(n8688) );
  NAND4_X1 U9856 ( .A1(n7566), .A2(n7564), .A3(P1_DATAO_REG_13__SCAN_IN), .A4(
        n7562), .ZN(n8690) );
  NAND2_X1 U9857 ( .A1(n7568), .A2(n8418), .ZN(n7567) );
  INV_X1 U9858 ( .A(n8420), .ZN(n7570) );
  NAND2_X1 U9859 ( .A1(n7569), .A2(n8420), .ZN(n8526) );
  NAND2_X1 U9860 ( .A1(n8516), .A2(n8515), .ZN(n7569) );
  NAND2_X1 U9861 ( .A1(n8737), .A2(n7574), .ZN(n7571) );
  NAND2_X1 U9862 ( .A1(n7571), .A2(n7572), .ZN(n8769) );
  NAND3_X1 U9863 ( .A1(n11964), .A2(n11965), .A3(n11959), .ZN(n7583) );
  OAI21_X1 U9864 ( .B1(n8467), .B2(n7601), .A(n7600), .ZN(n8861) );
  NAND2_X1 U9865 ( .A1(n12829), .A2(n7622), .ZN(n12816) );
  NAND3_X1 U9866 ( .A1(n7627), .A2(n6741), .A3(n7626), .ZN(n7625) );
  CLKBUF_X1 U9867 ( .A(n8612), .Z(n7630) );
  NAND2_X1 U9868 ( .A1(n7635), .A2(n7633), .ZN(n11732) );
  INV_X1 U9869 ( .A(n7636), .ZN(n8478) );
  NAND2_X1 U9870 ( .A1(n9443), .A2(n7640), .ZN(n7639) );
  OAI21_X2 U9871 ( .B1(n7863), .B2(n7663), .A(n7661), .ZN(n7779) );
  INV_X1 U9872 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7662) );
  INV_X1 U9873 ( .A(n12156), .ZN(n12161) );
  NAND3_X1 U9874 ( .A1(n12091), .A2(n12090), .A3(n6800), .ZN(n7675) );
  NAND3_X1 U9875 ( .A1(n7679), .A2(n12210), .A3(n7678), .ZN(n7677) );
  NAND2_X1 U9876 ( .A1(n7680), .A2(n12062), .ZN(n7678) );
  NAND3_X1 U9877 ( .A1(n12040), .A2(n12025), .A3(n12030), .ZN(n7681) );
  NAND2_X1 U9878 ( .A1(n12150), .A2(n12151), .ZN(n12149) );
  NOR2_X1 U9879 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7687) );
  NOR2_X1 U9880 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7686) );
  NOR2_X1 U9881 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7685) );
  XNOR2_X2 U9882 ( .A(n7688), .B(n8289), .ZN(n14071) );
  NAND2_X1 U9883 ( .A1(n11040), .A2(n7691), .ZN(n7690) );
  NAND2_X1 U9884 ( .A1(n11025), .A2(n7696), .ZN(n7695) );
  AND2_X2 U9885 ( .A1(n12213), .A2(n7697), .ZN(n7696) );
  INV_X1 U9886 ( .A(n11504), .ZN(n8114) );
  NAND2_X1 U9887 ( .A1(n10519), .A2(n6751), .ZN(n7701) );
  NAND3_X1 U9888 ( .A1(n7701), .A2(n7182), .A3(n7700), .ZN(n10511) );
  NAND2_X1 U9889 ( .A1(n14326), .A2(n7702), .ZN(n8144) );
  INV_X1 U9890 ( .A(n8322), .ZN(n7704) );
  NAND2_X1 U9891 ( .A1(n6724), .A2(n7709), .ZN(n7705) );
  NAND2_X1 U9892 ( .A1(n6724), .A2(n7707), .ZN(n7706) );
  NAND2_X1 U9893 ( .A1(n14246), .A2(n7712), .ZN(n7710) );
  NAND2_X1 U9894 ( .A1(n7714), .A2(n8260), .ZN(n14121) );
  NAND2_X1 U9895 ( .A1(n13971), .A2(n7728), .ZN(n7726) );
  NAND2_X1 U9896 ( .A1(n7732), .A2(n7733), .ZN(n12382) );
  NAND2_X1 U9897 ( .A1(n13989), .A2(n7734), .ZN(n7732) );
  NAND2_X1 U9898 ( .A1(n13989), .A2(n13990), .ZN(n13988) );
  INV_X1 U9899 ( .A(n10792), .ZN(n7742) );
  OAI211_X2 U9900 ( .C1(n6690), .C2(n14874), .A(n9134), .B(n9133), .ZN(n9974)
         );
  OR2_X1 U9901 ( .A1(n9142), .A2(n9771), .ZN(n9133) );
  OR2_X2 U9902 ( .A1(n9377), .A2(n9376), .ZN(n7767) );
  AND2_X1 U9903 ( .A1(n10499), .A2(n10668), .ZN(n10502) );
  AND2_X1 U9904 ( .A1(n11268), .A2(n9094), .ZN(n9562) );
  XNOR2_X1 U9905 ( .A(n13486), .B(n13485), .ZN(n13690) );
  NAND2_X1 U9906 ( .A1(n8848), .A2(n8847), .ZN(n12819) );
  AOI21_X1 U9907 ( .B1(n9319), .B2(n9318), .A(n9317), .ZN(n9320) );
  NAND2_X1 U9908 ( .A1(n13501), .A2(n13481), .ZN(n13484) );
  AOI21_X2 U9909 ( .B1(n12574), .B2(n12832), .A(n12463), .ZN(n12548) );
  OR2_X1 U9910 ( .A1(n12388), .A2(n8905), .ZN(n10957) );
  INV_X1 U9911 ( .A(n8905), .ZN(n8894) );
  NAND2_X1 U9912 ( .A1(n8629), .A2(n8437), .ZN(n8439) );
  NAND2_X1 U9913 ( .A1(n8617), .A2(n8435), .ZN(n8629) );
  NAND2_X1 U9914 ( .A1(n8558), .A2(n8557), .ZN(n8429) );
  NAND2_X1 U9915 ( .A1(n8426), .A2(n8425), .ZN(n8558) );
  NAND2_X1 U9916 ( .A1(n8861), .A2(n8468), .ZN(n8470) );
  XNOR2_X1 U9917 ( .A(n12803), .B(n12806), .ZN(n12979) );
  OR2_X1 U9918 ( .A1(n8517), .A2(SI_10_), .ZN(n8649) );
  XNOR2_X1 U9919 ( .A(n8335), .B(n12224), .ZN(n14086) );
  NAND2_X1 U9920 ( .A1(n14086), .A2(n14688), .ZN(n8351) );
  XNOR2_X1 U9921 ( .A(n8263), .B(n8262), .ZN(n13828) );
  NAND2_X1 U9922 ( .A1(n8705), .A2(n8704), .ZN(n8707) );
  NAND2_X1 U9923 ( .A1(n8690), .A2(n8446), .ZN(n8705) );
  XNOR2_X1 U9924 ( .A(n8288), .B(n8287), .ZN(n14087) );
  INV_X1 U9925 ( .A(n9419), .ZN(n9422) );
  XNOR2_X1 U9926 ( .A(n9536), .B(n9535), .ZN(n13823) );
  INV_X1 U9927 ( .A(n8941), .ZN(n8944) );
  AND2_X1 U9928 ( .A1(n9411), .A2(n9412), .ZN(n9417) );
  INV_X1 U9929 ( .A(n7904), .ZN(n7898) );
  NAND2_X1 U9931 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  NAND2_X1 U9932 ( .A1(n8838), .A2(n8837), .ZN(n8466) );
  NOR2_X2 U9933 ( .A1(n11355), .A2(n11352), .ZN(n11522) );
  NAND2_X1 U9934 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  NAND2_X1 U9935 ( .A1(n8406), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8408) );
  INV_X1 U9936 ( .A(n13479), .ZN(n13516) );
  NAND2_X1 U9937 ( .A1(n11749), .A2(n11750), .ZN(n11768) );
  INV_X1 U9938 ( .A(n14261), .ZN(n8325) );
  NAND2_X1 U9939 ( .A1(n9303), .A2(n9302), .ZN(n9305) );
  XNOR2_X1 U9940 ( .A(n11843), .B(n11995), .ZN(n12966) );
  NAND2_X1 U9941 ( .A1(n7829), .A2(SI_18_), .ZN(n7830) );
  NAND2_X1 U9942 ( .A1(n8114), .A2(n12218), .ZN(n8116) );
  XNOR2_X1 U9943 ( .A(n8251), .B(n8250), .ZN(n13832) );
  XNOR2_X1 U9944 ( .A(n12760), .B(n12762), .ZN(n13037) );
  NAND2_X1 U9945 ( .A1(n9152), .A2(n9153), .ZN(n9157) );
  NAND2_X1 U9946 ( .A1(n6690), .A2(n13840), .ZN(n9098) );
  NOR3_X1 U9947 ( .A1(n13653), .A2(n13652), .A3(n13651), .ZN(n7756) );
  INV_X1 U9948 ( .A(n15067), .ZN(n13643) );
  AND2_X1 U9949 ( .A1(n12496), .A2(n8989), .ZN(n7757) );
  AND2_X1 U9950 ( .A1(n9054), .A2(n9053), .ZN(n7758) );
  AND2_X1 U9951 ( .A1(n9649), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7759) );
  CLKBUF_X2 U9952 ( .A(P1_U4016), .Z(n14042) );
  AND2_X2 U9953 ( .A1(n8977), .A2(n10413), .ZN(n15382) );
  INV_X1 U9954 ( .A(n14111), .ZN(n14132) );
  INV_X1 U9955 ( .A(n14127), .ZN(n14124) );
  INV_X1 U9956 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8481) );
  INV_X1 U9957 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8621) );
  NOR2_X1 U9958 ( .A1(n8988), .A2(n11492), .ZN(n7761) );
  AND2_X1 U9959 ( .A1(n9607), .A2(n7770), .ZN(n7763) );
  INV_X1 U9960 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9143) );
  AND2_X1 U9961 ( .A1(n14641), .A2(n12562), .ZN(n7764) );
  AOI22_X1 U9962 ( .A1(n13372), .A2(n9170), .B1(n9974), .B2(n9593), .ZN(n9135)
         );
  NOR2_X1 U9963 ( .A1(n8622), .A2(n8605), .ZN(n7765) );
  AND2_X2 U9964 ( .A1(n9671), .A2(n9670), .ZN(n14857) );
  INV_X1 U9965 ( .A(n14857), .ZN(n9673) );
  INV_X1 U9966 ( .A(n12021), .ZN(n14040) );
  INV_X1 U9967 ( .A(n11980), .ZN(n8635) );
  AND2_X1 U9968 ( .A1(n9008), .A2(n9007), .ZN(n7766) );
  AND2_X1 U9969 ( .A1(n8336), .A2(n12009), .ZN(n14352) );
  AND2_X1 U9970 ( .A1(n13799), .A2(n13465), .ZN(n7768) );
  AND2_X1 U9971 ( .A1(n11767), .A2(n11769), .ZN(n7769) );
  AND2_X1 U9972 ( .A1(n9600), .A2(n9599), .ZN(n7770) );
  NAND2_X1 U9973 ( .A1(n14040), .A2(n7127), .ZN(n12031) );
  NAND2_X1 U9974 ( .A1(n9170), .A2(n13374), .ZN(n9114) );
  INV_X1 U9975 ( .A(n9151), .ZN(n9156) );
  NAND2_X1 U9976 ( .A1(n9211), .A2(n9210), .ZN(n9212) );
  OAI22_X1 U9977 ( .A1(n15103), .A2(n6685), .B1(n9435), .B2(n10823), .ZN(n9229) );
  NAND2_X1 U9978 ( .A1(n9250), .A2(n9249), .ZN(n9269) );
  OAI21_X1 U9979 ( .B1(n9303), .B2(n9302), .A(n9301), .ZN(n9304) );
  INV_X1 U9980 ( .A(n11979), .ZN(n11881) );
  NAND2_X1 U9981 ( .A1(n9378), .A2(n7767), .ZN(n9393) );
  INV_X1 U9982 ( .A(n9410), .ZN(n9416) );
  OAI22_X1 U9983 ( .A1(n13617), .A2(n9435), .B1(n13462), .B2(n6685), .ZN(n9420) );
  INV_X1 U9984 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9010) );
  INV_X1 U9985 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U9986 ( .A1(n9609), .A2(n9610), .ZN(n9611) );
  AND2_X1 U9987 ( .A1(n9027), .A2(n9649), .ZN(n9028) );
  INV_X1 U9988 ( .A(n12776), .ZN(n8895) );
  AND2_X1 U9989 ( .A1(n12898), .A2(n12897), .ZN(n8781) );
  INV_X1 U9990 ( .A(n11870), .ZN(n8567) );
  INV_X1 U9991 ( .A(n14262), .ZN(n8324) );
  NOR2_X1 U9992 ( .A1(n8187), .A2(SI_21_), .ZN(n7837) );
  INV_X1 U9993 ( .A(n8130), .ZN(n7828) );
  INV_X1 U9994 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12392) );
  INV_X1 U9995 ( .A(n8864), .ZN(n8396) );
  INV_X1 U9996 ( .A(n8696), .ZN(n8387) );
  NAND2_X1 U9997 ( .A1(n11895), .A2(n11894), .ZN(n11984) );
  INV_X1 U9998 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9221) );
  NOR2_X1 U9999 ( .A1(n9328), .A2(n9327), .ZN(n9326) );
  AND2_X1 U10000 ( .A1(n9383), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9050) );
  AND2_X1 U10001 ( .A1(n11655), .A2(n11673), .ZN(n11657) );
  OR2_X1 U10002 ( .A1(n9356), .A2(n13257), .ZN(n9367) );
  OR2_X1 U10003 ( .A1(n9310), .A2(n9309), .ZN(n9328) );
  INV_X1 U10004 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9182) );
  INV_X1 U10005 ( .A(n9643), .ZN(n9645) );
  INV_X1 U10006 ( .A(n14435), .ZN(n8338) );
  NOR2_X1 U10007 ( .A1(n8047), .A2(n8046), .ZN(n8064) );
  INV_X1 U10008 ( .A(n8013), .ZN(n7807) );
  AND2_X1 U10009 ( .A1(n8604), .A2(n15749), .ZN(n8622) );
  NOR2_X1 U10010 ( .A1(n12462), .A2(n12461), .ZN(n12463) );
  INV_X4 U10011 ( .A(n8494), .ZN(n10948) );
  INV_X1 U10012 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15749) );
  NAND2_X1 U10013 ( .A1(n8396), .A2(n8395), .ZN(n8876) );
  INV_X1 U10014 ( .A(n8830), .ZN(n8394) );
  OR2_X1 U10015 ( .A1(n8747), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8775) );
  AND2_X1 U10016 ( .A1(n15268), .A2(n8987), .ZN(n11492) );
  OAI21_X1 U10017 ( .B1(n12390), .B2(n13114), .A(n9005), .ZN(n9006) );
  AOI21_X1 U10018 ( .B1(n11723), .B2(n8703), .A(n7764), .ZN(n12945) );
  NAND2_X1 U10019 ( .A1(n8540), .A2(n8539), .ZN(n8426) );
  INV_X1 U10020 ( .A(n13217), .ZN(n13153) );
  NOR2_X1 U10021 ( .A1(n9469), .A2(n13285), .ZN(n9493) );
  AND2_X1 U10022 ( .A1(n9050), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9426) );
  OR2_X1 U10023 ( .A1(n14976), .A2(n14975), .ZN(n14978) );
  OR2_X1 U10024 ( .A1(n15015), .A2(n15014), .ZN(n15011) );
  NAND2_X1 U10025 ( .A1(n9258), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9294) );
  INV_X1 U10026 ( .A(n15103), .ZN(n10850) );
  INV_X1 U10027 ( .A(n13355), .ZN(n11571) );
  INV_X1 U10028 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9014) );
  OR2_X1 U10029 ( .A1(n8078), .A2(n8077), .ZN(n8108) );
  NOR2_X1 U10030 ( .A1(n8108), .A2(n8107), .ZN(n8123) );
  INV_X1 U10031 ( .A(n8193), .ZN(n8206) );
  NAND2_X1 U10032 ( .A1(n7966), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7993) );
  INV_X1 U10033 ( .A(n12188), .ZN(n12014) );
  OR2_X1 U10034 ( .A1(n8154), .A2(n8153), .ZN(n8166) );
  INV_X1 U10035 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8030) );
  NOR2_X1 U10036 ( .A1(n14088), .A2(n8349), .ZN(n8350) );
  OR2_X1 U10037 ( .A1(n9904), .A2(n8374), .ZN(n10348) );
  AND2_X1 U10038 ( .A1(n7817), .A2(n7816), .ZN(n8038) );
  NAND2_X1 U10039 ( .A1(n14550), .A2(n14551), .ZN(n14510) );
  NAND2_X1 U10040 ( .A1(n8622), .A2(n8621), .ZN(n8636) );
  OR2_X1 U10041 ( .A1(n10291), .A2(n12003), .ZN(n15143) );
  OR2_X1 U10042 ( .A1(n8818), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U10043 ( .A1(n11968), .A2(n11969), .ZN(n11995) );
  INV_X1 U10044 ( .A(n9006), .ZN(n9007) );
  NAND2_X1 U10045 ( .A1(n13054), .A2(n12833), .ZN(n11952) );
  AND2_X1 U10046 ( .A1(n11919), .A2(n11920), .ZN(n12921) );
  AND2_X1 U10047 ( .A1(n9003), .A2(n10411), .ZN(n15289) );
  AND2_X1 U10048 ( .A1(n8943), .A2(n11416), .ZN(n8948) );
  NAND2_X1 U10049 ( .A1(n8707), .A2(n8448), .ZN(n8721) );
  AND2_X1 U10050 ( .A1(n8443), .A2(n8442), .ZN(n8662) );
  AND2_X1 U10051 ( .A1(n8425), .A2(n8424), .ZN(n8539) );
  NAND2_X2 U10052 ( .A1(n11332), .A2(n9924), .ZN(n10229) );
  XNOR2_X1 U10053 ( .A(n9925), .B(n10229), .ZN(n9973) );
  OR2_X1 U10054 ( .A1(n10457), .A2(n15071), .ZN(n9966) );
  OR2_X1 U10055 ( .A1(n9896), .A2(n9895), .ZN(n10000) );
  OR2_X1 U10056 ( .A1(n14961), .A2(n14960), .ZN(n14963) );
  OR2_X1 U10057 ( .A1(n9993), .A2(n9994), .ZN(n10166) );
  INV_X1 U10058 ( .A(n13482), .ZN(n13447) );
  INV_X1 U10059 ( .A(n11700), .ZN(n11698) );
  INV_X1 U10060 ( .A(n11541), .ZN(n11558) );
  AND2_X1 U10061 ( .A1(n13866), .A2(n12328), .ZN(n13968) );
  AND3_X1 U10062 ( .A1(n10349), .A2(n10881), .A3(n10348), .ZN(n10355) );
  OR2_X1 U10063 ( .A1(n8166), .A2(n8165), .ZN(n8175) );
  OR2_X1 U10064 ( .A1(n14409), .A2(n14024), .ZN(n8322) );
  AND2_X1 U10065 ( .A1(n10884), .A2(n10883), .ZN(n10888) );
  INV_X1 U10066 ( .A(n14238), .ZN(n14316) );
  AND2_X1 U10067 ( .A1(n8342), .A2(n10891), .ZN(n14852) );
  INV_X1 U10068 ( .A(n7933), .ZN(n12034) );
  AND2_X1 U10069 ( .A1(n8846), .A2(n8845), .ZN(n12579) );
  OR2_X1 U10070 ( .A1(n8636), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8652) );
  INV_X1 U10071 ( .A(n15143), .ZN(n15149) );
  AND2_X1 U10072 ( .A1(n10278), .A2(n10277), .ZN(n15140) );
  NAND2_X1 U10073 ( .A1(n8882), .A2(n8881), .ZN(n12523) );
  INV_X1 U10074 ( .A(n12474), .ZN(n12505) );
  INV_X1 U10075 ( .A(n12562), .ZN(n12947) );
  OR2_X1 U10076 ( .A1(n8652), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8669) );
  INV_X1 U10077 ( .A(n11375), .ZN(n15295) );
  AND2_X1 U10078 ( .A1(n10677), .A2(n10772), .ZN(n15328) );
  INV_X1 U10079 ( .A(n12971), .ZN(n15380) );
  OR2_X2 U10080 ( .A1(n8802), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8804) );
  INV_X1 U10081 ( .A(n13312), .ZN(n13409) );
  AND4_X1 U10082 ( .A1(n9466), .A2(n9465), .A3(n9464), .A4(n9463), .ZN(n13469)
         );
  AND3_X1 U10083 ( .A1(n9360), .A2(n9359), .A3(n9358), .ZN(n13451) );
  INV_X1 U10084 ( .A(n15013), .ZN(n15032) );
  AND2_X1 U10085 ( .A1(n9898), .A2(n9875), .ZN(n15028) );
  NAND2_X1 U10086 ( .A1(n9965), .A2(n15072), .ZN(n15052) );
  INV_X1 U10087 ( .A(n15111), .ZN(n15079) );
  AND2_X1 U10088 ( .A1(n10045), .A2(n10044), .ZN(n10338) );
  AND2_X1 U10089 ( .A1(n9254), .A2(n9270), .ZN(n10002) );
  NAND2_X1 U10090 ( .A1(n10354), .A2(n14323), .ZN(n14012) );
  AND4_X1 U10091 ( .A1(n8223), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n14179)
         );
  AND4_X1 U10092 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n8110), .ZN(n14315)
         );
  OR2_X1 U10093 ( .A1(n14731), .A2(n14727), .ZN(n14785) );
  INV_X1 U10094 ( .A(n14785), .ZN(n14819) );
  NAND2_X1 U10095 ( .A1(n12237), .A2(n10353), .ZN(n14323) );
  NAND2_X1 U10096 ( .A1(n14319), .A2(n10892), .ZN(n14300) );
  AOI21_X1 U10097 ( .B1(n8384), .B2(n9906), .A(n9905), .ZN(n10881) );
  AND2_X1 U10098 ( .A1(n14857), .A2(n14680), .ZN(n14436) );
  INV_X1 U10099 ( .A(n14352), .ZN(n14688) );
  NOR2_X1 U10100 ( .A1(n8382), .A2(n10882), .ZN(n9671) );
  AND2_X1 U10101 ( .A1(n8026), .A2(n8042), .ZN(n11176) );
  AND2_X1 U10102 ( .A1(n9759), .A2(n9758), .ZN(n15232) );
  AND2_X1 U10103 ( .A1(n10294), .A2(n10293), .ZN(n15159) );
  NAND2_X1 U10104 ( .A1(n10276), .A2(n10413), .ZN(n15146) );
  NOR2_X1 U10105 ( .A1(n10284), .A2(n11797), .ZN(n10932) );
  CLKBUF_X1 U10106 ( .A(n10932), .Z(n10958) );
  INV_X1 U10107 ( .A(n15232), .ZN(n15251) );
  INV_X1 U10108 ( .A(n15262), .ZN(n15241) );
  NAND2_X1 U10109 ( .A1(n10477), .A2(n15328), .ZN(n15307) );
  INV_X1 U10110 ( .A(n13016), .ZN(n13024) );
  OR2_X1 U10111 ( .A1(n10426), .A2(n10425), .ZN(n15394) );
  INV_X1 U10112 ( .A(n15382), .ZN(n9009) );
  INV_X1 U10113 ( .A(n13109), .ZN(n13105) );
  OR2_X1 U10114 ( .A1(n11798), .A2(n11797), .ZN(n11799) );
  INV_X1 U10115 ( .A(SI_13_), .ZN(n15723) );
  INV_X1 U10116 ( .A(n13334), .ZN(n13348) );
  INV_X1 U10117 ( .A(n9967), .ZN(n13354) );
  INV_X1 U10118 ( .A(n9626), .ZN(n13428) );
  INV_X1 U10119 ( .A(n11279), .ZN(n13364) );
  INV_X1 U10120 ( .A(n14864), .ZN(n15044) );
  INV_X1 U10121 ( .A(n15055), .ZN(n13678) );
  INV_X1 U10122 ( .A(n13609), .ZN(n15063) );
  INV_X1 U10123 ( .A(n13503), .ZN(n13780) );
  NAND2_X1 U10124 ( .A1(n10338), .A2(n10337), .ZN(n15117) );
  AND2_X1 U10125 ( .A1(n9960), .A2(n9660), .ZN(n15072) );
  INV_X1 U10126 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9921) );
  INV_X1 U10127 ( .A(n14012), .ZN(n14002) );
  INV_X1 U10128 ( .A(n14305), .ZN(n14023) );
  OR2_X1 U10129 ( .A1(n14731), .A2(n10268), .ZN(n14828) );
  INV_X1 U10130 ( .A(n14729), .ZN(n14832) );
  INV_X1 U10131 ( .A(n14086), .ZN(n14100) );
  INV_X1 U10132 ( .A(n14329), .ZN(n14313) );
  AND2_X1 U10133 ( .A1(n14091), .A2(n14323), .ZN(n14309) );
  INV_X1 U10134 ( .A(n14345), .ZN(n14419) );
  INV_X1 U10135 ( .A(n14133), .ZN(n14440) );
  AND2_X1 U10136 ( .A1(n9986), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9909) );
  INV_X1 U10137 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10016) );
  INV_X1 U10138 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9919) );
  NOR2_X1 U10139 ( .A1(P2_U3088), .A2(n9871), .ZN(P2_U3947) );
  NAND2_X1 U10140 ( .A1(n7779), .A2(SI_1_), .ZN(n7780) );
  INV_X1 U10141 ( .A(SI_1_), .ZN(n9782) );
  OAI21_X1 U10142 ( .B1(SI_2_), .B2(n9782), .A(n7779), .ZN(n7774) );
  INV_X1 U10143 ( .A(SI_2_), .ZN(n15689) );
  OAI21_X1 U10144 ( .B1(SI_1_), .B2(n15689), .A(n7772), .ZN(n7773) );
  NAND2_X1 U10145 ( .A1(n7774), .A2(n7773), .ZN(n7777) );
  OAI211_X1 U10146 ( .C1(SI_1_), .C2(n7779), .A(n7775), .B(n15689), .ZN(n7776)
         );
  NAND3_X1 U10147 ( .A1(n7778), .A2(n7777), .A3(n7776), .ZN(n7917) );
  MUX2_X1 U10148 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7863), .Z(n7916) );
  NAND2_X1 U10149 ( .A1(n7917), .A2(n7916), .ZN(n7783) );
  NAND2_X1 U10150 ( .A1(n7781), .A2(SI_2_), .ZN(n7782) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7863), .Z(n7785) );
  NAND2_X1 U10152 ( .A1(n7785), .A2(SI_3_), .ZN(n7786) );
  MUX2_X1 U10153 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7845), .Z(n7788) );
  INV_X1 U10154 ( .A(n7939), .ZN(n7787) );
  NAND2_X1 U10155 ( .A1(n7788), .A2(SI_4_), .ZN(n7789) );
  MUX2_X1 U10156 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7845), .Z(n7792) );
  NAND2_X1 U10157 ( .A1(n7792), .A2(SI_5_), .ZN(n7793) );
  MUX2_X1 U10158 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7845), .Z(n7795) );
  NAND2_X1 U10159 ( .A1(n7795), .A2(SI_6_), .ZN(n7796) );
  MUX2_X1 U10160 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n7845), .Z(n7798) );
  NAND2_X1 U10161 ( .A1(n7798), .A2(SI_7_), .ZN(n7799) );
  MUX2_X1 U10162 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n7845), .Z(n7801) );
  NAND2_X1 U10163 ( .A1(n7801), .A2(SI_8_), .ZN(n7802) );
  MUX2_X1 U10164 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n7845), .Z(n7804) );
  NAND2_X1 U10165 ( .A1(n7804), .A2(SI_9_), .ZN(n7805) );
  MUX2_X1 U10166 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n7845), .Z(n7808) );
  INV_X1 U10167 ( .A(n7810), .ZN(n7811) );
  NAND2_X1 U10168 ( .A1(n7811), .A2(SI_11_), .ZN(n7812) );
  MUX2_X1 U10169 ( .A(n9919), .B(n9921), .S(n7845), .Z(n7814) );
  NAND2_X1 U10170 ( .A1(n7814), .A2(n15480), .ZN(n7817) );
  INV_X1 U10171 ( .A(n7814), .ZN(n7815) );
  NAND2_X1 U10172 ( .A1(n7815), .A2(SI_12_), .ZN(n7816) );
  MUX2_X1 U10173 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9773), .Z(n8055) );
  INV_X1 U10174 ( .A(SI_14_), .ZN(n15542) );
  MUX2_X1 U10175 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n7845), .Z(n8072) );
  INV_X1 U10176 ( .A(n8072), .ZN(n8087) );
  MUX2_X1 U10177 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n7845), .Z(n8092) );
  NAND2_X1 U10178 ( .A1(n8092), .A2(SI_15_), .ZN(n7821) );
  OAI21_X1 U10179 ( .B1(n15542), .B2(n8087), .A(n7821), .ZN(n7818) );
  INV_X1 U10180 ( .A(n7818), .ZN(n7819) );
  NOR2_X1 U10181 ( .A1(n8072), .A2(SI_14_), .ZN(n7822) );
  INV_X1 U10182 ( .A(SI_15_), .ZN(n9852) );
  INV_X1 U10183 ( .A(n8092), .ZN(n7820) );
  AOI22_X1 U10184 ( .A1(n7822), .A2(n7821), .B1(n9852), .B2(n7820), .ZN(n7823)
         );
  MUX2_X1 U10185 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n7845), .Z(n7825) );
  XNOR2_X1 U10186 ( .A(n7825), .B(n15453), .ZN(n8117) );
  INV_X1 U10187 ( .A(n7825), .ZN(n7826) );
  NAND2_X1 U10188 ( .A1(n7826), .A2(n15453), .ZN(n7827) );
  INV_X1 U10189 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10314) );
  MUX2_X1 U10190 ( .A(n10300), .B(n10314), .S(n7845), .Z(n8130) );
  MUX2_X1 U10191 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9773), .Z(n8145) );
  INV_X1 U10192 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10909) );
  INV_X1 U10193 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10907) );
  MUX2_X1 U10194 ( .A(n10909), .B(n10907), .S(n9773), .Z(n7831) );
  INV_X1 U10195 ( .A(SI_19_), .ZN(n10164) );
  NAND2_X1 U10196 ( .A1(n7831), .A2(n10164), .ZN(n7834) );
  INV_X1 U10197 ( .A(n7831), .ZN(n7832) );
  NAND2_X1 U10198 ( .A1(n7832), .A2(SI_19_), .ZN(n7833) );
  NAND2_X1 U10199 ( .A1(n7834), .A2(n7833), .ZN(n8159) );
  MUX2_X1 U10200 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9773), .Z(n8187) );
  MUX2_X1 U10201 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9773), .Z(n8182) );
  NOR2_X1 U10202 ( .A1(n8182), .A2(SI_20_), .ZN(n7835) );
  INV_X1 U10203 ( .A(n8182), .ZN(n7836) );
  INV_X1 U10204 ( .A(SI_20_), .ZN(n10454) );
  NOR2_X1 U10205 ( .A1(n7836), .A2(n10454), .ZN(n7839) );
  INV_X1 U10206 ( .A(n7837), .ZN(n7838) );
  AOI22_X1 U10207 ( .A1(n7839), .A2(n7838), .B1(n8187), .B2(SI_21_), .ZN(n7840) );
  INV_X1 U10208 ( .A(SI_22_), .ZN(n15742) );
  XNOR2_X2 U10209 ( .A(n7841), .B(n15742), .ZN(n9443) );
  MUX2_X1 U10210 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9773), .Z(n9442) );
  MUX2_X1 U10211 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9773), .Z(n8212) );
  INV_X1 U10212 ( .A(n8212), .ZN(n7843) );
  INV_X1 U10213 ( .A(SI_23_), .ZN(n15478) );
  NAND2_X1 U10214 ( .A1(n8212), .A2(SI_23_), .ZN(n7844) );
  MUX2_X1 U10215 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9773), .Z(n8226) );
  INV_X1 U10216 ( .A(n8226), .ZN(n7848) );
  NAND2_X1 U10217 ( .A1(n7846), .A2(SI_24_), .ZN(n7847) );
  INV_X1 U10218 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11822) );
  INV_X1 U10219 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13838) );
  MUX2_X1 U10220 ( .A(n11822), .B(n13838), .S(n9773), .Z(n7849) );
  INV_X1 U10221 ( .A(SI_25_), .ZN(n15715) );
  NAND2_X1 U10222 ( .A1(n7849), .A2(n15715), .ZN(n7852) );
  INV_X1 U10223 ( .A(n7849), .ZN(n7850) );
  NAND2_X1 U10224 ( .A1(n7850), .A2(SI_25_), .ZN(n7851) );
  NAND2_X1 U10225 ( .A1(n7852), .A2(n7851), .ZN(n8238) );
  INV_X1 U10226 ( .A(SI_26_), .ZN(n15673) );
  INV_X1 U10227 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14491) );
  INV_X1 U10228 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13833) );
  MUX2_X1 U10229 ( .A(n14491), .B(n13833), .S(n9773), .Z(n8249) );
  INV_X1 U10230 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14487) );
  INV_X1 U10231 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8473) );
  MUX2_X1 U10232 ( .A(n14487), .B(n8473), .S(n9773), .Z(n8261) );
  INV_X1 U10233 ( .A(n8261), .ZN(n7854) );
  NOR2_X1 U10234 ( .A1(n7854), .A2(SI_27_), .ZN(n7853) );
  INV_X1 U10235 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14485) );
  INV_X1 U10236 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8900) );
  MUX2_X1 U10237 ( .A(n14485), .B(n8900), .S(n9773), .Z(n7855) );
  INV_X1 U10238 ( .A(SI_28_), .ZN(n15660) );
  NAND2_X1 U10239 ( .A1(n7855), .A2(n15660), .ZN(n8277) );
  INV_X1 U10240 ( .A(n7855), .ZN(n7856) );
  NAND2_X1 U10241 ( .A1(n7856), .A2(SI_28_), .ZN(n7857) );
  NAND2_X1 U10242 ( .A1(n8277), .A2(n7857), .ZN(n8278) );
  INV_X2 U10243 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8101) );
  NOR2_X1 U10244 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n7860) );
  NOR2_X1 U10245 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n7859) );
  NOR2_X1 U10246 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n7858) );
  XNOR2_X2 U10247 ( .A(n7861), .B(n7866), .ZN(n14483) );
  NAND2_X4 U10248 ( .A1(n8204), .A2(n9773), .ZN(n7930) );
  OR2_X1 U10249 ( .A1(n7930), .A2(n14485), .ZN(n7864) );
  INV_X1 U10250 ( .A(n7872), .ZN(n14477) );
  INV_X1 U10251 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7869) );
  NAND2_X2 U10252 ( .A1(n14477), .A2(n14481), .ZN(n7921) );
  NAND2_X1 U10253 ( .A1(n6687), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U10254 ( .A1(n6943), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7883) );
  NOR2_X2 U10255 ( .A1(n7872), .A2(n14481), .ZN(n7885) );
  NAND2_X1 U10256 ( .A1(n7922), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7882) );
  INV_X1 U10257 ( .A(n14481), .ZN(n7871) );
  NAND2_X1 U10259 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n7873) );
  INV_X1 U10260 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8029) );
  INV_X1 U10261 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10262 ( .A1(n8064), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8078) );
  INV_X1 U10263 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8077) );
  INV_X1 U10264 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U10265 ( .A1(n8137), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8154) );
  INV_X1 U10266 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8153) );
  INV_X1 U10267 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8165) );
  INV_X1 U10268 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U10269 ( .A1(n8192), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U10270 ( .A1(n8206), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8205) );
  NAND2_X1 U10271 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n8218), .ZN(n8231) );
  INV_X1 U10272 ( .A(n8231), .ZN(n7874) );
  NAND2_X1 U10273 ( .A1(n7874), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8242) );
  INV_X1 U10274 ( .A(n8242), .ZN(n7875) );
  NAND2_X1 U10275 ( .A1(n7875), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8254) );
  INV_X1 U10276 ( .A(n8254), .ZN(n7876) );
  NAND2_X1 U10277 ( .A1(n7876), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8266) );
  INV_X1 U10278 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13847) );
  INV_X1 U10279 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7877) );
  OAI21_X1 U10280 ( .B1(n8266), .B2(n13847), .A(n7877), .ZN(n7880) );
  INV_X1 U10281 ( .A(n8266), .ZN(n7879) );
  AND2_X1 U10282 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n7878) );
  NAND2_X1 U10283 ( .A1(n7879), .A2(n7878), .ZN(n14089) );
  NAND2_X1 U10284 ( .A1(n7880), .A2(n14089), .ZN(n14115) );
  OR2_X1 U10285 ( .A1(n8282), .A2(n14115), .ZN(n7881) );
  NAND4_X1 U10286 ( .A1(n7884), .A2(n7883), .A3(n7882), .A4(n7881), .ZN(n14018) );
  INV_X1 U10287 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11003) );
  NAND2_X1 U10288 ( .A1(n11810), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7889) );
  INV_X1 U10289 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10094) );
  OR2_X1 U10290 ( .A1(n11814), .A2(n10094), .ZN(n7888) );
  INV_X1 U10291 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10292 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n7891) );
  INV_X1 U10293 ( .A(n7892), .ZN(n7893) );
  XNOR2_X1 U10294 ( .A(n7895), .B(n7894), .ZN(n9818) );
  OR2_X1 U10295 ( .A1(n11805), .A2(n9818), .ZN(n7897) );
  OR2_X1 U10296 ( .A1(n7930), .A2(n7663), .ZN(n7896) );
  NAND2_X1 U10297 ( .A1(n7904), .A2(n6967), .ZN(n12025) );
  NAND2_X1 U10298 ( .A1(n7923), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10299 ( .A1(n7885), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7900) );
  NAND4_X4 U10300 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n14043) );
  INV_X1 U10301 ( .A(SI_0_), .ZN(n9808) );
  XNOR2_X1 U10302 ( .A(n7903), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14497) );
  MUX2_X1 U10303 ( .A(n7684), .B(n14497), .S(n8204), .Z(n12017) );
  INV_X1 U10304 ( .A(n12017), .ZN(n10446) );
  NAND2_X1 U10305 ( .A1(n14043), .A2(n10446), .ZN(n10520) );
  NAND2_X1 U10306 ( .A1(n7904), .A2(n11001), .ZN(n7905) );
  INV_X1 U10307 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7906) );
  OR2_X1 U10308 ( .A1(n7921), .A2(n7906), .ZN(n7910) );
  INV_X1 U10309 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10899) );
  OR2_X1 U10310 ( .A1(n8267), .A2(n10899), .ZN(n7909) );
  NAND2_X1 U10311 ( .A1(n7885), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U10312 ( .A1(n11810), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7907) );
  AND4_X2 U10313 ( .A1(n7909), .A2(n7910), .A3(n7908), .A4(n7907), .ZN(n12021)
         );
  NOR2_X1 U10314 ( .A1(n7892), .A2(n8290), .ZN(n7911) );
  INV_X1 U10315 ( .A(n7912), .ZN(n7915) );
  INV_X1 U10316 ( .A(n7913), .ZN(n7914) );
  XNOR2_X1 U10317 ( .A(n7917), .B(n7916), .ZN(n9796) );
  OAI211_X1 U10318 ( .C1(n8204), .C2(n10097), .A(n7919), .B(n7918), .ZN(n12022) );
  NAND2_X1 U10319 ( .A1(n12021), .A2(n7127), .ZN(n7920) );
  INV_X2 U10320 ( .A(n7921), .ZN(n8345) );
  NAND2_X1 U10321 ( .A1(n7885), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U10322 ( .A1(n11810), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7925) );
  OR2_X1 U10323 ( .A1(n7913), .A2(n8290), .ZN(n7928) );
  XNOR2_X1 U10324 ( .A(n7928), .B(n15757), .ZN(n10098) );
  NAND2_X1 U10325 ( .A1(n9767), .A2(n7941), .ZN(n7932) );
  OR2_X1 U10326 ( .A1(n7930), .A2(n9768), .ZN(n7931) );
  OAI211_X1 U10327 ( .C1(n8204), .C2(n10098), .A(n7932), .B(n7931), .ZN(n7933)
         );
  XNOR2_X2 U10328 ( .A(n14039), .B(n12033), .ZN(n12202) );
  NAND2_X1 U10329 ( .A1(n10788), .A2(n12034), .ZN(n7934) );
  NAND2_X1 U10330 ( .A1(n10511), .A2(n7934), .ZN(n10547) );
  NAND2_X1 U10331 ( .A1(n8345), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7938) );
  INV_X1 U10332 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7935) );
  OR2_X1 U10333 ( .A1(n8217), .A2(n7935), .ZN(n7937) );
  XNOR2_X1 U10334 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11267) );
  INV_X1 U10335 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10107) );
  OR2_X1 U10336 ( .A1(n6899), .A2(n10107), .ZN(n7936) );
  XNOR2_X1 U10337 ( .A(n7940), .B(n7939), .ZN(n9792) );
  NAND2_X1 U10338 ( .A1(n9792), .A2(n7941), .ZN(n7944) );
  INV_X2 U10339 ( .A(n7930), .ZN(n8162) );
  INV_X2 U10340 ( .A(n8204), .ZN(n9985) );
  NAND2_X1 U10341 ( .A1(n7913), .A2(n15757), .ZN(n7948) );
  NAND2_X1 U10342 ( .A1(n7948), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7942) );
  XNOR2_X1 U10343 ( .A(n7942), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U10344 ( .A1(n8162), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9985), .B2(
        n10116), .ZN(n7943) );
  AND2_X2 U10345 ( .A1(n7944), .A2(n7943), .ZN(n12038) );
  XNOR2_X1 U10346 ( .A(n14038), .B(n12038), .ZN(n12204) );
  NAND2_X1 U10347 ( .A1(n10547), .A2(n12204), .ZN(n10546) );
  NAND2_X1 U10348 ( .A1(n12039), .A2(n12038), .ZN(n7945) );
  XNOR2_X1 U10349 ( .A(n7947), .B(n7946), .ZN(n9814) );
  NAND2_X1 U10350 ( .A1(n9814), .A2(n11804), .ZN(n7951) );
  NAND2_X1 U10351 ( .A1(n7960), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7949) );
  XNOR2_X1 U10352 ( .A(n7949), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U10353 ( .A1(n8162), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9985), .B2(
        n10117), .ZN(n7950) );
  NAND2_X1 U10354 ( .A1(n7923), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U10355 ( .A1(n6687), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7955) );
  AOI21_X1 U10356 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7952) );
  NOR2_X1 U10357 ( .A1(n7952), .A2(n7966), .ZN(n11253) );
  NAND2_X1 U10358 ( .A1(n8195), .A2(n11253), .ZN(n7954) );
  NAND2_X1 U10359 ( .A1(n7922), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7953) );
  NAND4_X1 U10360 ( .A1(n7956), .A2(n7955), .A3(n7954), .A4(n7953), .ZN(n14037) );
  XNOR2_X1 U10361 ( .A(n12047), .B(n11408), .ZN(n12205) );
  OR2_X1 U10362 ( .A1(n12047), .A2(n14037), .ZN(n7957) );
  NAND2_X1 U10363 ( .A1(n9820), .A2(n11804), .ZN(n7965) );
  INV_X1 U10364 ( .A(n7960), .ZN(n7962) );
  INV_X1 U10365 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U10366 ( .A1(n7962), .A2(n7961), .ZN(n7973) );
  NAND2_X1 U10367 ( .A1(n7973), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7963) );
  XNOR2_X1 U10368 ( .A(n7963), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U10369 ( .A1(n8162), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9985), .B2(
        n10156), .ZN(n7964) );
  NAND2_X1 U10370 ( .A1(n7923), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10371 ( .A1(n7922), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7969) );
  OAI21_X1 U10372 ( .B1(n7966), .B2(P1_REG3_REG_6__SCAN_IN), .A(n7993), .ZN(
        n11228) );
  OR2_X1 U10373 ( .A1(n8267), .A2(n11228), .ZN(n7968) );
  NAND2_X1 U10374 ( .A1(n6687), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7967) );
  NAND4_X1 U10375 ( .A1(n7970), .A2(n7969), .A3(n7968), .A4(n7967), .ZN(n14036) );
  XNOR2_X1 U10376 ( .A(n12052), .B(n14036), .ZN(n12207) );
  INV_X1 U10377 ( .A(n12207), .ZN(n10681) );
  XNOR2_X1 U10378 ( .A(n7972), .B(n7971), .ZN(n9827) );
  NAND2_X1 U10379 ( .A1(n9827), .A2(n11804), .ZN(n7979) );
  OAI21_X1 U10380 ( .B1(n7973), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7974) );
  MUX2_X1 U10381 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7974), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n7977) );
  AOI22_X1 U10382 ( .A1(n8162), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9985), .B2(
        n10144), .ZN(n7978) );
  INV_X1 U10383 ( .A(n14846), .ZN(n12060) );
  NAND2_X1 U10384 ( .A1(n8345), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7986) );
  INV_X1 U10385 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7980) );
  OR2_X1 U10386 ( .A1(n8217), .A2(n7980), .ZN(n7985) );
  INV_X1 U10387 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7981) );
  XNOR2_X1 U10388 ( .A(n7993), .B(n7981), .ZN(n11097) );
  OR2_X1 U10389 ( .A1(n8282), .A2(n11097), .ZN(n7984) );
  INV_X1 U10390 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7982) );
  OR2_X1 U10391 ( .A1(n6899), .A2(n7982), .ZN(n7983) );
  XNOR2_X1 U10392 ( .A(n12060), .B(n14035), .ZN(n12208) );
  INV_X1 U10393 ( .A(n12208), .ZN(n11087) );
  NAND2_X1 U10394 ( .A1(n14846), .A2(n12059), .ZN(n7987) );
  XNOR2_X1 U10395 ( .A(n7989), .B(n7988), .ZN(n9832) );
  NAND2_X1 U10396 ( .A1(n9832), .A2(n11804), .ZN(n7992) );
  OR2_X1 U10397 ( .A1(n7976), .A2(n8290), .ZN(n7990) );
  XNOR2_X1 U10398 ( .A(n7990), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U10399 ( .A1(n8162), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9985), .B2(
        n10437), .ZN(n7991) );
  NAND2_X1 U10400 ( .A1(n8345), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U10401 ( .A1(n7923), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7998) );
  INV_X1 U10402 ( .A(n7993), .ZN(n7994) );
  AOI21_X1 U10403 ( .B1(n7994), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n7995) );
  OR2_X1 U10404 ( .A1(n7995), .A2(n8006), .ZN(n11200) );
  OR2_X1 U10405 ( .A1(n8282), .A2(n11200), .ZN(n7997) );
  NAND2_X1 U10406 ( .A1(n7922), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7996) );
  NAND4_X1 U10407 ( .A1(n7999), .A2(n7998), .A3(n7997), .A4(n7996), .ZN(n14034) );
  XNOR2_X1 U10408 ( .A(n12063), .B(n14034), .ZN(n12210) );
  INV_X1 U10409 ( .A(n12210), .ZN(n10870) );
  OR2_X1 U10410 ( .A1(n12063), .A2(n14034), .ZN(n8000) );
  NAND2_X1 U10411 ( .A1(n7976), .A2(n8003), .ZN(n8098) );
  NAND2_X1 U10412 ( .A1(n8098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8015) );
  XNOR2_X1 U10413 ( .A(n8015), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U10414 ( .A1(n8162), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9985), .B2(
        n10732), .ZN(n8004) );
  NAND2_X1 U10415 ( .A1(n8345), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8011) );
  INV_X1 U10416 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8005) );
  OR2_X1 U10417 ( .A1(n8217), .A2(n8005), .ZN(n8010) );
  OR2_X1 U10418 ( .A1(n8006), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U10419 ( .A1(n8031), .A2(n8007), .ZN(n11033) );
  OR2_X1 U10420 ( .A1(n8282), .A2(n11033), .ZN(n8009) );
  INV_X1 U10421 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10429) );
  OR2_X1 U10422 ( .A1(n6899), .A2(n10429), .ZN(n8008) );
  XNOR2_X1 U10423 ( .A(n12070), .B(n12069), .ZN(n12212) );
  NAND2_X1 U10424 ( .A1(n12068), .A2(n12069), .ZN(n8012) );
  NAND2_X1 U10425 ( .A1(n8015), .A2(n15553), .ZN(n8024) );
  NAND2_X1 U10426 ( .A1(n8024), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8016) );
  XNOR2_X1 U10427 ( .A(n8016), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11174) );
  AOI22_X1 U10428 ( .A1(n8162), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9985), 
        .B2(n11174), .ZN(n8017) );
  NAND2_X1 U10429 ( .A1(n6943), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U10430 ( .A1(n7922), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U10431 ( .A1(n8345), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8019) );
  XNOR2_X1 U10432 ( .A(n8031), .B(n8030), .ZN(n11771) );
  OR2_X1 U10433 ( .A1(n8282), .A2(n11771), .ZN(n8018) );
  NAND4_X1 U10434 ( .A1(n8021), .A2(n8020), .A3(n8019), .A4(n8018), .ZN(n14032) );
  INV_X1 U10435 ( .A(n14032), .ZN(n11765) );
  NAND2_X1 U10436 ( .A1(n8025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8060) );
  INV_X1 U10437 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n15541) );
  OR2_X1 U10438 ( .A1(n8060), .A2(n15541), .ZN(n8026) );
  NAND2_X1 U10439 ( .A1(n8060), .A2(n15541), .ZN(n8042) );
  AOI22_X1 U10440 ( .A1(n8162), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9985), 
        .B2(n11176), .ZN(n8027) );
  NAND2_X1 U10441 ( .A1(n8345), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10442 ( .A1(n6943), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8035) );
  OAI21_X1 U10443 ( .B1(n8031), .B2(n8030), .A(n8029), .ZN(n8032) );
  NAND2_X1 U10444 ( .A1(n8032), .A2(n8047), .ZN(n11792) );
  OR2_X1 U10445 ( .A1(n8282), .A2(n11792), .ZN(n8034) );
  NAND2_X1 U10446 ( .A1(n7922), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8033) );
  NAND4_X1 U10447 ( .A1(n8036), .A2(n8035), .A3(n8034), .A4(n8033), .ZN(n14031) );
  INV_X1 U10448 ( .A(n12215), .ZN(n11190) );
  OR2_X1 U10449 ( .A1(n12080), .A2(n14031), .ZN(n8037) );
  OR2_X1 U10450 ( .A1(n8039), .A2(n8038), .ZN(n8040) );
  NAND2_X1 U10451 ( .A1(n8041), .A2(n8040), .ZN(n9918) );
  NAND2_X1 U10452 ( .A1(n9918), .A2(n7941), .ZN(n8045) );
  NAND2_X1 U10453 ( .A1(n8042), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8043) );
  XNOR2_X1 U10454 ( .A(n8043), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14058) );
  AOI22_X1 U10455 ( .A1(n8162), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9985), 
        .B2(n14058), .ZN(n8044) );
  NAND2_X1 U10456 ( .A1(n7923), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8053) );
  NAND2_X1 U10457 ( .A1(n6687), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8052) );
  INV_X1 U10458 ( .A(n8064), .ZN(n8049) );
  NAND2_X1 U10459 ( .A1(n8047), .A2(n8046), .ZN(n8048) );
  NAND2_X1 U10460 ( .A1(n8049), .A2(n8048), .ZN(n13895) );
  OR2_X1 U10461 ( .A1(n8282), .A2(n13895), .ZN(n8051) );
  NAND2_X1 U10462 ( .A1(n7922), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8050) );
  NAND4_X1 U10463 ( .A1(n8053), .A2(n8052), .A3(n8051), .A4(n8050), .ZN(n14029) );
  INV_X1 U10464 ( .A(n14029), .ZN(n12244) );
  XNOR2_X1 U10465 ( .A(n12246), .B(n12244), .ZN(n12214) );
  OR2_X1 U10466 ( .A1(n12246), .A2(n14029), .ZN(n8054) );
  XNOR2_X1 U10467 ( .A(n8055), .B(n15723), .ZN(n8056) );
  XNOR2_X1 U10468 ( .A(n8057), .B(n8056), .ZN(n10012) );
  NAND2_X1 U10469 ( .A1(n10012), .A2(n7941), .ZN(n8063) );
  OR2_X1 U10470 ( .A1(n8058), .A2(n8290), .ZN(n8059) );
  NAND2_X1 U10471 ( .A1(n8060), .A2(n8059), .ZN(n8073) );
  XNOR2_X1 U10472 ( .A(n8073), .B(n8061), .ZN(n14754) );
  AOI22_X1 U10473 ( .A1(n8162), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9985), 
        .B2(n14754), .ZN(n8062) );
  NAND2_X1 U10474 ( .A1(n8345), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U10475 ( .A1(n6943), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8068) );
  OR2_X1 U10476 ( .A1(n8064), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10477 ( .A1(n8078), .A2(n8065), .ZN(n13962) );
  OR2_X1 U10478 ( .A1(n8282), .A2(n13962), .ZN(n8067) );
  NAND2_X1 U10479 ( .A1(n7922), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8066) );
  NAND4_X1 U10480 ( .A1(n8069), .A2(n8068), .A3(n8067), .A4(n8066), .ZN(n14028) );
  XNOR2_X1 U10481 ( .A(n13964), .B(n14028), .ZN(n12216) );
  OR2_X1 U10482 ( .A1(n13964), .A2(n14028), .ZN(n8070) );
  XNOR2_X1 U10483 ( .A(n8089), .B(n15542), .ZN(n8086) );
  XNOR2_X1 U10484 ( .A(n8086), .B(n8072), .ZN(n10244) );
  NAND2_X1 U10485 ( .A1(n10244), .A2(n7941), .ZN(n8076) );
  OAI21_X1 U10486 ( .B1(n8073), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8074) );
  XNOR2_X1 U10487 ( .A(n8074), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14060) );
  AOI22_X1 U10488 ( .A1(n8162), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n14060), 
        .B2(n9985), .ZN(n8075) );
  NAND2_X1 U10489 ( .A1(n8345), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8083) );
  INV_X1 U10490 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14047) );
  OR2_X1 U10491 ( .A1(n8217), .A2(n14047), .ZN(n8082) );
  NAND2_X1 U10492 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  NAND2_X1 U10493 ( .A1(n8108), .A2(n8079), .ZN(n13857) );
  OR2_X1 U10494 ( .A1(n8267), .A2(n13857), .ZN(n8081) );
  INV_X1 U10495 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14056) );
  OR2_X1 U10496 ( .A1(n6899), .A2(n14056), .ZN(n8080) );
  OR2_X1 U10497 ( .A1(n14681), .A2(n13959), .ZN(n12096) );
  NAND2_X1 U10498 ( .A1(n14681), .A2(n13959), .ZN(n12095) );
  INV_X1 U10499 ( .A(n13959), .ZN(n14027) );
  NAND2_X1 U10500 ( .A1(n14681), .A2(n14027), .ZN(n8085) );
  INV_X1 U10501 ( .A(n8086), .ZN(n8088) );
  NAND2_X1 U10502 ( .A1(n8088), .A2(n8087), .ZN(n8091) );
  NAND2_X1 U10503 ( .A1(n8089), .A2(n15542), .ZN(n8090) );
  NAND2_X1 U10504 ( .A1(n8091), .A2(n8090), .ZN(n8094) );
  XNOR2_X1 U10505 ( .A(n8092), .B(n9852), .ZN(n8093) );
  NAND2_X1 U10506 ( .A1(n10334), .A2(n7941), .ZN(n8106) );
  NOR2_X1 U10507 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8096) );
  NAND4_X1 U10508 ( .A1(n8058), .A2(n8096), .A3(n8095), .A4(n15539), .ZN(n8097) );
  OR2_X1 U10509 ( .A1(n8098), .A2(n8097), .ZN(n8100) );
  NAND2_X1 U10510 ( .A1(n8100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8099) );
  MUX2_X1 U10511 ( .A(n8099), .B(P1_IR_REG_31__SCAN_IN), .S(n8101), .Z(n8103)
         );
  INV_X1 U10512 ( .A(n8100), .ZN(n8102) );
  NAND2_X1 U10513 ( .A1(n8102), .A2(n8101), .ZN(n8119) );
  NAND2_X1 U10514 ( .A1(n8103), .A2(n8119), .ZN(n14780) );
  INV_X1 U10515 ( .A(n14780), .ZN(n8104) );
  AOI22_X1 U10516 ( .A1(n8162), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9985), 
        .B2(n8104), .ZN(n8105) );
  NAND2_X1 U10517 ( .A1(n6687), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8113) );
  INV_X1 U10518 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11510) );
  OR2_X1 U10519 ( .A1(n8217), .A2(n11510), .ZN(n8112) );
  AND2_X1 U10520 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  OR2_X1 U10521 ( .A1(n8109), .A2(n8123), .ZN(n14009) );
  OR2_X1 U10522 ( .A1(n8282), .A2(n14009), .ZN(n8111) );
  INV_X1 U10523 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14772) );
  OR2_X1 U10524 ( .A1(n6899), .A2(n14772), .ZN(n8110) );
  NAND2_X1 U10525 ( .A1(n14421), .A2(n14315), .ZN(n12101) );
  INV_X1 U10526 ( .A(n14315), .ZN(n14026) );
  OR2_X1 U10527 ( .A1(n14421), .A2(n14026), .ZN(n8115) );
  XNOR2_X1 U10528 ( .A(n8118), .B(n8117), .ZN(n10241) );
  NAND2_X1 U10529 ( .A1(n10241), .A2(n7941), .ZN(n8122) );
  NAND2_X1 U10530 ( .A1(n8119), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8120) );
  XNOR2_X1 U10531 ( .A(n8120), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14795) );
  AOI22_X1 U10532 ( .A1(n8162), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9985), 
        .B2(n14795), .ZN(n8121) );
  NAND2_X2 U10533 ( .A1(n8122), .A2(n8121), .ZN(n14413) );
  NOR2_X1 U10534 ( .A1(n8123), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8124) );
  OR2_X1 U10535 ( .A1(n8137), .A2(n8124), .ZN(n14322) );
  OR2_X1 U10536 ( .A1(n14322), .A2(n8282), .ZN(n8128) );
  NAND2_X1 U10537 ( .A1(n6687), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U10538 ( .A1(n7923), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U10539 ( .A1(n7922), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8125) );
  NAND4_X1 U10540 ( .A1(n8128), .A2(n8127), .A3(n8126), .A4(n8125), .ZN(n14025) );
  XNOR2_X1 U10541 ( .A(n14413), .B(n14304), .ZN(n14327) );
  OR2_X1 U10542 ( .A1(n14413), .A2(n14025), .ZN(n8129) );
  XNOR2_X1 U10543 ( .A(n8130), .B(SI_17_), .ZN(n8131) );
  XNOR2_X1 U10544 ( .A(n8132), .B(n8131), .ZN(n10299) );
  NAND2_X1 U10545 ( .A1(n10299), .A2(n7941), .ZN(n8136) );
  NAND2_X1 U10546 ( .A1(n8133), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8134) );
  XNOR2_X1 U10547 ( .A(n8134), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U10548 ( .A1(n8162), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9985), 
        .B2(n14063), .ZN(n8135) );
  NAND2_X1 U10549 ( .A1(n6687), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8143) );
  OR2_X1 U10550 ( .A1(n8137), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8138) );
  AND2_X1 U10551 ( .A1(n8154), .A2(n8138), .ZN(n14298) );
  NAND2_X1 U10552 ( .A1(n14298), .A2(n8195), .ZN(n8142) );
  INV_X1 U10553 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8139) );
  OR2_X1 U10554 ( .A1(n8217), .A2(n8139), .ZN(n8141) );
  NAND2_X1 U10555 ( .A1(n7922), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8140) );
  NAND4_X1 U10556 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n14024) );
  NAND2_X1 U10557 ( .A1(n14409), .A2(n14024), .ZN(n8321) );
  XNOR2_X1 U10558 ( .A(n8146), .B(n8145), .ZN(n10776) );
  NAND2_X1 U10559 ( .A1(n10776), .A2(n7941), .ZN(n8150) );
  NAND2_X1 U10560 ( .A1(n8161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8147) );
  XNOR2_X1 U10561 ( .A(n8147), .B(n7754), .ZN(n14827) );
  INV_X1 U10562 ( .A(n14827), .ZN(n8148) );
  AOI22_X1 U10563 ( .A1(n8162), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9985), 
        .B2(n8148), .ZN(n8149) );
  NAND2_X1 U10564 ( .A1(n6687), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8152) );
  INV_X1 U10565 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14821) );
  OR2_X1 U10566 ( .A1(n8217), .A2(n14821), .ZN(n8151) );
  AND2_X1 U10567 ( .A1(n8152), .A2(n8151), .ZN(n8158) );
  NAND2_X1 U10568 ( .A1(n8154), .A2(n8153), .ZN(n8155) );
  NAND2_X1 U10569 ( .A1(n8166), .A2(n8155), .ZN(n14286) );
  OR2_X1 U10570 ( .A1(n14286), .A2(n8282), .ZN(n8157) );
  INV_X1 U10571 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14816) );
  OR2_X1 U10572 ( .A1(n6899), .A2(n14816), .ZN(n8156) );
  AND2_X1 U10573 ( .A1(n14290), .A2(n14023), .ZN(n12128) );
  OR2_X1 U10574 ( .A1(n14290), .A2(n14023), .ZN(n12127) );
  OAI21_X2 U10575 ( .B1(n14276), .B2(n12128), .A(n12127), .ZN(n14258) );
  XNOR2_X1 U10576 ( .A(n8160), .B(n8159), .ZN(n10906) );
  NAND2_X1 U10577 ( .A1(n10906), .A2(n7941), .ZN(n8164) );
  AOI22_X1 U10578 ( .A1(n8162), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14287), 
        .B2(n9985), .ZN(n8163) );
  NAND2_X1 U10579 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  NAND2_X1 U10580 ( .A1(n8175), .A2(n8167), .ZN(n14266) );
  AOI22_X1 U10581 ( .A1(n7922), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n7923), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10582 ( .A1(n8345), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8168) );
  OAI211_X1 U10583 ( .C1(n14266), .C2(n8282), .A(n8169), .B(n8168), .ZN(n14237) );
  INV_X1 U10584 ( .A(n14237), .ZN(n14279) );
  OR2_X1 U10585 ( .A1(n14265), .A2(n14279), .ZN(n12132) );
  NAND2_X1 U10586 ( .A1(n14265), .A2(n14279), .ZN(n12133) );
  NAND2_X1 U10587 ( .A1(n12132), .A2(n12133), .ZN(n14262) );
  NAND2_X1 U10588 ( .A1(n14258), .A2(n14262), .ZN(n8171) );
  OR2_X1 U10589 ( .A1(n14265), .A2(n14237), .ZN(n8170) );
  NAND2_X1 U10590 ( .A1(n11256), .A2(n11804), .ZN(n8173) );
  INV_X1 U10591 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11257) );
  OR2_X1 U10592 ( .A1(n7930), .A2(n11257), .ZN(n8172) );
  AND2_X1 U10593 ( .A1(n8175), .A2(n8174), .ZN(n8176) );
  OR2_X1 U10594 ( .A1(n8176), .A2(n8192), .ZN(n13953) );
  INV_X1 U10595 ( .A(n13953), .ZN(n14243) );
  INV_X1 U10596 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14393) );
  NAND2_X1 U10597 ( .A1(n6943), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U10598 ( .A1(n6687), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8177) );
  OAI211_X1 U10599 ( .C1(n14393), .C2(n6899), .A(n8178), .B(n8177), .ZN(n8179)
         );
  AOI21_X1 U10600 ( .B1(n14243), .B2(n8195), .A(n8179), .ZN(n14396) );
  INV_X1 U10601 ( .A(n14396), .ZN(n14269) );
  XNOR2_X1 U10602 ( .A(n14251), .B(n14269), .ZN(n14247) );
  OR2_X1 U10603 ( .A1(n6897), .A2(n14396), .ZN(n8180) );
  INV_X1 U10604 ( .A(n8181), .ZN(n8183) );
  NAND2_X1 U10605 ( .A1(n8183), .A2(n8182), .ZN(n8186) );
  OR2_X1 U10606 ( .A1(n8184), .A2(n10454), .ZN(n8185) );
  XNOR2_X1 U10607 ( .A(n8187), .B(SI_21_), .ZN(n8188) );
  NAND2_X1 U10608 ( .A1(n11341), .A2(n11804), .ZN(n8191) );
  INV_X1 U10609 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11345) );
  OR2_X1 U10610 ( .A1(n7930), .A2(n11345), .ZN(n8190) );
  NAND2_X2 U10611 ( .A1(n8191), .A2(n8190), .ZN(n14386) );
  OR2_X1 U10612 ( .A1(n8192), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8194) );
  AND2_X1 U10613 ( .A1(n8194), .A2(n8193), .ZN(n14229) );
  NAND2_X1 U10614 ( .A1(n14229), .A2(n8195), .ZN(n8201) );
  INV_X1 U10615 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10616 ( .A1(n7923), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10617 ( .A1(n8345), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8196) );
  OAI211_X1 U10618 ( .C1(n8198), .C2(n6899), .A(n8197), .B(n8196), .ZN(n8199)
         );
  INV_X1 U10619 ( .A(n8199), .ZN(n8200) );
  NAND2_X1 U10620 ( .A1(n8201), .A2(n8200), .ZN(n14240) );
  INV_X1 U10621 ( .A(n14240), .ZN(n8326) );
  XNOR2_X1 U10622 ( .A(n14386), .B(n8326), .ZN(n14225) );
  INV_X1 U10623 ( .A(n14225), .ZN(n8202) );
  NAND2_X1 U10624 ( .A1(n9443), .A2(n9766), .ZN(n8203) );
  NAND2_X1 U10625 ( .A1(n6687), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U10626 ( .A1(n7923), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8209) );
  OAI21_X1 U10627 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8206), .A(n8205), .ZN(
        n14214) );
  OR2_X1 U10628 ( .A1(n8282), .A2(n14214), .ZN(n8208) );
  NAND2_X1 U10629 ( .A1(n7922), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8207) );
  NAND4_X1 U10630 ( .A1(n8210), .A2(n8209), .A3(n8208), .A4(n8207), .ZN(n14224) );
  NAND2_X1 U10631 ( .A1(n14210), .A2(n14209), .ZN(n14208) );
  OR2_X1 U10632 ( .A1(n14211), .A2(n14224), .ZN(n8211) );
  XNOR2_X1 U10633 ( .A(n8212), .B(SI_23_), .ZN(n8213) );
  XNOR2_X1 U10634 ( .A(n8214), .B(n8213), .ZN(n11432) );
  NAND2_X1 U10635 ( .A1(n11432), .A2(n11804), .ZN(n8216) );
  INV_X1 U10636 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11434) );
  OR2_X1 U10637 ( .A1(n7930), .A2(n11434), .ZN(n8215) );
  NAND2_X1 U10638 ( .A1(n8345), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8223) );
  INV_X1 U10639 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14197) );
  OR2_X1 U10640 ( .A1(n8217), .A2(n14197), .ZN(n8222) );
  OAI21_X1 U10641 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8218), .A(n8231), .ZN(
        n14199) );
  OR2_X1 U10642 ( .A1(n8282), .A2(n14199), .ZN(n8221) );
  INV_X1 U10643 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8219) );
  OR2_X1 U10644 ( .A1(n6899), .A2(n8219), .ZN(n8220) );
  NAND2_X1 U10645 ( .A1(n14202), .A2(n14179), .ZN(n8328) );
  OR2_X1 U10646 ( .A1(n14202), .A2(n14179), .ZN(n8224) );
  NAND2_X1 U10647 ( .A1(n8328), .A2(n8224), .ZN(n14192) );
  NAND2_X2 U10648 ( .A1(n6722), .A2(n14192), .ZN(n14191) );
  OR2_X1 U10649 ( .A1(n14372), .A2(n14179), .ZN(n8225) );
  NAND2_X1 U10650 ( .A1(n11635), .A2(n11804), .ZN(n8229) );
  OR2_X1 U10651 ( .A1(n7930), .A2(n7602), .ZN(n8228) );
  NAND2_X1 U10652 ( .A1(n6687), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U10653 ( .A1(n6943), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8235) );
  INV_X1 U10654 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8230) );
  NAND2_X1 U10655 ( .A1(n8231), .A2(n8230), .ZN(n8232) );
  NAND2_X1 U10656 ( .A1(n8242), .A2(n8232), .ZN(n13942) );
  OR2_X1 U10657 ( .A1(n8267), .A2(n13942), .ZN(n8234) );
  NAND2_X1 U10658 ( .A1(n7922), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8233) );
  NAND4_X1 U10659 ( .A1(n8236), .A2(n8235), .A3(n8234), .A4(n8233), .ZN(n14021) );
  XNOR2_X1 U10660 ( .A(n14185), .B(n14021), .ZN(n14177) );
  OR2_X1 U10661 ( .A1(n14185), .A2(n14021), .ZN(n8237) );
  XNOR2_X1 U10662 ( .A(n8239), .B(n8238), .ZN(n11821) );
  NAND2_X1 U10663 ( .A1(n11821), .A2(n11804), .ZN(n8241) );
  OR2_X1 U10664 ( .A1(n7930), .A2(n11822), .ZN(n8240) );
  NAND2_X1 U10665 ( .A1(n6687), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8247) );
  NAND2_X1 U10666 ( .A1(n7923), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8246) );
  INV_X1 U10667 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U10668 ( .A1(n8242), .A2(n13909), .ZN(n8243) );
  NAND2_X1 U10669 ( .A1(n8254), .A2(n8243), .ZN(n14162) );
  OR2_X1 U10670 ( .A1(n8282), .A2(n14162), .ZN(n8245) );
  NAND2_X1 U10671 ( .A1(n7922), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8244) );
  NAND4_X1 U10672 ( .A1(n8247), .A2(n8246), .A3(n8245), .A4(n8244), .ZN(n14020) );
  XNOR2_X1 U10673 ( .A(n14167), .B(n14020), .ZN(n14157) );
  NAND2_X1 U10674 ( .A1(n14167), .A2(n14020), .ZN(n8248) );
  XNOR2_X1 U10675 ( .A(n8249), .B(SI_26_), .ZN(n8250) );
  NAND2_X1 U10676 ( .A1(n13832), .A2(n11804), .ZN(n8253) );
  OR2_X1 U10677 ( .A1(n7930), .A2(n14491), .ZN(n8252) );
  NAND2_X1 U10678 ( .A1(n6687), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10679 ( .A1(n7923), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8258) );
  INV_X1 U10680 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13995) );
  NAND2_X1 U10681 ( .A1(n8254), .A2(n13995), .ZN(n8255) );
  NAND2_X1 U10682 ( .A1(n8266), .A2(n8255), .ZN(n14148) );
  OR2_X1 U10683 ( .A1(n8282), .A2(n14148), .ZN(n8257) );
  NAND2_X1 U10684 ( .A1(n7922), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8256) );
  NAND4_X1 U10685 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n14019) );
  XNOR2_X1 U10686 ( .A(n13987), .B(n14019), .ZN(n14144) );
  INV_X1 U10687 ( .A(n14144), .ZN(n14142) );
  NAND2_X1 U10688 ( .A1(n6884), .A2(n14019), .ZN(n8260) );
  XNOR2_X1 U10689 ( .A(n8261), .B(SI_27_), .ZN(n8262) );
  OR2_X1 U10690 ( .A1(n7930), .A2(n14487), .ZN(n8264) );
  NAND2_X1 U10691 ( .A1(n8345), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U10692 ( .A1(n6943), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8270) );
  XNOR2_X1 U10693 ( .A(n8266), .B(n13847), .ZN(n13844) );
  OR2_X1 U10694 ( .A1(n8267), .A2(n13844), .ZN(n8269) );
  NAND2_X1 U10695 ( .A1(n7922), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8268) );
  NAND4_X1 U10696 ( .A1(n8271), .A2(n8270), .A3(n8269), .A4(n8268), .ZN(n14104) );
  INV_X1 U10697 ( .A(n14104), .ZN(n8272) );
  NAND2_X1 U10698 ( .A1(n14133), .A2(n8272), .ZN(n8333) );
  OR2_X1 U10699 ( .A1(n14133), .A2(n14104), .ZN(n8274) );
  INV_X1 U10700 ( .A(n14018), .ZN(n8275) );
  NAND2_X1 U10701 ( .A1(n14435), .A2(n8275), .ZN(n8334) );
  OR2_X1 U10702 ( .A1(n14435), .A2(n8275), .ZN(n8276) );
  NAND2_X1 U10703 ( .A1(n8334), .A2(n8276), .ZN(n12223) );
  INV_X1 U10704 ( .A(n12223), .ZN(n14107) );
  MUX2_X1 U10705 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n9773), .Z(n9537) );
  INV_X1 U10706 ( .A(SI_29_), .ZN(n13129) );
  XNOR2_X1 U10707 ( .A(n9537), .B(n13129), .ZN(n9535) );
  NAND2_X1 U10708 ( .A1(n13823), .A2(n11804), .ZN(n8281) );
  INV_X1 U10709 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14480) );
  OR2_X1 U10710 ( .A1(n7930), .A2(n14480), .ZN(n8280) );
  NAND2_X1 U10711 ( .A1(n6687), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8286) );
  NAND2_X1 U10712 ( .A1(n6943), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8285) );
  OR2_X1 U10713 ( .A1(n8282), .A2(n14089), .ZN(n8284) );
  NAND2_X1 U10714 ( .A1(n7922), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8283) );
  NAND4_X1 U10715 ( .A1(n8286), .A2(n8285), .A3(n8284), .A4(n8283), .ZN(n14105) );
  OR2_X1 U10716 ( .A1(n8293), .A2(n8290), .ZN(n8291) );
  MUX2_X1 U10717 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8291), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8294) );
  INV_X1 U10718 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U10719 ( .A1(n8295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10720 ( .A1(n6772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8298) );
  NAND2_X2 U10721 ( .A1(n12012), .A2(n12016), .ZN(n12376) );
  OAI21_X1 U10722 ( .B1(n12012), .B2(n12016), .A(n12376), .ZN(n10885) );
  OR2_X1 U10723 ( .A1(n10885), .A2(n14287), .ZN(n14283) );
  AND2_X1 U10724 ( .A1(n12188), .A2(n14287), .ZN(n8299) );
  NAND2_X1 U10725 ( .A1(n12189), .A2(n8299), .ZN(n10623) );
  NAND2_X1 U10726 ( .A1(n14283), .A2(n10623), .ZN(n14855) );
  INV_X1 U10727 ( .A(n12204), .ZN(n8304) );
  NAND2_X1 U10728 ( .A1(n12025), .A2(n12019), .ZN(n8300) );
  AND2_X1 U10729 ( .A1(n8300), .A2(n12023), .ZN(n10616) );
  NAND2_X1 U10730 ( .A1(n10616), .A2(n12201), .ZN(n8301) );
  NAND2_X1 U10731 ( .A1(n12021), .A2(n12022), .ZN(n12030) );
  NAND2_X1 U10732 ( .A1(n8301), .A2(n12030), .ZN(n10515) );
  NAND2_X1 U10733 ( .A1(n10515), .A2(n12202), .ZN(n8303) );
  NAND2_X1 U10734 ( .A1(n10788), .A2(n12033), .ZN(n8302) );
  NAND2_X1 U10735 ( .A1(n8303), .A2(n8302), .ZN(n10552) );
  NAND2_X1 U10736 ( .A1(n8304), .A2(n10552), .ZN(n8306) );
  INV_X1 U10737 ( .A(n12038), .ZN(n12041) );
  NAND2_X1 U10738 ( .A1(n12039), .A2(n12041), .ZN(n8305) );
  NAND2_X1 U10739 ( .A1(n8306), .A2(n8305), .ZN(n11039) );
  INV_X1 U10740 ( .A(n12205), .ZN(n8307) );
  NAND2_X1 U10741 ( .A1(n11039), .A2(n8307), .ZN(n8309) );
  NAND2_X1 U10742 ( .A1(n11408), .A2(n12047), .ZN(n8308) );
  NAND2_X1 U10743 ( .A1(n8309), .A2(n8308), .ZN(n10679) );
  INV_X1 U10744 ( .A(n14036), .ZN(n11405) );
  NAND2_X1 U10745 ( .A1(n12052), .A2(n11405), .ZN(n8310) );
  NOR2_X1 U10746 ( .A1(n14846), .A2(n14035), .ZN(n8311) );
  NAND2_X1 U10747 ( .A1(n14846), .A2(n14035), .ZN(n8312) );
  NAND2_X1 U10748 ( .A1(n10873), .A2(n12210), .ZN(n8314) );
  INV_X1 U10749 ( .A(n14034), .ZN(n11754) );
  OR2_X1 U10750 ( .A1(n12063), .A2(n11754), .ZN(n8313) );
  NAND2_X1 U10751 ( .A1(n8314), .A2(n8313), .ZN(n11028) );
  INV_X1 U10752 ( .A(n12069), .ZN(n14033) );
  OR2_X1 U10753 ( .A1(n12068), .A2(n14033), .ZN(n8315) );
  INV_X1 U10754 ( .A(n14031), .ZN(n11783) );
  OR2_X1 U10755 ( .A1(n12080), .A2(n11783), .ZN(n8316) );
  INV_X1 U10756 ( .A(n12214), .ZN(n11420) );
  NAND2_X1 U10757 ( .A1(n11451), .A2(n12216), .ZN(n8318) );
  INV_X1 U10758 ( .A(n14028), .ZN(n12256) );
  OR2_X1 U10759 ( .A1(n13964), .A2(n12256), .ZN(n8317) );
  NAND2_X1 U10760 ( .A1(n8318), .A2(n8317), .ZN(n11468) );
  INV_X1 U10761 ( .A(n12218), .ZN(n8319) );
  NAND2_X1 U10762 ( .A1(n14413), .A2(n14304), .ZN(n8320) );
  NAND2_X1 U10763 ( .A1(n8322), .A2(n8321), .ZN(n14294) );
  INV_X1 U10764 ( .A(n14294), .ZN(n14302) );
  NAND2_X1 U10765 ( .A1(n14301), .A2(n14024), .ZN(n8323) );
  XNOR2_X1 U10766 ( .A(n14290), .B(n14023), .ZN(n14278) );
  OR2_X1 U10767 ( .A1(n8326), .A2(n14386), .ZN(n8327) );
  INV_X1 U10768 ( .A(n14224), .ZN(n12321) );
  NAND2_X1 U10769 ( .A1(n14193), .A2(n8328), .ZN(n14178) );
  NAND2_X1 U10770 ( .A1(n14178), .A2(n14177), .ZN(n14176) );
  INV_X1 U10771 ( .A(n14021), .ZN(n8329) );
  NAND2_X1 U10772 ( .A1(n14185), .A2(n8329), .ZN(n8330) );
  NAND2_X1 U10773 ( .A1(n14176), .A2(n8330), .ZN(n14156) );
  INV_X1 U10774 ( .A(n14020), .ZN(n14180) );
  NAND2_X1 U10775 ( .A1(n14167), .A2(n14180), .ZN(n8331) );
  INV_X1 U10776 ( .A(n14019), .ZN(n8332) );
  NAND2_X1 U10777 ( .A1(n13987), .A2(n8332), .ZN(n14126) );
  NAND2_X1 U10778 ( .A1(n14102), .A2(n14107), .ZN(n14101) );
  NAND2_X1 U10779 ( .A1(n14101), .A2(n8334), .ZN(n8335) );
  NAND2_X1 U10780 ( .A1(n14496), .A2(n14287), .ZN(n8336) );
  NAND2_X1 U10781 ( .A1(n12183), .A2(n12014), .ZN(n12009) );
  INV_X1 U10782 ( .A(n12063), .ZN(n11634) );
  NAND2_X1 U10783 ( .A1(n11095), .A2(n11634), .ZN(n11032) );
  INV_X1 U10784 ( .A(n12080), .ZN(n14694) );
  INV_X1 U10785 ( .A(n12246), .ZN(n13902) );
  INV_X1 U10786 ( .A(n14421), .ZN(n8337) );
  NAND2_X1 U10787 ( .A1(n6897), .A2(n14264), .ZN(n14250) );
  OR2_X1 U10788 ( .A1(n14250), .A2(n14386), .ZN(n14227) );
  OR2_X2 U10789 ( .A1(n6884), .A2(n14160), .ZN(n14146) );
  INV_X1 U10790 ( .A(n12183), .ZN(n12013) );
  AOI21_X1 U10791 ( .B1(n12178), .B2(n14112), .A(n14423), .ZN(n8339) );
  INV_X1 U10792 ( .A(n12178), .ZN(n14097) );
  INV_X1 U10793 ( .A(n8340), .ZN(n10447) );
  NAND2_X1 U10794 ( .A1(n10447), .A2(n14287), .ZN(n8342) );
  NAND2_X1 U10795 ( .A1(n12013), .A2(n12014), .ZN(n12225) );
  INV_X1 U10796 ( .A(n12225), .ZN(n8341) );
  NAND2_X1 U10797 ( .A1(n8341), .A2(n12189), .ZN(n10891) );
  NAND2_X1 U10798 ( .A1(n14496), .A2(n12183), .ZN(n12191) );
  INV_X1 U10799 ( .A(n14483), .ZN(n10268) );
  NOR2_X2 U10800 ( .A1(n12191), .A2(n10268), .ZN(n14239) );
  INV_X1 U10801 ( .A(P1_B_REG_SCAN_IN), .ZN(n8343) );
  OR2_X1 U10802 ( .A1(n14488), .A2(n8343), .ZN(n8344) );
  AND2_X1 U10803 ( .A1(n14239), .A2(n8344), .ZN(n11815) );
  INV_X1 U10804 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10805 ( .A1(n7923), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10806 ( .A1(n8345), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8346) );
  OAI211_X1 U10807 ( .C1(n6899), .C2(n8348), .A(n8347), .B(n8346), .ZN(n14017)
         );
  NAND2_X1 U10808 ( .A1(n11815), .A2(n14017), .ZN(n14090) );
  INV_X1 U10809 ( .A(n12191), .ZN(n9987) );
  NAND2_X1 U10810 ( .A1(n14018), .A2(n14238), .ZN(n14092) );
  OAI211_X1 U10811 ( .C1(n14097), .C2(n14852), .A(n14090), .B(n14092), .ZN(
        n8349) );
  INV_X1 U10812 ( .A(n8352), .ZN(n8354) );
  INV_X1 U10813 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10814 ( .A1(n8354), .A2(n8353), .ZN(n8356) );
  OAI21_X2 U10815 ( .B1(n8356), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U10816 ( .A1(n8375), .A2(P1_B_REG_SCAN_IN), .ZN(n8358) );
  MUX2_X1 U10817 ( .A(n8358), .B(P1_B_REG_SCAN_IN), .S(n8376), .Z(n8361) );
  NAND2_X1 U10818 ( .A1(n8359), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8360) );
  OR2_X1 U10819 ( .A1(n9904), .A2(P1_D_REG_1__SCAN_IN), .ZN(n8362) );
  INV_X1 U10820 ( .A(n8383), .ZN(n14492) );
  NAND2_X1 U10821 ( .A1(n8375), .A2(n14492), .ZN(n9907) );
  NAND2_X1 U10822 ( .A1(n8362), .A2(n9907), .ZN(n10880) );
  NAND2_X1 U10823 ( .A1(n14248), .A2(n14287), .ZN(n10356) );
  NAND2_X1 U10824 ( .A1(n10880), .A2(n10356), .ZN(n8382) );
  NOR4_X1 U10825 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8367) );
  NOR4_X1 U10826 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8366) );
  NOR4_X1 U10827 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8365) );
  NOR4_X1 U10828 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8364) );
  NAND4_X1 U10829 ( .A1(n8367), .A2(n8366), .A3(n8365), .A4(n8364), .ZN(n8373)
         );
  NOR2_X1 U10830 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n8371) );
  NOR4_X1 U10831 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n8370) );
  NOR4_X1 U10832 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8369) );
  NOR4_X1 U10833 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8368) );
  NAND4_X1 U10834 ( .A1(n8371), .A2(n8370), .A3(n8369), .A4(n8368), .ZN(n8372)
         );
  NOR2_X1 U10835 ( .A1(n8373), .A2(n8372), .ZN(n8374) );
  INV_X1 U10836 ( .A(n8375), .ZN(n8378) );
  NAND2_X1 U10837 ( .A1(n8352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8379) );
  XNOR2_X1 U10838 ( .A(n8379), .B(n8353), .ZN(n9986) );
  NAND2_X1 U10839 ( .A1(n12188), .A2(n14071), .ZN(n8380) );
  NAND2_X1 U10840 ( .A1(n9987), .A2(n8380), .ZN(n12236) );
  AND2_X1 U10841 ( .A1(n12237), .A2(n12236), .ZN(n8381) );
  NAND2_X1 U10842 ( .A1(n10348), .A2(n8381), .ZN(n10882) );
  INV_X1 U10843 ( .A(n9904), .ZN(n8384) );
  INV_X1 U10844 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9906) );
  NOR2_X1 U10845 ( .A1(n8376), .A2(n8383), .ZN(n9905) );
  AND2_X2 U10846 ( .A1(n9671), .A2(n10881), .ZN(n14863) );
  NAND2_X1 U10847 ( .A1(n8551), .A2(n8550), .ZN(n8571) );
  INV_X1 U10848 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n15481) );
  INV_X1 U10849 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8386) );
  INV_X1 U10850 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8388) );
  NOR2_X1 U10851 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_REG3_REG_18__SCAN_IN), 
        .ZN(n8390) );
  INV_X1 U10852 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15658) );
  INV_X1 U10853 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n8393) );
  INV_X1 U10854 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8395) );
  INV_X1 U10855 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15555) );
  INV_X1 U10856 ( .A(n8890), .ZN(n8398) );
  INV_X1 U10857 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n15556) );
  NAND2_X1 U10858 ( .A1(n8398), .A2(n15556), .ZN(n12388) );
  NAND2_X1 U10859 ( .A1(n8890), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U10860 ( .A1(n12388), .A2(n8399), .ZN(n12773) );
  INV_X1 U10861 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13117) );
  INV_X1 U10862 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8407) );
  XNOR2_X2 U10863 ( .A(n8408), .B(n8407), .ZN(n13127) );
  INV_X1 U10864 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8414) );
  NAND2_X4 U10865 ( .A1(n8410), .A2(n13127), .ZN(n10950) );
  NAND2_X1 U10866 ( .A1(n8507), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U10867 ( .A1(n10948), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8412) );
  OAI211_X1 U10868 ( .C1(n10953), .C2(n8414), .A(n8413), .B(n8412), .ZN(n8415)
         );
  INV_X1 U10869 ( .A(n8502), .ZN(n8416) );
  NAND2_X1 U10870 ( .A1(n8491), .A2(n8416), .ZN(n8418) );
  NAND2_X1 U10871 ( .A1(n7662), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8417) );
  INV_X1 U10872 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U10873 ( .A1(n9797), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8419) );
  NAND2_X1 U10874 ( .A1(n9768), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U10875 ( .A1(n9793), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U10876 ( .A1(n9817), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U10877 ( .A1(n9824), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10878 ( .A1(n9821), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U10879 ( .A1(n9831), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U10880 ( .A1(n8433), .A2(n8432), .ZN(n8593) );
  NAND2_X1 U10881 ( .A1(n9835), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10882 ( .A1(n9833), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10883 ( .A1(n9838), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10884 ( .A1(n9840), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10885 ( .A1(n8438), .A2(n8436), .ZN(n8628) );
  INV_X1 U10886 ( .A(n8628), .ZN(n8437) );
  NAND2_X1 U10887 ( .A1(n9842), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8441) );
  INV_X1 U10888 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U10889 ( .A1(n9844), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U10890 ( .A1(n9848), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10891 ( .A1(n9850), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10892 ( .A1(n9919), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10893 ( .A1(n9921), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8444) );
  INV_X1 U10894 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10013) );
  INV_X1 U10895 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U10896 ( .A1(n10245), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8448) );
  INV_X1 U10897 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10297) );
  NAND2_X1 U10898 ( .A1(n10297), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8447) );
  AND2_X1 U10899 ( .A1(n8448), .A2(n8447), .ZN(n8704) );
  INV_X1 U10900 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U10901 ( .A1(n10335), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8450) );
  INV_X1 U10902 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U10903 ( .A1(n10368), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8449) );
  AND2_X1 U10904 ( .A1(n8450), .A2(n8449), .ZN(n8720) );
  INV_X1 U10905 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U10906 ( .A1(n10242), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8452) );
  INV_X1 U10907 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U10908 ( .A1(n10271), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8451) );
  AND2_X1 U10909 ( .A1(n8452), .A2(n8451), .ZN(n8736) );
  NAND2_X1 U10910 ( .A1(n10300), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10911 ( .A1(n10314), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10912 ( .A1(n8455), .A2(n8453), .ZN(n8754) );
  INV_X1 U10913 ( .A(n8754), .ZN(n8454) );
  INV_X1 U10914 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10779) );
  NAND2_X1 U10915 ( .A1(n10779), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8457) );
  INV_X1 U10916 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10777) );
  NAND2_X1 U10917 ( .A1(n10777), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8456) );
  AND2_X1 U10918 ( .A1(n8457), .A2(n8456), .ZN(n8768) );
  NAND2_X1 U10919 ( .A1(n10909), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10920 ( .A1(n10907), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8458) );
  AND2_X1 U10921 ( .A1(n8459), .A2(n8458), .ZN(n8782) );
  NAND2_X1 U10922 ( .A1(n11345), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8463) );
  INV_X1 U10923 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11343) );
  NAND2_X1 U10924 ( .A1(n11343), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8462) );
  AND2_X1 U10925 ( .A1(n8463), .A2(n8462), .ZN(n8811) );
  INV_X1 U10926 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11829) );
  XNOR2_X1 U10927 ( .A(n11829), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8826) );
  XNOR2_X1 U10928 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8837) );
  INV_X1 U10929 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U10930 ( .A1(n8464), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8465) );
  INV_X1 U10931 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11637) );
  NAND2_X1 U10932 ( .A1(n13838), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10933 ( .A1(n11822), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8469) );
  AND2_X1 U10934 ( .A1(n14491), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10935 ( .A1(n13833), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8472) );
  AND2_X1 U10936 ( .A1(n8473), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U10937 ( .A1(n14487), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8475) );
  XNOR2_X1 U10938 ( .A(n8900), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8477) );
  XNOR2_X1 U10939 ( .A(n8899), .B(n8477), .ZN(n11823) );
  XNOR2_X2 U10940 ( .A(n8482), .B(n8481), .ZN(n8927) );
  NAND2_X4 U10941 ( .A1(n8926), .A2(n8927), .ZN(n9692) );
  NAND2_X1 U10942 ( .A1(n11823), .A2(n11840), .ZN(n8484) );
  NAND2_X2 U10943 ( .A1(n9692), .A2(n9773), .ZN(n8517) );
  OR2_X1 U10944 ( .A1(n8517), .A2(n15660), .ZN(n8483) );
  INV_X1 U10945 ( .A(n13035), .ZN(n8897) );
  INV_X1 U10946 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9710) );
  OR2_X1 U10947 ( .A1(n8795), .A2(n9710), .ZN(n8488) );
  INV_X1 U10948 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10509) );
  OR2_X1 U10949 ( .A1(n8905), .A2(n10509), .ZN(n8487) );
  INV_X1 U10950 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9711) );
  OR2_X1 U10951 ( .A1(n10950), .A2(n9711), .ZN(n8486) );
  NAND2_X1 U10952 ( .A1(n10948), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8485) );
  INV_X1 U10953 ( .A(n15312), .ZN(n10280) );
  INV_X1 U10954 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8490) );
  OR2_X1 U10955 ( .A1(n8517), .A2(n9782), .ZN(n8492) );
  XNOR2_X1 U10956 ( .A(n8491), .B(n8502), .ZN(n9781) );
  NAND2_X1 U10957 ( .A1(n8832), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8499) );
  INV_X1 U10958 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9716) );
  OR2_X1 U10959 ( .A1(n10950), .A2(n9716), .ZN(n8498) );
  INV_X1 U10960 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n8493) );
  OR2_X1 U10961 ( .A1(n8905), .A2(n8493), .ZN(n8497) );
  INV_X1 U10962 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8495) );
  OR2_X1 U10963 ( .A1(n8494), .A2(n8495), .ZN(n8496) );
  NAND4_X2 U10964 ( .A1(n8499), .A2(n8498), .A3(n8497), .A4(n8496), .ZN(n10504) );
  OR2_X1 U10965 ( .A1(n8517), .A2(n9808), .ZN(n8504) );
  INV_X1 U10966 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U10967 ( .A1(n8500), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8501) );
  AND2_X1 U10968 ( .A1(n8502), .A2(n8501), .ZN(n9809) );
  OR2_X1 U10969 ( .A1(n8815), .A2(n9809), .ZN(n8503) );
  OAI211_X1 U10970 ( .C1(n9810), .C2(n9692), .A(n8504), .B(n8503), .ZN(n10279)
         );
  NAND2_X1 U10971 ( .A1(n10504), .A2(n10279), .ZN(n15320) );
  NAND2_X1 U10972 ( .A1(n15324), .A2(n15320), .ZN(n8506) );
  NAND2_X1 U10973 ( .A1(n15312), .A2(n15340), .ZN(n8505) );
  NAND2_X1 U10974 ( .A1(n8506), .A2(n8505), .ZN(n15309) );
  NAND2_X1 U10975 ( .A1(n8507), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8513) );
  INV_X1 U10976 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n8508) );
  OR2_X1 U10977 ( .A1(n8905), .A2(n8508), .ZN(n8512) );
  INV_X1 U10978 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9717) );
  OR2_X1 U10979 ( .A1(n8795), .A2(n9717), .ZN(n8511) );
  INV_X1 U10980 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8509) );
  NOR2_X1 U10981 ( .A1(n9678), .A2(n8681), .ZN(n8514) );
  XNOR2_X1 U10982 ( .A(n8516), .B(n8515), .ZN(n9787) );
  OR2_X1 U10983 ( .A1(n8517), .A2(SI_2_), .ZN(n8518) );
  INV_X1 U10984 ( .A(n11853), .ZN(n11012) );
  NAND2_X1 U10985 ( .A1(n11012), .A2(n6682), .ZN(n8520) );
  NAND2_X1 U10986 ( .A1(n10948), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8524) );
  INV_X1 U10987 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11018) );
  OR2_X1 U10988 ( .A1(n10950), .A2(n11018), .ZN(n8523) );
  OR2_X1 U10989 ( .A1(n8905), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8522) );
  INV_X1 U10990 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9723) );
  OR2_X1 U10991 ( .A1(n8795), .A2(n9723), .ZN(n8521) );
  AND4_X2 U10992 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n15314)
         );
  OR2_X1 U10993 ( .A1(n8517), .A2(SI_3_), .ZN(n8531) );
  XNOR2_X1 U10994 ( .A(n8526), .B(n8525), .ZN(n9777) );
  OR2_X1 U10995 ( .A1(n8815), .A2(n9777), .ZN(n8530) );
  NAND2_X1 U10996 ( .A1(n7311), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8527) );
  MUX2_X1 U10997 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8527), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n8528) );
  OR2_X1 U10998 ( .A1(n9692), .A2(n10611), .ZN(n8529) );
  NAND2_X1 U10999 ( .A1(n15314), .A2(n10764), .ZN(n11865) );
  INV_X1 U11000 ( .A(n15314), .ZN(n12623) );
  INV_X1 U11001 ( .A(n10764), .ZN(n11019) );
  NAND2_X1 U11002 ( .A1(n12623), .A2(n11019), .ZN(n11862) );
  NAND2_X1 U11003 ( .A1(n12623), .A2(n10764), .ZN(n8533) );
  NAND2_X1 U11004 ( .A1(n11013), .A2(n8533), .ZN(n11153) );
  NAND2_X1 U11005 ( .A1(n10948), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8538) );
  INV_X1 U11006 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11157) );
  OR2_X1 U11007 ( .A1(n10950), .A2(n11157), .ZN(n8537) );
  AND2_X1 U11008 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8534) );
  NOR2_X1 U11009 ( .A1(n8551), .A2(n8534), .ZN(n10995) );
  OR2_X1 U11010 ( .A1(n8905), .A2(n10995), .ZN(n8536) );
  INV_X1 U11011 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15386) );
  OR2_X1 U11012 ( .A1(n8795), .A2(n15386), .ZN(n8535) );
  OR2_X1 U11013 ( .A1(n8517), .A2(SI_4_), .ZN(n8548) );
  XNOR2_X1 U11014 ( .A(n8540), .B(n8539), .ZN(n9784) );
  OR2_X1 U11015 ( .A1(n8815), .A2(n9784), .ZN(n8547) );
  NAND2_X1 U11016 ( .A1(n8543), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8542) );
  MUX2_X1 U11017 ( .A(n8542), .B(P3_IR_REG_31__SCAN_IN), .S(n8541), .Z(n8545)
         );
  INV_X1 U11018 ( .A(n8561), .ZN(n8544) );
  OR2_X1 U11019 ( .A1(n9692), .A2(n9728), .ZN(n8546) );
  NAND2_X1 U11020 ( .A1(n11317), .A2(n11158), .ZN(n11866) );
  INV_X1 U11021 ( .A(n11317), .ZN(n10023) );
  INV_X1 U11022 ( .A(n11158), .ZN(n10996) );
  NAND2_X1 U11023 ( .A1(n10023), .A2(n10996), .ZN(n11869) );
  NAND2_X1 U11024 ( .A1(n11866), .A2(n11869), .ZN(n11152) );
  NAND2_X1 U11025 ( .A1(n11153), .A2(n11152), .ZN(n11151) );
  NAND2_X1 U11026 ( .A1(n10023), .A2(n11158), .ZN(n8549) );
  NAND2_X1 U11027 ( .A1(n11151), .A2(n8549), .ZN(n11313) );
  INV_X1 U11028 ( .A(n11313), .ZN(n8568) );
  NAND2_X1 U11029 ( .A1(n10948), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8556) );
  INV_X1 U11030 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9734) );
  OR2_X1 U11031 ( .A1(n10950), .A2(n9734), .ZN(n8555) );
  OR2_X1 U11032 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  AND2_X1 U11033 ( .A1(n8571), .A2(n8552), .ZN(n11312) );
  OR2_X1 U11034 ( .A1(n8905), .A2(n11312), .ZN(n8554) );
  INV_X1 U11035 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9733) );
  OR2_X1 U11036 ( .A1(n8795), .A2(n9733), .ZN(n8553) );
  OR2_X1 U11037 ( .A1(n8517), .A2(SI_5_), .ZN(n8566) );
  XNOR2_X1 U11038 ( .A(n8558), .B(n8557), .ZN(n9772) );
  OR2_X1 U11039 ( .A1(n8815), .A2(n9772), .ZN(n8565) );
  NOR2_X1 U11040 ( .A1(n8561), .A2(n8681), .ZN(n8559) );
  MUX2_X1 U11041 ( .A(n8681), .B(n8559), .S(P3_IR_REG_5__SCAN_IN), .Z(n8563)
         );
  NAND2_X1 U11042 ( .A1(n8561), .A2(n8560), .ZN(n8590) );
  INV_X1 U11043 ( .A(n8590), .ZN(n8562) );
  OR2_X1 U11044 ( .A1(n9692), .A2(n10570), .ZN(n8564) );
  NAND2_X1 U11045 ( .A1(n11303), .A2(n11311), .ZN(n11872) );
  INV_X1 U11046 ( .A(n11303), .ZN(n10028) );
  INV_X1 U11047 ( .A(n11311), .ZN(n8569) );
  NAND2_X1 U11048 ( .A1(n10028), .A2(n8569), .ZN(n11867) );
  NAND2_X1 U11049 ( .A1(n11303), .A2(n8569), .ZN(n8570) );
  NAND2_X1 U11050 ( .A1(n10948), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8576) );
  INV_X1 U11051 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15297) );
  OR2_X1 U11052 ( .A1(n10950), .A2(n15297), .ZN(n8575) );
  NAND2_X1 U11053 ( .A1(n8571), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8572) );
  AND2_X1 U11054 ( .A1(n8584), .A2(n8572), .ZN(n15293) );
  OR2_X1 U11055 ( .A1(n8905), .A2(n15293), .ZN(n8574) );
  INV_X1 U11056 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15389) );
  OR2_X1 U11057 ( .A1(n10953), .A2(n15389), .ZN(n8573) );
  AND4_X2 U11058 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n15130)
         );
  NAND2_X1 U11059 ( .A1(n8590), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8578) );
  INV_X1 U11060 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8577) );
  XNOR2_X1 U11061 ( .A(n8578), .B(n8577), .ZN(n9813) );
  INV_X1 U11062 ( .A(SI_6_), .ZN(n9811) );
  OR2_X1 U11063 ( .A1(n8517), .A2(n9811), .ZN(n8582) );
  XNOR2_X1 U11064 ( .A(n9821), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8579) );
  XNOR2_X1 U11065 ( .A(n8580), .B(n8579), .ZN(n9812) );
  OR2_X1 U11066 ( .A1(n8815), .A2(n9812), .ZN(n8581) );
  OAI211_X1 U11067 ( .C1(n9692), .C2(n9813), .A(n8582), .B(n8581), .ZN(n15292)
         );
  NAND2_X1 U11068 ( .A1(n15130), .A2(n15292), .ZN(n11877) );
  INV_X1 U11069 ( .A(n15130), .ZN(n10037) );
  INV_X1 U11070 ( .A(n15292), .ZN(n8583) );
  NAND2_X1 U11071 ( .A1(n10037), .A2(n8583), .ZN(n11874) );
  NAND2_X1 U11072 ( .A1(n10948), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8589) );
  INV_X1 U11073 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9744) );
  OR2_X1 U11074 ( .A1(n10950), .A2(n9744), .ZN(n8588) );
  AND2_X1 U11075 ( .A1(n8584), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8585) );
  NOR2_X1 U11076 ( .A1(n8604), .A2(n8585), .ZN(n15277) );
  OR2_X1 U11077 ( .A1(n8905), .A2(n15277), .ZN(n8587) );
  INV_X1 U11078 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9743) );
  OR2_X1 U11079 ( .A1(n8795), .A2(n9743), .ZN(n8586) );
  OAI21_X1 U11080 ( .B1(n8590), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8592) );
  INV_X1 U11081 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8591) );
  XNOR2_X1 U11082 ( .A(n8592), .B(n8591), .ZN(n10631) );
  INV_X1 U11083 ( .A(n10631), .ZN(n9745) );
  NAND2_X1 U11084 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  OR2_X1 U11085 ( .A1(n8815), .A2(n9789), .ZN(n8598) );
  OR2_X1 U11086 ( .A1(n8517), .A2(SI_7_), .ZN(n8597) );
  OAI211_X1 U11087 ( .C1(n9745), .C2(n9692), .A(n8598), .B(n8597), .ZN(n15276)
         );
  INV_X1 U11088 ( .A(n15276), .ZN(n15139) );
  NAND2_X1 U11089 ( .A1(n12497), .A2(n15139), .ZN(n8600) );
  INV_X1 U11090 ( .A(n8600), .ZN(n8599) );
  NOR2_X1 U11091 ( .A1(n8599), .A2(n15272), .ZN(n8602) );
  NAND2_X1 U11092 ( .A1(n10037), .A2(n15292), .ZN(n15270) );
  AND2_X1 U11093 ( .A1(n15270), .A2(n8600), .ZN(n8601) );
  NAND2_X1 U11094 ( .A1(n10948), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8609) );
  INV_X1 U11095 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n8603) );
  OR2_X1 U11096 ( .A1(n10950), .A2(n8603), .ZN(n8608) );
  NOR2_X1 U11097 ( .A1(n8604), .A2(n15749), .ZN(n8605) );
  OR2_X1 U11098 ( .A1(n8905), .A2(n7765), .ZN(n8607) );
  INV_X1 U11099 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15392) );
  INV_X1 U11100 ( .A(n15131), .ZN(n11497) );
  NAND2_X1 U11101 ( .A1(n8610), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8611) );
  MUX2_X1 U11102 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8611), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8613) );
  INV_X1 U11103 ( .A(n8612), .ZN(n8630) );
  NAND2_X1 U11104 ( .A1(n8613), .A2(n8630), .ZN(n9804) );
  INV_X1 U11105 ( .A(SI_8_), .ZN(n9803) );
  OR2_X1 U11106 ( .A1(n8517), .A2(n9803), .ZN(n8619) );
  OR2_X1 U11107 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  NAND2_X1 U11108 ( .A1(n8617), .A2(n8616), .ZN(n9802) );
  OR2_X1 U11109 ( .A1(n8815), .A2(n9802), .ZN(n8618) );
  OAI211_X1 U11110 ( .C1(n9692), .C2(n9804), .A(n8619), .B(n8618), .ZN(n12495)
         );
  INV_X1 U11111 ( .A(n12495), .ZN(n8620) );
  NAND2_X1 U11112 ( .A1(n11497), .A2(n8620), .ZN(n11883) );
  NAND2_X1 U11113 ( .A1(n15131), .A2(n12495), .ZN(n11882) );
  NAND2_X1 U11114 ( .A1(n11369), .A2(n11979), .ZN(n11368) );
  NAND2_X1 U11115 ( .A1(n10948), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8627) );
  INV_X1 U11116 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11500) );
  OR2_X1 U11117 ( .A1(n10950), .A2(n11500), .ZN(n8626) );
  INV_X1 U11118 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11058) );
  OR2_X1 U11119 ( .A1(n8622), .A2(n8621), .ZN(n8623) );
  AND2_X1 U11120 ( .A1(n8636), .A2(n8623), .ZN(n11591) );
  OR2_X1 U11121 ( .A1(n8905), .A2(n11591), .ZN(n8624) );
  XNOR2_X1 U11122 ( .A(n8629), .B(n8628), .ZN(n9805) );
  OR2_X1 U11123 ( .A1(n8815), .A2(n9805), .ZN(n8634) );
  OR2_X1 U11124 ( .A1(n8517), .A2(SI_9_), .ZN(n8633) );
  OR2_X1 U11125 ( .A1(n8612), .A2(n8681), .ZN(n8631) );
  XNOR2_X1 U11126 ( .A(n8631), .B(P3_IR_REG_9__SCAN_IN), .ZN(n15180) );
  OR2_X1 U11127 ( .A1(n9692), .A2(n15180), .ZN(n8632) );
  NAND2_X1 U11128 ( .A1(n12496), .A2(n11885), .ZN(n11599) );
  OAI21_X1 U11129 ( .B1(n12496), .B2(n11885), .A(n11599), .ZN(n11980) );
  NAND2_X1 U11130 ( .A1(n10948), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8641) );
  INV_X1 U11131 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11707) );
  OR2_X1 U11132 ( .A1(n10950), .A2(n11707), .ZN(n8640) );
  NAND2_X1 U11133 ( .A1(n8636), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8637) );
  AND2_X1 U11134 ( .A1(n8652), .A2(n8637), .ZN(n15160) );
  OR2_X1 U11135 ( .A1(n8905), .A2(n15160), .ZN(n8639) );
  INV_X1 U11136 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11076) );
  INV_X1 U11137 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8642) );
  OR2_X1 U11138 ( .A1(n8741), .A2(n8681), .ZN(n8643) );
  XNOR2_X1 U11139 ( .A(n8643), .B(P3_IR_REG_10__SCAN_IN), .ZN(n11083) );
  OR2_X1 U11140 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  AND2_X1 U11141 ( .A1(n8647), .A2(n8646), .ZN(n9798) );
  OR2_X1 U11142 ( .A1(n8815), .A2(n9798), .ZN(n8648) );
  NAND2_X1 U11143 ( .A1(n8650), .A2(n11982), .ZN(n11606) );
  INV_X1 U11144 ( .A(n15153), .ZN(n11711) );
  NAND2_X1 U11145 ( .A1(n12401), .A2(n11711), .ZN(n8651) );
  NAND2_X1 U11146 ( .A1(n10948), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8658) );
  INV_X1 U11147 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14650) );
  OR2_X1 U11148 ( .A1(n10950), .A2(n14650), .ZN(n8657) );
  NAND2_X1 U11149 ( .A1(n8652), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8653) );
  AND2_X1 U11150 ( .A1(n8669), .A2(n8653), .ZN(n14656) );
  OR2_X1 U11151 ( .A1(n8905), .A2(n14656), .ZN(n8656) );
  INV_X1 U11152 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8654) );
  OR2_X1 U11153 ( .A1(n8795), .A2(n8654), .ZN(n8655) );
  INV_X1 U11154 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U11155 ( .A1(n8741), .A2(n8659), .ZN(n8680) );
  NAND2_X1 U11156 ( .A1(n8680), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8661) );
  INV_X1 U11157 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8660) );
  XNOR2_X1 U11158 ( .A(n8661), .B(n8660), .ZN(n15194) );
  AOI22_X1 U11159 ( .A1(n8790), .A2(n9800), .B1(n8789), .B2(n15194), .ZN(n8667) );
  OR2_X1 U11160 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  NAND2_X1 U11161 ( .A1(n8665), .A2(n8664), .ZN(n9801) );
  NAND2_X1 U11162 ( .A1(n9801), .A2(n11840), .ZN(n8666) );
  NAND2_X1 U11163 ( .A1(n12583), .A2(n12587), .ZN(n11895) );
  INV_X1 U11164 ( .A(n12583), .ZN(n10030) );
  NAND2_X1 U11165 ( .A1(n10030), .A2(n14651), .ZN(n11894) );
  NAND2_X1 U11166 ( .A1(n12583), .A2(n14651), .ZN(n8668) );
  NAND2_X1 U11167 ( .A1(n8507), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11168 ( .A1(n8669), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8670) );
  AND2_X1 U11169 ( .A1(n8696), .A2(n8670), .ZN(n12515) );
  OR2_X1 U11170 ( .A1(n8905), .A2(n12515), .ZN(n8674) );
  INV_X1 U11171 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12646) );
  OR2_X1 U11172 ( .A1(n10953), .A2(n12646), .ZN(n8673) );
  INV_X1 U11173 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8671) );
  OR2_X1 U11174 ( .A1(n8494), .A2(n8671), .ZN(n8672) );
  OR2_X1 U11175 ( .A1(n8677), .A2(n8676), .ZN(n8678) );
  NAND2_X1 U11176 ( .A1(n8679), .A2(n8678), .ZN(n9819) );
  OR2_X1 U11177 ( .A1(n9819), .A2(n8815), .ZN(n8687) );
  NOR2_X1 U11178 ( .A1(n8680), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8684) );
  OR2_X1 U11179 ( .A1(n8684), .A2(n8681), .ZN(n8682) );
  MUX2_X1 U11180 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8682), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8685) );
  INV_X1 U11181 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U11182 ( .A1(n8684), .A2(n8683), .ZN(n8708) );
  AOI22_X1 U11183 ( .A1(n8790), .A2(SI_12_), .B1(n8789), .B2(n15214), .ZN(
        n8686) );
  NAND2_X1 U11184 ( .A1(n8687), .A2(n8686), .ZN(n12517) );
  NAND2_X1 U11185 ( .A1(n14639), .A2(n12517), .ZN(n11899) );
  INV_X1 U11186 ( .A(n12517), .ZN(n11727) );
  NAND2_X1 U11187 ( .A1(n11727), .A2(n12566), .ZN(n11900) );
  NAND2_X1 U11188 ( .A1(n11899), .A2(n11900), .ZN(n11985) );
  NAND2_X1 U11189 ( .A1(n12517), .A2(n12566), .ZN(n14635) );
  NAND2_X1 U11190 ( .A1(n8688), .A2(n10013), .ZN(n8689) );
  NAND2_X1 U11191 ( .A1(n8690), .A2(n8689), .ZN(n9836) );
  NAND2_X1 U11192 ( .A1(n9836), .A2(n11840), .ZN(n8693) );
  NAND2_X1 U11193 ( .A1(n8708), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8691) );
  XNOR2_X1 U11194 ( .A(n8691), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12668) );
  INV_X1 U11195 ( .A(n12668), .ZN(n15234) );
  AOI22_X1 U11196 ( .A1(n8790), .A2(n15723), .B1(n8789), .B2(n15234), .ZN(
        n8692) );
  NAND2_X1 U11197 ( .A1(n8693), .A2(n8692), .ZN(n14641) );
  NAND2_X1 U11198 ( .A1(n10948), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8701) );
  INV_X1 U11199 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8694) );
  OR2_X1 U11200 ( .A1(n10950), .A2(n8694), .ZN(n8700) );
  INV_X1 U11201 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8695) );
  OR2_X1 U11202 ( .A1(n10953), .A2(n8695), .ZN(n8699) );
  NAND2_X1 U11203 ( .A1(n8696), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8697) );
  AND2_X1 U11204 ( .A1(n8713), .A2(n8697), .ZN(n14642) );
  OR2_X1 U11205 ( .A1(n8905), .A2(n14642), .ZN(n8698) );
  OR2_X1 U11206 ( .A1(n14641), .A2(n12562), .ZN(n8702) );
  AND2_X1 U11207 ( .A1(n14635), .A2(n8702), .ZN(n8703) );
  OR2_X1 U11208 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  NAND2_X1 U11209 ( .A1(n8707), .A2(n8706), .ZN(n9845) );
  NAND2_X1 U11210 ( .A1(n9845), .A2(n11840), .ZN(n8712) );
  OR2_X1 U11211 ( .A1(n8708), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U11212 ( .A1(n8724), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8710) );
  INV_X1 U11213 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8709) );
  XNOR2_X1 U11214 ( .A(n8710), .B(n8709), .ZN(n15248) );
  AOI22_X1 U11215 ( .A1(n8790), .A2(n15542), .B1(n8789), .B2(n15248), .ZN(
        n8711) );
  NAND2_X1 U11216 ( .A1(n8507), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8718) );
  INV_X1 U11217 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13020) );
  OR2_X1 U11218 ( .A1(n8795), .A2(n13020), .ZN(n8717) );
  NAND2_X1 U11219 ( .A1(n8713), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8714) );
  AND2_X1 U11220 ( .A1(n8728), .A2(n8714), .ZN(n12455) );
  OR2_X1 U11221 ( .A1(n8905), .A2(n12455), .ZN(n8716) );
  INV_X1 U11222 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13108) );
  OR2_X1 U11223 ( .A1(n8494), .A2(n13108), .ZN(n8715) );
  NAND4_X1 U11224 ( .A1(n8718), .A2(n8717), .A3(n8716), .A4(n8715), .ZN(n12936) );
  OR2_X1 U11225 ( .A1(n13113), .A2(n12936), .ZN(n11910) );
  NAND2_X1 U11226 ( .A1(n13113), .A2(n12936), .ZN(n11908) );
  NAND2_X1 U11227 ( .A1(n11910), .A2(n11908), .ZN(n12942) );
  OR2_X1 U11228 ( .A1(n13113), .A2(n14640), .ZN(n8719) );
  OR2_X1 U11229 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  NAND2_X1 U11230 ( .A1(n8723), .A2(n8722), .ZN(n9853) );
  OR2_X1 U11231 ( .A1(n9853), .A2(n8815), .ZN(n8727) );
  OAI21_X1 U11232 ( .B1(n8724), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U11233 ( .A(n8725), .B(P3_IR_REG_15__SCAN_IN), .ZN(n14626) );
  AOI22_X1 U11234 ( .A1(n8790), .A2(SI_15_), .B1(n8789), .B2(n14626), .ZN(
        n8726) );
  NAND2_X1 U11235 ( .A1(n10948), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8733) );
  INV_X1 U11236 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14616) );
  OR2_X1 U11237 ( .A1(n10950), .A2(n14616), .ZN(n8732) );
  NAND2_X1 U11238 ( .A1(n8728), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8729) );
  AND2_X1 U11239 ( .A1(n8747), .A2(n8729), .ZN(n12614) );
  OR2_X1 U11240 ( .A1(n8905), .A2(n12614), .ZN(n8731) );
  INV_X1 U11241 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14628) );
  OR2_X1 U11242 ( .A1(n10953), .A2(n14628), .ZN(n8730) );
  NAND4_X1 U11243 ( .A1(n8733), .A2(n8732), .A3(n8731), .A4(n8730), .ZN(n12949) );
  AND2_X1 U11244 ( .A1(n13102), .A2(n12949), .ZN(n8734) );
  OR2_X1 U11245 ( .A1(n13102), .A2(n12949), .ZN(n8735) );
  OR2_X1 U11246 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  NAND2_X1 U11247 ( .A1(n8739), .A2(n8738), .ZN(n9917) );
  OR2_X1 U11248 ( .A1(n9917), .A2(n8815), .ZN(n8746) );
  NAND2_X1 U11249 ( .A1(n8743), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8742) );
  MUX2_X1 U11250 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8742), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8744) );
  AND2_X1 U11251 ( .A1(n8744), .A2(n8757), .ZN(n12673) );
  AOI22_X1 U11252 ( .A1(n8790), .A2(SI_16_), .B1(n8789), .B2(n12673), .ZN(
        n8745) );
  NAND2_X1 U11253 ( .A1(n10948), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8752) );
  INV_X1 U11254 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12927) );
  OR2_X1 U11255 ( .A1(n10950), .A2(n12927), .ZN(n8751) );
  NAND2_X1 U11256 ( .A1(n8747), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8748) );
  AND2_X1 U11257 ( .A1(n8775), .A2(n8748), .ZN(n12928) );
  OR2_X1 U11258 ( .A1(n8905), .A2(n12928), .ZN(n8750) );
  INV_X1 U11259 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13013) );
  OR2_X1 U11260 ( .A1(n8795), .A2(n13013), .ZN(n8749) );
  OR2_X1 U11261 ( .A1(n13095), .A2(n12528), .ZN(n11919) );
  NAND2_X1 U11262 ( .A1(n13095), .A2(n12528), .ZN(n11920) );
  NAND2_X1 U11263 ( .A1(n13095), .A2(n12937), .ZN(n8753) );
  XNOR2_X1 U11264 ( .A(n8755), .B(n8754), .ZN(n10010) );
  NAND2_X1 U11265 ( .A1(n10010), .A2(n11840), .ZN(n8762) );
  NAND2_X1 U11266 ( .A1(n8757), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8756) );
  MUX2_X1 U11267 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8756), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8759) );
  INV_X1 U11268 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11269 ( .A1(n8759), .A2(n8786), .ZN(n12718) );
  INV_X1 U11270 ( .A(n12718), .ZN(n8760) );
  AOI22_X1 U11271 ( .A1(n8790), .A2(SI_17_), .B1(n8789), .B2(n8760), .ZN(n8761) );
  NAND2_X1 U11272 ( .A1(n10948), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8767) );
  INV_X1 U11273 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12915) );
  OR2_X1 U11274 ( .A1(n10950), .A2(n12915), .ZN(n8766) );
  INV_X1 U11275 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8763) );
  XNOR2_X1 U11276 ( .A(n8775), .B(n8763), .ZN(n12541) );
  OR2_X1 U11277 ( .A1(n8905), .A2(n12541), .ZN(n8765) );
  INV_X1 U11278 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13010) );
  OR2_X1 U11279 ( .A1(n10953), .A2(n13010), .ZN(n8764) );
  OR2_X1 U11280 ( .A1(n13089), .A2(n12596), .ZN(n11927) );
  NAND2_X1 U11281 ( .A1(n13089), .A2(n12596), .ZN(n11923) );
  NAND2_X1 U11282 ( .A1(n11927), .A2(n11923), .ZN(n12911) );
  NAND2_X1 U11283 ( .A1(n12910), .A2(n12911), .ZN(n12909) );
  OR2_X1 U11284 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  NAND2_X1 U11285 ( .A1(n8771), .A2(n8770), .ZN(n10018) );
  OR2_X1 U11286 ( .A1(n10018), .A2(n8815), .ZN(n8774) );
  NAND2_X1 U11287 ( .A1(n8786), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8772) );
  XNOR2_X1 U11288 ( .A(n8772), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U11289 ( .A1(n8790), .A2(SI_18_), .B1(n8789), .B2(n12715), .ZN(
        n8773) );
  NAND2_X1 U11290 ( .A1(n10948), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8780) );
  INV_X1 U11291 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12902) );
  OR2_X1 U11292 ( .A1(n10950), .A2(n12902), .ZN(n8779) );
  OAI21_X1 U11293 ( .B1(n8775), .B2(P3_REG3_REG_17__SCAN_IN), .A(
        P3_REG3_REG_18__SCAN_IN), .ZN(n8776) );
  AND2_X1 U11294 ( .A1(n8793), .A2(n8776), .ZN(n12595) );
  OR2_X1 U11295 ( .A1(n8905), .A2(n12595), .ZN(n8778) );
  INV_X1 U11296 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13007) );
  OR2_X1 U11297 ( .A1(n8795), .A2(n13007), .ZN(n8777) );
  NAND2_X1 U11298 ( .A1(n13083), .A2(n12543), .ZN(n11929) );
  INV_X1 U11299 ( .A(n12596), .ZN(n12423) );
  NAND2_X1 U11300 ( .A1(n13089), .A2(n12423), .ZN(n12897) );
  OR2_X1 U11301 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  NAND2_X1 U11302 ( .A1(n8785), .A2(n8784), .ZN(n10163) );
  NAND2_X1 U11303 ( .A1(n10163), .A2(n11840), .ZN(n8792) );
  INV_X1 U11304 ( .A(n8912), .ZN(n8787) );
  NAND2_X1 U11305 ( .A1(n8787), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8788) );
  AOI22_X1 U11306 ( .A1(n8790), .A2(n10164), .B1(n8789), .B2(n7624), .ZN(n8791) );
  NAND2_X1 U11307 ( .A1(n8793), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11308 ( .A1(n8807), .A2(n8794), .ZN(n12475) );
  NAND2_X1 U11309 ( .A1(n8894), .A2(n12475), .ZN(n8799) );
  INV_X1 U11310 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13076) );
  OR2_X1 U11311 ( .A1(n8494), .A2(n13076), .ZN(n8798) );
  INV_X1 U11312 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12888) );
  OR2_X1 U11313 ( .A1(n10950), .A2(n12888), .ZN(n8797) );
  INV_X1 U11314 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13004) );
  OR2_X1 U11315 ( .A1(n8795), .A2(n13004), .ZN(n8796) );
  NAND4_X1 U11316 ( .A1(n8799), .A2(n8798), .A3(n8797), .A4(n8796), .ZN(n12868) );
  NAND2_X1 U11317 ( .A1(n13080), .A2(n12868), .ZN(n11934) );
  NAND2_X1 U11318 ( .A1(n11933), .A2(n11934), .ZN(n12889) );
  OR2_X1 U11319 ( .A1(n13083), .A2(n12912), .ZN(n12883) );
  AND2_X1 U11320 ( .A1(n12889), .A2(n12883), .ZN(n8800) );
  INV_X1 U11321 ( .A(n12868), .ZN(n12597) );
  OR2_X1 U11322 ( .A1(n13080), .A2(n12597), .ZN(n8801) );
  NAND2_X1 U11323 ( .A1(n8802), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U11324 ( .A1(n8804), .A2(n8803), .ZN(n10453) );
  OR2_X1 U11325 ( .A1(n8517), .A2(n10454), .ZN(n8805) );
  NAND2_X1 U11326 ( .A1(n8807), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U11327 ( .A1(n8818), .A2(n8808), .ZN(n12872) );
  AOI22_X1 U11328 ( .A1(n12872), .A2(n8894), .B1(n8832), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n8810) );
  AOI22_X1 U11329 ( .A1(n10948), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n8507), 
        .B2(P3_REG2_REG_20__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U11330 ( .A1(n12876), .A2(n12474), .ZN(n11938) );
  NAND2_X2 U11331 ( .A1(n12867), .A2(n12877), .ZN(n12856) );
  OR2_X1 U11332 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  NAND2_X1 U11333 ( .A1(n8814), .A2(n8813), .ZN(n10675) );
  INV_X1 U11334 ( .A(SI_21_), .ZN(n10676) );
  OR2_X1 U11335 ( .A1(n8517), .A2(n10676), .ZN(n8816) );
  NAND2_X1 U11336 ( .A1(n8818), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U11337 ( .A1(n8830), .A2(n8819), .ZN(n12864) );
  NAND2_X1 U11338 ( .A1(n12864), .A2(n8894), .ZN(n8822) );
  AOI22_X1 U11339 ( .A1(n10948), .A2(P3_REG0_REG_21__SCAN_IN), .B1(n8507), 
        .B2(P3_REG2_REG_21__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11340 ( .A1(n8832), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U11341 ( .A1(n13070), .A2(n8824), .ZN(n11941) );
  NAND2_X1 U11342 ( .A1(n11942), .A2(n11941), .ZN(n12857) );
  NAND2_X1 U11343 ( .A1(n12876), .A2(n12505), .ZN(n12858) );
  AND2_X1 U11344 ( .A1(n12857), .A2(n12858), .ZN(n8823) );
  OR2_X1 U11345 ( .A1(n13070), .A2(n12869), .ZN(n8825) );
  XNOR2_X1 U11346 ( .A(n8827), .B(n8826), .ZN(n10774) );
  NAND2_X1 U11347 ( .A1(n10774), .A2(n11840), .ZN(n8829) );
  OR2_X1 U11348 ( .A1(n8517), .A2(n15742), .ZN(n8828) );
  NAND2_X2 U11349 ( .A1(n8829), .A2(n8828), .ZN(n13064) );
  INV_X1 U11350 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13063) );
  NAND2_X1 U11351 ( .A1(n8830), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U11352 ( .A1(n8841), .A2(n8831), .ZN(n12849) );
  NAND2_X1 U11353 ( .A1(n12849), .A2(n8894), .ZN(n8834) );
  AOI22_X1 U11354 ( .A1(n8832), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n8507), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n8833) );
  OAI211_X1 U11355 ( .C1(n8494), .C2(n13063), .A(n8834), .B(n8833), .ZN(n12573) );
  NOR2_X1 U11356 ( .A1(n13064), .A2(n12573), .ZN(n8836) );
  NAND2_X1 U11357 ( .A1(n13064), .A2(n12573), .ZN(n8835) );
  XNOR2_X1 U11358 ( .A(n8838), .B(n8837), .ZN(n10946) );
  NAND2_X1 U11359 ( .A1(n10946), .A2(n11840), .ZN(n8840) );
  OR2_X1 U11360 ( .A1(n8517), .A2(n15478), .ZN(n8839) );
  XNOR2_X1 U11361 ( .A(n8841), .B(P3_REG3_REG_23__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U11362 ( .A1(n12837), .A2(n8894), .ZN(n8846) );
  INV_X1 U11363 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U11364 ( .A1(n10948), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11365 ( .A1(n8507), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8842) );
  OAI211_X1 U11366 ( .C1(n12991), .C2(n10953), .A(n8843), .B(n8842), .ZN(n8844) );
  INV_X1 U11367 ( .A(n8844), .ZN(n8845) );
  NAND2_X1 U11368 ( .A1(n12987), .A2(n12846), .ZN(n8847) );
  XNOR2_X1 U11369 ( .A(n8849), .B(n7602), .ZN(n11271) );
  NAND2_X1 U11370 ( .A1(n11271), .A2(n11840), .ZN(n8851) );
  INV_X1 U11371 ( .A(SI_24_), .ZN(n11272) );
  OR2_X1 U11372 ( .A1(n8517), .A2(n11272), .ZN(n8850) );
  NAND2_X2 U11373 ( .A1(n8851), .A2(n8850), .ZN(n13054) );
  NAND2_X1 U11374 ( .A1(n8852), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U11375 ( .A1(n8864), .A2(n8853), .ZN(n12824) );
  NAND2_X1 U11376 ( .A1(n12824), .A2(n8894), .ZN(n8858) );
  INV_X1 U11377 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12984) );
  NAND2_X1 U11378 ( .A1(n10948), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11379 ( .A1(n8507), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8854) );
  OAI211_X1 U11380 ( .C1(n12984), .C2(n10953), .A(n8855), .B(n8854), .ZN(n8856) );
  INV_X1 U11381 ( .A(n8856), .ZN(n8857) );
  AND2_X1 U11382 ( .A1(n13054), .A2(n12522), .ZN(n8859) );
  OAI22_X1 U11383 ( .A1(n12819), .A2(n8859), .B1(n12522), .B2(n13054), .ZN(
        n12804) );
  XNOR2_X1 U11384 ( .A(n13838), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8860) );
  XNOR2_X1 U11385 ( .A(n8861), .B(n8860), .ZN(n11414) );
  NAND2_X1 U11386 ( .A1(n11414), .A2(n11840), .ZN(n8863) );
  OR2_X1 U11387 ( .A1(n8517), .A2(n15715), .ZN(n8862) );
  NAND2_X1 U11388 ( .A1(n8864), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U11389 ( .A1(n8876), .A2(n8865), .ZN(n12810) );
  NAND2_X1 U11390 ( .A1(n12810), .A2(n8894), .ZN(n8870) );
  INV_X1 U11391 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12982) );
  NAND2_X1 U11392 ( .A1(n10948), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U11393 ( .A1(n8507), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8866) );
  OAI211_X1 U11394 ( .C1(n12982), .C2(n10953), .A(n8867), .B(n8866), .ZN(n8868) );
  INV_X1 U11395 ( .A(n8868), .ZN(n8869) );
  NAND2_X1 U11396 ( .A1(n12811), .A2(n12821), .ZN(n8871) );
  NAND2_X2 U11397 ( .A1(n12805), .A2(n8871), .ZN(n12795) );
  XNOR2_X1 U11398 ( .A(n13833), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8872) );
  XNOR2_X1 U11399 ( .A(n8873), .B(n8872), .ZN(n11479) );
  NAND2_X1 U11400 ( .A1(n11479), .A2(n11840), .ZN(n8875) );
  OR2_X1 U11401 ( .A1(n8517), .A2(n15673), .ZN(n8874) );
  NAND2_X1 U11402 ( .A1(n8876), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11403 ( .A1(n8888), .A2(n8877), .ZN(n12799) );
  NAND2_X1 U11404 ( .A1(n12799), .A2(n8894), .ZN(n8882) );
  INV_X1 U11405 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12976) );
  NAND2_X1 U11406 ( .A1(n8507), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U11407 ( .A1(n10948), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8878) );
  OAI211_X1 U11408 ( .C1(n12976), .C2(n10953), .A(n8879), .B(n8878), .ZN(n8880) );
  INV_X1 U11409 ( .A(n8880), .ZN(n8881) );
  OR2_X1 U11410 ( .A1(n13044), .A2(n12523), .ZN(n8883) );
  XNOR2_X1 U11411 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8884) );
  XNOR2_X1 U11412 ( .A(n8885), .B(n8884), .ZN(n11800) );
  NAND2_X1 U11413 ( .A1(n11800), .A2(n11840), .ZN(n8887) );
  INV_X1 U11414 ( .A(SI_27_), .ZN(n15494) );
  OR2_X1 U11415 ( .A1(n8517), .A2(n15494), .ZN(n8886) );
  NAND2_X1 U11416 ( .A1(n8888), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U11417 ( .A1(n8890), .A2(n8889), .ZN(n12788) );
  INV_X1 U11418 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12974) );
  NAND2_X1 U11419 ( .A1(n8507), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11420 ( .A1(n10948), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8891) );
  OAI211_X1 U11421 ( .C1(n12974), .C2(n10953), .A(n8892), .B(n8891), .ZN(n8893) );
  NAND2_X1 U11422 ( .A1(n12787), .A2(n12766), .ZN(n12758) );
  OR2_X2 U11423 ( .A1(n13035), .A2(n12782), .ZN(n11965) );
  NAND2_X1 U11424 ( .A1(n13035), .A2(n12782), .ZN(n9001) );
  INV_X1 U11425 ( .A(n12766), .ZN(n10780) );
  OR2_X1 U11426 ( .A1(n12787), .A2(n10780), .ZN(n12761) );
  AND2_X1 U11427 ( .A1(n12762), .A2(n12761), .ZN(n8896) );
  OAI21_X1 U11428 ( .B1(n12782), .B2(n8897), .A(n12764), .ZN(n8910) );
  AND2_X1 U11429 ( .A1(n14485), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U11430 ( .A1(n8900), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8901) );
  XNOR2_X1 U11431 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11830) );
  XNOR2_X1 U11432 ( .A(n11832), .B(n11830), .ZN(n13126) );
  NAND2_X1 U11433 ( .A1(n13126), .A2(n11840), .ZN(n8904) );
  OR2_X1 U11434 ( .A1(n8517), .A2(n13129), .ZN(n8903) );
  INV_X1 U11435 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n12964) );
  NAND2_X1 U11436 ( .A1(n10948), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U11437 ( .A1(n8507), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8906) );
  OAI211_X1 U11438 ( .C1(n10953), .C2(n12964), .A(n8907), .B(n8906), .ZN(n8908) );
  INV_X1 U11439 ( .A(n8908), .ZN(n8909) );
  NAND2_X1 U11440 ( .A1(n12965), .A2(n12767), .ZN(n11969) );
  XNOR2_X1 U11441 ( .A(n8910), .B(n11995), .ZN(n8934) );
  INV_X1 U11442 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11443 ( .A1(n8918), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8913) );
  MUX2_X1 U11444 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8913), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8915) );
  NAND2_X1 U11445 ( .A1(n8916), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8917) );
  MUX2_X1 U11446 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8917), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8919) );
  NAND2_X1 U11447 ( .A1(n11855), .A2(n9002), .ZN(n11851) );
  NAND2_X1 U11448 ( .A1(n8914), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8920) );
  XNOR2_X1 U11449 ( .A(n8920), .B(n7632), .ZN(n10772) );
  NAND2_X1 U11450 ( .A1(n12742), .A2(n12004), .ZN(n8935) );
  INV_X1 U11451 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U11452 ( .A1(n10948), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U11453 ( .A1(n8507), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8921) );
  OAI211_X1 U11454 ( .C1(n8923), .C2(n10953), .A(n8922), .B(n8921), .ZN(n8924)
         );
  INV_X1 U11455 ( .A(n8924), .ZN(n8925) );
  INV_X1 U11456 ( .A(n8926), .ZN(n9755) );
  NAND2_X1 U11457 ( .A1(n9755), .A2(n12651), .ZN(n9694) );
  NAND2_X1 U11458 ( .A1(n9692), .A2(n9694), .ZN(n8929) );
  AND2_X1 U11459 ( .A1(n9755), .A2(P3_B_REG_SCAN_IN), .ZN(n8928) );
  OR2_X1 U11460 ( .A1(n15315), .A2(n8928), .ZN(n12750) );
  NOR2_X1 U11461 ( .A1(n11845), .A2(n12750), .ZN(n8932) );
  INV_X1 U11462 ( .A(n8929), .ZN(n8930) );
  NOR2_X1 U11463 ( .A1(n12782), .A2(n15313), .ZN(n8931) );
  OAI21_X1 U11464 ( .B1(n8934), .B2(n15311), .A(n8933), .ZN(n12391) );
  INV_X1 U11465 ( .A(n12391), .ZN(n12963) );
  NAND2_X1 U11466 ( .A1(n6680), .A2(n7624), .ZN(n10421) );
  INV_X1 U11467 ( .A(n10421), .ZN(n11974) );
  NAND2_X1 U11468 ( .A1(n11959), .A2(n11974), .ZN(n10407) );
  INV_X1 U11469 ( .A(n8935), .ZN(n8936) );
  NAND2_X1 U11470 ( .A1(n6833), .A2(n8936), .ZN(n10285) );
  AND2_X1 U11471 ( .A1(n10407), .A2(n10285), .ZN(n8972) );
  NAND2_X1 U11472 ( .A1(n6779), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8937) );
  MUX2_X1 U11473 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8937), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8939) );
  NAND2_X1 U11474 ( .A1(n8939), .A2(n8938), .ZN(n11274) );
  XNOR2_X1 U11475 ( .A(n11274), .B(P3_B_REG_SCAN_IN), .ZN(n8943) );
  NAND2_X1 U11476 ( .A1(n8938), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8940) );
  MUX2_X1 U11477 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8940), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8942) );
  NAND2_X1 U11478 ( .A1(n8942), .A2(n8944), .ZN(n11416) );
  NAND2_X1 U11479 ( .A1(n8944), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8945) );
  MUX2_X1 U11480 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8945), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8947) );
  NAND2_X1 U11481 ( .A1(n8947), .A2(n8946), .ZN(n11481) );
  INV_X1 U11482 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U11483 ( .A1(n11798), .A2(n9826), .ZN(n8950) );
  NAND2_X1 U11484 ( .A1(n11481), .A2(n11416), .ZN(n8949) );
  NAND2_X1 U11485 ( .A1(n8950), .A2(n8949), .ZN(n10470) );
  INV_X1 U11486 ( .A(n10470), .ZN(n10423) );
  INV_X1 U11487 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U11488 ( .A1(n11798), .A2(n8951), .ZN(n8953) );
  NAND2_X1 U11489 ( .A1(n11481), .A2(n11274), .ZN(n8952) );
  NAND2_X1 U11490 ( .A1(n10423), .A2(n13116), .ZN(n10416) );
  NOR2_X1 U11491 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8957) );
  NOR4_X1 U11492 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8956) );
  NOR4_X1 U11493 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8955) );
  NOR4_X1 U11494 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8954) );
  NAND4_X1 U11495 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n8963)
         );
  NOR4_X1 U11496 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8961) );
  NOR4_X1 U11497 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8960) );
  NOR4_X1 U11498 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8959) );
  NOR4_X1 U11499 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8958) );
  NAND4_X1 U11500 ( .A1(n8961), .A2(n8960), .A3(n8959), .A4(n8958), .ZN(n8962)
         );
  OAI21_X1 U11501 ( .B1(n8963), .B2(n8962), .A(n11798), .ZN(n10412) );
  INV_X1 U11502 ( .A(n10412), .ZN(n8970) );
  OR2_X1 U11503 ( .A1(n10416), .A2(n8970), .ZN(n10282) );
  NAND2_X1 U11504 ( .A1(n10677), .A2(n6680), .ZN(n8964) );
  NAND2_X1 U11505 ( .A1(n8964), .A2(n10772), .ZN(n8968) );
  NAND2_X1 U11506 ( .A1(n6680), .A2(n12004), .ZN(n8965) );
  NAND2_X1 U11507 ( .A1(n8965), .A2(n12742), .ZN(n8966) );
  NAND2_X1 U11508 ( .A1(n8966), .A2(n10677), .ZN(n8967) );
  NAND2_X1 U11509 ( .A1(n8968), .A2(n8967), .ZN(n10281) );
  INV_X1 U11510 ( .A(n10281), .ZN(n8971) );
  INV_X1 U11511 ( .A(n13116), .ZN(n8969) );
  NAND2_X1 U11512 ( .A1(n10470), .A2(n8969), .ZN(n10473) );
  OAI22_X1 U11513 ( .A1(n8972), .A2(n10282), .B1(n8971), .B2(n10291), .ZN(
        n8977) );
  INV_X1 U11514 ( .A(n11481), .ZN(n8974) );
  NOR2_X1 U11515 ( .A1(n11416), .A2(n11274), .ZN(n8973) );
  NAND2_X1 U11516 ( .A1(n8974), .A2(n8973), .ZN(n10284) );
  NAND2_X1 U11517 ( .A1(n6840), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8976) );
  XNOR2_X1 U11518 ( .A(n8976), .B(n8975), .ZN(n10283) );
  NAND2_X1 U11519 ( .A1(n10284), .A2(n13115), .ZN(n10476) );
  INV_X1 U11520 ( .A(n15301), .ZN(n8979) );
  NOR2_X1 U11521 ( .A1(n11853), .A2(n6682), .ZN(n8978) );
  AOI21_X2 U11522 ( .B1(n6999), .B2(n8979), .A(n8978), .ZN(n11861) );
  INV_X1 U11523 ( .A(n10279), .ZN(n10481) );
  NOR2_X2 U11524 ( .A1(n10504), .A2(n10481), .ZN(n11856) );
  NAND2_X1 U11525 ( .A1(n15299), .A2(n6999), .ZN(n15303) );
  NAND2_X1 U11526 ( .A1(n11861), .A2(n15303), .ZN(n11011) );
  NAND2_X1 U11527 ( .A1(n11011), .A2(n11977), .ZN(n11010) );
  NAND2_X1 U11528 ( .A1(n11149), .A2(n11976), .ZN(n8980) );
  NAND2_X1 U11529 ( .A1(n8980), .A2(n11866), .ZN(n11310) );
  NAND2_X1 U11530 ( .A1(n11310), .A2(n11870), .ZN(n8981) );
  NAND2_X1 U11531 ( .A1(n15282), .A2(n15283), .ZN(n11364) );
  INV_X1 U11532 ( .A(n8987), .ZN(n8983) );
  INV_X1 U11533 ( .A(n12497), .ZN(n11370) );
  NAND2_X1 U11534 ( .A1(n11370), .A2(n15139), .ZN(n11365) );
  AND2_X1 U11535 ( .A1(n11365), .A2(n11882), .ZN(n8982) );
  INV_X1 U11536 ( .A(n11885), .ZN(n8989) );
  OR2_X1 U11537 ( .A1(n12496), .A2(n8989), .ZN(n8984) );
  AND2_X1 U11538 ( .A1(n11877), .A2(n8985), .ZN(n8986) );
  NAND2_X1 U11539 ( .A1(n11364), .A2(n8986), .ZN(n8991) );
  NOR2_X1 U11540 ( .A1(n7761), .A2(n7757), .ZN(n8990) );
  NAND2_X1 U11541 ( .A1(n12401), .A2(n15153), .ZN(n11890) );
  INV_X1 U11542 ( .A(n11985), .ZN(n11721) );
  NAND2_X1 U11543 ( .A1(n11722), .A2(n11721), .ZN(n8992) );
  INV_X1 U11544 ( .A(n14641), .ZN(n12570) );
  NAND2_X1 U11545 ( .A1(n14641), .A2(n12947), .ZN(n11905) );
  INV_X1 U11546 ( .A(n11908), .ZN(n8993) );
  INV_X1 U11547 ( .A(n12949), .ZN(n12532) );
  OR2_X1 U11548 ( .A1(n13102), .A2(n12532), .ZN(n11918) );
  NAND2_X1 U11549 ( .A1(n13102), .A2(n12532), .ZN(n11912) );
  NAND2_X1 U11550 ( .A1(n8994), .A2(n11912), .ZN(n12922) );
  NAND2_X1 U11551 ( .A1(n12922), .A2(n12921), .ZN(n12920) );
  INV_X1 U11552 ( .A(n12911), .ZN(n12907) );
  NAND2_X1 U11553 ( .A1(n12908), .A2(n12907), .ZN(n8995) );
  INV_X1 U11554 ( .A(n12898), .ZN(n8996) );
  INV_X1 U11555 ( .A(n12890), .ZN(n8997) );
  NAND2_X1 U11556 ( .A1(n8997), .A2(n11934), .ZN(n8998) );
  NAND2_X1 U11557 ( .A1(n8998), .A2(n11933), .ZN(n12878) );
  NAND2_X1 U11558 ( .A1(n13064), .A2(n12832), .ZN(n11946) );
  NAND2_X1 U11559 ( .A1(n12843), .A2(n11946), .ZN(n8999) );
  NAND2_X1 U11560 ( .A1(n8999), .A2(n11945), .ZN(n12827) );
  NAND2_X1 U11561 ( .A1(n12803), .A2(n12802), .ZN(n9000) );
  NAND2_X1 U11562 ( .A1(n12811), .A2(n12605), .ZN(n11957) );
  NAND2_X1 U11563 ( .A1(n9000), .A2(n11957), .ZN(n12793) );
  NAND2_X1 U11564 ( .A1(n13044), .A2(n12781), .ZN(n11960) );
  AND2_X2 U11565 ( .A1(n12777), .A2(n12776), .ZN(n12779) );
  NAND2_X1 U11566 ( .A1(n9001), .A2(n12758), .ZN(n11964) );
  OAI21_X2 U11567 ( .B1(n12779), .B2(n11964), .A(n11965), .ZN(n11843) );
  NAND3_X1 U11568 ( .A1(n15339), .A2(n10281), .A3(n11974), .ZN(n9003) );
  NOR2_X1 U11569 ( .A1(n12742), .A2(n10772), .ZN(n10418) );
  NAND2_X1 U11570 ( .A1(n9002), .A2(n10418), .ZN(n10411) );
  NAND2_X1 U11571 ( .A1(n6680), .A2(n12742), .ZN(n15327) );
  OR2_X1 U11572 ( .A1(n15327), .A2(n12004), .ZN(n12971) );
  AND2_X1 U11573 ( .A1(n15289), .A2(n12971), .ZN(n11610) );
  INV_X1 U11574 ( .A(n11610), .ZN(n15368) );
  NAND2_X1 U11575 ( .A1(n12966), .A2(n13109), .ZN(n9008) );
  INV_X1 U11576 ( .A(n12965), .ZN(n12390) );
  NAND2_X1 U11577 ( .A1(n15382), .A2(n15328), .ZN(n13114) );
  INV_X1 U11578 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9004) );
  OR2_X1 U11579 ( .A1(n15382), .A2(n9004), .ZN(n9005) );
  OAI21_X1 U11580 ( .B1(n12963), .B2(n9009), .A(n7766), .ZN(P3_U3456) );
  NOR2_X1 U11581 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n9013) );
  NAND4_X1 U11582 ( .A1(n9013), .A2(n9012), .A3(n9011), .A4(n9010), .ZN(n9286)
         );
  NOR3_X2 U11583 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .A3(
        P2_IR_REG_3__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U11584 ( .A1(n9019), .A2(n9039), .ZN(n9026) );
  NOR2_X2 U11585 ( .A1(n9037), .A2(n9026), .ZN(n9033) );
  INV_X1 U11586 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9045) );
  OAI21_X1 U11587 ( .B1(n9649), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9022) );
  OAI21_X1 U11588 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_27__SCAN_IN), 
        .A(n9022), .ZN(n9023) );
  INV_X1 U11589 ( .A(n9023), .ZN(n9024) );
  AOI21_X1 U11590 ( .B1(n9025), .B2(n7759), .A(n9024), .ZN(n9031) );
  NOR2_X1 U11591 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n9027) );
  INV_X1 U11592 ( .A(n9555), .ZN(n9063) );
  NAND2_X1 U11593 ( .A1(n9398), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9032) );
  INV_X1 U11594 ( .A(n9047), .ZN(n9034) );
  NAND2_X1 U11595 ( .A1(n9034), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9035) );
  INV_X1 U11596 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9038) );
  NAND3_X1 U11597 ( .A1(n9335), .A2(n9039), .A3(n9038), .ZN(n9040) );
  XNOR2_X1 U11598 ( .A(n9041), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11599 ( .A1(n9042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9043) );
  INV_X1 U11600 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9044) );
  AND2_X1 U11601 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  INV_X1 U11602 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9644) );
  INV_X4 U11603 ( .A(n9617), .ZN(n9593) );
  AND2_X1 U11604 ( .A1(n9095), .A2(n9661), .ZN(n9113) );
  INV_X1 U11605 ( .A(n9113), .ZN(n9170) );
  AND2_X1 U11606 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9071) );
  NAND2_X1 U11607 ( .A1(n9071), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U11608 ( .A1(n9181), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9222) );
  INV_X1 U11609 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9236) );
  INV_X1 U11610 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9293) );
  INV_X1 U11611 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9309) );
  INV_X1 U11612 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U11613 ( .A1(n9326), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9356) );
  INV_X1 U11614 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13257) );
  INV_X1 U11615 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13277) );
  INV_X1 U11616 ( .A(n9426), .ZN(n9052) );
  INV_X1 U11617 ( .A(n9050), .ZN(n9404) );
  INV_X1 U11618 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13304) );
  NAND2_X1 U11619 ( .A1(n9404), .A2(n13304), .ZN(n9051) );
  AND2_X1 U11620 ( .A1(n9052), .A2(n9051), .ZN(n13615) );
  INV_X1 U11621 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9053) );
  NAND2_X2 U11622 ( .A1(n13818), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9078) );
  INV_X1 U11623 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9085) );
  XNOR2_X2 U11624 ( .A(n9078), .B(n9085), .ZN(n9058) );
  NAND2_X1 U11625 ( .A1(n9055), .A2(n9054), .ZN(n9056) );
  INV_X1 U11626 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9061) );
  INV_X2 U11627 ( .A(n9558), .ZN(n9582) );
  NAND2_X1 U11628 ( .A1(n9582), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9060) );
  NAND2_X1 U11629 ( .A1(n9587), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9059) );
  OAI211_X1 U11630 ( .C1(n9567), .C2(n9061), .A(n9060), .B(n9059), .ZN(n9062)
         );
  AOI21_X1 U11631 ( .B1(n13615), .B2(n9428), .A(n9062), .ZN(n13462) );
  OAI22_X1 U11632 ( .A1(n13617), .A2(n6685), .B1(n9435), .B2(n13462), .ZN(
        n9418) );
  INV_X1 U11633 ( .A(n9418), .ZN(n9423) );
  NAND2_X1 U11634 ( .A1(n9814), .A2(n9579), .ZN(n9070) );
  INV_X1 U11635 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U11636 ( .A1(n9144), .A2(n9064), .ZN(n9158) );
  NAND2_X1 U11637 ( .A1(n9288), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9065) );
  MUX2_X1 U11638 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9065), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9068) );
  INV_X1 U11639 ( .A(n9288), .ZN(n9067) );
  INV_X1 U11640 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9066) );
  NAND2_X1 U11641 ( .A1(n9067), .A2(n9066), .ZN(n9196) );
  NAND2_X1 U11642 ( .A1(n9068), .A2(n9196), .ZN(n14913) );
  INV_X1 U11643 ( .A(n14913), .ZN(n9886) );
  AOI22_X1 U11644 ( .A1(n9255), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7283), .B2(
        n9886), .ZN(n9069) );
  NAND2_X1 U11645 ( .A1(n9582), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U11646 ( .A1(n9109), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9076) );
  INV_X1 U11647 ( .A(n9071), .ZN(n9164) );
  INV_X1 U11648 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11649 ( .A1(n9164), .A2(n9072), .ZN(n9073) );
  NAND2_X1 U11650 ( .A1(n9183), .A2(n9073), .ZN(n13265) );
  OR2_X1 U11651 ( .A1(n9569), .A2(n13265), .ZN(n9075) );
  NAND2_X1 U11652 ( .A1(n9587), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9074) );
  NAND4_X1 U11653 ( .A1(n9077), .A2(n9076), .A3(n9075), .A4(n9074), .ZN(n13369) );
  AOI22_X1 U11654 ( .A1(n15078), .A2(n9594), .B1(n9593), .B2(n13369), .ZN(
        n9176) );
  INV_X1 U11655 ( .A(n9617), .ZN(n9096) );
  AOI22_X1 U11656 ( .A1(n9085), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n9083) );
  INV_X1 U11657 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11658 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9079) );
  OAI21_X1 U11659 ( .B1(n9080), .B2(P2_IR_REG_30__SCAN_IN), .A(n9079), .ZN(
        n9081) );
  NAND2_X1 U11660 ( .A1(n9078), .A2(n9081), .ZN(n9082) );
  OAI21_X1 U11661 ( .B1(n9078), .B2(n9083), .A(n9082), .ZN(n9084) );
  NAND2_X1 U11662 ( .A1(n9084), .A2(n7378), .ZN(n9093) );
  AOI22_X1 U11663 ( .A1(n9085), .A2(P2_REG3_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n9089) );
  INV_X1 U11664 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U11665 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .ZN(n9086) );
  OAI21_X1 U11666 ( .B1(n9911), .B2(P2_IR_REG_30__SCAN_IN), .A(n9086), .ZN(
        n9087) );
  NAND2_X1 U11667 ( .A1(n9078), .A2(n9087), .ZN(n9088) );
  OAI21_X1 U11668 ( .B1(n9078), .B2(n9089), .A(n9088), .ZN(n9091) );
  NAND2_X1 U11669 ( .A1(n9091), .A2(n9090), .ZN(n9092) );
  INV_X1 U11670 ( .A(n11827), .ZN(n9667) );
  OAI21_X1 U11671 ( .B1(n9667), .B2(n13400), .A(n9922), .ZN(n9101) );
  NAND3_X1 U11672 ( .A1(n9095), .A2(n9661), .A3(n13375), .ZN(n9100) );
  OAI211_X1 U11673 ( .C1(n9096), .C2(n13375), .A(n9101), .B(n9100), .ZN(n9104)
         );
  NAND2_X1 U11674 ( .A1(n7845), .A2(SI_0_), .ZN(n9097) );
  XNOR2_X1 U11675 ( .A(n9097), .B(n7158), .ZN(n13840) );
  INV_X1 U11676 ( .A(n9926), .ZN(n9099) );
  NAND3_X1 U11677 ( .A1(n9099), .A2(n9095), .A3(n13375), .ZN(n9103) );
  OAI211_X1 U11678 ( .C1(n13375), .C2(n9101), .A(n9926), .B(n9100), .ZN(n9102)
         );
  NAND2_X1 U11679 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9105) );
  MUX2_X1 U11680 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9105), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9108) );
  INV_X1 U11681 ( .A(n9106), .ZN(n9107) );
  NAND2_X1 U11682 ( .A1(n9108), .A2(n9107), .ZN(n13377) );
  NAND2_X1 U11683 ( .A1(n9109), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9112) );
  INV_X1 U11684 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9110) );
  INV_X1 U11685 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13376) );
  OAI22_X1 U11686 ( .A1(n9925), .A2(n9113), .B1(n10196), .B2(n9617), .ZN(n9119) );
  NAND2_X1 U11687 ( .A1(n9115), .A2(n9114), .ZN(n9116) );
  NAND2_X1 U11688 ( .A1(n9117), .A2(n9116), .ZN(n9123) );
  INV_X1 U11689 ( .A(n9118), .ZN(n9121) );
  INV_X1 U11690 ( .A(n9119), .ZN(n9120) );
  NAND2_X1 U11691 ( .A1(n9121), .A2(n9120), .ZN(n9122) );
  NAND2_X1 U11692 ( .A1(n9428), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U11693 ( .A1(n9109), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9127) );
  INV_X1 U11694 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9124) );
  NAND4_X2 U11695 ( .A1(n9128), .A2(n9127), .A3(n9126), .A4(n9125), .ZN(n13372) );
  NOR2_X1 U11696 ( .A1(n6677), .A2(n9143), .ZN(n9129) );
  MUX2_X1 U11697 ( .A(n9143), .B(n9129), .S(P2_IR_REG_2__SCAN_IN), .Z(n9130)
         );
  INV_X1 U11698 ( .A(n9130), .ZN(n9132) );
  INV_X1 U11699 ( .A(n9144), .ZN(n9131) );
  NAND2_X1 U11700 ( .A1(n9132), .A2(n9131), .ZN(n14874) );
  AOI22_X1 U11701 ( .A1(n13372), .A2(n9593), .B1(n9974), .B2(n9170), .ZN(n9136) );
  NAND2_X1 U11702 ( .A1(n9109), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9141) );
  OR2_X1 U11703 ( .A1(n9569), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9140) );
  INV_X1 U11704 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9137) );
  OR2_X1 U11705 ( .A1(n9571), .A2(n9137), .ZN(n9139) );
  INV_X1 U11706 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9855) );
  OR2_X1 U11707 ( .A1(n9558), .A2(n9855), .ZN(n9138) );
  AND4_X2 U11708 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n10206)
         );
  NAND2_X1 U11709 ( .A1(n9063), .A2(n9767), .ZN(n9150) );
  OR2_X1 U11710 ( .A1(n9142), .A2(n9770), .ZN(n9149) );
  NOR2_X1 U11711 ( .A1(n9144), .A2(n9143), .ZN(n9145) );
  MUX2_X1 U11712 ( .A(n9143), .B(n9145), .S(P2_IR_REG_3__SCAN_IN), .Z(n9146)
         );
  INV_X1 U11713 ( .A(n9146), .ZN(n9147) );
  NAND2_X1 U11714 ( .A1(n9147), .A2(n9158), .ZN(n14887) );
  OR2_X1 U11715 ( .A1(n6690), .A2(n14887), .ZN(n9148) );
  OAI22_X1 U11716 ( .A1(n10206), .A2(n6685), .B1(n10339), .B2(n9344), .ZN(
        n9153) );
  INV_X1 U11717 ( .A(n10206), .ZN(n13371) );
  AOI22_X1 U11718 ( .A1(n9170), .A2(n13371), .B1(n10963), .B2(n9593), .ZN(
        n9151) );
  INV_X1 U11719 ( .A(n9153), .ZN(n9154) );
  NAND2_X1 U11720 ( .A1(n9792), .A2(n9063), .ZN(n9162) );
  NAND2_X1 U11721 ( .A1(n9158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9159) );
  MUX2_X1 U11722 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9159), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9160) );
  AND2_X1 U11723 ( .A1(n9160), .A2(n9288), .ZN(n9884) );
  AOI22_X1 U11724 ( .A1(n9255), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7283), .B2(
        n9884), .ZN(n9161) );
  NAND2_X1 U11725 ( .A1(n9582), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9169) );
  INV_X1 U11726 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9163) );
  OR2_X1 U11727 ( .A1(n9567), .A2(n9163), .ZN(n9168) );
  OAI21_X1 U11728 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9164), .ZN(n13293) );
  OR2_X1 U11729 ( .A1(n9586), .A2(n13293), .ZN(n9167) );
  INV_X1 U11730 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9165) );
  OR2_X1 U11731 ( .A1(n9571), .A2(n9165), .ZN(n9166) );
  INV_X1 U11732 ( .A(n9170), .ZN(n9344) );
  OAI22_X1 U11733 ( .A1(n10661), .A2(n6685), .B1(n10664), .B2(n9344), .ZN(
        n9171) );
  OAI22_X1 U11734 ( .A1(n10661), .A2(n9344), .B1(n10664), .B2(n6685), .ZN(
        n9174) );
  INV_X1 U11735 ( .A(n9171), .ZN(n9172) );
  INV_X1 U11736 ( .A(n15078), .ZN(n10798) );
  INV_X1 U11737 ( .A(n13369), .ZN(n10812) );
  OAI22_X1 U11738 ( .A1(n10798), .A2(n6685), .B1(n9435), .B2(n10812), .ZN(
        n9175) );
  NAND2_X1 U11739 ( .A1(n9820), .A2(n9063), .ZN(n9180) );
  NAND2_X1 U11740 ( .A1(n9196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9178) );
  XNOR2_X1 U11741 ( .A(n9178), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U11742 ( .A1(n9255), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7283), .B2(
        n9888), .ZN(n9179) );
  NAND2_X1 U11743 ( .A1(n9109), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9189) );
  INV_X1 U11744 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9861) );
  OR2_X1 U11745 ( .A1(n9558), .A2(n9861), .ZN(n9188) );
  INV_X1 U11746 ( .A(n9181), .ZN(n9203) );
  NAND2_X1 U11747 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  NAND2_X1 U11748 ( .A1(n9203), .A2(n9184), .ZN(n15051) );
  OR2_X1 U11749 ( .A1(n9586), .A2(n15051), .ZN(n9187) );
  INV_X1 U11750 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9185) );
  OR2_X1 U11751 ( .A1(n9571), .A2(n9185), .ZN(n9186) );
  OAI22_X1 U11752 ( .A1(n15089), .A2(n6685), .B1(n9435), .B2(n10814), .ZN(
        n9191) );
  NAND2_X1 U11753 ( .A1(n9190), .A2(n9191), .ZN(n9195) );
  OAI22_X1 U11754 ( .A1(n15089), .A2(n9344), .B1(n10814), .B2(n6685), .ZN(
        n9194) );
  INV_X1 U11755 ( .A(n9190), .ZN(n9193) );
  INV_X1 U11756 ( .A(n9191), .ZN(n9192) );
  NAND2_X1 U11757 ( .A1(n9827), .A2(n9579), .ZN(n9201) );
  INV_X1 U11758 ( .A(n9196), .ZN(n9198) );
  INV_X1 U11759 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U11760 ( .A1(n9198), .A2(n9197), .ZN(n9214) );
  NAND2_X1 U11761 ( .A1(n9214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9199) );
  XNOR2_X1 U11762 ( .A(n9199), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9890) );
  AOI22_X1 U11763 ( .A1(n9255), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7283), .B2(
        n9890), .ZN(n9200) );
  NAND2_X1 U11764 ( .A1(n9201), .A2(n9200), .ZN(n10817) );
  NAND2_X1 U11765 ( .A1(n9582), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U11766 ( .A1(n9109), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9207) );
  INV_X1 U11767 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U11768 ( .A1(n9203), .A2(n9202), .ZN(n9204) );
  NAND2_X1 U11769 ( .A1(n9222), .A2(n9204), .ZN(n10830) );
  OR2_X1 U11770 ( .A1(n9569), .A2(n10830), .ZN(n9206) );
  NAND2_X1 U11771 ( .A1(n9587), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9205) );
  NAND4_X1 U11772 ( .A1(n9208), .A2(n9207), .A3(n9206), .A4(n9205), .ZN(n13368) );
  AOI22_X1 U11773 ( .A1(n10817), .A2(n9594), .B1(n9593), .B2(n13368), .ZN(
        n9210) );
  INV_X1 U11774 ( .A(n10817), .ZN(n15096) );
  INV_X1 U11775 ( .A(n13368), .ZN(n10816) );
  OAI22_X1 U11776 ( .A1(n15096), .A2(n6685), .B1(n9435), .B2(n10816), .ZN(
        n9209) );
  OAI21_X1 U11777 ( .B1(n9211), .B2(n9210), .A(n9209), .ZN(n9213) );
  NAND2_X1 U11778 ( .A1(n9832), .A2(n9579), .ZN(n9219) );
  NAND2_X1 U11779 ( .A1(n9216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9215) );
  MUX2_X1 U11780 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9215), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9217) );
  NAND2_X1 U11781 ( .A1(n9217), .A2(n9251), .ZN(n14951) );
  INV_X1 U11782 ( .A(n14951), .ZN(n9892) );
  AOI22_X1 U11783 ( .A1(n9398), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7283), .B2(
        n9892), .ZN(n9218) );
  NAND2_X1 U11784 ( .A1(n9582), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9228) );
  INV_X1 U11785 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9220) );
  OR2_X1 U11786 ( .A1(n9567), .A2(n9220), .ZN(n9227) );
  NAND2_X1 U11787 ( .A1(n9222), .A2(n9221), .ZN(n9223) );
  NAND2_X1 U11788 ( .A1(n9237), .A2(n9223), .ZN(n10755) );
  OR2_X1 U11789 ( .A1(n9586), .A2(n10755), .ZN(n9226) );
  INV_X1 U11790 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9224) );
  OR2_X1 U11791 ( .A1(n9571), .A2(n9224), .ZN(n9225) );
  OAI22_X1 U11792 ( .A1(n15103), .A2(n9344), .B1(n10823), .B2(n6685), .ZN(
        n9231) );
  INV_X1 U11793 ( .A(n9229), .ZN(n9230) );
  NAND2_X1 U11794 ( .A1(n9837), .A2(n9579), .ZN(n9234) );
  NAND2_X1 U11795 ( .A1(n9251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9232) );
  XNOR2_X1 U11796 ( .A(n9232), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9894) );
  AOI22_X1 U11797 ( .A1(n9255), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7283), .B2(
        n9894), .ZN(n9233) );
  NAND2_X1 U11798 ( .A1(n9587), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9242) );
  INV_X1 U11799 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10805) );
  OR2_X1 U11800 ( .A1(n9558), .A2(n10805), .ZN(n9241) );
  INV_X1 U11801 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9997) );
  OR2_X1 U11802 ( .A1(n9567), .A2(n9997), .ZN(n9240) );
  INV_X1 U11803 ( .A(n9235), .ZN(n9260) );
  NAND2_X1 U11804 ( .A1(n9237), .A2(n9236), .ZN(n9238) );
  NAND2_X1 U11805 ( .A1(n9260), .A2(n9238), .ZN(n10920) );
  OR2_X1 U11806 ( .A1(n9569), .A2(n10920), .ZN(n9239) );
  OAI22_X1 U11807 ( .A1(n11120), .A2(n9344), .B1(n11115), .B2(n6685), .ZN(
        n9247) );
  NAND2_X1 U11808 ( .A1(n9243), .A2(n9247), .ZN(n9245) );
  OAI22_X1 U11809 ( .A1(n11120), .A2(n6685), .B1(n9435), .B2(n11115), .ZN(
        n9244) );
  NAND2_X1 U11810 ( .A1(n9245), .A2(n9244), .ZN(n9250) );
  INV_X1 U11811 ( .A(n9247), .ZN(n9248) );
  NAND2_X1 U11812 ( .A1(n9246), .A2(n9248), .ZN(n9249) );
  NAND2_X1 U11813 ( .A1(n9841), .A2(n9579), .ZN(n9257) );
  OAI21_X1 U11814 ( .B1(n9251), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9253) );
  INV_X1 U11815 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9252) );
  OR2_X1 U11816 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  NAND2_X1 U11817 ( .A1(n9253), .A2(n9252), .ZN(n9270) );
  AOI22_X1 U11818 ( .A1(n7283), .A2(n10002), .B1(n9398), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U11819 ( .A1(n9582), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9265) );
  NAND2_X1 U11820 ( .A1(n9109), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9264) );
  INV_X1 U11821 ( .A(n9258), .ZN(n9276) );
  INV_X1 U11822 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U11823 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  NAND2_X1 U11824 ( .A1(n9276), .A2(n9261), .ZN(n11130) );
  OR2_X1 U11825 ( .A1(n9586), .A2(n11130), .ZN(n9263) );
  NAND2_X1 U11826 ( .A1(n9587), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9262) );
  NAND4_X1 U11827 ( .A1(n9265), .A2(n9264), .A3(n9263), .A4(n9262), .ZN(n13365) );
  AOI22_X1 U11828 ( .A1(n11283), .A2(n9576), .B1(n9594), .B2(n13365), .ZN(
        n9268) );
  INV_X1 U11829 ( .A(n9268), .ZN(n9267) );
  AOI22_X1 U11830 ( .A1(n11283), .A2(n9594), .B1(n9593), .B2(n13365), .ZN(
        n9266) );
  NAND2_X1 U11831 ( .A1(n9847), .A2(n9579), .ZN(n9273) );
  NAND2_X1 U11832 ( .A1(n9270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9271) );
  XNOR2_X1 U11833 ( .A(n9271), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U11834 ( .A1(n10167), .A2(n7283), .B1(n9398), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11835 ( .A1(n9109), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9281) );
  INV_X1 U11836 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9274) );
  OR2_X1 U11837 ( .A1(n9571), .A2(n9274), .ZN(n9280) );
  INV_X1 U11838 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11839 ( .A1(n9276), .A2(n9275), .ZN(n9277) );
  NAND2_X1 U11840 ( .A1(n9294), .A2(n9277), .ZN(n11334) );
  OR2_X1 U11841 ( .A1(n9569), .A2(n11334), .ZN(n9279) );
  INV_X1 U11842 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11335) );
  OR2_X1 U11843 ( .A1(n9558), .A2(n11335), .ZN(n9278) );
  OAI22_X1 U11844 ( .A1(n11486), .A2(n6685), .B1(n9435), .B2(n11279), .ZN(
        n9284) );
  INV_X1 U11845 ( .A(n9282), .ZN(n9283) );
  NAND2_X1 U11846 ( .A1(n9918), .A2(n9579), .ZN(n9292) );
  OAI21_X1 U11847 ( .B1(n9288), .B2(n9287), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9289) );
  MUX2_X1 U11848 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9289), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9290) );
  AND2_X1 U11849 ( .A1(n9285), .A2(n9290), .ZN(n10170) );
  AOI22_X1 U11850 ( .A1(n9398), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7283), 
        .B2(n10170), .ZN(n9291) );
  NAND2_X1 U11851 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  NAND2_X1 U11852 ( .A1(n9310), .A2(n9295), .ZN(n11360) );
  OR2_X1 U11853 ( .A1(n9586), .A2(n11360), .ZN(n9299) );
  NAND2_X1 U11854 ( .A1(n9109), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U11855 ( .A1(n9587), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11856 ( .A1(n9582), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9296) );
  NAND4_X1 U11857 ( .A1(n9299), .A2(n9298), .A3(n9297), .A4(n9296), .ZN(n13363) );
  AOI22_X1 U11858 ( .A1(n11384), .A2(n9576), .B1(n9594), .B2(n13363), .ZN(
        n9302) );
  AOI22_X1 U11859 ( .A1(n11384), .A2(n9594), .B1(n9576), .B2(n13363), .ZN(
        n9300) );
  INV_X1 U11860 ( .A(n9300), .ZN(n9301) );
  NAND2_X1 U11861 ( .A1(n9305), .A2(n9304), .ZN(n9319) );
  NAND2_X1 U11862 ( .A1(n10012), .A2(n9579), .ZN(n9308) );
  NAND2_X1 U11863 ( .A1(n9285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9306) );
  XNOR2_X1 U11864 ( .A(n9306), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U11865 ( .A1(n9255), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7283), 
        .B2(n11669), .ZN(n9307) );
  NAND2_X1 U11866 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  AND2_X1 U11867 ( .A1(n9328), .A2(n9311), .ZN(n11387) );
  NAND2_X1 U11868 ( .A1(n9428), .A2(n11387), .ZN(n9316) );
  INV_X1 U11869 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11668) );
  OR2_X1 U11870 ( .A1(n9567), .A2(n11668), .ZN(n9315) );
  INV_X1 U11871 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11388) );
  OR2_X1 U11872 ( .A1(n9558), .A2(n11388), .ZN(n9314) );
  INV_X1 U11873 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9312) );
  OR2_X1 U11874 ( .A1(n9571), .A2(n9312), .ZN(n9313) );
  OAI22_X1 U11875 ( .A1(n14668), .A2(n9344), .B1(n11531), .B2(n6685), .ZN(
        n9318) );
  INV_X1 U11876 ( .A(n11531), .ZN(n13362) );
  AOI22_X1 U11877 ( .A1(n7230), .A2(n9576), .B1(n9594), .B2(n13362), .ZN(n9317) );
  NAND2_X1 U11878 ( .A1(n10244), .A2(n9579), .ZN(n9323) );
  NAND2_X1 U11879 ( .A1(n9037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9321) );
  XNOR2_X1 U11880 ( .A(n9321), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U11881 ( .A1(n9255), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7283), 
        .B2(n11673), .ZN(n9322) );
  NAND2_X1 U11882 ( .A1(n9582), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11883 ( .A1(n9109), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9324) );
  AND2_X1 U11884 ( .A1(n9325), .A2(n9324), .ZN(n9332) );
  INV_X1 U11885 ( .A(n9326), .ZN(n9339) );
  NAND2_X1 U11886 ( .A1(n9328), .A2(n9327), .ZN(n9329) );
  NAND2_X1 U11887 ( .A1(n9339), .A2(n9329), .ZN(n11551) );
  OR2_X1 U11888 ( .A1(n11551), .A2(n9569), .ZN(n9331) );
  NAND2_X1 U11889 ( .A1(n9587), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9330) );
  OAI22_X1 U11890 ( .A1(n11648), .A2(n6685), .B1(n9435), .B2(n11560), .ZN(
        n9334) );
  AOI22_X1 U11891 ( .A1(n11553), .A2(n9594), .B1(n9576), .B2(n13361), .ZN(
        n9333) );
  NAND2_X1 U11892 ( .A1(n10334), .A2(n9579), .ZN(n9338) );
  OR2_X1 U11893 ( .A1(n9335), .A2(n9143), .ZN(n9336) );
  INV_X1 U11894 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9350) );
  XNOR2_X1 U11895 ( .A(n9336), .B(n9350), .ZN(n11674) );
  INV_X1 U11896 ( .A(n11674), .ZN(n15007) );
  AOI22_X1 U11897 ( .A1(n9255), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7283), 
        .B2(n15007), .ZN(n9337) );
  INV_X1 U11898 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n13346) );
  NAND2_X1 U11899 ( .A1(n9339), .A2(n13346), .ZN(n9340) );
  NAND2_X1 U11900 ( .A1(n9356), .A2(n9340), .ZN(n11572) );
  OR2_X1 U11901 ( .A1(n11572), .A2(n9569), .ZN(n9343) );
  AOI22_X1 U11902 ( .A1(n9109), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n9582), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11903 ( .A1(n9587), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9341) );
  OAI22_X1 U11904 ( .A1(n13355), .A2(n9344), .B1(n13137), .B2(n6685), .ZN(
        n9346) );
  INV_X1 U11905 ( .A(n13137), .ZN(n13360) );
  AOI22_X1 U11906 ( .A1(n11571), .A2(n9576), .B1(n9594), .B2(n13360), .ZN(
        n9345) );
  AOI21_X1 U11907 ( .B1(n9347), .B2(n9346), .A(n9345), .ZN(n9349) );
  NAND2_X1 U11908 ( .A1(n10241), .A2(n9579), .ZN(n9355) );
  NAND2_X1 U11909 ( .A1(n9335), .A2(n9350), .ZN(n9352) );
  NAND2_X1 U11910 ( .A1(n9352), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9351) );
  MUX2_X1 U11911 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9351), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9353) );
  OR2_X1 U11912 ( .A1(n9352), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n9379) );
  AND2_X1 U11913 ( .A1(n9353), .A2(n9379), .ZN(n15023) );
  AOI22_X1 U11914 ( .A1(n9255), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7283), 
        .B2(n15023), .ZN(n9354) );
  NAND2_X1 U11915 ( .A1(n9356), .A2(n13257), .ZN(n9357) );
  AND2_X1 U11916 ( .A1(n9367), .A2(n9357), .ZN(n13254) );
  NAND2_X1 U11917 ( .A1(n13254), .A2(n9428), .ZN(n9360) );
  AOI22_X1 U11918 ( .A1(n9109), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9582), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U11919 ( .A1(n9587), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9358) );
  OAI22_X1 U11920 ( .A1(n13452), .A2(n6685), .B1(n9435), .B2(n13451), .ZN(
        n9362) );
  INV_X1 U11921 ( .A(n13451), .ZN(n13359) );
  AOI22_X1 U11922 ( .A1(n13813), .A2(n9594), .B1(n9593), .B2(n13359), .ZN(
        n9361) );
  NAND2_X1 U11923 ( .A1(n10299), .A2(n9579), .ZN(n9365) );
  NAND2_X1 U11924 ( .A1(n9379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9363) );
  XNOR2_X1 U11925 ( .A(n9363), .B(P2_IR_REG_17__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U11926 ( .A1(n9255), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7283), 
        .B2(n11678), .ZN(n9364) );
  INV_X1 U11927 ( .A(n9366), .ZN(n9385) );
  NAND2_X1 U11928 ( .A1(n9367), .A2(n13277), .ZN(n9368) );
  NAND2_X1 U11929 ( .A1(n9385), .A2(n9368), .ZN(n13275) );
  OR2_X1 U11930 ( .A1(n13275), .A2(n9569), .ZN(n9373) );
  INV_X1 U11931 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13756) );
  NAND2_X1 U11932 ( .A1(n9582), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U11933 ( .A1(n9587), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9369) );
  OAI211_X1 U11934 ( .C1(n9567), .C2(n13756), .A(n9370), .B(n9369), .ZN(n9371)
         );
  INV_X1 U11935 ( .A(n9371), .ZN(n9372) );
  OAI22_X1 U11936 ( .A1(n13810), .A2(n9435), .B1(n13455), .B2(n6685), .ZN(
        n9376) );
  INV_X1 U11937 ( .A(n13455), .ZN(n13421) );
  AOI22_X1 U11938 ( .A1(n13672), .A2(n9576), .B1(n9594), .B2(n13421), .ZN(
        n9374) );
  INV_X1 U11939 ( .A(n9375), .ZN(n9378) );
  NAND2_X1 U11940 ( .A1(n10776), .A2(n9579), .ZN(n9382) );
  OAI21_X1 U11941 ( .B1(n9379), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9380) );
  XNOR2_X1 U11942 ( .A(n9380), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U11943 ( .A1(n9255), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7283), 
        .B2(n13388), .ZN(n9381) );
  INV_X1 U11944 ( .A(n9383), .ZN(n9402) );
  INV_X1 U11945 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11946 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  AND2_X1 U11947 ( .A1(n9402), .A2(n9386), .ZN(n13654) );
  NAND2_X1 U11948 ( .A1(n13654), .A2(n9428), .ZN(n9392) );
  INV_X1 U11949 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11950 ( .A1(n9587), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U11951 ( .A1(n9109), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9387) );
  OAI211_X1 U11952 ( .C1(n9558), .C2(n9389), .A(n9388), .B(n9387), .ZN(n9390)
         );
  INV_X1 U11953 ( .A(n9390), .ZN(n9391) );
  OAI22_X1 U11954 ( .A1(n13656), .A2(n6685), .B1(n9435), .B2(n13457), .ZN(
        n9394) );
  INV_X1 U11955 ( .A(n13656), .ZN(n13749) );
  INV_X1 U11956 ( .A(n13457), .ZN(n13424) );
  AOI22_X1 U11957 ( .A1(n13749), .A2(n9594), .B1(n9593), .B2(n13424), .ZN(
        n9395) );
  OAI22_X1 U11958 ( .A1(n9396), .A2(n9395), .B1(n9394), .B2(n9393), .ZN(n9411)
         );
  NAND2_X1 U11959 ( .A1(n10906), .A2(n9579), .ZN(n9400) );
  AOI22_X1 U11960 ( .A1(n9398), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7283), 
        .B2(n9094), .ZN(n9399) );
  INV_X1 U11961 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11962 ( .A1(n9402), .A2(n9401), .ZN(n9403) );
  NAND2_X1 U11963 ( .A1(n9404), .A2(n9403), .ZN(n13638) );
  OR2_X1 U11964 ( .A1(n13638), .A2(n9569), .ZN(n9409) );
  INV_X1 U11965 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13747) );
  NAND2_X1 U11966 ( .A1(n9587), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U11967 ( .A1(n9582), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9405) );
  OAI211_X1 U11968 ( .C1(n9567), .C2(n13747), .A(n9406), .B(n9405), .ZN(n9407)
         );
  INV_X1 U11969 ( .A(n9407), .ZN(n9408) );
  OAI22_X1 U11970 ( .A1(n13804), .A2(n9435), .B1(n9626), .B2(n6685), .ZN(n9412) );
  OAI22_X1 U11971 ( .A1(n13804), .A2(n6685), .B1(n9435), .B2(n9626), .ZN(n9410) );
  INV_X1 U11972 ( .A(n9411), .ZN(n9414) );
  INV_X1 U11973 ( .A(n9412), .ZN(n9413) );
  NAND2_X1 U11974 ( .A1(n9414), .A2(n9413), .ZN(n9415) );
  NAND2_X1 U11975 ( .A1(n9419), .A2(n9418), .ZN(n9421) );
  INV_X1 U11976 ( .A(n9438), .ZN(n9434) );
  NAND2_X1 U11977 ( .A1(n11341), .A2(n9579), .ZN(n9425) );
  NAND2_X1 U11978 ( .A1(n9398), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9424) );
  OR2_X1 U11979 ( .A1(n9426), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9427) );
  AND2_X1 U11980 ( .A1(n9446), .A2(n9427), .ZN(n13605) );
  NAND2_X1 U11981 ( .A1(n13605), .A2(n9428), .ZN(n9433) );
  INV_X1 U11982 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13738) );
  NAND2_X1 U11983 ( .A1(n9582), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U11984 ( .A1(n9587), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9429) );
  OAI211_X1 U11985 ( .C1(n9567), .C2(n13738), .A(n9430), .B(n9429), .ZN(n9431)
         );
  INV_X1 U11986 ( .A(n9431), .ZN(n9432) );
  OAI22_X1 U11987 ( .A1(n13799), .A2(n9435), .B1(n13465), .B2(n6685), .ZN(
        n9436) );
  NAND2_X1 U11988 ( .A1(n9434), .A2(n9436), .ZN(n9441) );
  OAI22_X1 U11989 ( .A1(n13799), .A2(n6685), .B1(n9435), .B2(n13465), .ZN(
        n9440) );
  INV_X1 U11990 ( .A(n9436), .ZN(n9437) );
  XNOR2_X1 U11991 ( .A(n9443), .B(n7642), .ZN(n11826) );
  NAND2_X1 U11992 ( .A1(n11826), .A2(n9579), .ZN(n9445) );
  NAND2_X1 U11993 ( .A1(n9398), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9444) );
  INV_X1 U11994 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13313) );
  NAND2_X1 U11995 ( .A1(n9446), .A2(n13313), .ZN(n9448) );
  INV_X1 U11996 ( .A(n9462), .ZN(n9447) );
  NAND2_X1 U11997 ( .A1(n9448), .A2(n9447), .ZN(n13311) );
  OR2_X1 U11998 ( .A1(n13311), .A2(n9569), .ZN(n9454) );
  INV_X1 U11999 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U12000 ( .A1(n9587), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9450) );
  NAND2_X1 U12001 ( .A1(n9582), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9449) );
  OAI211_X1 U12002 ( .C1(n9567), .C2(n9451), .A(n9450), .B(n9449), .ZN(n9452)
         );
  INV_X1 U12003 ( .A(n9452), .ZN(n9453) );
  NAND2_X1 U12004 ( .A1(n9454), .A2(n9453), .ZN(n13467) );
  AOI22_X1 U12005 ( .A1(n13730), .A2(n9576), .B1(n9594), .B2(n13467), .ZN(
        n9456) );
  INV_X1 U12006 ( .A(n13730), .ZN(n13595) );
  INV_X1 U12007 ( .A(n13467), .ZN(n13435) );
  OAI22_X1 U12008 ( .A1(n13595), .A2(n9435), .B1(n13435), .B2(n6685), .ZN(
        n9455) );
  OAI21_X1 U12009 ( .B1(n9457), .B2(n9456), .A(n9455), .ZN(n9459) );
  NAND2_X1 U12010 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  NAND2_X1 U12011 ( .A1(n11432), .A2(n9579), .ZN(n9461) );
  NAND2_X1 U12012 ( .A1(n9398), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U12013 ( .A1(n9109), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9466) );
  INV_X1 U12014 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13792) );
  OR2_X1 U12015 ( .A1(n9571), .A2(n13792), .ZN(n9465) );
  NAND2_X1 U12016 ( .A1(n9462), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9469) );
  OAI21_X1 U12017 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n9462), .A(n9469), .ZN(
        n13211) );
  OR2_X1 U12018 ( .A1(n9586), .A2(n13211), .ZN(n9464) );
  INV_X1 U12019 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13576) );
  OR2_X1 U12020 ( .A1(n9558), .A2(n13576), .ZN(n9463) );
  OAI22_X1 U12021 ( .A1(n13794), .A2(n9435), .B1(n13469), .B2(n6685), .ZN(
        n9504) );
  NAND2_X1 U12022 ( .A1(n11635), .A2(n9579), .ZN(n9468) );
  NAND2_X1 U12023 ( .A1(n9398), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U12024 ( .A1(n9109), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9475) );
  INV_X1 U12025 ( .A(n9469), .ZN(n9471) );
  INV_X1 U12026 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13285) );
  INV_X1 U12027 ( .A(n9493), .ZN(n9470) );
  OAI21_X1 U12028 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n9471), .A(n9470), .ZN(
        n13284) );
  OR2_X1 U12029 ( .A1(n9586), .A2(n13284), .ZN(n9474) );
  NAND2_X1 U12030 ( .A1(n9587), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U12031 ( .A1(n9582), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9472) );
  NAND4_X1 U12032 ( .A1(n9475), .A2(n9474), .A3(n9473), .A4(n9472), .ZN(n13473) );
  AND2_X1 U12033 ( .A1(n13473), .A2(n9593), .ZN(n9476) );
  AOI21_X1 U12034 ( .B1(n13718), .B2(n9594), .A(n9476), .ZN(n9529) );
  NAND2_X1 U12035 ( .A1(n13718), .A2(n9593), .ZN(n9478) );
  NAND2_X1 U12036 ( .A1(n13473), .A2(n9594), .ZN(n9477) );
  NAND2_X1 U12037 ( .A1(n9478), .A2(n9477), .ZN(n9528) );
  NAND2_X1 U12038 ( .A1(n13832), .A2(n9579), .ZN(n9480) );
  NAND2_X1 U12039 ( .A1(n9398), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U12040 ( .A1(n9109), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9487) );
  NAND3_X1 U12041 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .A3(n9493), .ZN(n9509) );
  INV_X1 U12042 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U12043 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(n9493), .ZN(n9481) );
  NAND2_X1 U12044 ( .A1(n9482), .A2(n9481), .ZN(n9483) );
  NAND2_X1 U12045 ( .A1(n9509), .A2(n9483), .ZN(n13531) );
  OR2_X1 U12046 ( .A1(n9586), .A2(n13531), .ZN(n9486) );
  NAND2_X1 U12047 ( .A1(n9582), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U12048 ( .A1(n9587), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9484) );
  NAND4_X1 U12049 ( .A1(n9487), .A2(n9486), .A3(n9485), .A4(n9484), .ZN(n13476) );
  AND2_X1 U12050 ( .A1(n13476), .A2(n9593), .ZN(n9488) );
  AOI21_X1 U12051 ( .B1(n13707), .B2(n9594), .A(n9488), .ZN(n9523) );
  NAND2_X1 U12052 ( .A1(n13707), .A2(n9593), .ZN(n9490) );
  NAND2_X1 U12053 ( .A1(n13476), .A2(n9594), .ZN(n9489) );
  NAND2_X1 U12054 ( .A1(n9490), .A2(n9489), .ZN(n9522) );
  NAND2_X1 U12055 ( .A1(n9523), .A2(n9522), .ZN(n9527) );
  NAND2_X1 U12056 ( .A1(n11821), .A2(n9579), .ZN(n9492) );
  NAND2_X1 U12057 ( .A1(n9398), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9491) );
  NAND2_X2 U12058 ( .A1(n9492), .A2(n9491), .ZN(n13788) );
  NAND2_X1 U12059 ( .A1(n9109), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9497) );
  XNOR2_X1 U12060 ( .A(P2_REG3_REG_25__SCAN_IN), .B(n9493), .ZN(n13550) );
  OR2_X1 U12061 ( .A1(n9569), .A2(n13550), .ZN(n9496) );
  NAND2_X1 U12062 ( .A1(n9587), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U12063 ( .A1(n9582), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9494) );
  NAND4_X1 U12064 ( .A1(n9497), .A2(n9496), .A3(n9495), .A4(n9494), .ZN(n13475) );
  AND2_X1 U12065 ( .A1(n13475), .A2(n9593), .ZN(n9498) );
  AOI21_X1 U12066 ( .B1(n13788), .B2(n9594), .A(n9498), .ZN(n9519) );
  NAND2_X1 U12067 ( .A1(n13788), .A2(n9576), .ZN(n9500) );
  NAND2_X1 U12068 ( .A1(n13475), .A2(n9594), .ZN(n9499) );
  NAND2_X1 U12069 ( .A1(n9500), .A2(n9499), .ZN(n9518) );
  NAND2_X1 U12070 ( .A1(n9519), .A2(n9518), .ZN(n9501) );
  NAND2_X1 U12071 ( .A1(n9527), .A2(n9501), .ZN(n9530) );
  AOI21_X1 U12072 ( .B1(n9529), .B2(n9528), .A(n9530), .ZN(n9502) );
  INV_X1 U12073 ( .A(n13469), .ZN(n13470) );
  AOI22_X1 U12074 ( .A1(n13471), .A2(n9576), .B1(n9594), .B2(n13470), .ZN(
        n9503) );
  NAND2_X1 U12075 ( .A1(n9398), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9505) );
  NAND2_X1 U12076 ( .A1(n9582), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U12077 ( .A1(n9109), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9513) );
  INV_X1 U12078 ( .A(n9509), .ZN(n9507) );
  NAND2_X1 U12079 ( .A1(n9507), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9584) );
  INV_X1 U12080 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9508) );
  NAND2_X1 U12081 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  NAND2_X1 U12082 ( .A1(n9584), .A2(n9510), .ZN(n13520) );
  OR2_X1 U12083 ( .A1(n9586), .A2(n13520), .ZN(n9512) );
  NAND2_X1 U12084 ( .A1(n9587), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9511) );
  NAND4_X1 U12085 ( .A1(n9514), .A2(n9513), .A3(n9512), .A4(n9511), .ZN(n13358) );
  AND2_X1 U12086 ( .A1(n13358), .A2(n9593), .ZN(n9515) );
  AOI21_X1 U12087 ( .B1(n13522), .B2(n9594), .A(n9515), .ZN(n9598) );
  NAND2_X1 U12088 ( .A1(n13522), .A2(n9593), .ZN(n9517) );
  NAND2_X1 U12089 ( .A1(n13358), .A2(n9594), .ZN(n9516) );
  NAND2_X1 U12090 ( .A1(n9517), .A2(n9516), .ZN(n9597) );
  INV_X1 U12091 ( .A(n9518), .ZN(n9521) );
  INV_X1 U12092 ( .A(n9519), .ZN(n9520) );
  AND2_X1 U12093 ( .A1(n9521), .A2(n9520), .ZN(n9526) );
  INV_X1 U12094 ( .A(n9522), .ZN(n9525) );
  INV_X1 U12095 ( .A(n9523), .ZN(n9524) );
  AOI22_X1 U12096 ( .A1(n9527), .A2(n9526), .B1(n9525), .B2(n9524), .ZN(n9532)
         );
  OR3_X1 U12097 ( .A1(n9530), .A2(n9529), .A3(n9528), .ZN(n9531) );
  OAI211_X1 U12098 ( .C1(n9598), .C2(n9597), .A(n9532), .B(n9531), .ZN(n9533)
         );
  INV_X1 U12099 ( .A(n9533), .ZN(n9534) );
  INV_X1 U12100 ( .A(n9537), .ZN(n9538) );
  NAND2_X1 U12101 ( .A1(n9538), .A2(n13129), .ZN(n9539) );
  MUX2_X1 U12102 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9773), .Z(n9541) );
  NAND2_X1 U12103 ( .A1(n9541), .A2(SI_30_), .ZN(n9542) );
  OAI21_X1 U12104 ( .B1(SI_30_), .B2(n9541), .A(n9542), .ZN(n9551) );
  MUX2_X1 U12105 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9773), .Z(n9543) );
  XNOR2_X1 U12106 ( .A(n9543), .B(SI_31_), .ZN(n9544) );
  NAND2_X1 U12107 ( .A1(n13816), .A2(n9579), .ZN(n9547) );
  NAND2_X1 U12108 ( .A1(n9398), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9546) );
  INV_X1 U12109 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13684) );
  NAND2_X1 U12110 ( .A1(n9582), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U12111 ( .A1(n9587), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9548) );
  OAI211_X1 U12112 ( .C1(n9567), .C2(n13684), .A(n9549), .B(n9548), .ZN(n13410) );
  INV_X1 U12113 ( .A(n13410), .ZN(n9550) );
  OAI22_X1 U12114 ( .A1(n13771), .A2(n9435), .B1(n9550), .B2(n6685), .ZN(n9578) );
  NAND2_X1 U12115 ( .A1(n9552), .A2(n9551), .ZN(n9553) );
  NAND2_X1 U12116 ( .A1(n9398), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9556) );
  INV_X1 U12117 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13688) );
  OR2_X1 U12118 ( .A1(n9567), .A2(n13688), .ZN(n9561) );
  INV_X1 U12119 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13415) );
  OR2_X1 U12120 ( .A1(n9558), .A2(n13415), .ZN(n9560) );
  INV_X1 U12121 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13773) );
  OR2_X1 U12122 ( .A1(n9571), .A2(n13773), .ZN(n9559) );
  AND3_X1 U12123 ( .A1(n9561), .A2(n9560), .A3(n9559), .ZN(n13449) );
  OAI22_X1 U12124 ( .A1(n13775), .A2(n9435), .B1(n13449), .B2(n6685), .ZN(
        n9610) );
  INV_X1 U12125 ( .A(n13449), .ZN(n13356) );
  NAND2_X1 U12126 ( .A1(n13410), .A2(n9594), .ZN(n9616) );
  NAND2_X1 U12127 ( .A1(n13400), .A2(n11268), .ZN(n9957) );
  NAND2_X1 U12128 ( .A1(n10460), .A2(n9667), .ZN(n9622) );
  NAND4_X1 U12129 ( .A1(n9616), .A2(n9661), .A3(n9957), .A4(n9622), .ZN(n9563)
         );
  AOI22_X1 U12130 ( .A1(n13418), .A2(n9576), .B1(n13356), .B2(n9563), .ZN(
        n9609) );
  NAND2_X1 U12131 ( .A1(n13823), .A2(n9579), .ZN(n9565) );
  NAND2_X1 U12132 ( .A1(n9398), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U12133 ( .A1(n9582), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9575) );
  INV_X1 U12134 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9566) );
  OR2_X1 U12135 ( .A1(n9567), .A2(n9566), .ZN(n9574) );
  INV_X1 U12136 ( .A(n9584), .ZN(n9568) );
  NAND2_X1 U12137 ( .A1(n9568), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13489) );
  OR2_X1 U12138 ( .A1(n9569), .A2(n13489), .ZN(n9573) );
  INV_X1 U12139 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9570) );
  OR2_X1 U12140 ( .A1(n9571), .A2(n9570), .ZN(n9572) );
  AOI22_X1 U12141 ( .A1(n13491), .A2(n9576), .B1(n9594), .B2(n13357), .ZN(
        n9601) );
  OAI22_X1 U12142 ( .A1(n13692), .A2(n9435), .B1(n13230), .B2(n6685), .ZN(
        n9602) );
  OAI22_X1 U12143 ( .A1(n9610), .A2(n9609), .B1(n9601), .B2(n9602), .ZN(n9577)
         );
  OAI21_X1 U12144 ( .B1(n9578), .B2(n9614), .A(n9577), .ZN(n9607) );
  NAND2_X1 U12145 ( .A1(n13825), .A2(n9579), .ZN(n9581) );
  NAND2_X1 U12146 ( .A1(n9398), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9580) );
  NAND2_X1 U12147 ( .A1(n9582), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U12148 ( .A1(n9109), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9590) );
  INV_X1 U12149 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U12150 ( .A1(n9584), .A2(n9583), .ZN(n9585) );
  NAND2_X1 U12151 ( .A1(n13489), .A2(n9585), .ZN(n13504) );
  OR2_X1 U12152 ( .A1(n9586), .A2(n13504), .ZN(n9589) );
  NAND2_X1 U12153 ( .A1(n9587), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9588) );
  NAND4_X1 U12154 ( .A1(n9591), .A2(n9590), .A3(n9589), .A4(n9588), .ZN(n13482) );
  AND2_X1 U12155 ( .A1(n13482), .A2(n9593), .ZN(n9592) );
  AOI21_X1 U12156 ( .B1(n13503), .B2(n9594), .A(n9592), .ZN(n9604) );
  NAND2_X1 U12157 ( .A1(n13503), .A2(n9593), .ZN(n9596) );
  NAND2_X1 U12158 ( .A1(n13482), .A2(n9594), .ZN(n9595) );
  NAND2_X1 U12159 ( .A1(n9596), .A2(n9595), .ZN(n9603) );
  NAND2_X1 U12160 ( .A1(n9604), .A2(n9603), .ZN(n9600) );
  NAND2_X1 U12161 ( .A1(n9598), .A2(n9597), .ZN(n9599) );
  INV_X1 U12162 ( .A(n9601), .ZN(n9606) );
  INV_X1 U12163 ( .A(n9602), .ZN(n9605) );
  OAI22_X1 U12164 ( .A1(n9606), .A2(n9605), .B1(n9604), .B2(n9603), .ZN(n9608)
         );
  OAI21_X1 U12165 ( .B1(n9641), .B2(n9608), .A(n9607), .ZN(n9612) );
  INV_X1 U12166 ( .A(n9614), .ZN(n9615) );
  INV_X1 U12167 ( .A(n9922), .ZN(n9924) );
  NAND2_X1 U12168 ( .A1(n9661), .A2(n13400), .ZN(n9620) );
  OAI211_X1 U12169 ( .C1(n9924), .C2(n9667), .A(n9957), .B(n9620), .ZN(n9621)
         );
  INV_X1 U12170 ( .A(n11268), .ZN(n9963) );
  NAND2_X1 U12171 ( .A1(n9661), .A2(n9963), .ZN(n10047) );
  OAI21_X1 U12172 ( .B1(n10047), .B2(n13400), .A(n9622), .ZN(n9623) );
  XNOR2_X1 U12173 ( .A(n13418), .B(n13356), .ZN(n9640) );
  NAND2_X1 U12174 ( .A1(n13503), .A2(n13447), .ZN(n9624) );
  INV_X1 U12175 ( .A(n13476), .ZN(n9625) );
  OR2_X1 U12176 ( .A1(n13707), .A2(n9625), .ZN(n13441) );
  NAND2_X1 U12177 ( .A1(n13707), .A2(n9625), .ZN(n13442) );
  NAND2_X1 U12178 ( .A1(n13441), .A2(n13442), .ZN(n13535) );
  INV_X1 U12179 ( .A(n13475), .ZN(n13440) );
  XNOR2_X1 U12180 ( .A(n13788), .B(n13440), .ZN(n13545) );
  INV_X1 U12181 ( .A(n13473), .ZN(n13438) );
  XNOR2_X1 U12182 ( .A(n13471), .B(n13469), .ZN(n13579) );
  NAND2_X1 U12183 ( .A1(n13741), .A2(n13462), .ZN(n13429) );
  NAND2_X1 U12184 ( .A1(n13637), .A2(n13428), .ZN(n13458) );
  XNOR2_X1 U12185 ( .A(n13749), .B(n13457), .ZN(n13646) );
  NAND2_X1 U12186 ( .A1(n13813), .A2(n13451), .ZN(n9627) );
  NAND2_X1 U12187 ( .A1(n13664), .A2(n9627), .ZN(n11700) );
  XNOR2_X1 U12188 ( .A(n7230), .B(n13362), .ZN(n11386) );
  INV_X1 U12189 ( .A(n13365), .ZN(n11275) );
  XNOR2_X1 U12190 ( .A(n11283), .B(n11275), .ZN(n11121) );
  INV_X1 U12191 ( .A(n11120), .ZN(n10809) );
  INV_X1 U12192 ( .A(n11115), .ZN(n13366) );
  XNOR2_X1 U12193 ( .A(n10809), .B(n13366), .ZN(n10821) );
  INV_X1 U12194 ( .A(n15089), .ZN(n15054) );
  XNOR2_X1 U12195 ( .A(n15078), .B(n13369), .ZN(n10810) );
  NAND2_X1 U12196 ( .A1(n9099), .A2(n13375), .ZN(n10178) );
  INV_X1 U12197 ( .A(n13375), .ZN(n9628) );
  NAND2_X1 U12198 ( .A1(n9926), .A2(n9628), .ZN(n9629) );
  NAND2_X1 U12199 ( .A1(n10178), .A2(n9629), .ZN(n10469) );
  AND4_X1 U12200 ( .A1(n10214), .A2(n10182), .A3(n9963), .A4(n10469), .ZN(
        n9630) );
  INV_X1 U12201 ( .A(n10661), .ZN(n13295) );
  INV_X1 U12202 ( .A(n10664), .ZN(n13370) );
  XNOR2_X1 U12203 ( .A(n13295), .B(n13370), .ZN(n10659) );
  XNOR2_X1 U12204 ( .A(n13371), .B(n10963), .ZN(n10203) );
  NAND4_X1 U12205 ( .A1(n10810), .A2(n9630), .A3(n10659), .A4(n10203), .ZN(
        n9631) );
  NOR2_X1 U12206 ( .A1(n10801), .A2(n9631), .ZN(n9632) );
  INV_X1 U12207 ( .A(n10823), .ZN(n13367) );
  XNOR2_X1 U12208 ( .A(n10850), .B(n13367), .ZN(n10852) );
  XNOR2_X1 U12209 ( .A(n10817), .B(n13368), .ZN(n10815) );
  NAND4_X1 U12210 ( .A1(n10821), .A2(n9632), .A3(n10852), .A4(n10815), .ZN(
        n9633) );
  NOR2_X1 U12211 ( .A1(n11121), .A2(n9633), .ZN(n9634) );
  XNOR2_X1 U12212 ( .A(n11489), .B(n13364), .ZN(n11327) );
  XNOR2_X1 U12213 ( .A(n11384), .B(n13363), .ZN(n11288) );
  NAND4_X1 U12214 ( .A1(n11386), .A2(n9634), .A3(n11327), .A4(n11288), .ZN(
        n9635) );
  NOR2_X1 U12215 ( .A1(n11700), .A2(n9635), .ZN(n9636) );
  XNOR2_X1 U12216 ( .A(n11553), .B(n13361), .ZN(n11541) );
  XNOR2_X1 U12217 ( .A(n13672), .B(n13421), .ZN(n13662) );
  NAND4_X1 U12218 ( .A1(n11688), .A2(n9636), .A3(n11541), .A4(n13662), .ZN(
        n9637) );
  XNOR2_X1 U12219 ( .A(n13730), .B(n13435), .ZN(n13588) );
  INV_X1 U12220 ( .A(n13799), .ZN(n13237) );
  XNOR2_X1 U12221 ( .A(n13237), .B(n13465), .ZN(n13602) );
  NOR2_X1 U12222 ( .A1(n13481), .A2(n9638), .ZN(n9639) );
  INV_X1 U12223 ( .A(n9661), .ZN(n11342) );
  NAND2_X1 U12224 ( .A1(n9645), .A2(n9644), .ZN(n9651) );
  NAND2_X1 U12225 ( .A1(n9651), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9647) );
  INV_X1 U12226 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9646) );
  XNOR2_X1 U12227 ( .A(n9647), .B(n9646), .ZN(n9960) );
  INV_X1 U12228 ( .A(n9960), .ZN(n9648) );
  AND2_X1 U12229 ( .A1(n9648), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11395) );
  INV_X1 U12230 ( .A(n11395), .ZN(n9666) );
  XNOR2_X1 U12231 ( .A(n9650), .B(n9649), .ZN(n13834) );
  INV_X1 U12232 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9652) );
  NAND2_X1 U12233 ( .A1(n9653), .A2(n9652), .ZN(n9658) );
  NAND2_X1 U12234 ( .A1(n9658), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9655) );
  XNOR2_X1 U12235 ( .A(n9655), .B(n9654), .ZN(n13835) );
  NAND2_X1 U12236 ( .A1(n9656), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9657) );
  MUX2_X1 U12237 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9657), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9659) );
  NAND2_X1 U12238 ( .A1(n9659), .A2(n9658), .ZN(n11636) );
  NOR3_X1 U12239 ( .A1(n13834), .A2(n13835), .A3(n11636), .ZN(n9677) );
  INV_X1 U12240 ( .A(n9677), .ZN(n9959) );
  AND2_X1 U12241 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9959), .ZN(n9660) );
  INV_X1 U12242 ( .A(n9957), .ZN(n9948) );
  INV_X1 U12243 ( .A(n9662), .ZN(n9873) );
  OAI21_X1 U12244 ( .B1(n9663), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9664) );
  XNOR2_X1 U12245 ( .A(n9664), .B(P2_IR_REG_27__SCAN_IN), .ZN(n13830) );
  NAND4_X1 U12246 ( .A1(n15072), .A2(n9948), .A3(n13331), .A4(n13830), .ZN(
        n9665) );
  OAI211_X1 U12247 ( .C1(n9667), .C2(n9666), .A(n9665), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9668) );
  NAND2_X1 U12248 ( .A1(n9669), .A2(n9668), .ZN(P2_U3328) );
  INV_X1 U12249 ( .A(n10881), .ZN(n9670) );
  NAND2_X1 U12250 ( .A1(n9672), .A2(n14857), .ZN(n9675) );
  NAND2_X1 U12251 ( .A1(n9673), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U12252 ( .A1(n9675), .A2(n9674), .ZN(P1_U3525) );
  INV_X1 U12253 ( .A(n9909), .ZN(n9676) );
  NOR2_X1 U12254 ( .A1(n10259), .A2(n9676), .ZN(P1_U4016) );
  NAND2_X1 U12255 ( .A1(n9960), .A2(n9677), .ZN(n9871) );
  INV_X1 U12256 ( .A(n13115), .ZN(n11797) );
  NAND2_X1 U12257 ( .A1(n9813), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9686) );
  OAI21_X1 U12258 ( .B1(n9813), .B2(P3_REG2_REG_6__SCAN_IN), .A(n9686), .ZN(
        n10578) );
  NAND2_X1 U12259 ( .A1(n9678), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9680) );
  OAI21_X1 U12260 ( .B1(n9783), .B2(n9679), .A(n9680), .ZN(n10397) );
  NAND2_X1 U12261 ( .A1(n10399), .A2(n9680), .ZN(n10691) );
  OR2_X1 U12262 ( .A1(n9719), .A2(n15319), .ZN(n9681) );
  NAND2_X1 U12263 ( .A1(n10690), .A2(n9681), .ZN(n9682) );
  NAND2_X1 U12264 ( .A1(n9682), .A2(n9778), .ZN(n10533) );
  NAND2_X1 U12265 ( .A1(n10533), .A2(n9683), .ZN(n10593) );
  XNOR2_X1 U12266 ( .A(n9728), .B(n11157), .ZN(n10534) );
  NOR2_X1 U12267 ( .A1(n9685), .A2(n10560), .ZN(n10579) );
  INV_X1 U12268 ( .A(n9686), .ZN(n9687) );
  NOR2_X1 U12269 ( .A1(n10577), .A2(n9687), .ZN(n9688) );
  NOR2_X1 U12270 ( .A1(n9745), .A2(n9688), .ZN(n9689) );
  NAND2_X1 U12271 ( .A1(n9804), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11061) );
  OAI21_X1 U12272 ( .B1(n9804), .B2(P3_REG2_REG_8__SCAN_IN), .A(n11061), .ZN(
        n9690) );
  NAND2_X1 U12273 ( .A1(n9691), .A2(n9690), .ZN(n9696) );
  INV_X1 U12274 ( .A(n10283), .ZN(n9693) );
  OAI21_X1 U12275 ( .B1(n11967), .B2(n9693), .A(n9692), .ZN(n9759) );
  OR2_X1 U12276 ( .A1(n10283), .A2(P3_U3151), .ZN(n12007) );
  AND2_X1 U12277 ( .A1(n10476), .A2(n12007), .ZN(n9757) );
  OR2_X1 U12278 ( .A1(n9759), .A2(n9757), .ZN(n9708) );
  INV_X1 U12279 ( .A(n9708), .ZN(n9756) );
  INV_X1 U12280 ( .A(n9694), .ZN(n9695) );
  NAND2_X1 U12281 ( .A1(n9756), .A2(n9695), .ZN(n15266) );
  AOI21_X1 U12282 ( .B1(n11062), .B2(n9696), .A(n15266), .ZN(n9765) );
  NAND2_X1 U12283 ( .A1(n9813), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9702) );
  OAI21_X1 U12284 ( .B1(n9813), .B2(P3_REG1_REG_6__SCAN_IN), .A(n9702), .ZN(
        n10582) );
  XNOR2_X1 U12285 ( .A(n9719), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n10695) );
  NAND2_X1 U12286 ( .A1(n10695), .A2(n10694), .ZN(n10693) );
  OR2_X1 U12287 ( .A1(n9719), .A2(n9717), .ZN(n9697) );
  NAND2_X1 U12288 ( .A1(n10693), .A2(n9697), .ZN(n9698) );
  NAND2_X1 U12289 ( .A1(n9698), .A2(n9778), .ZN(n10527) );
  NAND2_X1 U12290 ( .A1(n10527), .A2(n9699), .ZN(n10596) );
  OR2_X2 U12291 ( .A1(n10596), .A2(n9723), .ZN(n10598) );
  XNOR2_X1 U12292 ( .A(n9728), .B(n15386), .ZN(n10528) );
  NOR2_X1 U12293 ( .A1(n9700), .A2(n10570), .ZN(n9701) );
  INV_X1 U12294 ( .A(n9702), .ZN(n9703) );
  NOR2_X1 U12295 ( .A1(n9745), .A2(n9704), .ZN(n9705) );
  NAND2_X1 U12296 ( .A1(n9804), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11072) );
  OAI21_X1 U12297 ( .B1(n9804), .B2(P3_REG1_REG_8__SCAN_IN), .A(n11072), .ZN(
        n9706) );
  NAND2_X1 U12298 ( .A1(n9707), .A2(n9706), .ZN(n9709) );
  NOR2_X1 U12299 ( .A1(n9708), .A2(n12651), .ZN(n15262) );
  AOI21_X1 U12300 ( .B1(n11073), .B2(n9709), .A(n15241), .ZN(n9764) );
  MUX2_X1 U12301 ( .A(n9711), .B(n9710), .S(n6684), .Z(n9712) );
  INV_X1 U12302 ( .A(n9783), .ZN(n10403) );
  NAND2_X1 U12303 ( .A1(n9712), .A2(n10403), .ZN(n10701) );
  INV_X1 U12304 ( .A(n9712), .ZN(n9713) );
  NAND2_X1 U12305 ( .A1(n9713), .A2(n9783), .ZN(n9714) );
  NAND2_X1 U12306 ( .A1(n10701), .A2(n9714), .ZN(n10393) );
  INV_X1 U12307 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9715) );
  INV_X4 U12308 ( .A(n12651), .ZN(n12735) );
  MUX2_X1 U12309 ( .A(n9716), .B(n9715), .S(n12735), .Z(n15162) );
  NAND2_X1 U12310 ( .A1(n10392), .A2(n10701), .ZN(n9722) );
  MUX2_X1 U12311 ( .A(n15319), .B(n9717), .S(n12735), .Z(n9718) );
  NAND2_X1 U12312 ( .A1(n9718), .A2(n9719), .ZN(n10606) );
  INV_X1 U12313 ( .A(n9718), .ZN(n9720) );
  INV_X1 U12314 ( .A(n9719), .ZN(n10710) );
  NAND2_X1 U12315 ( .A1(n9720), .A2(n10710), .ZN(n9721) );
  AND2_X1 U12316 ( .A1(n10606), .A2(n9721), .ZN(n10702) );
  NAND2_X1 U12317 ( .A1(n9722), .A2(n10702), .ZN(n10705) );
  NAND2_X1 U12318 ( .A1(n10705), .A2(n10606), .ZN(n9727) );
  MUX2_X1 U12319 ( .A(n11018), .B(n9723), .S(n12735), .Z(n9724) );
  NAND2_X1 U12320 ( .A1(n9724), .A2(n10611), .ZN(n10542) );
  INV_X1 U12321 ( .A(n9724), .ZN(n9725) );
  NAND2_X1 U12322 ( .A1(n9725), .A2(n9778), .ZN(n9726) );
  AND2_X1 U12323 ( .A1(n10542), .A2(n9726), .ZN(n10604) );
  NAND2_X1 U12324 ( .A1(n10608), .A2(n10542), .ZN(n9732) );
  MUX2_X1 U12325 ( .A(n11157), .B(n15386), .S(n12735), .Z(n9729) );
  NAND2_X1 U12326 ( .A1(n9729), .A2(n9728), .ZN(n10557) );
  INV_X1 U12327 ( .A(n9729), .ZN(n9730) );
  NAND2_X1 U12328 ( .A1(n9730), .A2(n10539), .ZN(n9731) );
  AND2_X1 U12329 ( .A1(n10557), .A2(n9731), .ZN(n10540) );
  NAND2_X1 U12330 ( .A1(n9732), .A2(n10540), .ZN(n10558) );
  NAND2_X1 U12331 ( .A1(n10558), .A2(n10557), .ZN(n9738) );
  MUX2_X1 U12332 ( .A(n9734), .B(n9733), .S(n12735), .Z(n9735) );
  NAND2_X1 U12333 ( .A1(n9735), .A2(n10570), .ZN(n10574) );
  INV_X1 U12334 ( .A(n9735), .ZN(n9736) );
  NAND2_X1 U12335 ( .A1(n9736), .A2(n9774), .ZN(n9737) );
  AND2_X1 U12336 ( .A1(n10574), .A2(n9737), .ZN(n10555) );
  NAND2_X1 U12337 ( .A1(n10575), .A2(n10574), .ZN(n9742) );
  MUX2_X1 U12338 ( .A(n15297), .B(n15389), .S(n12735), .Z(n9739) );
  INV_X1 U12339 ( .A(n9813), .ZN(n10591) );
  NAND2_X1 U12340 ( .A1(n9739), .A2(n10591), .ZN(n10634) );
  INV_X1 U12341 ( .A(n9739), .ZN(n9740) );
  NAND2_X1 U12342 ( .A1(n9740), .A2(n9813), .ZN(n9741) );
  AND2_X1 U12343 ( .A1(n10634), .A2(n9741), .ZN(n10572) );
  NAND2_X1 U12344 ( .A1(n9742), .A2(n10572), .ZN(n10635) );
  NAND2_X1 U12345 ( .A1(n10635), .A2(n10634), .ZN(n9749) );
  MUX2_X1 U12346 ( .A(n9744), .B(n9743), .S(n12735), .Z(n9746) );
  NAND2_X1 U12347 ( .A1(n9746), .A2(n9745), .ZN(n9752) );
  INV_X1 U12348 ( .A(n9746), .ZN(n9747) );
  NAND2_X1 U12349 ( .A1(n9747), .A2(n10631), .ZN(n9748) );
  AND2_X1 U12350 ( .A1(n9752), .A2(n9748), .ZN(n10632) );
  NAND2_X1 U12351 ( .A1(n10637), .A2(n9752), .ZN(n9750) );
  MUX2_X1 U12352 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12735), .Z(n11053) );
  INV_X1 U12353 ( .A(n9804), .ZN(n11054) );
  XNOR2_X1 U12354 ( .A(n11053), .B(n11054), .ZN(n9751) );
  INV_X1 U12355 ( .A(n9751), .ZN(n9753) );
  NAND3_X1 U12356 ( .A1(n10637), .A2(n9753), .A3(n9752), .ZN(n9754) );
  NAND2_X1 U12357 ( .A1(n10958), .A2(n8926), .ZN(n15253) );
  AOI21_X1 U12358 ( .B1(n11057), .B2(n9754), .A(n15253), .ZN(n9763) );
  MUX2_X1 U12359 ( .A(n9756), .B(P3_U3897), .S(n9755), .Z(n15259) );
  INV_X1 U12360 ( .A(n15259), .ZN(n15235) );
  INV_X1 U12361 ( .A(n9757), .ZN(n9758) );
  NOR2_X1 U12362 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15749), .ZN(n9760) );
  AOI21_X1 U12363 ( .B1(n15232), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n9760), .ZN(
        n9761) );
  OAI21_X1 U12364 ( .B1(n15235), .B2(n9804), .A(n9761), .ZN(n9762) );
  OR4_X1 U12365 ( .A1(n9765), .A2(n9764), .A3(n9763), .A4(n9762), .ZN(P3_U3190) );
  NAND2_X1 U12366 ( .A1(n9773), .A2(P1_U3086), .ZN(n14490) );
  AND2_X1 U12367 ( .A1(n9766), .A2(P1_U3086), .ZN(n11431) );
  INV_X2 U12368 ( .A(n11431), .ZN(n14494) );
  INV_X1 U12369 ( .A(n9767), .ZN(n9769) );
  OAI222_X1 U12370 ( .A1(n14490), .A2(n9768), .B1(n14494), .B2(n9769), .C1(
        P1_U3086), .C2(n10098), .ZN(P1_U3352) );
  NOR2_X1 U12371 ( .A1(n9773), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13829) );
  INV_X1 U12372 ( .A(n13829), .ZN(n13839) );
  OAI222_X1 U12373 ( .A1(n13839), .A2(n9770), .B1(n13837), .B2(n9769), .C1(
        P2_U3088), .C2(n14887), .ZN(P2_U3324) );
  OAI222_X1 U12374 ( .A1(n13839), .A2(n9771), .B1(n13837), .B2(n9796), .C1(
        P2_U3088), .C2(n14874), .ZN(P2_U3325) );
  NOR2_X1 U12375 ( .A1(n9773), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13123) );
  INV_X1 U12376 ( .A(n9772), .ZN(n9776) );
  INV_X1 U12377 ( .A(SI_5_), .ZN(n9775) );
  OAI222_X1 U12378 ( .A1(n11825), .A2(n9776), .B1(n13130), .B2(n9775), .C1(
        n9774), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12379 ( .A(n9777), .ZN(n9780) );
  INV_X1 U12380 ( .A(SI_3_), .ZN(n9779) );
  OAI222_X1 U12381 ( .A1(n11825), .A2(n9780), .B1(n13130), .B2(n9779), .C1(
        n9778), .C2(P3_U3151), .ZN(P3_U3292) );
  INV_X1 U12382 ( .A(n9784), .ZN(n9786) );
  INV_X1 U12383 ( .A(SI_4_), .ZN(n9785) );
  OAI222_X1 U12384 ( .A1(n11825), .A2(n9786), .B1(n13130), .B2(n9785), .C1(
        n10539), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12385 ( .A(n9787), .ZN(n9788) );
  OAI222_X1 U12386 ( .A1(n11825), .A2(n9788), .B1(n13130), .B2(n15689), .C1(
        n10710), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12387 ( .A(n9789), .ZN(n9791) );
  INV_X1 U12388 ( .A(SI_7_), .ZN(n9790) );
  OAI222_X1 U12389 ( .A1(n11825), .A2(n9791), .B1(n13130), .B2(n9790), .C1(
        n10631), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12390 ( .A(n9792), .ZN(n9794) );
  INV_X1 U12391 ( .A(n10116), .ZN(n10308) );
  OAI222_X1 U12392 ( .A1(n14490), .A2(n9793), .B1(n14494), .B2(n9794), .C1(
        P1_U3086), .C2(n10308), .ZN(P1_U3351) );
  INV_X1 U12393 ( .A(n9884), .ZN(n14900) );
  OAI222_X1 U12394 ( .A1(n13839), .A2(n9795), .B1(n13837), .B2(n9794), .C1(
        P2_U3088), .C2(n14900), .ZN(P2_U3323) );
  INV_X1 U12395 ( .A(n14490), .ZN(n14474) );
  INV_X1 U12396 ( .A(n14474), .ZN(n14486) );
  OAI222_X1 U12397 ( .A1(n14486), .A2(n9797), .B1(n14494), .B2(n9796), .C1(
        P1_U3086), .C2(n10097), .ZN(P1_U3353) );
  OAI222_X1 U12398 ( .A1(n14494), .A2(n9818), .B1(n10095), .B2(P1_U3086), .C1(
        n7663), .C2(n14486), .ZN(P1_U3354) );
  INV_X1 U12399 ( .A(n9798), .ZN(n9799) );
  INV_X1 U12400 ( .A(SI_10_), .ZN(n15503) );
  INV_X1 U12401 ( .A(n11083), .ZN(n12640) );
  OAI222_X1 U12402 ( .A1(n11825), .A2(n9799), .B1(n13130), .B2(n15503), .C1(
        n12640), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U12403 ( .A1(n11825), .A2(n9801), .B1(n13130), .B2(n9800), .C1(
        n15194), .C2(P3_U3151), .ZN(P3_U3284) );
  OAI222_X1 U12404 ( .A1(P3_U3151), .A2(n9804), .B1(n13130), .B2(n9803), .C1(
        n11825), .C2(n9802), .ZN(P3_U3287) );
  INV_X1 U12405 ( .A(n9805), .ZN(n9807) );
  INV_X1 U12406 ( .A(SI_9_), .ZN(n9806) );
  OAI222_X1 U12407 ( .A1(n7217), .A2(P3_U3151), .B1(n11825), .B2(n9807), .C1(
        n9806), .C2(n13130), .ZN(P3_U3286) );
  OAI222_X1 U12408 ( .A1(n9810), .A2(P3_U3151), .B1(n11825), .B2(n9809), .C1(
        n9808), .C2(n13130), .ZN(P3_U3295) );
  OAI222_X1 U12409 ( .A1(n9813), .A2(P3_U3151), .B1(n11825), .B2(n9812), .C1(
        n9811), .C2(n13130), .ZN(P3_U3289) );
  INV_X1 U12410 ( .A(n9814), .ZN(n9816) );
  OAI222_X1 U12411 ( .A1(n13839), .A2(n9815), .B1(n13837), .B2(n9816), .C1(
        P2_U3088), .C2(n14913), .ZN(P2_U3322) );
  INV_X1 U12412 ( .A(n10117), .ZN(n10137) );
  OAI222_X1 U12413 ( .A1(n14490), .A2(n9817), .B1(n14494), .B2(n9816), .C1(
        P1_U3086), .C2(n10137), .ZN(P1_U3350) );
  OAI222_X1 U12414 ( .A1(P2_U3088), .A2(n13377), .B1(n13837), .B2(n9818), .C1(
        n7662), .C2(n13839), .ZN(P2_U3326) );
  INV_X1 U12415 ( .A(n15214), .ZN(n12663) );
  OAI222_X1 U12416 ( .A1(n11825), .A2(n9819), .B1(n13130), .B2(n15480), .C1(
        n12663), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12417 ( .A(n9820), .ZN(n9823) );
  INV_X1 U12418 ( .A(n9888), .ZN(n14926) );
  OAI222_X1 U12419 ( .A1(n13839), .A2(n9821), .B1(n13837), .B2(n9823), .C1(
        P2_U3088), .C2(n14926), .ZN(P2_U3321) );
  INV_X1 U12420 ( .A(n10156), .ZN(n9822) );
  OAI222_X1 U12421 ( .A1(n14490), .A2(n9824), .B1(n14494), .B2(n9823), .C1(
        P1_U3086), .C2(n9822), .ZN(P1_U3349) );
  NAND2_X1 U12422 ( .A1(n10423), .A2(n13115), .ZN(n9825) );
  OAI21_X1 U12423 ( .B1(n13115), .B2(n9826), .A(n9825), .ZN(P3_U3377) );
  INV_X1 U12424 ( .A(n9827), .ZN(n9830) );
  INV_X1 U12425 ( .A(n10144), .ZN(n9828) );
  OAI222_X1 U12426 ( .A1(n14490), .A2(n9829), .B1(n14494), .B2(n9830), .C1(
        P1_U3086), .C2(n9828), .ZN(P1_U3348) );
  INV_X1 U12427 ( .A(n9890), .ZN(n14938) );
  OAI222_X1 U12428 ( .A1(n13839), .A2(n9831), .B1(n13837), .B2(n9830), .C1(
        P2_U3088), .C2(n14938), .ZN(P2_U3320) );
  INV_X1 U12429 ( .A(n9832), .ZN(n9834) );
  OAI222_X1 U12430 ( .A1(n13839), .A2(n9833), .B1(n13837), .B2(n9834), .C1(
        P2_U3088), .C2(n14951), .ZN(P2_U3319) );
  INV_X1 U12431 ( .A(n10437), .ZN(n10112) );
  OAI222_X1 U12432 ( .A1(n14490), .A2(n9835), .B1(n14494), .B2(n9834), .C1(
        P1_U3086), .C2(n10112), .ZN(P1_U3347) );
  OAI222_X1 U12433 ( .A1(n11825), .A2(n9836), .B1(n13130), .B2(n15723), .C1(
        n15234), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12434 ( .A(n9837), .ZN(n9839) );
  INV_X1 U12435 ( .A(n10732), .ZN(n10435) );
  OAI222_X1 U12436 ( .A1(n14490), .A2(n9838), .B1(n14494), .B2(n9839), .C1(
        P1_U3086), .C2(n10435), .ZN(P1_U3346) );
  INV_X1 U12437 ( .A(n9894), .ZN(n9998) );
  OAI222_X1 U12438 ( .A1(n13839), .A2(n9840), .B1(n13837), .B2(n9839), .C1(
        P2_U3088), .C2(n9998), .ZN(P2_U3318) );
  INV_X1 U12439 ( .A(n9841), .ZN(n9843) );
  INV_X1 U12440 ( .A(n11174), .ZN(n10737) );
  OAI222_X1 U12441 ( .A1(n14490), .A2(n9842), .B1(n14494), .B2(n9843), .C1(
        P1_U3086), .C2(n10737), .ZN(P1_U3345) );
  INV_X1 U12442 ( .A(n10002), .ZN(n14966) );
  OAI222_X1 U12443 ( .A1(n13839), .A2(n9844), .B1(n13837), .B2(n9843), .C1(
        P2_U3088), .C2(n14966), .ZN(P2_U3317) );
  OAI222_X1 U12444 ( .A1(n11825), .A2(n9845), .B1(n13130), .B2(n15542), .C1(
        n15248), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X2 U12445 ( .A(P2_U3947), .ZN(n13373) );
  NAND2_X1 U12446 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n13373), .ZN(n9846) );
  OAI21_X1 U12447 ( .B1(n13462), .B2(n13373), .A(n9846), .ZN(P2_U3551) );
  INV_X1 U12448 ( .A(n9847), .ZN(n9849) );
  INV_X1 U12449 ( .A(n11176), .ZN(n14736) );
  OAI222_X1 U12450 ( .A1(n14490), .A2(n9848), .B1(n14494), .B2(n9849), .C1(
        P1_U3086), .C2(n14736), .ZN(P1_U3344) );
  INV_X1 U12451 ( .A(n10167), .ZN(n9995) );
  OAI222_X1 U12452 ( .A1(n13839), .A2(n9850), .B1(n13837), .B2(n9849), .C1(
        P2_U3088), .C2(n9995), .ZN(P2_U3316) );
  INV_X1 U12453 ( .A(n14626), .ZN(n9851) );
  OAI222_X1 U12454 ( .A1(n11825), .A2(n9853), .B1(n13130), .B2(n9852), .C1(
        n9851), .C2(P3_U3151), .ZN(P3_U3280) );
  MUX2_X1 U12455 ( .A(n10805), .B(P2_REG2_REG_9__SCAN_IN), .S(n9894), .Z(n9869) );
  MUX2_X1 U12456 ( .A(n9124), .B(P2_REG2_REG_2__SCAN_IN), .S(n14874), .Z(
        n14867) );
  INV_X1 U12457 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10925) );
  MUX2_X1 U12458 ( .A(n10925), .B(P2_REG2_REG_1__SCAN_IN), .S(n13377), .Z(
        n13381) );
  AND2_X1 U12459 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n13380) );
  NAND2_X1 U12460 ( .A1(n13381), .A2(n13380), .ZN(n13379) );
  OAI21_X1 U12461 ( .B1(n10925), .B2(n13377), .A(n13379), .ZN(n14866) );
  NAND2_X1 U12462 ( .A1(n14867), .A2(n14866), .ZN(n14865) );
  OR2_X1 U12463 ( .A1(n14874), .A2(n9124), .ZN(n9854) );
  NAND2_X1 U12464 ( .A1(n14865), .A2(n9854), .ZN(n14879) );
  MUX2_X1 U12465 ( .A(n9855), .B(P2_REG2_REG_3__SCAN_IN), .S(n14887), .Z(
        n14880) );
  NAND2_X1 U12466 ( .A1(n14879), .A2(n14880), .ZN(n14878) );
  OR2_X1 U12467 ( .A1(n14887), .A2(n9855), .ZN(n9856) );
  NAND2_X1 U12468 ( .A1(n14878), .A2(n9856), .ZN(n14892) );
  INV_X1 U12469 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9857) );
  MUX2_X1 U12470 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9857), .S(n9884), .Z(n14893) );
  NAND2_X1 U12471 ( .A1(n14892), .A2(n14893), .ZN(n14891) );
  NAND2_X1 U12472 ( .A1(n9884), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U12473 ( .A1(n14891), .A2(n9858), .ZN(n14909) );
  INV_X1 U12474 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9859) );
  MUX2_X1 U12475 ( .A(n9859), .B(P2_REG2_REG_5__SCAN_IN), .S(n14913), .Z(
        n14910) );
  NAND2_X1 U12476 ( .A1(n14909), .A2(n14910), .ZN(n14908) );
  NAND2_X1 U12477 ( .A1(n9886), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12478 ( .A1(n14908), .A2(n9860), .ZN(n14922) );
  XNOR2_X1 U12479 ( .A(n9888), .B(n9861), .ZN(n14923) );
  NAND2_X1 U12480 ( .A1(n14922), .A2(n14923), .ZN(n14921) );
  NAND2_X1 U12481 ( .A1(n9888), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U12482 ( .A1(n14921), .A2(n9862), .ZN(n14935) );
  INV_X1 U12483 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9863) );
  MUX2_X1 U12484 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9863), .S(n9890), .Z(n14934) );
  NAND2_X1 U12485 ( .A1(n14935), .A2(n14934), .ZN(n14933) );
  NAND2_X1 U12486 ( .A1(n9890), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U12487 ( .A1(n14933), .A2(n9864), .ZN(n14945) );
  INV_X1 U12488 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9865) );
  MUX2_X1 U12489 ( .A(n9865), .B(P2_REG2_REG_8__SCAN_IN), .S(n14951), .Z(
        n14944) );
  NAND2_X1 U12490 ( .A1(n14945), .A2(n14944), .ZN(n14943) );
  NAND2_X1 U12491 ( .A1(n9892), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U12492 ( .A1(n14943), .A2(n9866), .ZN(n9868) );
  OR2_X1 U12493 ( .A1(n9868), .A2(n9869), .ZN(n9990) );
  INV_X1 U12494 ( .A(n9990), .ZN(n9867) );
  AOI21_X1 U12495 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9903) );
  NAND2_X1 U12496 ( .A1(n9960), .A2(n9958), .ZN(n9870) );
  NAND2_X1 U12497 ( .A1(n9870), .A2(n6690), .ZN(n9872) );
  AND2_X1 U12498 ( .A1(n9872), .A2(n9871), .ZN(n9876) );
  INV_X1 U12499 ( .A(n9876), .ZN(n9898) );
  OR2_X1 U12500 ( .A1(n9662), .A2(P2_U3088), .ZN(n13827) );
  INV_X1 U12501 ( .A(n13827), .ZN(n9874) );
  AND2_X1 U12502 ( .A1(n13830), .A2(n9874), .ZN(n9875) );
  INV_X1 U12503 ( .A(n15028), .ZN(n15018) );
  AND2_X1 U12504 ( .A1(n9876), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14864) );
  AND2_X1 U12505 ( .A1(n9662), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9877) );
  NAND2_X1 U12506 ( .A1(n9898), .A2(n9877), .ZN(n15035) );
  NAND2_X1 U12507 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10918) );
  OAI21_X1 U12508 ( .B1(n15035), .B2(n9998), .A(n10918), .ZN(n9901) );
  INV_X1 U12509 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9878) );
  MUX2_X1 U12510 ( .A(n9878), .B(P2_REG1_REG_2__SCAN_IN), .S(n14874), .Z(
        n14870) );
  INV_X1 U12511 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10186) );
  MUX2_X1 U12512 ( .A(n10186), .B(P2_REG1_REG_1__SCAN_IN), .S(n13377), .Z(
        n13384) );
  AND2_X1 U12513 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13383) );
  NAND2_X1 U12514 ( .A1(n13384), .A2(n13383), .ZN(n13382) );
  INV_X1 U12515 ( .A(n13377), .ZN(n9879) );
  NAND2_X1 U12516 ( .A1(n9879), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U12517 ( .A1(n13382), .A2(n9880), .ZN(n14869) );
  NAND2_X1 U12518 ( .A1(n14870), .A2(n14869), .ZN(n14868) );
  OR2_X1 U12519 ( .A1(n14874), .A2(n9878), .ZN(n9881) );
  NAND2_X1 U12520 ( .A1(n14868), .A2(n9881), .ZN(n14882) );
  INV_X1 U12521 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9882) );
  MUX2_X1 U12522 ( .A(n9882), .B(P2_REG1_REG_3__SCAN_IN), .S(n14887), .Z(
        n14883) );
  NAND2_X1 U12523 ( .A1(n14882), .A2(n14883), .ZN(n14881) );
  OR2_X1 U12524 ( .A1(n14887), .A2(n9882), .ZN(n9883) );
  NAND2_X1 U12525 ( .A1(n14881), .A2(n9883), .ZN(n14895) );
  MUX2_X1 U12526 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9163), .S(n9884), .Z(n14896) );
  NAND2_X1 U12527 ( .A1(n14895), .A2(n14896), .ZN(n14894) );
  NAND2_X1 U12528 ( .A1(n9884), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U12529 ( .A1(n14894), .A2(n9885), .ZN(n14906) );
  INV_X1 U12530 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15120) );
  MUX2_X1 U12531 ( .A(n15120), .B(P2_REG1_REG_5__SCAN_IN), .S(n14913), .Z(
        n14907) );
  NAND2_X1 U12532 ( .A1(n14906), .A2(n14907), .ZN(n14905) );
  NAND2_X1 U12533 ( .A1(n9886), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U12534 ( .A1(n14905), .A2(n9887), .ZN(n14919) );
  INV_X1 U12535 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15122) );
  MUX2_X1 U12536 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15122), .S(n9888), .Z(
        n14920) );
  NAND2_X1 U12537 ( .A1(n14919), .A2(n14920), .ZN(n14918) );
  NAND2_X1 U12538 ( .A1(n9888), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U12539 ( .A1(n14918), .A2(n9889), .ZN(n14932) );
  INV_X1 U12540 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15124) );
  MUX2_X1 U12541 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n15124), .S(n9890), .Z(
        n14931) );
  NAND2_X1 U12542 ( .A1(n14932), .A2(n14931), .ZN(n14930) );
  NAND2_X1 U12543 ( .A1(n9890), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U12544 ( .A1(n14930), .A2(n9891), .ZN(n14948) );
  MUX2_X1 U12545 ( .A(n9220), .B(P2_REG1_REG_8__SCAN_IN), .S(n14951), .Z(
        n14947) );
  NAND2_X1 U12546 ( .A1(n14948), .A2(n14947), .ZN(n14946) );
  NAND2_X1 U12547 ( .A1(n9892), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U12548 ( .A1(n14946), .A2(n9893), .ZN(n9896) );
  MUX2_X1 U12549 ( .A(n9997), .B(P2_REG1_REG_9__SCAN_IN), .S(n9894), .Z(n9895)
         );
  NAND2_X1 U12550 ( .A1(n9896), .A2(n9895), .ZN(n9899) );
  NOR2_X1 U12551 ( .A1(n13830), .A2(n13827), .ZN(n9897) );
  NAND2_X1 U12552 ( .A1(n9898), .A2(n9897), .ZN(n15013) );
  AOI21_X1 U12553 ( .B1(n10000), .B2(n9899), .A(n15013), .ZN(n9900) );
  AOI211_X1 U12554 ( .C1(n14864), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n9901), .B(
        n9900), .ZN(n9902) );
  OAI21_X1 U12555 ( .B1(n9903), .B2(n15018), .A(n9902), .ZN(P2_U3223) );
  NAND2_X1 U12556 ( .A1(n9904), .A2(n12237), .ZN(n14833) );
  AOI22_X1 U12557 ( .A1(n14833), .A2(n9906), .B1(n9909), .B2(n9905), .ZN(
        P1_U3445) );
  INV_X1 U12558 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9910) );
  INV_X1 U12559 ( .A(n9907), .ZN(n9908) );
  AOI22_X1 U12560 ( .A1(n14833), .A2(n9910), .B1(n9909), .B2(n9908), .ZN(
        P1_U3446) );
  OAI211_X1 U12561 ( .C1(n15018), .C2(P2_REG2_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .B(n15035), .ZN(n9912) );
  AOI21_X1 U12562 ( .B1(n15032), .B2(n9911), .A(n9912), .ZN(n9916) );
  AOI21_X1 U12563 ( .B1(n15028), .B2(P2_REG2_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U12564 ( .A1(n14864), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9914) );
  NAND3_X1 U12565 ( .A1(n9912), .A2(n15032), .A3(P2_REG1_REG_0__SCAN_IN), .ZN(
        n9913) );
  OAI211_X1 U12566 ( .C1(n9916), .C2(n9915), .A(n9914), .B(n9913), .ZN(
        P2_U3214) );
  INV_X1 U12567 ( .A(n12673), .ZN(n12692) );
  OAI222_X1 U12568 ( .A1(n11825), .A2(n9917), .B1(n12692), .B2(P3_U3151), .C1(
        n15453), .C2(n13130), .ZN(P3_U3279) );
  INV_X1 U12569 ( .A(n9918), .ZN(n9920) );
  INV_X1 U12570 ( .A(n14058), .ZN(n11180) );
  OAI222_X1 U12571 ( .A1(n14486), .A2(n9919), .B1(n14494), .B2(n9920), .C1(
        P1_U3086), .C2(n11180), .ZN(P1_U3343) );
  INV_X1 U12572 ( .A(n10170), .ZN(n11665) );
  OAI222_X1 U12573 ( .A1(n13839), .A2(n9921), .B1(n13837), .B2(n9920), .C1(
        P2_U3088), .C2(n11665), .ZN(P2_U3315) );
  XNOR2_X1 U12574 ( .A(n9922), .B(n11827), .ZN(n9923) );
  NAND2_X1 U12575 ( .A1(n11342), .A2(n11827), .ZN(n10051) );
  NAND2_X1 U12576 ( .A1(n13374), .A2(n13651), .ZN(n9972) );
  XNOR2_X1 U12577 ( .A(n9973), .B(n9972), .ZN(n9928) );
  OR2_X1 U12578 ( .A1(n9926), .A2(n13375), .ZN(n10181) );
  OAI21_X1 U12579 ( .B1(n9926), .B2(n13651), .A(n10181), .ZN(n10060) );
  AOI21_X1 U12580 ( .B1(n9926), .B2(n10229), .A(n10060), .ZN(n9927) );
  AOI21_X1 U12581 ( .B1(n9928), .B2(n9927), .A(n9971), .ZN(n9970) );
  INV_X1 U12582 ( .A(P2_B_REG_SCAN_IN), .ZN(n9929) );
  XNOR2_X1 U12583 ( .A(n11636), .B(n9929), .ZN(n9932) );
  INV_X1 U12584 ( .A(n13835), .ZN(n9931) );
  INV_X1 U12585 ( .A(n13834), .ZN(n9930) );
  OR2_X1 U12586 ( .A1(n15068), .A2(P2_D_REG_1__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U12587 ( .A1(n13835), .A2(n13834), .ZN(n9933) );
  NAND2_X1 U12588 ( .A1(n9934), .A2(n9933), .ZN(n10045) );
  INV_X1 U12589 ( .A(n15072), .ZN(n15074) );
  NOR2_X1 U12590 ( .A1(n10045), .A2(n15074), .ZN(n15073) );
  NOR4_X1 U12591 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9938) );
  NOR4_X1 U12592 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9937) );
  NOR4_X1 U12593 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9936) );
  NOR4_X1 U12594 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9935) );
  NAND4_X1 U12595 ( .A1(n9938), .A2(n9937), .A3(n9936), .A4(n9935), .ZN(n9945)
         );
  NOR2_X1 U12596 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9942) );
  NOR4_X1 U12597 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9941) );
  NOR4_X1 U12598 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9940) );
  NOR4_X1 U12599 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9939) );
  NAND4_X1 U12600 ( .A1(n9942), .A2(n9941), .A3(n9940), .A4(n9939), .ZN(n9944)
         );
  INV_X1 U12601 ( .A(n15068), .ZN(n9943) );
  OAI21_X1 U12602 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n10336) );
  NAND2_X1 U12603 ( .A1(n15073), .A2(n10336), .ZN(n10457) );
  OR2_X1 U12604 ( .A1(n15068), .A2(P2_D_REG_0__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U12605 ( .A1(n11636), .A2(n13834), .ZN(n9946) );
  NAND2_X1 U12606 ( .A1(n9947), .A2(n9946), .ZN(n15071) );
  INV_X1 U12607 ( .A(n9966), .ZN(n9951) );
  OR2_X1 U12608 ( .A1(n10051), .A2(n9948), .ZN(n15111) );
  INV_X1 U12609 ( .A(n9958), .ZN(n9949) );
  AND2_X1 U12610 ( .A1(n15111), .A2(n9949), .ZN(n9950) );
  NAND2_X1 U12611 ( .A1(n9951), .A2(n9950), .ZN(n13339) );
  NOR2_X2 U12612 ( .A1(n9966), .A2(n9957), .ZN(n13334) );
  NAND2_X1 U12613 ( .A1(n9958), .A2(n9662), .ZN(n13312) );
  NAND2_X1 U12614 ( .A1(n13372), .A2(n13409), .ZN(n9953) );
  NAND2_X1 U12615 ( .A1(n13331), .A2(n13375), .ZN(n9952) );
  NAND2_X1 U12616 ( .A1(n9953), .A2(n9952), .ZN(n10184) );
  INV_X1 U12617 ( .A(n10336), .ZN(n9954) );
  NOR2_X1 U12618 ( .A1(n15071), .A2(n9954), .ZN(n10046) );
  INV_X1 U12619 ( .A(n10045), .ZN(n9955) );
  NAND2_X1 U12620 ( .A1(n10046), .A2(n9955), .ZN(n9956) );
  INV_X1 U12621 ( .A(n10051), .ZN(n9964) );
  NAND2_X1 U12622 ( .A1(n9964), .A2(n10460), .ZN(n10043) );
  NAND2_X1 U12623 ( .A1(n9956), .A2(n10043), .ZN(n9962) );
  NAND2_X1 U12624 ( .A1(n9958), .A2(n9957), .ZN(n10455) );
  AND3_X1 U12625 ( .A1(n10455), .A2(n9960), .A3(n9959), .ZN(n9961) );
  NAND2_X1 U12626 ( .A1(n9962), .A2(n9961), .ZN(n10235) );
  OR2_X1 U12627 ( .A1(n10235), .A2(P2_U3088), .ZN(n10059) );
  AOI22_X1 U12628 ( .A1(n13334), .A2(n10184), .B1(n10059), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U12629 ( .A1(n9964), .A2(n9963), .ZN(n10645) );
  INV_X1 U12630 ( .A(n10043), .ZN(n9965) );
  NAND2_X1 U12631 ( .A1(n9967), .A2(n10197), .ZN(n9968) );
  OAI211_X1 U12632 ( .C1(n9970), .C2(n13339), .A(n9969), .B(n9968), .ZN(
        P2_U3194) );
  AOI21_X1 U12633 ( .B1(n9973), .B2(n9972), .A(n9971), .ZN(n9978) );
  INV_X1 U12634 ( .A(n9974), .ZN(n10344) );
  XNOR2_X1 U12635 ( .A(n10344), .B(n10229), .ZN(n9976) );
  NAND2_X1 U12636 ( .A1(n13372), .A2(n13651), .ZN(n9975) );
  NAND2_X1 U12637 ( .A1(n9976), .A2(n9975), .ZN(n10230) );
  OAI21_X1 U12638 ( .B1(n9976), .B2(n9975), .A(n10230), .ZN(n9977) );
  NOR2_X1 U12639 ( .A1(n9978), .A2(n9977), .ZN(n10232) );
  AOI21_X1 U12640 ( .B1(n9978), .B2(n9977), .A(n10232), .ZN(n9983) );
  NOR2_X1 U12641 ( .A1(n10206), .A2(n13312), .ZN(n9980) );
  NOR2_X1 U12642 ( .A1(n10196), .A2(n13448), .ZN(n9979) );
  OR2_X1 U12643 ( .A1(n9980), .A2(n9979), .ZN(n10216) );
  AOI22_X1 U12644 ( .A1(n13334), .A2(n10216), .B1(n10059), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U12645 ( .A1(n9967), .A2(n9974), .ZN(n9981) );
  OAI211_X1 U12646 ( .C1(n9983), .C2(n13339), .A(n9982), .B(n9981), .ZN(
        P2_U3209) );
  INV_X1 U12647 ( .A(n12237), .ZN(n10359) );
  INV_X1 U12648 ( .A(n9986), .ZN(n9984) );
  NAND2_X1 U12649 ( .A1(n9984), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12240) );
  NAND2_X1 U12650 ( .A1(n10359), .A2(n12240), .ZN(n10071) );
  AOI21_X1 U12651 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(n10070) );
  INV_X1 U12652 ( .A(n10070), .ZN(n9988) );
  AND2_X1 U12653 ( .A1(n10071), .A2(n9988), .ZN(n14729) );
  NOR2_X1 U12654 ( .A1(n14729), .A2(n14042), .ZN(P1_U3085) );
  XNOR2_X1 U12655 ( .A(n10167), .B(P2_REG2_REG_11__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U12656 ( .A1(n9998), .A2(n10805), .ZN(n9989) );
  NAND2_X1 U12657 ( .A1(n9990), .A2(n9989), .ZN(n14957) );
  INV_X1 U12658 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11131) );
  MUX2_X1 U12659 ( .A(n11131), .B(P2_REG2_REG_10__SCAN_IN), .S(n10002), .Z(
        n14956) );
  OR2_X1 U12660 ( .A1(n14957), .A2(n14956), .ZN(n14959) );
  NAND2_X1 U12661 ( .A1(n10002), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U12662 ( .A1(n14959), .A2(n9991), .ZN(n9993) );
  INV_X1 U12663 ( .A(n10166), .ZN(n9992) );
  AOI21_X1 U12664 ( .B1(n9994), .B2(n9993), .A(n9992), .ZN(n10009) );
  NAND2_X1 U12665 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11144)
         );
  OAI21_X1 U12666 ( .B1(n15035), .B2(n9995), .A(n11144), .ZN(n9996) );
  AOI21_X1 U12667 ( .B1(n14864), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9996), .ZN(
        n10008) );
  NAND2_X1 U12668 ( .A1(n9998), .A2(n9997), .ZN(n9999) );
  NAND2_X1 U12669 ( .A1(n10000), .A2(n9999), .ZN(n14961) );
  INV_X1 U12670 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10001) );
  MUX2_X1 U12671 ( .A(n10001), .B(P2_REG1_REG_10__SCAN_IN), .S(n10002), .Z(
        n14960) );
  NAND2_X1 U12672 ( .A1(n10002), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U12673 ( .A1(n14963), .A2(n10003), .ZN(n10006) );
  INV_X1 U12674 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10004) );
  MUX2_X1 U12675 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10004), .S(n10167), .Z(
        n10005) );
  NAND2_X1 U12676 ( .A1(n10006), .A2(n10005), .ZN(n10169) );
  OAI211_X1 U12677 ( .C1(n10006), .C2(n10005), .A(n10169), .B(n15032), .ZN(
        n10007) );
  OAI211_X1 U12678 ( .C1(n10009), .C2(n15018), .A(n10008), .B(n10007), .ZN(
        P2_U3225) );
  INV_X1 U12679 ( .A(n10010), .ZN(n10011) );
  INV_X1 U12680 ( .A(SI_17_), .ZN(n15545) );
  OAI222_X1 U12681 ( .A1(n12718), .A2(P3_U3151), .B1(n11825), .B2(n10011), 
        .C1(n15545), .C2(n13130), .ZN(P3_U3278) );
  INV_X1 U12682 ( .A(n11669), .ZN(n14981) );
  INV_X1 U12683 ( .A(n10012), .ZN(n10014) );
  OAI222_X1 U12684 ( .A1(P2_U3088), .A2(n14981), .B1(n13837), .B2(n10014), 
        .C1(n10013), .C2(n13839), .ZN(P2_U3314) );
  INV_X1 U12685 ( .A(n14754), .ZN(n10015) );
  OAI222_X1 U12686 ( .A1(n14490), .A2(n10016), .B1(P1_U3086), .B2(n10015), 
        .C1(n10014), .C2(n14494), .ZN(P1_U3342) );
  INV_X1 U12687 ( .A(SI_18_), .ZN(n10017) );
  INV_X1 U12688 ( .A(n12715), .ZN(n12719) );
  OAI222_X1 U12689 ( .A1(n11825), .A2(n10018), .B1(n13130), .B2(n10017), .C1(
        n12719), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U12690 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n10020) );
  NAND2_X1 U12691 ( .A1(n12496), .A2(n10958), .ZN(n10019) );
  OAI21_X1 U12692 ( .B1(n10958), .B2(n10020), .A(n10019), .ZN(P3_U3500) );
  INV_X1 U12693 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n15671) );
  NAND2_X1 U12694 ( .A1(n12947), .A2(n10958), .ZN(n10021) );
  OAI21_X1 U12695 ( .B1(n10958), .B2(n15671), .A(n10021), .ZN(P3_U3504) );
  INV_X1 U12696 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n15731) );
  NAND2_X1 U12697 ( .A1(n12949), .A2(n10958), .ZN(n10022) );
  OAI21_X1 U12698 ( .B1(P3_U3897), .B2(n15731), .A(n10022), .ZN(P3_U3506) );
  INV_X1 U12699 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n15744) );
  NAND2_X1 U12700 ( .A1(n10023), .A2(P3_U3897), .ZN(n10024) );
  OAI21_X1 U12701 ( .B1(n10958), .B2(n15744), .A(n10024), .ZN(P3_U3495) );
  INV_X1 U12702 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U12703 ( .A1(n12423), .A2(P3_U3897), .ZN(n10025) );
  OAI21_X1 U12704 ( .B1(n10958), .B2(n10026), .A(n10025), .ZN(P3_U3508) );
  INV_X1 U12705 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n15717) );
  NAND2_X1 U12706 ( .A1(n12497), .A2(P3_U3897), .ZN(n10027) );
  OAI21_X1 U12707 ( .B1(n10958), .B2(n15717), .A(n10027), .ZN(P3_U3498) );
  INV_X1 U12708 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n15530) );
  NAND2_X1 U12709 ( .A1(n10028), .A2(P3_U3897), .ZN(n10029) );
  OAI21_X1 U12710 ( .B1(n10958), .B2(n15530), .A(n10029), .ZN(P3_U3496) );
  INV_X1 U12711 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15685) );
  NAND2_X1 U12712 ( .A1(n10030), .A2(P3_U3897), .ZN(n10031) );
  OAI21_X1 U12713 ( .B1(P3_U3897), .B2(n15685), .A(n10031), .ZN(P3_U3502) );
  INV_X1 U12714 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n15706) );
  NAND2_X1 U12715 ( .A1(n12937), .A2(P3_U3897), .ZN(n10032) );
  OAI21_X1 U12716 ( .B1(n10958), .B2(n15706), .A(n10032), .ZN(P3_U3507) );
  INV_X1 U12717 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n15716) );
  NAND2_X1 U12718 ( .A1(n12912), .A2(P3_U3897), .ZN(n10033) );
  OAI21_X1 U12719 ( .B1(n10932), .B2(n15716), .A(n10033), .ZN(P3_U3509) );
  INV_X1 U12720 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n10035) );
  NAND2_X1 U12721 ( .A1(n12936), .A2(P3_U3897), .ZN(n10034) );
  OAI21_X1 U12722 ( .B1(n10932), .B2(n10035), .A(n10034), .ZN(P3_U3505) );
  INV_X1 U12723 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n15724) );
  NAND2_X1 U12724 ( .A1(n12868), .A2(P3_U3897), .ZN(n10036) );
  OAI21_X1 U12725 ( .B1(P3_U3897), .B2(n15724), .A(n10036), .ZN(P3_U3510) );
  INV_X1 U12726 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n15696) );
  NAND2_X1 U12727 ( .A1(n10037), .A2(P3_U3897), .ZN(n10038) );
  OAI21_X1 U12728 ( .B1(n10958), .B2(n15696), .A(n10038), .ZN(P3_U3497) );
  INV_X1 U12729 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U12730 ( .A1(n12401), .A2(P3_U3897), .ZN(n10039) );
  OAI21_X1 U12731 ( .B1(P3_U3897), .B2(n10040), .A(n10039), .ZN(P3_U3501) );
  INV_X1 U12732 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U12733 ( .A1(n11497), .A2(P3_U3897), .ZN(n10041) );
  OAI21_X1 U12734 ( .B1(n10958), .B2(n10042), .A(n10041), .ZN(P3_U3499) );
  AND3_X1 U12735 ( .A1(n15072), .A2(n10043), .A3(n10455), .ZN(n10044) );
  AND2_X2 U12736 ( .A1(n10046), .A2(n10338), .ZN(n15129) );
  NAND2_X1 U12737 ( .A1(n13374), .A2(n13409), .ZN(n10064) );
  OR2_X1 U12738 ( .A1(n11827), .A2(n13400), .ZN(n10048) );
  NAND2_X1 U12739 ( .A1(n10048), .A2(n10047), .ZN(n15048) );
  INV_X1 U12740 ( .A(n15048), .ZN(n13622) );
  AND2_X1 U12741 ( .A1(n6873), .A2(n13622), .ZN(n10049) );
  OR2_X1 U12742 ( .A1(n10049), .A2(n10469), .ZN(n10050) );
  NAND2_X1 U12743 ( .A1(n10064), .A2(n10050), .ZN(n10463) );
  INV_X1 U12744 ( .A(n9095), .ZN(n15083) );
  OR2_X1 U12745 ( .A1(n9926), .A2(n10051), .ZN(n10461) );
  OAI21_X1 U12746 ( .B1(n10469), .B2(n15083), .A(n10461), .ZN(n10052) );
  NOR2_X1 U12747 ( .A1(n10463), .A2(n10052), .ZN(n15076) );
  NAND2_X1 U12748 ( .A1(n15127), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10053) );
  OAI21_X1 U12749 ( .B1(n15127), .B2(n15076), .A(n10053), .ZN(P2_U3499) );
  INV_X1 U12750 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n15489) );
  NAND2_X1 U12751 ( .A1(n10504), .A2(P3_U3897), .ZN(n10054) );
  OAI21_X1 U12752 ( .B1(P3_U3897), .B2(n15489), .A(n10054), .ZN(P3_U3491) );
  INV_X1 U12753 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U12754 ( .A1(n11853), .A2(P3_U3897), .ZN(n10055) );
  OAI21_X1 U12755 ( .B1(P3_U3897), .B2(n10056), .A(n10055), .ZN(P3_U3493) );
  INV_X1 U12756 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U12757 ( .A1(n10280), .A2(P3_U3897), .ZN(n10057) );
  OAI21_X1 U12758 ( .B1(n10958), .B2(n10058), .A(n10057), .ZN(P3_U3492) );
  AOI22_X1 U12759 ( .A1(n9967), .A2(n9099), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10059), .ZN(n10063) );
  AND3_X1 U12760 ( .A1(n9926), .A2(n13375), .A3(n13191), .ZN(n10061) );
  OAI21_X1 U12761 ( .B1(n10061), .B2(n10060), .A(n13343), .ZN(n10062) );
  OAI211_X1 U12762 ( .C1(n10064), .C2(n13348), .A(n10063), .B(n10062), .ZN(
        P2_U3204) );
  INV_X1 U12763 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U12764 ( .A1(n12505), .A2(P3_U3897), .ZN(n10065) );
  OAI21_X1 U12765 ( .B1(n10932), .B2(n10066), .A(n10065), .ZN(P3_U3511) );
  INV_X1 U12766 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15690) );
  NAND2_X1 U12767 ( .A1(n12566), .A2(n10958), .ZN(n10067) );
  OAI21_X1 U12768 ( .B1(P3_U3897), .B2(n15690), .A(n10067), .ZN(P3_U3503) );
  INV_X1 U12769 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n15697) );
  NAND2_X1 U12770 ( .A1(n12869), .A2(n10958), .ZN(n10068) );
  OAI21_X1 U12771 ( .B1(P3_U3897), .B2(n15697), .A(n10068), .ZN(P3_U3512) );
  INV_X1 U12772 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n15674) );
  NAND2_X1 U12773 ( .A1(n12573), .A2(P3_U3897), .ZN(n10069) );
  OAI21_X1 U12774 ( .B1(n10932), .B2(n15674), .A(n10069), .ZN(P3_U3513) );
  NAND2_X1 U12775 ( .A1(n10071), .A2(n10070), .ZN(n14731) );
  NAND2_X1 U12776 ( .A1(n6889), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10075) );
  INV_X1 U12777 ( .A(n10072), .ZN(n10074) );
  INV_X1 U12778 ( .A(n10093), .ZN(n10073) );
  INV_X1 U12779 ( .A(n14488), .ZN(n14727) );
  AOI211_X1 U12780 ( .C1(n10075), .C2(n10074), .A(n10073), .B(n14785), .ZN(
        n10080) );
  NAND2_X1 U12781 ( .A1(n6889), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10264) );
  INV_X1 U12782 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10076) );
  OR2_X1 U12783 ( .A1(n14483), .A2(n14488), .ZN(n10077) );
  AOI211_X1 U12784 ( .C1(n10264), .C2(n10078), .A(n10086), .B(n14789), .ZN(
        n10079) );
  NOR2_X1 U12785 ( .A1(n10080), .A2(n10079), .ZN(n10082) );
  AOI22_X1 U12786 ( .A1(n14729), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10081) );
  OAI211_X1 U12787 ( .C1(n10095), .C2(n14828), .A(n10082), .B(n10081), .ZN(
        P1_U3244) );
  INV_X1 U12788 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10085) );
  INV_X1 U12789 ( .A(n14828), .ZN(n14796) );
  INV_X1 U12790 ( .A(n10098), .ZN(n10114) );
  NAND2_X1 U12791 ( .A1(n14796), .A2(n10114), .ZN(n10084) );
  NAND2_X1 U12792 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n10083) );
  OAI211_X1 U12793 ( .C1(n10085), .C2(n14832), .A(n10084), .B(n10083), .ZN(
        n10105) );
  INV_X1 U12794 ( .A(n10097), .ZN(n10250) );
  INV_X1 U12795 ( .A(n10095), .ZN(n10087) );
  AOI21_X1 U12796 ( .B1(n10087), .B2(P1_REG2_REG_1__SCAN_IN), .A(n10086), .ZN(
        n10248) );
  INV_X1 U12797 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10088) );
  INV_X1 U12798 ( .A(n10089), .ZN(n10247) );
  INV_X1 U12799 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10090) );
  MUX2_X1 U12800 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10090), .S(n10098), .Z(
        n10091) );
  AOI211_X1 U12801 ( .C1(n10092), .C2(n10091), .A(n10113), .B(n14789), .ZN(
        n10104) );
  INV_X1 U12802 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10096) );
  OAI21_X1 U12803 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(n10252) );
  NAND2_X1 U12804 ( .A1(n10252), .A2(n10253), .ZN(n10251) );
  OAI21_X1 U12805 ( .B1(n10097), .B2(n10096), .A(n10251), .ZN(n10101) );
  INV_X1 U12806 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10099) );
  MUX2_X1 U12807 ( .A(n10099), .B(P1_REG1_REG_3__SCAN_IN), .S(n10098), .Z(
        n10100) );
  NOR2_X1 U12808 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  NOR3_X1 U12809 ( .A1(n14785), .A2(n10106), .A3(n10102), .ZN(n10103) );
  OR3_X1 U12810 ( .A1(n10105), .A2(n10104), .A3(n10103), .ZN(P1_U3246) );
  MUX2_X1 U12811 ( .A(n10107), .B(P1_REG1_REG_4__SCAN_IN), .S(n10116), .Z(
        n10302) );
  NOR2_X1 U12812 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  AOI21_X1 U12813 ( .B1(n10116), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10301), .ZN(
        n10127) );
  XOR2_X1 U12814 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10117), .Z(n10128) );
  NAND2_X1 U12815 ( .A1(n10127), .A2(n10128), .ZN(n10126) );
  OAI21_X1 U12816 ( .B1(n10117), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10126), .ZN(
        n10154) );
  XNOR2_X1 U12817 ( .A(n10156), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10155) );
  XNOR2_X1 U12818 ( .A(n10144), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n10142) );
  NOR2_X1 U12819 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  INV_X1 U12820 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10108) );
  MUX2_X1 U12821 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10108), .S(n10437), .Z(
        n10109) );
  OAI21_X1 U12822 ( .B1(n10110), .B2(n10109), .A(n10430), .ZN(n10124) );
  AND2_X1 U12823 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11628) );
  AOI21_X1 U12824 ( .B1(n14729), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11628), .ZN(
        n10111) );
  OAI21_X1 U12825 ( .B1(n14828), .B2(n10112), .A(n10111), .ZN(n10123) );
  MUX2_X1 U12826 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7935), .S(n10116), .Z(
        n10115) );
  INV_X1 U12827 ( .A(n10115), .ZN(n10305) );
  XNOR2_X1 U12828 ( .A(n10117), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n10130) );
  XNOR2_X1 U12829 ( .A(n10156), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n10151) );
  NOR2_X1 U12830 ( .A1(n10152), .A2(n10151), .ZN(n10150) );
  XNOR2_X1 U12831 ( .A(n10144), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n10139) );
  INV_X1 U12832 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10118) );
  MUX2_X1 U12833 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10118), .S(n10437), .Z(
        n10119) );
  INV_X1 U12834 ( .A(n10119), .ZN(n10120) );
  AOI211_X1 U12835 ( .C1(n10121), .C2(n10120), .A(n14789), .B(n10436), .ZN(
        n10122) );
  AOI211_X1 U12836 ( .C1(n14819), .C2(n10124), .A(n10123), .B(n10122), .ZN(
        n10125) );
  INV_X1 U12837 ( .A(n10125), .ZN(P1_U3251) );
  OAI21_X1 U12838 ( .B1(n10128), .B2(n10127), .A(n10126), .ZN(n10133) );
  AOI211_X1 U12839 ( .C1(n10131), .C2(n10130), .A(n14789), .B(n10129), .ZN(
        n10132) );
  AOI21_X1 U12840 ( .B1(n14819), .B2(n10133), .A(n10132), .ZN(n10136) );
  NAND2_X1 U12841 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11250) );
  INV_X1 U12842 ( .A(n11250), .ZN(n10134) );
  AOI21_X1 U12843 ( .B1(n14729), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10134), .ZN(
        n10135) );
  OAI211_X1 U12844 ( .C1(n10137), .C2(n14828), .A(n10136), .B(n10135), .ZN(
        P1_U3248) );
  AOI211_X1 U12845 ( .C1(n10140), .C2(n10139), .A(n14789), .B(n10138), .ZN(
        n10149) );
  AOI211_X1 U12846 ( .C1(n10143), .C2(n10142), .A(n14785), .B(n10141), .ZN(
        n10148) );
  INV_X1 U12847 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10146) );
  NAND2_X1 U12848 ( .A1(n14796), .A2(n10144), .ZN(n10145) );
  NAND2_X1 U12849 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11445) );
  OAI211_X1 U12850 ( .C1(n10146), .C2(n14832), .A(n10145), .B(n11445), .ZN(
        n10147) );
  OR3_X1 U12851 ( .A1(n10149), .A2(n10148), .A3(n10147), .ZN(P1_U3250) );
  AOI211_X1 U12852 ( .C1(n10152), .C2(n10151), .A(n14789), .B(n10150), .ZN(
        n10162) );
  AOI211_X1 U12853 ( .C1(n10155), .C2(n10154), .A(n10153), .B(n14785), .ZN(
        n10161) );
  INV_X1 U12854 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U12855 ( .A1(n14796), .A2(n10156), .ZN(n10158) );
  NAND2_X1 U12856 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10157) );
  OAI211_X1 U12857 ( .C1(n10159), .C2(n14832), .A(n10158), .B(n10157), .ZN(
        n10160) );
  OR3_X1 U12858 ( .A1(n10162), .A2(n10161), .A3(n10160), .ZN(P1_U3249) );
  OAI222_X1 U12859 ( .A1(P3_U3151), .A2(n7624), .B1(n13130), .B2(n10164), .C1(
        n11825), .C2(n10163), .ZN(P3_U3276) );
  INV_X1 U12860 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11651) );
  XNOR2_X1 U12861 ( .A(n10170), .B(n11651), .ZN(n11649) );
  OR2_X1 U12862 ( .A1(n10167), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10165) );
  NAND2_X1 U12863 ( .A1(n10166), .A2(n10165), .ZN(n11650) );
  XOR2_X1 U12864 ( .A(n11649), .B(n11650), .Z(n10177) );
  NAND2_X1 U12865 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11358)
         );
  OAI21_X1 U12866 ( .B1(n15035), .B2(n11665), .A(n11358), .ZN(n10175) );
  NAND2_X1 U12867 ( .A1(n10167), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10168) );
  NAND2_X1 U12868 ( .A1(n10169), .A2(n10168), .ZN(n10172) );
  INV_X1 U12869 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14675) );
  MUX2_X1 U12870 ( .A(n14675), .B(P2_REG1_REG_12__SCAN_IN), .S(n10170), .Z(
        n10171) );
  NAND2_X1 U12871 ( .A1(n10172), .A2(n10171), .ZN(n10173) );
  AOI21_X1 U12872 ( .B1(n11667), .B2(n10173), .A(n15013), .ZN(n10174) );
  AOI211_X1 U12873 ( .C1(n14864), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n10175), 
        .B(n10174), .ZN(n10176) );
  OAI21_X1 U12874 ( .B1(n15018), .B2(n10177), .A(n10176), .ZN(P2_U3226) );
  INV_X1 U12875 ( .A(n10178), .ZN(n10180) );
  INV_X1 U12876 ( .A(n10190), .ZN(n10179) );
  AOI21_X1 U12877 ( .B1(n10180), .B2(n10182), .A(n10179), .ZN(n10931) );
  NAND2_X1 U12878 ( .A1(n6873), .A2(n15083), .ZN(n15099) );
  INV_X1 U12879 ( .A(n15099), .ZN(n13759) );
  INV_X1 U12880 ( .A(n10181), .ZN(n10183) );
  NAND2_X1 U12881 ( .A1(n10182), .A2(n10183), .ZN(n10199) );
  OAI21_X1 U12882 ( .B1(n10183), .B2(n10182), .A(n10199), .ZN(n10185) );
  AOI21_X1 U12883 ( .B1(n10185), .B2(n15048), .A(n10184), .ZN(n10926) );
  NAND2_X1 U12884 ( .A1(n9925), .A2(n9926), .ZN(n10212) );
  OAI211_X1 U12885 ( .C1(n9925), .C2(n9926), .A(n10749), .B(n10212), .ZN(
        n10927) );
  OAI211_X1 U12886 ( .C1(n10931), .C2(n13759), .A(n10926), .B(n10927), .ZN(
        n10365) );
  NAND2_X1 U12887 ( .A1(n15129), .A2(n15079), .ZN(n13758) );
  OAI22_X1 U12888 ( .A1(n13758), .A2(n9925), .B1(n15129), .B2(n10186), .ZN(
        n10187) );
  AOI21_X1 U12889 ( .B1(n15129), .B2(n10365), .A(n10187), .ZN(n10188) );
  INV_X1 U12890 ( .A(n10188), .ZN(P2_U3500) );
  NAND2_X1 U12891 ( .A1(n10196), .A2(n9925), .ZN(n10189) );
  INV_X1 U12892 ( .A(n10214), .ZN(n10210) );
  INV_X1 U12893 ( .A(n13372), .ZN(n10200) );
  NAND2_X1 U12894 ( .A1(n10200), .A2(n10344), .ZN(n10191) );
  INV_X1 U12895 ( .A(n10203), .ZN(n10225) );
  NAND2_X1 U12896 ( .A1(n10206), .A2(n10339), .ZN(n10192) );
  INV_X1 U12897 ( .A(n10659), .ZN(n10193) );
  NAND2_X1 U12898 ( .A1(n10194), .A2(n10193), .ZN(n10654) );
  OAI21_X1 U12899 ( .B1(n10194), .B2(n10193), .A(n10654), .ZN(n10195) );
  INV_X1 U12900 ( .A(n10195), .ZN(n10652) );
  NAND2_X1 U12901 ( .A1(n10197), .A2(n10196), .ZN(n10198) );
  NAND2_X1 U12902 ( .A1(n10199), .A2(n10198), .ZN(n10215) );
  NAND2_X1 U12903 ( .A1(n10215), .A2(n10214), .ZN(n10202) );
  NAND2_X1 U12904 ( .A1(n10200), .A2(n9974), .ZN(n10201) );
  NAND2_X1 U12905 ( .A1(n10202), .A2(n10201), .ZN(n10226) );
  NAND2_X1 U12906 ( .A1(n10226), .A2(n10203), .ZN(n10205) );
  NAND2_X1 U12907 ( .A1(n10963), .A2(n10206), .ZN(n10204) );
  NAND2_X1 U12908 ( .A1(n10205), .A2(n10204), .ZN(n10660) );
  XNOR2_X1 U12909 ( .A(n10660), .B(n10659), .ZN(n10207) );
  OAI22_X1 U12910 ( .A1(n10812), .A2(n13312), .B1(n10206), .B2(n13448), .ZN(
        n13296) );
  AOI21_X1 U12911 ( .B1(n10207), .B2(n15048), .A(n13296), .ZN(n10649) );
  OR2_X1 U12912 ( .A1(n10212), .A2(n9974), .ZN(n10224) );
  INV_X1 U12913 ( .A(n10655), .ZN(n10656) );
  OAI211_X1 U12914 ( .C1(n10661), .C2(n10223), .A(n10656), .B(n10749), .ZN(
        n10646) );
  OAI211_X1 U12915 ( .C1(n10652), .C2(n13759), .A(n10649), .B(n10646), .ZN(
        n10370) );
  OAI22_X1 U12916 ( .A1(n13758), .A2(n10661), .B1(n15129), .B2(n9163), .ZN(
        n10208) );
  AOI21_X1 U12917 ( .B1(n10370), .B2(n15129), .A(n10208), .ZN(n10209) );
  INV_X1 U12918 ( .A(n10209), .ZN(P2_U3503) );
  INV_X1 U12919 ( .A(n10212), .ZN(n10213) );
  OAI211_X1 U12920 ( .C1(n10213), .C2(n10344), .A(n10749), .B(n10224), .ZN(
        n10862) );
  INV_X1 U12921 ( .A(n10862), .ZN(n10219) );
  XNOR2_X1 U12922 ( .A(n10215), .B(n10214), .ZN(n10217) );
  AOI21_X1 U12923 ( .B1(n10217), .B2(n15048), .A(n10216), .ZN(n10866) );
  INV_X1 U12924 ( .A(n10866), .ZN(n10218) );
  AOI211_X1 U12925 ( .C1(n15099), .C2(n10864), .A(n10219), .B(n10218), .ZN(
        n10347) );
  INV_X1 U12926 ( .A(n13758), .ZN(n13766) );
  AOI22_X1 U12927 ( .A1(n13766), .A2(n9974), .B1(n15127), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10220) );
  OAI21_X1 U12928 ( .B1(n10347), .B2(n15127), .A(n10220), .ZN(P2_U3501) );
  OAI21_X1 U12929 ( .B1(n10222), .B2(n10225), .A(n10221), .ZN(n10968) );
  AOI211_X1 U12930 ( .C1(n10963), .C2(n10224), .A(n13191), .B(n10223), .ZN(
        n10962) );
  XNOR2_X1 U12931 ( .A(n10226), .B(n10225), .ZN(n10227) );
  AOI22_X1 U12932 ( .A1(n13370), .A2(n13409), .B1(n13331), .B2(n13372), .ZN(
        n10234) );
  OAI21_X1 U12933 ( .B1(n10227), .B2(n13622), .A(n10234), .ZN(n10961) );
  AOI211_X1 U12934 ( .C1(n15099), .C2(n10968), .A(n10962), .B(n10961), .ZN(
        n10342) );
  AOI22_X1 U12935 ( .A1(n13766), .A2(n10963), .B1(n15127), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10228) );
  OAI21_X1 U12936 ( .B1(n10342), .B2(n15127), .A(n10228), .ZN(P2_U3502) );
  XNOR2_X1 U12937 ( .A(n10963), .B(n13226), .ZN(n10316) );
  NAND2_X1 U12938 ( .A1(n13371), .A2(n13191), .ZN(n10315) );
  XNOR2_X1 U12939 ( .A(n10316), .B(n10315), .ZN(n10318) );
  INV_X1 U12940 ( .A(n10230), .ZN(n10231) );
  XOR2_X1 U12941 ( .A(n10319), .B(n10318), .Z(n10238) );
  INV_X1 U12942 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10233) );
  OAI22_X1 U12943 ( .A1(n13348), .A2(n10234), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10233), .ZN(n10237) );
  NAND2_X1 U12944 ( .A1(n10235), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13336) );
  OAI22_X1 U12945 ( .A1(n13354), .A2(n10339), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13336), .ZN(n10236) );
  AOI211_X1 U12946 ( .C1(n13343), .C2(n10238), .A(n10237), .B(n10236), .ZN(
        n10239) );
  INV_X1 U12947 ( .A(n10239), .ZN(P2_U3190) );
  INV_X1 U12948 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n15566) );
  NAND2_X1 U12949 ( .A1(n12846), .A2(P3_U3897), .ZN(n10240) );
  OAI21_X1 U12950 ( .B1(P3_U3897), .B2(n15566), .A(n10240), .ZN(P3_U3514) );
  INV_X1 U12951 ( .A(n10241), .ZN(n10272) );
  INV_X1 U12952 ( .A(n14795), .ZN(n10243) );
  OAI222_X1 U12953 ( .A1(n14494), .A2(n10272), .B1(n10243), .B2(P1_U3086), 
        .C1(n10242), .C2(n14486), .ZN(P1_U3339) );
  INV_X1 U12954 ( .A(n10244), .ZN(n10298) );
  INV_X1 U12955 ( .A(n14060), .ZN(n14761) );
  OAI222_X1 U12956 ( .A1(n14494), .A2(n10298), .B1(n14761), .B2(P1_U3086), 
        .C1(n10245), .C2(n14486), .ZN(P1_U3341) );
  AOI211_X1 U12957 ( .C1(n10248), .C2(n10247), .A(n10246), .B(n14789), .ZN(
        n10249) );
  INV_X1 U12958 ( .A(n10249), .ZN(n10257) );
  AOI22_X1 U12959 ( .A1(n14729), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10256) );
  NAND2_X1 U12960 ( .A1(n14796), .A2(n10250), .ZN(n10255) );
  OAI211_X1 U12961 ( .C1(n10253), .C2(n10252), .A(n14819), .B(n10251), .ZN(
        n10254) );
  NAND4_X1 U12962 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n10270) );
  NAND2_X4 U12963 ( .A1(n14423), .A2(n11247), .ZN(n12322) );
  INV_X1 U12964 ( .A(n14043), .ZN(n10261) );
  INV_X1 U12965 ( .A(n12016), .ZN(n10258) );
  INV_X1 U12966 ( .A(n10259), .ZN(n10782) );
  NAND2_X1 U12967 ( .A1(n12358), .A2(n14043), .ZN(n10263) );
  NAND2_X1 U12968 ( .A1(n10782), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10262) );
  XNOR2_X1 U12969 ( .A(n10373), .B(n10375), .ZN(n10362) );
  INV_X1 U12970 ( .A(n10264), .ZN(n10265) );
  MUX2_X1 U12971 ( .A(n10362), .B(n10265), .S(n14727), .Z(n10269) );
  INV_X1 U12972 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10266) );
  AOI21_X1 U12973 ( .B1(n14727), .B2(n10266), .A(n14483), .ZN(n14726) );
  OAI21_X1 U12974 ( .B1(n6889), .B2(n14726), .A(n14042), .ZN(n10267) );
  AOI21_X1 U12975 ( .B1(n10269), .B2(n10268), .A(n10267), .ZN(n10312) );
  OR2_X1 U12976 ( .A1(n10270), .A2(n10312), .ZN(P1_U3245) );
  INV_X1 U12977 ( .A(n15023), .ZN(n10273) );
  OAI222_X1 U12978 ( .A1(P2_U3088), .A2(n10273), .B1(n13837), .B2(n10272), 
        .C1(n10271), .C2(n13839), .ZN(P2_U3311) );
  NAND2_X1 U12979 ( .A1(n10504), .A2(n6935), .ZN(n11854) );
  INV_X1 U12980 ( .A(n11854), .ZN(n10274) );
  NOR2_X1 U12981 ( .A1(n11856), .A2(n10274), .ZN(n11975) );
  NAND2_X1 U12982 ( .A1(n15339), .A2(n10281), .ZN(n10275) );
  OAI22_X1 U12983 ( .A1(n10282), .A2(n10275), .B1(n10291), .B2(n10285), .ZN(
        n10276) );
  NAND2_X1 U12984 ( .A1(n10413), .A2(n11974), .ZN(n12003) );
  NOR2_X1 U12985 ( .A1(n15143), .A2(n15315), .ZN(n12615) );
  NAND2_X1 U12986 ( .A1(n10282), .A2(n15327), .ZN(n10278) );
  AND2_X1 U12987 ( .A1(n15328), .A2(n10413), .ZN(n10277) );
  AOI22_X1 U12988 ( .A1(n10280), .A2(n12615), .B1(n15140), .B2(n10279), .ZN(
        n10296) );
  NAND2_X1 U12989 ( .A1(n10282), .A2(n10281), .ZN(n10289) );
  AND2_X1 U12990 ( .A1(n10284), .A2(n10283), .ZN(n10288) );
  INV_X1 U12991 ( .A(n10285), .ZN(n10286) );
  NAND2_X1 U12992 ( .A1(n10291), .A2(n10286), .ZN(n10287) );
  NAND2_X1 U12993 ( .A1(n11959), .A2(n10421), .ZN(n10415) );
  NAND4_X1 U12994 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10415), .ZN(
        n10290) );
  NAND2_X1 U12995 ( .A1(n10290), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10294) );
  INV_X1 U12996 ( .A(n10407), .ZN(n10292) );
  NAND3_X1 U12997 ( .A1(n10292), .A2(n10413), .A3(n10291), .ZN(n10293) );
  NAND2_X1 U12998 ( .A1(n15159), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10672) );
  NAND2_X1 U12999 ( .A1(n10672), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10295) );
  OAI211_X1 U13000 ( .C1(n11975), .C2(n15146), .A(n10296), .B(n10295), .ZN(
        P3_U3172) );
  INV_X1 U13001 ( .A(n11673), .ZN(n14994) );
  OAI222_X1 U13002 ( .A1(P2_U3088), .A2(n14994), .B1(n13837), .B2(n10298), 
        .C1(n10297), .C2(n13839), .ZN(P2_U3313) );
  INV_X1 U13003 ( .A(n10299), .ZN(n10313) );
  INV_X1 U13004 ( .A(n14063), .ZN(n14810) );
  OAI222_X1 U13005 ( .A1(n14494), .A2(n10313), .B1(n14810), .B2(P1_U3086), 
        .C1(n10300), .C2(n14490), .ZN(P1_U3338) );
  AOI211_X1 U13006 ( .C1(n10303), .C2(n10302), .A(n10301), .B(n14785), .ZN(
        n10311) );
  AOI211_X1 U13007 ( .C1(n10306), .C2(n10305), .A(n10304), .B(n14789), .ZN(
        n10310) );
  NAND2_X1 U13008 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U13009 ( .A1(n14729), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10307) );
  OAI211_X1 U13010 ( .C1(n14828), .C2(n10308), .A(n11262), .B(n10307), .ZN(
        n10309) );
  OR4_X1 U13011 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        P1_U3247) );
  INV_X1 U13012 ( .A(n11678), .ZN(n15036) );
  OAI222_X1 U13013 ( .A1(n13839), .A2(n10314), .B1(n13837), .B2(n10313), .C1(
        n15036), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13014 ( .A(n10315), .ZN(n10317) );
  AOI22_X1 U13015 ( .A1(n10319), .A2(n10318), .B1(n10317), .B2(n10316), .ZN(
        n13291) );
  NOR2_X1 U13016 ( .A1(n10664), .A2(n10749), .ZN(n10321) );
  XNOR2_X1 U13017 ( .A(n13295), .B(n13226), .ZN(n10320) );
  NOR2_X1 U13018 ( .A1(n10320), .A2(n10321), .ZN(n10322) );
  AOI21_X1 U13019 ( .B1(n10321), .B2(n10320), .A(n10322), .ZN(n13290) );
  NAND2_X1 U13020 ( .A1(n13291), .A2(n13290), .ZN(n13289) );
  INV_X1 U13021 ( .A(n10322), .ZN(n10323) );
  NAND2_X1 U13022 ( .A1(n13289), .A2(n10323), .ZN(n13262) );
  AND2_X1 U13023 ( .A1(n13369), .A2(n13191), .ZN(n10325) );
  XNOR2_X1 U13024 ( .A(n15078), .B(n13226), .ZN(n10324) );
  NOR2_X1 U13025 ( .A1(n10324), .A2(n10325), .ZN(n10326) );
  AOI21_X1 U13026 ( .B1(n10325), .B2(n10324), .A(n10326), .ZN(n13263) );
  INV_X1 U13027 ( .A(n10326), .ZN(n10327) );
  NOR2_X1 U13028 ( .A1(n10814), .A2(n10749), .ZN(n10486) );
  XNOR2_X1 U13029 ( .A(n15089), .B(n13226), .ZN(n10487) );
  XOR2_X1 U13030 ( .A(n10486), .B(n10487), .Z(n10488) );
  XNOR2_X1 U13031 ( .A(n10489), .B(n10488), .ZN(n10333) );
  NAND2_X1 U13032 ( .A1(n13368), .A2(n13409), .ZN(n10329) );
  NAND2_X1 U13033 ( .A1(n13369), .A2(n13331), .ZN(n10328) );
  NAND2_X1 U13034 ( .A1(n10329), .A2(n10328), .ZN(n15047) );
  NAND2_X1 U13035 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14928) );
  INV_X1 U13036 ( .A(n14928), .ZN(n10331) );
  OAI22_X1 U13037 ( .A1(n13354), .A2(n15089), .B1(n15051), .B2(n13336), .ZN(
        n10330) );
  AOI211_X1 U13038 ( .C1(n13334), .C2(n15047), .A(n10331), .B(n10330), .ZN(
        n10332) );
  OAI21_X1 U13039 ( .B1(n10333), .B2(n13339), .A(n10332), .ZN(P2_U3211) );
  INV_X1 U13040 ( .A(n10334), .ZN(n10367) );
  OAI222_X1 U13041 ( .A1(n14494), .A2(n10367), .B1(n14780), .B2(P1_U3086), 
        .C1(n10335), .C2(n14486), .ZN(P1_U3340) );
  AND2_X1 U13042 ( .A1(n15071), .A2(n10336), .ZN(n10337) );
  INV_X2 U13043 ( .A(n15117), .ZN(n15119) );
  NAND2_X1 U13044 ( .A1(n15119), .A2(n15079), .ZN(n13809) );
  OAI22_X1 U13045 ( .A1(n13809), .A2(n10339), .B1(n15119), .B2(n9137), .ZN(
        n10340) );
  INV_X1 U13046 ( .A(n10340), .ZN(n10341) );
  OAI21_X1 U13047 ( .B1(n10342), .B2(n15117), .A(n10341), .ZN(P2_U3439) );
  INV_X1 U13048 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10343) );
  OAI22_X1 U13049 ( .A1(n13809), .A2(n10344), .B1(n15119), .B2(n10343), .ZN(
        n10345) );
  INV_X1 U13050 ( .A(n10345), .ZN(n10346) );
  OAI21_X1 U13051 ( .B1(n10347), .B2(n15117), .A(n10346), .ZN(P2_U3436) );
  INV_X1 U13052 ( .A(n10880), .ZN(n10349) );
  NAND2_X1 U13053 ( .A1(n10355), .A2(n12237), .ZN(n10352) );
  NAND2_X1 U13054 ( .A1(n14852), .A2(n12191), .ZN(n10350) );
  INV_X1 U13055 ( .A(n12236), .ZN(n10351) );
  NOR2_X2 U13056 ( .A1(n13996), .A2(n14395), .ZN(n13950) );
  INV_X1 U13057 ( .A(n7904), .ZN(n14041) );
  OR2_X1 U13058 ( .A1(n10352), .A2(n10891), .ZN(n10354) );
  INV_X1 U13059 ( .A(n10356), .ZN(n10353) );
  AOI22_X1 U13060 ( .A1(n13950), .A2(n14041), .B1(n10446), .B2(n14012), .ZN(
        n10361) );
  INV_X1 U13061 ( .A(n10355), .ZN(n10357) );
  NAND2_X1 U13062 ( .A1(n10357), .A2(n10356), .ZN(n10358) );
  NAND2_X1 U13063 ( .A1(n10358), .A2(n12236), .ZN(n10783) );
  OR2_X1 U13064 ( .A1(n10783), .A2(n10359), .ZN(n10388) );
  NAND2_X1 U13065 ( .A1(n10388), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10360) );
  OAI211_X1 U13066 ( .C1(n10362), .C2(n14014), .A(n10361), .B(n10360), .ZN(
        P1_U3232) );
  INV_X1 U13067 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n15732) );
  NAND2_X1 U13068 ( .A1(n12522), .A2(P3_U3897), .ZN(n10363) );
  OAI21_X1 U13069 ( .B1(n10958), .B2(n15732), .A(n10363), .ZN(P3_U3515) );
  OAI22_X1 U13070 ( .A1(n13809), .A2(n9925), .B1(n15119), .B2(n9110), .ZN(
        n10364) );
  AOI21_X1 U13071 ( .B1(n15119), .B2(n10365), .A(n10364), .ZN(n10366) );
  INV_X1 U13072 ( .A(n10366), .ZN(P2_U3433) );
  OAI222_X1 U13073 ( .A1(n13839), .A2(n10368), .B1(n13837), .B2(n10367), .C1(
        n11674), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI22_X1 U13074 ( .A1(n13809), .A2(n10661), .B1(n15119), .B2(n9165), .ZN(
        n10369) );
  AOI21_X1 U13075 ( .B1(n10370), .B2(n15119), .A(n10369), .ZN(n10371) );
  INV_X1 U13076 ( .A(n10371), .ZN(P2_U3442) );
  OAI22_X1 U13077 ( .A1(n12322), .A2(n7904), .B1(n11001), .B2(n6683), .ZN(
        n10383) );
  XNOR2_X1 U13078 ( .A(n10372), .B(n12376), .ZN(n10384) );
  AOI21_X1 U13079 ( .B1(n10377), .B2(n10376), .A(n10385), .ZN(n10380) );
  NOR2_X2 U13080 ( .A1(n13996), .A2(n14316), .ZN(n14007) );
  AOI22_X1 U13081 ( .A1(n14007), .A2(n14043), .B1(n13950), .B2(n14040), .ZN(
        n10379) );
  AOI22_X1 U13082 ( .A1(n14012), .A2(n6967), .B1(n10388), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10378) );
  OAI211_X1 U13083 ( .C1(n10380), .C2(n14014), .A(n10379), .B(n10378), .ZN(
        P1_U3222) );
  OAI22_X1 U13084 ( .A1(n7127), .A2(n10381), .B1(n6683), .B2(n12021), .ZN(
        n10382) );
  XNOR2_X1 U13085 ( .A(n10382), .B(n12376), .ZN(n10790) );
  OAI22_X1 U13086 ( .A1(n12322), .A2(n12021), .B1(n7127), .B2(n6683), .ZN(
        n10789) );
  XNOR2_X1 U13087 ( .A(n10790), .B(n10789), .ZN(n10791) );
  INV_X1 U13088 ( .A(n10383), .ZN(n10387) );
  INV_X1 U13089 ( .A(n10384), .ZN(n10386) );
  XOR2_X1 U13090 ( .A(n10791), .B(n10792), .Z(n10391) );
  AOI22_X1 U13091 ( .A1(n14012), .A2(n12022), .B1(n10388), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13092 ( .A1(n14007), .A2(n14041), .B1(n13950), .B2(n6871), .ZN(
        n10389) );
  OAI211_X1 U13093 ( .C1(n10391), .C2(n14014), .A(n10390), .B(n10389), .ZN(
        P1_U3237) );
  INV_X1 U13094 ( .A(n10392), .ZN(n10704) );
  AOI21_X1 U13095 ( .B1(n15161), .B2(n10393), .A(n10704), .ZN(n10406) );
  INV_X1 U13096 ( .A(n10394), .ZN(n10396) );
  OAI21_X1 U13097 ( .B1(n10396), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10395), .ZN(
        n10402) );
  OAI22_X1 U13098 ( .A1(n15251), .A2(n15475), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10509), .ZN(n10401) );
  NAND2_X1 U13099 ( .A1(n10397), .A2(n9711), .ZN(n10398) );
  AOI21_X1 U13100 ( .B1(n10399), .B2(n10398), .A(n15266), .ZN(n10400) );
  AOI211_X1 U13101 ( .C1(n15262), .C2(n10402), .A(n10401), .B(n10400), .ZN(
        n10405) );
  NAND2_X1 U13102 ( .A1(n15259), .A2(n10403), .ZN(n10404) );
  OAI211_X1 U13103 ( .C1(n10406), .C2(n15253), .A(n10405), .B(n10404), .ZN(
        P3_U3183) );
  NAND2_X1 U13104 ( .A1(n10407), .A2(n15339), .ZN(n10408) );
  OR2_X1 U13105 ( .A1(n11975), .A2(n10408), .ZN(n10410) );
  OR2_X1 U13106 ( .A1(n15312), .A2(n15315), .ZN(n10409) );
  NAND2_X1 U13107 ( .A1(n10410), .A2(n10409), .ZN(n10478) );
  NAND2_X1 U13108 ( .A1(n11967), .A2(n10411), .ZN(n10472) );
  AND2_X1 U13109 ( .A1(n10413), .A2(n10412), .ZN(n10414) );
  AND2_X1 U13110 ( .A1(n10416), .A2(n10473), .ZN(n10417) );
  OAI211_X1 U13111 ( .C1(n10470), .C2(n10472), .A(n10475), .B(n10417), .ZN(
        n10426) );
  NAND2_X1 U13112 ( .A1(n15328), .A2(n6680), .ZN(n10420) );
  INV_X1 U13113 ( .A(n10418), .ZN(n10419) );
  NAND2_X1 U13114 ( .A1(n10420), .A2(n10419), .ZN(n10422) );
  NAND2_X1 U13115 ( .A1(n10422), .A2(n10421), .ZN(n10424) );
  AOI21_X1 U13116 ( .B1(n10424), .B2(n11967), .A(n10423), .ZN(n10425) );
  OAI22_X1 U13117 ( .A1(n13024), .A2(n6935), .B1(n15396), .B2(n9715), .ZN(
        n10427) );
  AOI21_X1 U13118 ( .B1(n10478), .B2(n15396), .A(n10427), .ZN(n10428) );
  INV_X1 U13119 ( .A(n10428), .ZN(P3_U3459) );
  MUX2_X1 U13120 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10429), .S(n10732), .Z(
        n10432) );
  OAI21_X1 U13121 ( .B1(n10437), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10430), .ZN(
        n10431) );
  NAND2_X1 U13122 ( .A1(n10431), .A2(n10432), .ZN(n10731) );
  OAI21_X1 U13123 ( .B1(n10432), .B2(n10431), .A(n10731), .ZN(n10442) );
  INV_X1 U13124 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10433) );
  NOR2_X1 U13125 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10433), .ZN(n11752) );
  AOI21_X1 U13126 ( .B1(n14729), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n11752), .ZN(
        n10434) );
  OAI21_X1 U13127 ( .B1(n14828), .B2(n10435), .A(n10434), .ZN(n10441) );
  XNOR2_X1 U13128 ( .A(n10732), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n10438) );
  NOR2_X1 U13129 ( .A1(n10439), .A2(n10438), .ZN(n10726) );
  AOI211_X1 U13130 ( .C1(n10439), .C2(n10438), .A(n14789), .B(n10726), .ZN(
        n10440) );
  AOI211_X1 U13131 ( .C1(n14819), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        n10443) );
  INV_X1 U13132 ( .A(n10443), .ZN(P1_U3252) );
  NAND2_X1 U13133 ( .A1(n14043), .A2(n12017), .ZN(n10444) );
  AND2_X1 U13134 ( .A1(n12019), .A2(n10444), .ZN(n12203) );
  INV_X1 U13135 ( .A(n12203), .ZN(n10445) );
  OAI21_X1 U13136 ( .B1(n14688), .B2(n14855), .A(n10445), .ZN(n10449) );
  AOI22_X1 U13137 ( .A1(n14041), .A2(n14239), .B1(n10447), .B2(n10446), .ZN(
        n10448) );
  AND2_X1 U13138 ( .A1(n10449), .A2(n10448), .ZN(n14835) );
  NAND2_X1 U13139 ( .A1(n14861), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10450) );
  OAI21_X1 U13140 ( .B1(n14861), .B2(n14835), .A(n10450), .ZN(P1_U3528) );
  OAI22_X1 U13141 ( .A1(n13114), .A2(n6935), .B1(n15382), .B2(n8495), .ZN(
        n10451) );
  AOI21_X1 U13142 ( .B1(n10478), .B2(n15382), .A(n10451), .ZN(n10452) );
  INV_X1 U13143 ( .A(n10452), .ZN(P3_U3390) );
  OAI222_X1 U13144 ( .A1(P3_U3151), .A2(n6680), .B1(n13130), .B2(n10454), .C1(
        n11825), .C2(n10453), .ZN(P3_U3275) );
  NAND2_X1 U13145 ( .A1(n15071), .A2(n10455), .ZN(n10456) );
  OR2_X1 U13146 ( .A1(n10457), .A2(n10456), .ZN(n10458) );
  NAND2_X1 U13147 ( .A1(n13643), .A2(n10459), .ZN(n11340) );
  INV_X1 U13148 ( .A(n15052), .ZN(n13674) );
  NOR2_X1 U13149 ( .A1(n10461), .A2(n10460), .ZN(n10462) );
  NOR2_X1 U13150 ( .A1(n10463), .A2(n10462), .ZN(n10464) );
  NOR2_X1 U13151 ( .A1(n15067), .A2(n10464), .ZN(n10467) );
  INV_X1 U13152 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10465) );
  NOR2_X1 U13153 ( .A1(n13643), .A2(n10465), .ZN(n10466) );
  AOI211_X1 U13154 ( .C1(n13674), .C2(P2_REG3_REG_0__SCAN_IN), .A(n10467), .B(
        n10466), .ZN(n10468) );
  OAI21_X1 U13155 ( .B1(n10469), .B2(n11340), .A(n10468), .ZN(P2_U3265) );
  NAND2_X1 U13156 ( .A1(n10472), .A2(n10470), .ZN(n10471) );
  OAI21_X1 U13157 ( .B1(n10472), .B2(n13116), .A(n10471), .ZN(n10474) );
  NAND3_X1 U13158 ( .A1(n10475), .A2(n10474), .A3(n10473), .ZN(n10480) );
  NOR2_X1 U13159 ( .A1(n10476), .A2(n15327), .ZN(n10477) );
  MUX2_X1 U13160 ( .A(n10478), .B(P3_REG2_REG_0__SCAN_IN), .S(n15337), .Z(
        n10479) );
  INV_X1 U13161 ( .A(n10479), .ZN(n10484) );
  INV_X1 U13162 ( .A(n15327), .ZN(n11973) );
  OR2_X1 U13163 ( .A1(n10480), .A2(n11973), .ZN(n11375) );
  NAND2_X1 U13164 ( .A1(n15295), .A2(n15328), .ZN(n14652) );
  OAI22_X1 U13165 ( .A1(n14652), .A2(n6935), .B1(n8493), .B2(n15307), .ZN(
        n10482) );
  INV_X1 U13166 ( .A(n10482), .ZN(n10483) );
  NAND2_X1 U13167 ( .A1(n10484), .A2(n10483), .ZN(P3_U3233) );
  INV_X1 U13168 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n15565) );
  NAND2_X1 U13169 ( .A1(n12821), .A2(P3_U3897), .ZN(n10485) );
  OAI21_X1 U13170 ( .B1(P3_U3897), .B2(n15565), .A(n10485), .ZN(P3_U3516) );
  XNOR2_X1 U13171 ( .A(n10817), .B(n13226), .ZN(n10745) );
  NAND2_X1 U13172 ( .A1(n13368), .A2(n13651), .ZN(n10744) );
  XNOR2_X1 U13173 ( .A(n10745), .B(n10744), .ZN(n10747) );
  XNOR2_X1 U13174 ( .A(n10748), .B(n10747), .ZN(n10493) );
  OAI22_X1 U13175 ( .A1(n10823), .A2(n13312), .B1(n10814), .B2(n13448), .ZN(
        n10835) );
  AOI22_X1 U13176 ( .A1(n13334), .A2(n10835), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10490) );
  OAI21_X1 U13177 ( .B1(n10830), .B2(n13336), .A(n10490), .ZN(n10491) );
  AOI21_X1 U13178 ( .B1(n10817), .B2(n9967), .A(n10491), .ZN(n10492) );
  OAI21_X1 U13179 ( .B1(n10493), .B2(n13339), .A(n10492), .ZN(P2_U3185) );
  INV_X1 U13180 ( .A(n10672), .ZN(n10510) );
  NAND2_X1 U13181 ( .A1(n10677), .A2(n12742), .ZN(n10495) );
  NAND2_X1 U13182 ( .A1(n10495), .A2(n6680), .ZN(n10496) );
  OR2_X1 U13183 ( .A1(n15312), .A2(n10497), .ZN(n10499) );
  NAND2_X1 U13184 ( .A1(n15312), .A2(n10498), .ZN(n10668) );
  AND2_X1 U13185 ( .A1(n15320), .A2(n12484), .ZN(n10500) );
  OAI21_X1 U13186 ( .B1(n10500), .B2(n15299), .A(n10502), .ZN(n10669) );
  INV_X1 U13187 ( .A(n11856), .ZN(n15325) );
  NAND3_X1 U13188 ( .A1(n15325), .A2(n15324), .A3(n12435), .ZN(n10501) );
  OAI211_X1 U13189 ( .C1(n10502), .C2(n15320), .A(n10669), .B(n10501), .ZN(
        n10503) );
  NAND2_X1 U13190 ( .A1(n10503), .A2(n15134), .ZN(n10508) );
  NAND2_X1 U13191 ( .A1(n10504), .A2(n12946), .ZN(n10506) );
  NAND2_X1 U13192 ( .A1(n11853), .A2(n12948), .ZN(n10505) );
  NAND2_X1 U13193 ( .A1(n10506), .A2(n10505), .ZN(n15321) );
  AOI22_X1 U13194 ( .A1(n15321), .A2(n15149), .B1(n15140), .B2(n15329), .ZN(
        n10507) );
  OAI211_X1 U13195 ( .C1(n10510), .C2(n10509), .A(n10508), .B(n10507), .ZN(
        P3_U3162) );
  OAI21_X1 U13196 ( .B1(n10512), .B2(n7182), .A(n10511), .ZN(n10887) );
  NAND2_X1 U13197 ( .A1(n10622), .A2(n12033), .ZN(n10513) );
  NAND2_X1 U13198 ( .A1(n10513), .A2(n14248), .ZN(n10514) );
  NOR2_X1 U13199 ( .A1(n10548), .A2(n10514), .ZN(n10890) );
  XNOR2_X1 U13200 ( .A(n10515), .B(n12202), .ZN(n10516) );
  OAI22_X1 U13201 ( .A1(n12039), .A2(n14395), .B1(n12021), .B2(n14316), .ZN(
        n10785) );
  AOI21_X1 U13202 ( .B1(n10516), .B2(n14688), .A(n10785), .ZN(n10898) );
  INV_X1 U13203 ( .A(n10898), .ZN(n10517) );
  AOI211_X1 U13204 ( .C1(n14855), .C2(n10887), .A(n10890), .B(n10517), .ZN(
        n10721) );
  INV_X1 U13205 ( .A(n14852), .ZN(n14680) );
  AOI22_X1 U13206 ( .A1(n14345), .A2(n12033), .B1(n14861), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n10518) );
  OAI21_X1 U13207 ( .B1(n10721), .B2(n14861), .A(n10518), .ZN(P1_U3531) );
  INV_X1 U13208 ( .A(n10623), .ZN(n14842) );
  OAI21_X1 U13209 ( .B1(n12200), .B2(n10520), .A(n10519), .ZN(n11006) );
  OAI21_X1 U13210 ( .B1(n11001), .B2(n12017), .A(n10621), .ZN(n11002) );
  OAI22_X1 U13211 ( .A1(n14395), .A2(n12021), .B1(n11002), .B2(n14423), .ZN(
        n10524) );
  XNOR2_X1 U13212 ( .A(n14041), .B(n11002), .ZN(n10521) );
  MUX2_X1 U13213 ( .A(n10521), .B(n12200), .S(n14043), .Z(n10522) );
  INV_X1 U13214 ( .A(n14283), .ZN(n11421) );
  AOI222_X1 U13215 ( .A1(n10522), .A2(n14688), .B1(n11006), .B2(n11421), .C1(
        n14043), .C2(n14238), .ZN(n11007) );
  INV_X1 U13216 ( .A(n11007), .ZN(n10523) );
  AOI211_X1 U13217 ( .C1(n14842), .C2(n11006), .A(n10524), .B(n10523), .ZN(
        n10717) );
  AOI22_X1 U13218 ( .A1(n14345), .A2(n6967), .B1(n14861), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n10525) );
  OAI21_X1 U13219 ( .B1(n10717), .B2(n14861), .A(n10525), .ZN(P1_U3529) );
  INV_X1 U13220 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15750) );
  NOR2_X1 U13221 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15750), .ZN(n10532) );
  INV_X1 U13222 ( .A(n10526), .ZN(n10530) );
  NAND3_X1 U13223 ( .A1(n10598), .A2(n10528), .A3(n10527), .ZN(n10529) );
  AOI21_X1 U13224 ( .B1(n10530), .B2(n10529), .A(n15241), .ZN(n10531) );
  AOI211_X1 U13225 ( .C1(n15232), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n10532), .B(
        n10531), .ZN(n10538) );
  AND3_X1 U13226 ( .A1(n10595), .A2(n10534), .A3(n10533), .ZN(n10535) );
  INV_X1 U13227 ( .A(n15266), .ZN(n10700) );
  OAI21_X1 U13228 ( .B1(n10536), .B2(n10535), .A(n10700), .ZN(n10537) );
  OAI211_X1 U13229 ( .C1(n15235), .C2(n10539), .A(n10538), .B(n10537), .ZN(
        n10545) );
  INV_X1 U13230 ( .A(n10540), .ZN(n10541) );
  NAND3_X1 U13231 ( .A1(n10608), .A2(n10542), .A3(n10541), .ZN(n10543) );
  AOI21_X1 U13232 ( .B1(n10558), .B2(n10543), .A(n15253), .ZN(n10544) );
  OR2_X1 U13233 ( .A1(n10545), .A2(n10544), .ZN(P3_U3186) );
  OAI21_X1 U13234 ( .B1(n10547), .B2(n12204), .A(n10546), .ZN(n10985) );
  OAI211_X1 U13235 ( .C1(n10548), .C2(n12038), .A(n11045), .B(n14248), .ZN(
        n10551) );
  NAND2_X1 U13236 ( .A1(n14239), .A2(n14037), .ZN(n10550) );
  NAND2_X1 U13237 ( .A1(n6871), .A2(n14238), .ZN(n10549) );
  AND2_X1 U13238 ( .A1(n10550), .A2(n10549), .ZN(n11263) );
  NAND2_X1 U13239 ( .A1(n10551), .A2(n11263), .ZN(n10980) );
  XNOR2_X1 U13240 ( .A(n12204), .B(n10552), .ZN(n10553) );
  NOR2_X1 U13241 ( .A1(n10553), .A2(n14352), .ZN(n10979) );
  AOI211_X1 U13242 ( .C1(n14855), .C2(n10985), .A(n10980), .B(n10979), .ZN(
        n10725) );
  AOI22_X1 U13243 ( .A1(n14345), .A2(n12041), .B1(n14861), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n10554) );
  OAI21_X1 U13244 ( .B1(n10725), .B2(n14861), .A(n10554), .ZN(P1_U3532) );
  INV_X1 U13245 ( .A(n10555), .ZN(n10556) );
  NAND3_X1 U13246 ( .A1(n10558), .A2(n10557), .A3(n10556), .ZN(n10559) );
  AOI21_X1 U13247 ( .B1(n10575), .B2(n10559), .A(n15253), .ZN(n10569) );
  AOI21_X1 U13248 ( .B1(n10561), .B2(n9734), .A(n10560), .ZN(n10567) );
  NOR2_X1 U13249 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8550), .ZN(n10565) );
  AOI21_X1 U13250 ( .B1(n6725), .B2(n9733), .A(n10562), .ZN(n10563) );
  NOR2_X1 U13251 ( .A1(n10563), .A2(n15241), .ZN(n10564) );
  AOI211_X1 U13252 ( .C1(n15232), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n10565), .B(
        n10564), .ZN(n10566) );
  OAI21_X1 U13253 ( .B1(n10567), .B2(n15266), .A(n10566), .ZN(n10568) );
  AOI211_X1 U13254 ( .C1(n15259), .C2(n10570), .A(n10569), .B(n10568), .ZN(
        n10571) );
  INV_X1 U13255 ( .A(n10571), .ZN(P3_U3187) );
  INV_X1 U13256 ( .A(n10572), .ZN(n10573) );
  NAND3_X1 U13257 ( .A1(n10575), .A2(n10574), .A3(n10573), .ZN(n10576) );
  AOI21_X1 U13258 ( .B1(n10635), .B2(n10576), .A(n15253), .ZN(n10590) );
  AOI21_X1 U13259 ( .B1(n10579), .B2(n10578), .A(n10577), .ZN(n10588) );
  INV_X1 U13260 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10580) );
  NOR2_X1 U13261 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10580), .ZN(n10586) );
  AOI21_X1 U13262 ( .B1(n10583), .B2(n10582), .A(n10581), .ZN(n10584) );
  NOR2_X1 U13263 ( .A1(n15241), .A2(n10584), .ZN(n10585) );
  AOI211_X1 U13264 ( .C1(n15232), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n10586), .B(
        n10585), .ZN(n10587) );
  OAI21_X1 U13265 ( .B1(n10588), .B2(n15266), .A(n10587), .ZN(n10589) );
  AOI211_X1 U13266 ( .C1(n15259), .C2(n10591), .A(n10590), .B(n10589), .ZN(
        n10592) );
  INV_X1 U13267 ( .A(n10592), .ZN(P3_U3188) );
  NAND2_X1 U13268 ( .A1(n10593), .A2(n11018), .ZN(n10594) );
  AND2_X1 U13269 ( .A1(n10595), .A2(n10594), .ZN(n10603) );
  NAND2_X1 U13270 ( .A1(n10596), .A2(n9723), .ZN(n10597) );
  NAND2_X1 U13271 ( .A1(n10598), .A2(n10597), .ZN(n10599) );
  NAND2_X1 U13272 ( .A1(n15262), .A2(n10599), .ZN(n10602) );
  INV_X1 U13273 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11020) );
  NOR2_X1 U13274 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11020), .ZN(n10600) );
  AOI21_X1 U13275 ( .B1(n15232), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10600), .ZN(
        n10601) );
  OAI211_X1 U13276 ( .C1(n15266), .C2(n10603), .A(n10602), .B(n10601), .ZN(
        n10610) );
  INV_X1 U13277 ( .A(n10604), .ZN(n10605) );
  NAND3_X1 U13278 ( .A1(n10705), .A2(n10606), .A3(n10605), .ZN(n10607) );
  AOI21_X1 U13279 ( .B1(n10608), .B2(n10607), .A(n15253), .ZN(n10609) );
  AOI211_X1 U13280 ( .C1(n15259), .C2(n10611), .A(n10610), .B(n10609), .ZN(
        n10612) );
  INV_X1 U13281 ( .A(n10612), .ZN(P3_U3185) );
  OAI21_X1 U13282 ( .B1(n10614), .B2(n10615), .A(n10613), .ZN(n10620) );
  INV_X1 U13283 ( .A(n10620), .ZN(n10905) );
  OAI22_X1 U13284 ( .A1(n10788), .A2(n14395), .B1(n7904), .B2(n14316), .ZN(
        n10619) );
  XNOR2_X1 U13285 ( .A(n10616), .B(n10615), .ZN(n10617) );
  NOR2_X1 U13286 ( .A1(n10617), .A2(n14352), .ZN(n10618) );
  AOI211_X1 U13287 ( .C1(n11421), .C2(n10620), .A(n10619), .B(n10618), .ZN(
        n10902) );
  OAI211_X1 U13288 ( .C1(n7128), .C2(n7127), .A(n14248), .B(n10622), .ZN(
        n10900) );
  OAI211_X1 U13289 ( .C1(n10905), .C2(n10623), .A(n10902), .B(n10900), .ZN(
        n10742) );
  OAI22_X1 U13290 ( .A1(n14419), .A2(n7127), .B1(n14863), .B2(n10096), .ZN(
        n10624) );
  AOI21_X1 U13291 ( .B1(n14863), .B2(n10742), .A(n10624), .ZN(n10625) );
  INV_X1 U13292 ( .A(n10625), .ZN(P1_U3530) );
  AOI21_X1 U13293 ( .B1(n9744), .B2(n10627), .A(n10626), .ZN(n10628) );
  OR2_X1 U13294 ( .A1(n10628), .A2(n15266), .ZN(n10630) );
  INV_X1 U13295 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15730) );
  NOR2_X1 U13296 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15730), .ZN(n15138) );
  AOI21_X1 U13297 ( .B1(n15232), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n15138), .ZN(
        n10629) );
  OAI211_X1 U13298 ( .C1(n15235), .C2(n10631), .A(n10630), .B(n10629), .ZN(
        n10643) );
  INV_X1 U13299 ( .A(n10632), .ZN(n10633) );
  NAND3_X1 U13300 ( .A1(n10635), .A2(n10634), .A3(n10633), .ZN(n10636) );
  AOI21_X1 U13301 ( .B1(n10637), .B2(n10636), .A(n15253), .ZN(n10642) );
  AOI21_X1 U13302 ( .B1(n9743), .B2(n10639), .A(n10638), .ZN(n10640) );
  NOR2_X1 U13303 ( .A1(n10640), .A2(n15241), .ZN(n10641) );
  OR3_X1 U13304 ( .A1(n10643), .A2(n10642), .A3(n10641), .ZN(P3_U3189) );
  INV_X1 U13305 ( .A(n6873), .ZN(n15106) );
  NAND2_X1 U13306 ( .A1(n13643), .A2(n15106), .ZN(n10644) );
  NOR2_X2 U13307 ( .A1(n15067), .A2(n10645), .ZN(n15055) );
  NOR2_X1 U13308 ( .A1(n15052), .A2(n13293), .ZN(n10648) );
  NAND2_X1 U13309 ( .A1(n13643), .A2(n13400), .ZN(n15062) );
  NOR2_X1 U13310 ( .A1(n15062), .A2(n10646), .ZN(n10647) );
  AOI211_X1 U13311 ( .C1(n15055), .C2(n13295), .A(n10648), .B(n10647), .ZN(
        n10651) );
  MUX2_X1 U13312 ( .A(n10649), .B(n9857), .S(n15067), .Z(n10650) );
  OAI211_X1 U13313 ( .C1(n15063), .C2(n10652), .A(n10651), .B(n10650), .ZN(
        P2_U3261) );
  NAND2_X1 U13314 ( .A1(n10661), .A2(n10664), .ZN(n10653) );
  XNOR2_X1 U13315 ( .A(n10799), .B(n10810), .ZN(n15082) );
  AOI211_X1 U13316 ( .C1(n15078), .C2(n10656), .A(n13191), .B(n15061), .ZN(
        n15077) );
  NAND2_X1 U13317 ( .A1(n15055), .A2(n15078), .ZN(n10657) );
  OAI21_X1 U13318 ( .B1(n15052), .B2(n13265), .A(n10657), .ZN(n10658) );
  AOI21_X1 U13319 ( .B1(n13673), .B2(n15077), .A(n10658), .ZN(n10667) );
  NAND2_X1 U13320 ( .A1(n10660), .A2(n10659), .ZN(n10663) );
  OR2_X1 U13321 ( .A1(n13370), .A2(n10661), .ZN(n10662) );
  NAND2_X1 U13322 ( .A1(n10663), .A2(n10662), .ZN(n10811) );
  XNOR2_X1 U13323 ( .A(n10811), .B(n10810), .ZN(n10665) );
  OAI22_X1 U13324 ( .A1(n10814), .A2(n13312), .B1(n10664), .B2(n13448), .ZN(
        n13267) );
  AOI21_X1 U13325 ( .B1(n10665), .B2(n15048), .A(n13267), .ZN(n15080) );
  MUX2_X1 U13326 ( .A(n15080), .B(n9859), .S(n15067), .Z(n10666) );
  OAI211_X1 U13327 ( .C1(n15063), .C2(n15082), .A(n10667), .B(n10666), .ZN(
        P2_U3260) );
  XNOR2_X1 U13328 ( .A(n6682), .B(n12484), .ZN(n10759) );
  XNOR2_X1 U13329 ( .A(n10759), .B(n11853), .ZN(n10762) );
  NAND2_X1 U13330 ( .A1(n10669), .A2(n10668), .ZN(n10763) );
  XOR2_X1 U13331 ( .A(n10762), .B(n10763), .Z(n10674) );
  NAND2_X1 U13332 ( .A1(n15149), .A2(n12946), .ZN(n12617) );
  NOR2_X1 U13333 ( .A1(n15312), .A2(n12617), .ZN(n10671) );
  INV_X1 U13334 ( .A(n12615), .ZN(n12578) );
  INV_X1 U13335 ( .A(n15140), .ZN(n15154) );
  OAI22_X1 U13336 ( .A1(n12578), .A2(n15314), .B1(n15154), .B2(n6682), .ZN(
        n10670) );
  AOI211_X1 U13337 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n10672), .A(n10671), .B(
        n10670), .ZN(n10673) );
  OAI21_X1 U13338 ( .B1(n10674), .B2(n15146), .A(n10673), .ZN(P3_U3177) );
  OAI222_X1 U13339 ( .A1(P3_U3151), .A2(n10677), .B1(n13130), .B2(n10676), 
        .C1(n11825), .C2(n10675), .ZN(P3_U3274) );
  INV_X1 U13340 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n15533) );
  NAND2_X1 U13341 ( .A1(n12523), .A2(n10958), .ZN(n10678) );
  OAI21_X1 U13342 ( .B1(P3_U3897), .B2(n15533), .A(n10678), .ZN(P3_U3517) );
  XNOR2_X1 U13343 ( .A(n10679), .B(n7693), .ZN(n11235) );
  OAI21_X1 U13344 ( .B1(n10682), .B2(n10681), .A(n10680), .ZN(n10683) );
  INV_X1 U13345 ( .A(n10683), .ZN(n11238) );
  AOI22_X1 U13346 ( .A1(n14035), .A2(n14239), .B1(n14238), .B2(n14037), .ZN(
        n11231) );
  NAND2_X1 U13347 ( .A1(n11046), .A2(n12052), .ZN(n10684) );
  NAND2_X1 U13348 ( .A1(n10684), .A2(n14248), .ZN(n10685) );
  OR2_X1 U13349 ( .A1(n10685), .A2(n11094), .ZN(n11232) );
  OAI211_X1 U13350 ( .C1(n11238), .C2(n14684), .A(n11231), .B(n11232), .ZN(
        n10686) );
  AOI21_X1 U13351 ( .B1(n14688), .B2(n11235), .A(n10686), .ZN(n10714) );
  INV_X1 U13352 ( .A(n12052), .ZN(n11407) );
  INV_X1 U13353 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10687) );
  OAI22_X1 U13354 ( .A1(n14419), .A2(n11407), .B1(n14863), .B2(n10687), .ZN(
        n10688) );
  INV_X1 U13355 ( .A(n10688), .ZN(n10689) );
  OAI21_X1 U13356 ( .B1(n10714), .B2(n14861), .A(n10689), .ZN(P1_U3534) );
  OAI21_X1 U13357 ( .B1(n10692), .B2(n10691), .A(n10690), .ZN(n10699) );
  OAI21_X1 U13358 ( .B1(n10695), .B2(n10694), .A(n10693), .ZN(n10696) );
  AND2_X1 U13359 ( .A1(n15262), .A2(n10696), .ZN(n10698) );
  INV_X1 U13360 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14501) );
  OAI22_X1 U13361 ( .A1(n15251), .A2(n14501), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8508), .ZN(n10697) );
  AOI211_X1 U13362 ( .C1(n10700), .C2(n10699), .A(n10698), .B(n10697), .ZN(
        n10709) );
  INV_X1 U13363 ( .A(n10701), .ZN(n10703) );
  NOR3_X1 U13364 ( .A1(n10704), .A2(n10703), .A3(n10702), .ZN(n10707) );
  INV_X1 U13365 ( .A(n10705), .ZN(n10706) );
  INV_X1 U13366 ( .A(n15253), .ZN(n15237) );
  OAI21_X1 U13367 ( .B1(n10707), .B2(n10706), .A(n15237), .ZN(n10708) );
  OAI211_X1 U13368 ( .C1(n15235), .C2(n10710), .A(n10709), .B(n10708), .ZN(
        P3_U3184) );
  INV_X1 U13369 ( .A(n14436), .ZN(n14469) );
  INV_X1 U13370 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10711) );
  OAI22_X1 U13371 ( .A1(n14469), .A2(n11407), .B1(n14857), .B2(n10711), .ZN(
        n10712) );
  INV_X1 U13372 ( .A(n10712), .ZN(n10713) );
  OAI21_X1 U13373 ( .B1(n10714), .B2(n9673), .A(n10713), .ZN(P1_U3477) );
  OAI22_X1 U13374 ( .A1(n14469), .A2(n11001), .B1(n14857), .B2(n7886), .ZN(
        n10715) );
  INV_X1 U13375 ( .A(n10715), .ZN(n10716) );
  OAI21_X1 U13376 ( .B1(n10717), .B2(n9673), .A(n10716), .ZN(P1_U3462) );
  INV_X1 U13377 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10718) );
  OAI22_X1 U13378 ( .A1(n14469), .A2(n12034), .B1(n14857), .B2(n10718), .ZN(
        n10719) );
  INV_X1 U13379 ( .A(n10719), .ZN(n10720) );
  OAI21_X1 U13380 ( .B1(n10721), .B2(n9673), .A(n10720), .ZN(P1_U3468) );
  INV_X1 U13381 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10722) );
  OAI22_X1 U13382 ( .A1(n14469), .A2(n12038), .B1(n14857), .B2(n10722), .ZN(
        n10723) );
  INV_X1 U13383 ( .A(n10723), .ZN(n10724) );
  OAI21_X1 U13384 ( .B1(n10725), .B2(n9673), .A(n10724), .ZN(P1_U3471) );
  INV_X1 U13385 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10727) );
  MUX2_X1 U13386 ( .A(n10727), .B(P1_REG2_REG_10__SCAN_IN), .S(n11174), .Z(
        n10728) );
  AOI211_X1 U13387 ( .C1(n10729), .C2(n10728), .A(n14789), .B(n11168), .ZN(
        n10740) );
  INV_X1 U13388 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10730) );
  MUX2_X1 U13389 ( .A(n10730), .B(P1_REG1_REG_10__SCAN_IN), .S(n11174), .Z(
        n10734) );
  OAI21_X1 U13390 ( .B1(n10732), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10731), .ZN(
        n10733) );
  NOR2_X1 U13391 ( .A1(n10733), .A2(n10734), .ZN(n11173) );
  AOI211_X1 U13392 ( .C1(n10734), .C2(n10733), .A(n14785), .B(n11173), .ZN(
        n10739) );
  NAND2_X1 U13393 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10736)
         );
  NAND2_X1 U13394 ( .A1(n14729), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10735) );
  OAI211_X1 U13395 ( .C1(n14828), .C2(n10737), .A(n10736), .B(n10735), .ZN(
        n10738) );
  OR3_X1 U13396 ( .A1(n10740), .A2(n10739), .A3(n10738), .ZN(P1_U3253) );
  OAI22_X1 U13397 ( .A1(n14469), .A2(n7127), .B1(n14857), .B2(n7906), .ZN(
        n10741) );
  AOI21_X1 U13398 ( .B1(n14857), .B2(n10742), .A(n10741), .ZN(n10743) );
  INV_X1 U13399 ( .A(n10743), .ZN(P1_U3465) );
  INV_X1 U13400 ( .A(n10744), .ZN(n10746) );
  NOR2_X1 U13401 ( .A1(n10823), .A2(n10749), .ZN(n10751) );
  XNOR2_X1 U13402 ( .A(n15103), .B(n13186), .ZN(n10750) );
  NOR2_X1 U13403 ( .A1(n10750), .A2(n10751), .ZN(n10912) );
  AOI21_X1 U13404 ( .B1(n10751), .B2(n10750), .A(n10912), .ZN(n10752) );
  OAI21_X1 U13405 ( .B1(n10753), .B2(n10752), .A(n10914), .ZN(n10754) );
  NAND2_X1 U13406 ( .A1(n10754), .A2(n13343), .ZN(n10758) );
  INV_X1 U13407 ( .A(n10755), .ZN(n10849) );
  INV_X1 U13408 ( .A(n13336), .ZN(n13350) );
  AOI22_X1 U13409 ( .A1(n13366), .A2(n13409), .B1(n13331), .B2(n13368), .ZN(
        n10855) );
  NAND2_X1 U13410 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14953) );
  OAI21_X1 U13411 ( .B1(n13348), .B2(n10855), .A(n14953), .ZN(n10756) );
  AOI21_X1 U13412 ( .B1(n10849), .B2(n13350), .A(n10756), .ZN(n10757) );
  OAI211_X1 U13413 ( .C1(n15103), .C2(n13354), .A(n10758), .B(n10757), .ZN(
        P2_U3193) );
  INV_X1 U13414 ( .A(n10759), .ZN(n10760) );
  NOR2_X1 U13415 ( .A1(n10760), .A2(n11853), .ZN(n10761) );
  AOI21_X2 U13416 ( .B1(n10763), .B2(n10762), .A(n10761), .ZN(n10766) );
  XNOR2_X1 U13417 ( .A(n10764), .B(n12484), .ZN(n10987) );
  XNOR2_X1 U13418 ( .A(n10987), .B(n15314), .ZN(n10765) );
  NAND2_X1 U13419 ( .A1(n10766), .A2(n10765), .ZN(n10990) );
  OAI211_X1 U13420 ( .C1(n10766), .C2(n10765), .A(n10990), .B(n15134), .ZN(
        n10770) );
  INV_X1 U13421 ( .A(n12617), .ZN(n12575) );
  OAI22_X1 U13422 ( .A1(n12578), .A2(n11317), .B1(n15154), .B2(n11019), .ZN(
        n10768) );
  MUX2_X1 U13423 ( .A(n12619), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n10767) );
  AOI211_X1 U13424 ( .C1(n12575), .C2(n11853), .A(n10768), .B(n10767), .ZN(
        n10769) );
  NAND2_X1 U13425 ( .A1(n10770), .A2(n10769), .ZN(P3_U3158) );
  NOR2_X1 U13426 ( .A1(n13130), .A2(SI_22_), .ZN(n10771) );
  AOI21_X1 U13427 ( .B1(n10772), .B2(P3_STATE_REG_SCAN_IN), .A(n10771), .ZN(
        n10773) );
  OAI21_X1 U13428 ( .B1(n10774), .B2(n11825), .A(n10773), .ZN(n10775) );
  INV_X1 U13429 ( .A(n10775), .ZN(P3_U3273) );
  INV_X1 U13430 ( .A(n10776), .ZN(n10778) );
  INV_X1 U13431 ( .A(n13388), .ZN(n11679) );
  OAI222_X1 U13432 ( .A1(n13839), .A2(n10777), .B1(n13837), .B2(n10778), .C1(
        P2_U3088), .C2(n11679), .ZN(P2_U3309) );
  OAI222_X1 U13433 ( .A1(n14486), .A2(n10779), .B1(n14494), .B2(n10778), .C1(
        P1_U3086), .C2(n14827), .ZN(P1_U3337) );
  INV_X1 U13434 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n15477) );
  NAND2_X1 U13435 ( .A1(n10780), .A2(P3_U3897), .ZN(n10781) );
  OAI21_X1 U13436 ( .B1(P3_U3897), .B2(n15477), .A(n10781), .ZN(P3_U3518) );
  INV_X1 U13437 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10889) );
  OAI21_X1 U13438 ( .B1(n10783), .B2(n10782), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n10784) );
  INV_X1 U13439 ( .A(n14010), .ZN(n13999) );
  INV_X1 U13440 ( .A(n13996), .ZN(n13863) );
  AOI22_X1 U13441 ( .A1(n13863), .A2(n10785), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10786) );
  OAI21_X1 U13442 ( .B1(n12034), .B2(n14002), .A(n10786), .ZN(n10796) );
  OAI22_X1 U13443 ( .A1(n12322), .A2(n10788), .B1(n12034), .B2(n6683), .ZN(
        n11239) );
  AOI211_X1 U13444 ( .C1(n10794), .C2(n10793), .A(n14014), .B(n6835), .ZN(
        n10795) );
  AOI211_X1 U13445 ( .C1(n10889), .C2(n13999), .A(n10796), .B(n10795), .ZN(
        n10797) );
  INV_X1 U13446 ( .A(n10797), .ZN(P1_U3218) );
  OR2_X1 U13447 ( .A1(n15089), .A2(n10814), .ZN(n10802) );
  INV_X1 U13448 ( .A(n10815), .ZN(n10833) );
  NAND2_X1 U13449 ( .A1(n10817), .A2(n13368), .ZN(n10803) );
  NAND2_X1 U13450 ( .A1(n10827), .A2(n10803), .ZN(n10842) );
  INV_X1 U13451 ( .A(n10852), .ZN(n10841) );
  NAND2_X1 U13452 ( .A1(n10842), .A2(n10841), .ZN(n10844) );
  OR2_X1 U13453 ( .A1(n15103), .A2(n10823), .ZN(n10804) );
  INV_X1 U13454 ( .A(n10821), .ZN(n11113) );
  XNOR2_X1 U13455 ( .A(n11114), .B(n11113), .ZN(n10972) );
  OAI22_X1 U13456 ( .A1(n13643), .A2(n10805), .B1(n10920), .B2(n15052), .ZN(
        n10808) );
  INV_X1 U13457 ( .A(n11129), .ZN(n10806) );
  OAI211_X1 U13458 ( .C1(n11120), .C2(n10847), .A(n10806), .B(n10749), .ZN(
        n10970) );
  NOR2_X1 U13459 ( .A1(n10970), .A2(n15062), .ZN(n10807) );
  AOI211_X1 U13460 ( .C1(n15055), .C2(n10809), .A(n10808), .B(n10807), .ZN(
        n10826) );
  NAND2_X1 U13461 ( .A1(n15078), .A2(n10812), .ZN(n10813) );
  NAND2_X1 U13462 ( .A1(n10834), .A2(n10815), .ZN(n10819) );
  NAND2_X1 U13463 ( .A1(n10817), .A2(n10816), .ZN(n10818) );
  OR2_X1 U13464 ( .A1(n15103), .A2(n13367), .ZN(n10820) );
  XNOR2_X1 U13465 ( .A(n11119), .B(n10821), .ZN(n10824) );
  NAND2_X1 U13466 ( .A1(n13365), .A2(n13409), .ZN(n10822) );
  OAI21_X1 U13467 ( .B1(n10823), .B2(n13448), .A(n10822), .ZN(n10917) );
  AOI21_X1 U13468 ( .B1(n10824), .B2(n15048), .A(n10917), .ZN(n10971) );
  OR2_X1 U13469 ( .A1(n10971), .A2(n15067), .ZN(n10825) );
  OAI211_X1 U13470 ( .C1(n10972), .C2(n15063), .A(n10826), .B(n10825), .ZN(
        P2_U3256) );
  OAI21_X1 U13471 ( .B1(n10828), .B2(n10833), .A(n10827), .ZN(n15094) );
  INV_X1 U13472 ( .A(n15060), .ZN(n10829) );
  OAI211_X1 U13473 ( .C1(n15096), .C2(n10829), .A(n10845), .B(n10749), .ZN(
        n15095) );
  INV_X1 U13474 ( .A(n15095), .ZN(n10832) );
  OAI22_X1 U13475 ( .A1(n13678), .A2(n15096), .B1(n15052), .B2(n10830), .ZN(
        n10831) );
  AOI21_X1 U13476 ( .B1(n13673), .B2(n10832), .A(n10831), .ZN(n10840) );
  XNOR2_X1 U13477 ( .A(n10834), .B(n10833), .ZN(n10837) );
  INV_X1 U13478 ( .A(n10835), .ZN(n10836) );
  OAI21_X1 U13479 ( .B1(n10837), .B2(n13622), .A(n10836), .ZN(n15097) );
  INV_X1 U13480 ( .A(n15097), .ZN(n10838) );
  MUX2_X1 U13481 ( .A(n9863), .B(n10838), .S(n13643), .Z(n10839) );
  OAI211_X1 U13482 ( .C1(n15063), .C2(n15094), .A(n10840), .B(n10839), .ZN(
        P2_U3258) );
  OR2_X1 U13483 ( .A1(n10842), .A2(n10841), .ZN(n10843) );
  AND2_X1 U13484 ( .A1(n10844), .A2(n10843), .ZN(n15107) );
  NAND2_X1 U13485 ( .A1(n10845), .A2(n10850), .ZN(n10846) );
  NAND2_X1 U13486 ( .A1(n10846), .A2(n10749), .ZN(n10848) );
  OR2_X1 U13487 ( .A1(n10848), .A2(n10847), .ZN(n15102) );
  AOI22_X1 U13488 ( .A1(n15055), .A2(n10850), .B1(n10849), .B2(n13674), .ZN(
        n10851) );
  OAI21_X1 U13489 ( .B1(n15062), .B2(n15102), .A(n10851), .ZN(n10858) );
  XNOR2_X1 U13490 ( .A(n10853), .B(n10852), .ZN(n10854) );
  NAND2_X1 U13491 ( .A1(n10854), .A2(n15048), .ZN(n10856) );
  NAND2_X1 U13492 ( .A1(n10856), .A2(n10855), .ZN(n15105) );
  MUX2_X1 U13493 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n15105), .S(n13643), .Z(
        n10857) );
  AOI211_X1 U13494 ( .C1(n15107), .C2(n13609), .A(n10858), .B(n10857), .ZN(
        n10859) );
  INV_X1 U13495 ( .A(n10859), .ZN(P2_U3257) );
  NAND2_X1 U13496 ( .A1(n15055), .A2(n9974), .ZN(n10861) );
  AOI22_X1 U13497 ( .A1(n15067), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n13674), .ZN(n10860) );
  OAI211_X1 U13498 ( .C1(n15062), .C2(n10862), .A(n10861), .B(n10860), .ZN(
        n10863) );
  AOI21_X1 U13499 ( .B1(n13609), .B2(n10864), .A(n10863), .ZN(n10865) );
  OAI21_X1 U13500 ( .B1(n15067), .B2(n10866), .A(n10865), .ZN(P2_U3263) );
  INV_X1 U13501 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n15502) );
  INV_X1 U13502 ( .A(n12782), .ZN(n10867) );
  NAND2_X1 U13503 ( .A1(n10867), .A2(P3_U3897), .ZN(n10868) );
  OAI21_X1 U13504 ( .B1(P3_U3897), .B2(n15502), .A(n10868), .ZN(P3_U3519) );
  OAI21_X1 U13505 ( .B1(n10871), .B2(n10870), .A(n10869), .ZN(n11206) );
  OR2_X1 U13506 ( .A1(n11095), .A2(n11634), .ZN(n10872) );
  AND3_X1 U13507 ( .A1(n11032), .A2(n10872), .A3(n14248), .ZN(n11199) );
  XNOR2_X1 U13508 ( .A(n10873), .B(n12210), .ZN(n10874) );
  OAI222_X1 U13509 ( .A1(n14395), .A2(n12069), .B1(n10874), .B2(n14352), .C1(
        n14316), .C2(n12059), .ZN(n11203) );
  AOI211_X1 U13510 ( .C1(n14855), .C2(n11206), .A(n11199), .B(n11203), .ZN(
        n10879) );
  AOI22_X1 U13511 ( .A1(n14345), .A2(n12063), .B1(n14861), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n10875) );
  OAI21_X1 U13512 ( .B1(n10879), .B2(n14861), .A(n10875), .ZN(P1_U3536) );
  INV_X1 U13513 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10876) );
  OAI22_X1 U13514 ( .A1(n14469), .A2(n11634), .B1(n14857), .B2(n10876), .ZN(
        n10877) );
  INV_X1 U13515 ( .A(n10877), .ZN(n10878) );
  OAI21_X1 U13516 ( .B1(n10879), .B2(n9673), .A(n10878), .ZN(P1_U3483) );
  NOR2_X1 U13517 ( .A1(n10881), .A2(n10880), .ZN(n10884) );
  INV_X1 U13518 ( .A(n10882), .ZN(n10883) );
  INV_X1 U13519 ( .A(n10885), .ZN(n10886) );
  NAND2_X1 U13520 ( .A1(n14329), .A2(n10887), .ZN(n10896) );
  INV_X1 U13521 ( .A(n14323), .ZN(n14297) );
  AOI22_X1 U13522 ( .A1(n14333), .A2(n10890), .B1(n14297), .B2(n10889), .ZN(
        n10895) );
  INV_X1 U13523 ( .A(n10891), .ZN(n10892) );
  OR2_X1 U13524 ( .A1(n14300), .A2(n12034), .ZN(n10894) );
  INV_X1 U13525 ( .A(n14319), .ZN(n14320) );
  NAND2_X1 U13526 ( .A1(n14320), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10893) );
  AND4_X1 U13527 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n10897) );
  OAI21_X1 U13528 ( .B1(n14309), .B2(n10898), .A(n10897), .ZN(P1_U3290) );
  OR2_X1 U13529 ( .A1(n12016), .A2(n14071), .ZN(n12192) );
  OR2_X1 U13530 ( .A1(n14309), .A2(n12192), .ZN(n14293) );
  OAI22_X1 U13531 ( .A1(n14253), .A2(n10900), .B1(n10899), .B2(n14323), .ZN(
        n10901) );
  AOI21_X1 U13532 ( .B1(n14325), .B2(n12022), .A(n10901), .ZN(n10904) );
  MUX2_X1 U13533 ( .A(n10088), .B(n10902), .S(n14319), .Z(n10903) );
  OAI211_X1 U13534 ( .C1(n10905), .C2(n14293), .A(n10904), .B(n10903), .ZN(
        P1_U3291) );
  INV_X1 U13535 ( .A(n10906), .ZN(n10908) );
  OAI222_X1 U13536 ( .A1(n13839), .A2(n10907), .B1(n13837), .B2(n10908), .C1(
        P2_U3088), .C2(n13400), .ZN(P2_U3308) );
  OAI222_X1 U13537 ( .A1(n14486), .A2(n10909), .B1(n14494), .B2(n10908), .C1(
        P1_U3086), .C2(n14071), .ZN(P1_U3336) );
  NOR2_X1 U13538 ( .A1(n11115), .A2(n10749), .ZN(n10911) );
  XNOR2_X1 U13539 ( .A(n11120), .B(n13186), .ZN(n10910) );
  NOR2_X1 U13540 ( .A1(n10910), .A2(n10911), .ZN(n10937) );
  AOI21_X1 U13541 ( .B1(n10911), .B2(n10910), .A(n10937), .ZN(n10916) );
  INV_X1 U13542 ( .A(n10912), .ZN(n10913) );
  NAND2_X1 U13543 ( .A1(n10914), .A2(n10913), .ZN(n10915) );
  OAI21_X1 U13544 ( .B1(n10916), .B2(n10915), .A(n6898), .ZN(n10923) );
  NOR2_X1 U13545 ( .A1(n13354), .A2(n11120), .ZN(n10922) );
  NAND2_X1 U13546 ( .A1(n13334), .A2(n10917), .ZN(n10919) );
  OAI211_X1 U13547 ( .C1(n13336), .C2(n10920), .A(n10919), .B(n10918), .ZN(
        n10921) );
  AOI211_X1 U13548 ( .C1(n10923), .C2(n13343), .A(n10922), .B(n10921), .ZN(
        n10924) );
  INV_X1 U13549 ( .A(n10924), .ZN(P2_U3203) );
  OAI22_X1 U13550 ( .A1(n15067), .A2(n10926), .B1(n13376), .B2(n15052), .ZN(
        n10929) );
  OAI22_X1 U13551 ( .A1(n13678), .A2(n9925), .B1(n10927), .B2(n15062), .ZN(
        n10928) );
  AOI211_X1 U13552 ( .C1(n15067), .C2(P2_REG2_REG_1__SCAN_IN), .A(n10929), .B(
        n10928), .ZN(n10930) );
  OAI21_X1 U13553 ( .B1(n15063), .B2(n10931), .A(n10930), .ZN(P2_U3264) );
  INV_X1 U13554 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15684) );
  INV_X1 U13555 ( .A(n11845), .ZN(n10933) );
  NAND2_X1 U13556 ( .A1(n10933), .A2(n10932), .ZN(n10934) );
  OAI21_X1 U13557 ( .B1(P3_U3897), .B2(n15684), .A(n10934), .ZN(P3_U3521) );
  INV_X1 U13558 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n15491) );
  INV_X1 U13559 ( .A(n12767), .ZN(n10935) );
  NAND2_X1 U13560 ( .A1(n10935), .A2(n10958), .ZN(n10936) );
  OAI21_X1 U13561 ( .B1(P3_U3897), .B2(n15491), .A(n10936), .ZN(P3_U3520) );
  INV_X1 U13562 ( .A(n10937), .ZN(n10938) );
  NAND2_X1 U13563 ( .A1(n13365), .A2(n13651), .ZN(n11138) );
  XNOR2_X1 U13564 ( .A(n11283), .B(n13226), .ZN(n11137) );
  XOR2_X1 U13565 ( .A(n11138), .B(n11137), .Z(n11139) );
  XNOR2_X1 U13566 ( .A(n11140), .B(n11139), .ZN(n10945) );
  NOR2_X1 U13567 ( .A1(n11279), .A2(n13312), .ZN(n10941) );
  NOR2_X1 U13568 ( .A1(n11115), .A2(n13448), .ZN(n10940) );
  OR2_X1 U13569 ( .A1(n10941), .A2(n10940), .ZN(n11124) );
  NAND2_X1 U13570 ( .A1(n13334), .A2(n11124), .ZN(n10942) );
  NAND2_X1 U13571 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14968)
         );
  OAI211_X1 U13572 ( .C1(n13336), .C2(n11130), .A(n10942), .B(n14968), .ZN(
        n10943) );
  AOI21_X1 U13573 ( .B1(n11283), .B2(n9967), .A(n10943), .ZN(n10944) );
  OAI21_X1 U13574 ( .B1(n10945), .B2(n13339), .A(n10944), .ZN(P2_U3189) );
  NAND2_X1 U13575 ( .A1(n10946), .A2(n13123), .ZN(n10947) );
  OAI211_X1 U13576 ( .C1(n15478), .C2(n13130), .A(n10947), .B(n12007), .ZN(
        P3_U3272) );
  INV_X1 U13577 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n10960) );
  INV_X1 U13578 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U13579 ( .A1(n10948), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10952) );
  INV_X1 U13580 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n10949) );
  OR2_X1 U13581 ( .A1(n10950), .A2(n10949), .ZN(n10951) );
  OAI211_X1 U13582 ( .C1(n10954), .C2(n10953), .A(n10952), .B(n10951), .ZN(
        n10955) );
  INV_X1 U13583 ( .A(n10955), .ZN(n10956) );
  NAND2_X1 U13584 ( .A1(n12752), .A2(n10958), .ZN(n10959) );
  OAI21_X1 U13585 ( .B1(P3_U3897), .B2(n10960), .A(n10959), .ZN(P3_U3522) );
  MUX2_X1 U13586 ( .A(n10961), .B(P2_REG2_REG_3__SCAN_IN), .S(n15067), .Z(
        n10967) );
  NAND2_X1 U13587 ( .A1(n13673), .A2(n10962), .ZN(n10965) );
  NAND2_X1 U13588 ( .A1(n15055), .A2(n10963), .ZN(n10964) );
  OAI211_X1 U13589 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n15052), .A(n10965), .B(
        n10964), .ZN(n10966) );
  AOI211_X1 U13590 ( .C1(n13609), .C2(n10968), .A(n10967), .B(n10966), .ZN(
        n10969) );
  INV_X1 U13591 ( .A(n10969), .ZN(P2_U3262) );
  OAI211_X1 U13592 ( .C1(n10972), .C2(n13759), .A(n10971), .B(n10970), .ZN(
        n10977) );
  OAI22_X1 U13593 ( .A1(n13758), .A2(n11120), .B1(n15129), .B2(n9997), .ZN(
        n10973) );
  AOI21_X1 U13594 ( .B1(n10977), .B2(n15129), .A(n10973), .ZN(n10974) );
  INV_X1 U13595 ( .A(n10974), .ZN(P2_U3508) );
  INV_X1 U13596 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10975) );
  OAI22_X1 U13597 ( .A1(n13809), .A2(n11120), .B1(n15119), .B2(n10975), .ZN(
        n10976) );
  AOI21_X1 U13598 ( .B1(n10977), .B2(n15119), .A(n10976), .ZN(n10978) );
  INV_X1 U13599 ( .A(n10978), .ZN(P2_U3457) );
  MUX2_X1 U13600 ( .A(n10979), .B(P1_REG2_REG_4__SCAN_IN), .S(n14309), .Z(
        n10984) );
  NAND2_X1 U13601 ( .A1(n14319), .A2(n14071), .ZN(n11215) );
  INV_X1 U13602 ( .A(n11215), .ZN(n10981) );
  AOI22_X1 U13603 ( .A1(n10981), .A2(n10980), .B1(n7408), .B2(n14297), .ZN(
        n10982) );
  OAI21_X1 U13604 ( .B1(n12038), .B2(n14300), .A(n10982), .ZN(n10983) );
  AOI211_X1 U13605 ( .C1(n14329), .C2(n10985), .A(n10984), .B(n10983), .ZN(
        n10986) );
  INV_X1 U13606 ( .A(n10986), .ZN(P1_U3289) );
  XNOR2_X1 U13607 ( .A(n11158), .B(n12435), .ZN(n11104) );
  XNOR2_X1 U13608 ( .A(n11104), .B(n11317), .ZN(n10994) );
  INV_X1 U13609 ( .A(n10987), .ZN(n10988) );
  OR2_X1 U13610 ( .A1(n15314), .A2(n10988), .ZN(n10989) );
  INV_X1 U13611 ( .A(n11106), .ZN(n10992) );
  AOI21_X1 U13612 ( .B1(n10994), .B2(n10993), .A(n10992), .ZN(n11000) );
  INV_X1 U13613 ( .A(n10995), .ZN(n11159) );
  OAI22_X1 U13614 ( .A1(n15154), .A2(n10996), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15750), .ZN(n10998) );
  OAI22_X1 U13615 ( .A1(n12578), .A2(n11303), .B1(n15314), .B2(n12617), .ZN(
        n10997) );
  AOI211_X1 U13616 ( .C1(n11159), .C2(n12619), .A(n10998), .B(n10997), .ZN(
        n10999) );
  OAI21_X1 U13617 ( .B1(n11000), .B2(n15146), .A(n10999), .ZN(P3_U3170) );
  INV_X1 U13618 ( .A(n14293), .ZN(n11101) );
  NAND2_X1 U13619 ( .A1(n14333), .A2(n14248), .ZN(n11513) );
  OAI22_X1 U13620 ( .A1(n11513), .A2(n11002), .B1(n14300), .B2(n11001), .ZN(
        n11005) );
  NOR2_X1 U13621 ( .A1(n14309), .A2(n14395), .ZN(n14270) );
  INV_X1 U13622 ( .A(n14270), .ZN(n11164) );
  OAI22_X1 U13623 ( .A1(n11164), .A2(n12021), .B1(n11003), .B2(n14323), .ZN(
        n11004) );
  AOI211_X1 U13624 ( .C1(n11101), .C2(n11006), .A(n11005), .B(n11004), .ZN(
        n11009) );
  MUX2_X1 U13625 ( .A(n11007), .B(n10076), .S(n14320), .Z(n11008) );
  NAND2_X1 U13626 ( .A1(n11009), .A2(n11008), .ZN(P1_U3292) );
  OAI21_X1 U13627 ( .B1(n11011), .B2(n11977), .A(n11010), .ZN(n15350) );
  INV_X1 U13628 ( .A(n15350), .ZN(n11023) );
  NAND2_X1 U13629 ( .A1(n11855), .A2(n11973), .ZN(n15281) );
  NOR2_X1 U13630 ( .A1(n15337), .A2(n15281), .ZN(n15333) );
  INV_X1 U13631 ( .A(n15333), .ZN(n12840) );
  INV_X1 U13632 ( .A(n15289), .ZN(n15326) );
  OAI22_X1 U13633 ( .A1(n11012), .A2(n15313), .B1(n11317), .B2(n15315), .ZN(
        n11017) );
  INV_X1 U13634 ( .A(n11013), .ZN(n11014) );
  AOI211_X1 U13635 ( .C1(n11977), .C2(n11015), .A(n15311), .B(n11014), .ZN(
        n11016) );
  AOI211_X1 U13636 ( .C1(n15326), .C2(n15350), .A(n11017), .B(n11016), .ZN(
        n15347) );
  INV_X2 U13637 ( .A(n15337), .ZN(n15335) );
  MUX2_X1 U13638 ( .A(n11018), .B(n15347), .S(n15335), .Z(n11022) );
  NOR2_X1 U13639 ( .A1(n11019), .A2(n15339), .ZN(n15349) );
  AOI22_X1 U13640 ( .A1(n15295), .A2(n15349), .B1(n15332), .B2(n11020), .ZN(
        n11021) );
  OAI211_X1 U13641 ( .C1(n11023), .C2(n12840), .A(n11022), .B(n11021), .ZN(
        P3_U3230) );
  OAI21_X1 U13642 ( .B1(n11025), .B2(n7398), .A(n11024), .ZN(n11222) );
  INV_X1 U13643 ( .A(n11222), .ZN(n11038) );
  INV_X1 U13644 ( .A(n11026), .ZN(n11027) );
  AOI21_X1 U13645 ( .B1(n7398), .B2(n11028), .A(n11027), .ZN(n11031) );
  NAND2_X1 U13646 ( .A1(n11222), .A2(n11421), .ZN(n11030) );
  AOI22_X1 U13647 ( .A1(n14239), .A2(n14032), .B1(n14034), .B2(n14238), .ZN(
        n11029) );
  OAI211_X1 U13648 ( .C1(n11031), .C2(n14352), .A(n11030), .B(n11029), .ZN(
        n11220) );
  NAND2_X1 U13649 ( .A1(n11220), .A2(n14319), .ZN(n11037) );
  AOI211_X1 U13650 ( .C1(n12070), .C2(n11032), .A(n14423), .B(n7121), .ZN(
        n11221) );
  INV_X1 U13651 ( .A(n11033), .ZN(n11756) );
  AOI22_X1 U13652 ( .A1(n14320), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11756), 
        .B2(n14297), .ZN(n11034) );
  OAI21_X1 U13653 ( .B1(n12068), .B2(n14300), .A(n11034), .ZN(n11035) );
  AOI21_X1 U13654 ( .B1(n11221), .B2(n14333), .A(n11035), .ZN(n11036) );
  OAI211_X1 U13655 ( .C1(n11038), .C2(n14293), .A(n11037), .B(n11036), .ZN(
        P1_U3284) );
  XNOR2_X1 U13656 ( .A(n11039), .B(n12205), .ZN(n11044) );
  OAI21_X1 U13657 ( .B1(n11041), .B2(n12205), .A(n11040), .ZN(n14840) );
  OAI22_X1 U13658 ( .A1(n11405), .A2(n14395), .B1(n12039), .B2(n14316), .ZN(
        n11042) );
  AOI21_X1 U13659 ( .B1(n14840), .B2(n11421), .A(n11042), .ZN(n11043) );
  OAI21_X1 U13660 ( .B1(n14352), .B2(n11044), .A(n11043), .ZN(n14838) );
  INV_X1 U13661 ( .A(n14838), .ZN(n11052) );
  AOI21_X1 U13662 ( .B1(n11045), .B2(n12047), .A(n14423), .ZN(n11047) );
  NAND2_X1 U13663 ( .A1(n11047), .A2(n11046), .ZN(n14836) );
  NAND2_X1 U13664 ( .A1(n14325), .A2(n12047), .ZN(n11049) );
  AOI22_X1 U13665 ( .A1(n14309), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n11253), 
        .B2(n14297), .ZN(n11048) );
  OAI211_X1 U13666 ( .C1(n14253), .C2(n14836), .A(n11049), .B(n11048), .ZN(
        n11050) );
  AOI21_X1 U13667 ( .B1(n11101), .B2(n14840), .A(n11050), .ZN(n11051) );
  OAI21_X1 U13668 ( .B1(n11052), .B2(n14309), .A(n11051), .ZN(P1_U3288) );
  MUX2_X1 U13669 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12735), .Z(n12641) );
  XOR2_X1 U13670 ( .A(n11083), .B(n12641), .Z(n12642) );
  INV_X1 U13671 ( .A(n11053), .ZN(n11055) );
  NAND2_X1 U13672 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  MUX2_X1 U13673 ( .A(n11500), .B(n11058), .S(n12735), .Z(n11060) );
  INV_X1 U13674 ( .A(n11060), .ZN(n11059) );
  NAND2_X1 U13675 ( .A1(n11059), .A2(n7217), .ZN(n15174) );
  AND2_X1 U13676 ( .A1(n11060), .A2(n15180), .ZN(n15175) );
  XOR2_X1 U13677 ( .A(n12642), .B(n12643), .Z(n11085) );
  NOR2_X1 U13678 ( .A1(n15180), .A2(n11063), .ZN(n11064) );
  NAND2_X1 U13679 ( .A1(n12640), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n12658) );
  NAND2_X1 U13680 ( .A1(n11083), .A2(n11707), .ZN(n11065) );
  NAND2_X1 U13681 ( .A1(n12658), .A2(n11065), .ZN(n11067) );
  INV_X1 U13682 ( .A(n12659), .ZN(n11066) );
  AOI21_X1 U13683 ( .B1(n11068), .B2(n11067), .A(n11066), .ZN(n11071) );
  NAND2_X1 U13684 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n15151)
         );
  INV_X1 U13685 ( .A(n15151), .ZN(n11069) );
  AOI21_X1 U13686 ( .B1(n15232), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11069), 
        .ZN(n11070) );
  OAI21_X1 U13687 ( .B1(n15266), .B2(n11071), .A(n11070), .ZN(n11082) );
  NOR2_X1 U13688 ( .A1(n15180), .A2(n11074), .ZN(n11075) );
  NAND2_X1 U13689 ( .A1(n12640), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12624) );
  NAND2_X1 U13690 ( .A1(n11083), .A2(n11076), .ZN(n11077) );
  NAND2_X1 U13691 ( .A1(n12624), .A2(n11077), .ZN(n11078) );
  NAND2_X1 U13692 ( .A1(n11079), .A2(n11078), .ZN(n11080) );
  AOI21_X1 U13693 ( .B1(n12625), .B2(n11080), .A(n15241), .ZN(n11081) );
  AOI211_X1 U13694 ( .C1(n15259), .C2(n11083), .A(n11082), .B(n11081), .ZN(
        n11084) );
  OAI21_X1 U13695 ( .B1(n11085), .B2(n15253), .A(n11084), .ZN(P3_U3192) );
  XNOR2_X1 U13696 ( .A(n11086), .B(n11087), .ZN(n11093) );
  OR2_X1 U13697 ( .A1(n11088), .A2(n11087), .ZN(n11089) );
  NAND2_X1 U13698 ( .A1(n11090), .A2(n11089), .ZN(n14843) );
  NAND2_X1 U13699 ( .A1(n14843), .A2(n11421), .ZN(n11092) );
  AOI22_X1 U13700 ( .A1(n14239), .A2(n14034), .B1(n14036), .B2(n14238), .ZN(
        n11091) );
  OAI211_X1 U13701 ( .C1(n14352), .C2(n11093), .A(n11092), .B(n11091), .ZN(
        n14848) );
  INV_X1 U13702 ( .A(n14848), .ZN(n11103) );
  OAI21_X1 U13703 ( .B1(n11094), .B2(n14846), .A(n14248), .ZN(n11096) );
  OR2_X1 U13704 ( .A1(n11096), .A2(n11095), .ZN(n14844) );
  NAND2_X1 U13705 ( .A1(n14325), .A2(n12060), .ZN(n11099) );
  INV_X1 U13706 ( .A(n11097), .ZN(n11448) );
  AOI22_X1 U13707 ( .A1(n14320), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n11448), 
        .B2(n14297), .ZN(n11098) );
  OAI211_X1 U13708 ( .C1(n14253), .C2(n14844), .A(n11099), .B(n11098), .ZN(
        n11100) );
  AOI21_X1 U13709 ( .B1(n14843), .B2(n11101), .A(n11100), .ZN(n11102) );
  OAI21_X1 U13710 ( .B1(n11103), .B2(n14309), .A(n11102), .ZN(P1_U3286) );
  NAND2_X1 U13711 ( .A1(n11317), .A2(n11104), .ZN(n11105) );
  XNOR2_X1 U13712 ( .A(n11311), .B(n12484), .ZN(n11295) );
  XNOR2_X1 U13713 ( .A(n11295), .B(n11303), .ZN(n11293) );
  XNOR2_X1 U13714 ( .A(n11294), .B(n11293), .ZN(n11111) );
  OAI22_X1 U13715 ( .A1(n12578), .A2(n15130), .B1(n11317), .B2(n12617), .ZN(
        n11107) );
  INV_X1 U13716 ( .A(n11107), .ZN(n11109) );
  AOI22_X1 U13717 ( .A1(n15140), .A2(n11311), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11108) );
  OAI211_X1 U13718 ( .C1(n11312), .C2(n15159), .A(n11109), .B(n11108), .ZN(
        n11110) );
  AOI21_X1 U13719 ( .B1(n11111), .B2(n15134), .A(n11110), .ZN(n11112) );
  INV_X1 U13720 ( .A(n11112), .ZN(P3_U3167) );
  OR2_X1 U13721 ( .A1(n11116), .A2(n11121), .ZN(n11117) );
  NAND2_X1 U13722 ( .A1(n11285), .A2(n11117), .ZN(n11128) );
  OR2_X1 U13723 ( .A1(n11128), .A2(n6873), .ZN(n11127) );
  NOR2_X1 U13724 ( .A1(n11120), .A2(n13366), .ZN(n11118) );
  NAND2_X1 U13725 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  NAND2_X1 U13726 ( .A1(n11277), .A2(n11123), .ZN(n11125) );
  AOI21_X1 U13727 ( .B1(n11125), .B2(n7325), .A(n11124), .ZN(n11126) );
  AND2_X1 U13728 ( .A1(n11127), .A2(n11126), .ZN(n15116) );
  INV_X1 U13729 ( .A(n11128), .ZN(n15114) );
  INV_X1 U13730 ( .A(n11340), .ZN(n11135) );
  INV_X1 U13731 ( .A(n11283), .ZN(n15112) );
  OAI211_X1 U13732 ( .C1(n11129), .C2(n15112), .A(n10749), .B(n11333), .ZN(
        n15110) );
  OAI22_X1 U13733 ( .A1(n13643), .A2(n11131), .B1(n11130), .B2(n15052), .ZN(
        n11132) );
  AOI21_X1 U13734 ( .B1(n15055), .B2(n11283), .A(n11132), .ZN(n11133) );
  OAI21_X1 U13735 ( .B1(n15062), .B2(n15110), .A(n11133), .ZN(n11134) );
  AOI21_X1 U13736 ( .B1(n15114), .B2(n11135), .A(n11134), .ZN(n11136) );
  OAI21_X1 U13737 ( .B1(n15116), .B2(n15067), .A(n11136), .ZN(P2_U3255) );
  XNOR2_X1 U13738 ( .A(n11486), .B(n13226), .ZN(n11142) );
  NAND2_X1 U13739 ( .A1(n13364), .A2(n13191), .ZN(n11141) );
  NOR2_X1 U13740 ( .A1(n11142), .A2(n11141), .ZN(n11346) );
  NOR2_X1 U13741 ( .A1(n11346), .A2(n6832), .ZN(n11143) );
  XNOR2_X1 U13742 ( .A(n11347), .B(n11143), .ZN(n11148) );
  INV_X1 U13743 ( .A(n13363), .ZN(n11381) );
  OAI22_X1 U13744 ( .A1(n11275), .A2(n13448), .B1(n11381), .B2(n13312), .ZN(
        n11329) );
  NAND2_X1 U13745 ( .A1(n13334), .A2(n11329), .ZN(n11145) );
  OAI211_X1 U13746 ( .C1(n13336), .C2(n11334), .A(n11145), .B(n11144), .ZN(
        n11146) );
  AOI21_X1 U13747 ( .B1(n11489), .B2(n9967), .A(n11146), .ZN(n11147) );
  OAI21_X1 U13748 ( .B1(n11148), .B2(n13339), .A(n11147), .ZN(P2_U3208) );
  XNOR2_X1 U13749 ( .A(n11149), .B(n11976), .ZN(n15353) );
  INV_X1 U13750 ( .A(n15353), .ZN(n11162) );
  NAND2_X1 U13751 ( .A1(n15353), .A2(n15326), .ZN(n11156) );
  OAI22_X1 U13752 ( .A1(n11303), .A2(n15315), .B1(n15314), .B2(n15313), .ZN(
        n11150) );
  INV_X1 U13753 ( .A(n11150), .ZN(n11155) );
  OAI211_X1 U13754 ( .C1(n11153), .C2(n11152), .A(n11151), .B(n15322), .ZN(
        n11154) );
  AND3_X1 U13755 ( .A1(n11156), .A2(n11155), .A3(n11154), .ZN(n15355) );
  MUX2_X1 U13756 ( .A(n11157), .B(n15355), .S(n15335), .Z(n11161) );
  AND2_X1 U13757 ( .A1(n11158), .A2(n15328), .ZN(n15352) );
  AOI22_X1 U13758 ( .A1(n15295), .A2(n15352), .B1(n15332), .B2(n11159), .ZN(
        n11160) );
  OAI211_X1 U13759 ( .C1(n11162), .C2(n12840), .A(n11161), .B(n11160), .ZN(
        P3_U3229) );
  AOI22_X1 U13760 ( .A1(n14320), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14297), .ZN(n11163) );
  OAI21_X1 U13761 ( .B1(n11164), .B2(n7904), .A(n11163), .ZN(n11167) );
  NAND2_X1 U13762 ( .A1(n14319), .A2(n14688), .ZN(n14220) );
  AOI21_X1 U13763 ( .B1(n14313), .B2(n14220), .A(n12203), .ZN(n11166) );
  AOI21_X1 U13764 ( .B1(n11513), .B2(n14300), .A(n12017), .ZN(n11165) );
  OR3_X1 U13765 ( .A1(n11167), .A2(n11166), .A3(n11165), .ZN(P1_U3293) );
  INV_X1 U13766 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11425) );
  XNOR2_X1 U13767 ( .A(n14058), .B(n11425), .ZN(n11170) );
  XNOR2_X1 U13768 ( .A(n11176), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n14738) );
  OAI21_X1 U13769 ( .B1(n11170), .B2(n11169), .A(n14045), .ZN(n11171) );
  INV_X1 U13770 ( .A(n14789), .ZN(n14824) );
  NAND2_X1 U13771 ( .A1(n11171), .A2(n14824), .ZN(n11184) );
  INV_X1 U13772 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11172) );
  MUX2_X1 U13773 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n11172), .S(n14058), .Z(
        n11178) );
  INV_X1 U13774 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11175) );
  MUX2_X1 U13775 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11175), .S(n11176), .Z(
        n14734) );
  OAI21_X1 U13776 ( .B1(n11176), .B2(P1_REG1_REG_11__SCAN_IN), .A(n14733), 
        .ZN(n11177) );
  OAI21_X1 U13777 ( .B1(n11178), .B2(n11177), .A(n14057), .ZN(n11182) );
  NAND2_X1 U13778 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13896)
         );
  NAND2_X1 U13779 ( .A1(n14729), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11179) );
  OAI211_X1 U13780 ( .C1(n14828), .C2(n11180), .A(n13896), .B(n11179), .ZN(
        n11181) );
  AOI21_X1 U13781 ( .B1(n11182), .B2(n14819), .A(n11181), .ZN(n11183) );
  NAND2_X1 U13782 ( .A1(n11184), .A2(n11183), .ZN(P1_U3255) );
  XNOR2_X1 U13783 ( .A(n11190), .B(n11185), .ZN(n11186) );
  NAND2_X1 U13784 ( .A1(n11186), .A2(n14688), .ZN(n11188) );
  AOI22_X1 U13785 ( .A1(n14239), .A2(n14029), .B1(n14032), .B2(n14238), .ZN(
        n11187) );
  NAND2_X1 U13786 ( .A1(n11188), .A2(n11187), .ZN(n14695) );
  INV_X1 U13787 ( .A(n14695), .ZN(n11198) );
  OAI21_X1 U13788 ( .B1(n11191), .B2(n11190), .A(n11189), .ZN(n14697) );
  OAI211_X1 U13789 ( .C1(n14694), .C2(n11192), .A(n6717), .B(n14248), .ZN(
        n14693) );
  INV_X1 U13790 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11193) );
  OAI22_X1 U13791 ( .A1(n14319), .A2(n11193), .B1(n11792), .B2(n14323), .ZN(
        n11194) );
  AOI21_X1 U13792 ( .B1(n14325), .B2(n12080), .A(n11194), .ZN(n11195) );
  OAI21_X1 U13793 ( .B1(n14693), .B2(n14253), .A(n11195), .ZN(n11196) );
  AOI21_X1 U13794 ( .B1(n14697), .B2(n14329), .A(n11196), .ZN(n11197) );
  OAI21_X1 U13795 ( .B1(n14309), .B2(n11198), .A(n11197), .ZN(P1_U3282) );
  INV_X1 U13796 ( .A(n11199), .ZN(n11202) );
  INV_X1 U13797 ( .A(n11200), .ZN(n11631) );
  AOI22_X1 U13798 ( .A1(n14325), .A2(n12063), .B1(n14297), .B2(n11631), .ZN(
        n11201) );
  OAI21_X1 U13799 ( .B1(n11215), .B2(n11202), .A(n11201), .ZN(n11205) );
  MUX2_X1 U13800 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11203), .S(n14319), .Z(
        n11204) );
  AOI211_X1 U13801 ( .C1(n14329), .C2(n11206), .A(n11205), .B(n11204), .ZN(
        n11207) );
  INV_X1 U13802 ( .A(n11207), .ZN(P1_U3285) );
  AOI21_X1 U13803 ( .B1(n11208), .B2(n12213), .A(n14352), .ZN(n11210) );
  AOI22_X1 U13804 ( .A1(n11210), .A2(n11209), .B1(n14238), .B2(n14033), .ZN(
        n14851) );
  OAI21_X1 U13805 ( .B1(n11212), .B2(n12213), .A(n11211), .ZN(n14854) );
  NAND2_X1 U13806 ( .A1(n14854), .A2(n14329), .ZN(n11219) );
  OAI22_X1 U13807 ( .A1(n14319), .A2(n10727), .B1(n11771), .B2(n14323), .ZN(
        n11217) );
  XNOR2_X1 U13808 ( .A(n11213), .B(n7126), .ZN(n11214) );
  AOI22_X1 U13809 ( .A1(n11214), .A2(n14248), .B1(n14239), .B2(n14031), .ZN(
        n14850) );
  NOR2_X1 U13810 ( .A1(n14850), .A2(n11215), .ZN(n11216) );
  AOI211_X1 U13811 ( .C1(n14325), .C2(n12073), .A(n11217), .B(n11216), .ZN(
        n11218) );
  OAI211_X1 U13812 ( .C1(n14309), .C2(n14851), .A(n11219), .B(n11218), .ZN(
        P1_U3283) );
  AOI211_X1 U13813 ( .C1(n14842), .C2(n11222), .A(n11221), .B(n11220), .ZN(
        n11227) );
  INV_X1 U13814 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11223) );
  OAI22_X1 U13815 ( .A1(n14469), .A2(n12068), .B1(n14857), .B2(n11223), .ZN(
        n11224) );
  INV_X1 U13816 ( .A(n11224), .ZN(n11225) );
  OAI21_X1 U13817 ( .B1(n11227), .B2(n9673), .A(n11225), .ZN(P1_U3486) );
  AOI22_X1 U13818 ( .A1(n14345), .A2(n12070), .B1(n14861), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11226) );
  OAI21_X1 U13819 ( .B1(n11227), .B2(n14861), .A(n11226), .ZN(P1_U3537) );
  NAND2_X1 U13820 ( .A1(n14320), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11230) );
  INV_X1 U13821 ( .A(n11228), .ZN(n11411) );
  NAND2_X1 U13822 ( .A1(n14297), .A2(n11411), .ZN(n11229) );
  OAI211_X1 U13823 ( .C1(n14320), .C2(n11231), .A(n11230), .B(n11229), .ZN(
        n11234) );
  NOR2_X1 U13824 ( .A1(n14253), .A2(n11232), .ZN(n11233) );
  AOI211_X1 U13825 ( .C1(n14325), .C2(n12052), .A(n11234), .B(n11233), .ZN(
        n11237) );
  INV_X1 U13826 ( .A(n14220), .ZN(n14205) );
  NAND2_X1 U13827 ( .A1(n11235), .A2(n14205), .ZN(n11236) );
  OAI211_X1 U13828 ( .C1(n11238), .C2(n14313), .A(n11237), .B(n11236), .ZN(
        P1_U3287) );
  OAI22_X1 U13829 ( .A1(n12322), .A2(n12039), .B1(n12038), .B2(n6683), .ZN(
        n11244) );
  INV_X1 U13830 ( .A(n11244), .ZN(n11241) );
  OAI22_X1 U13831 ( .A1(n12038), .A2(n6878), .B1(n6683), .B2(n12039), .ZN(
        n11242) );
  XOR2_X1 U13832 ( .A(n12376), .B(n11242), .Z(n11260) );
  INV_X1 U13833 ( .A(n11243), .ZN(n11245) );
  AND2_X1 U13834 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  AOI22_X1 U13835 ( .A1(n12378), .A2(n14037), .B1(n6688), .B2(n12047), .ZN(
        n11248) );
  XNOR2_X1 U13836 ( .A(n11248), .B(n12376), .ZN(n11398) );
  AOI22_X1 U13837 ( .A1(n12375), .A2(n14037), .B1(n12378), .B2(n12047), .ZN(
        n11399) );
  XNOR2_X1 U13838 ( .A(n11398), .B(n11399), .ZN(n11249) );
  XNOR2_X1 U13839 ( .A(n11400), .B(n11249), .ZN(n11255) );
  INV_X1 U13840 ( .A(n12047), .ZN(n14837) );
  AOI22_X1 U13841 ( .A1(n13950), .A2(n14036), .B1(n14007), .B2(n14038), .ZN(
        n11251) );
  OAI211_X1 U13842 ( .C1(n14837), .C2(n14002), .A(n11251), .B(n11250), .ZN(
        n11252) );
  AOI21_X1 U13843 ( .B1(n11253), .B2(n13999), .A(n11252), .ZN(n11254) );
  OAI21_X1 U13844 ( .B1(n11255), .B2(n14014), .A(n11254), .ZN(P1_U3227) );
  INV_X1 U13845 ( .A(n11256), .ZN(n11269) );
  OAI222_X1 U13846 ( .A1(n14494), .A2(n11269), .B1(n12188), .B2(P1_U3086), 
        .C1(n11257), .C2(n14486), .ZN(P1_U3335) );
  AOI211_X1 U13847 ( .C1(n11260), .C2(n11259), .A(n14014), .B(n11258), .ZN(
        n11261) );
  INV_X1 U13848 ( .A(n11261), .ZN(n11266) );
  OAI21_X1 U13849 ( .B1(n13996), .B2(n11263), .A(n11262), .ZN(n11264) );
  AOI21_X1 U13850 ( .B1(n12041), .B2(n14012), .A(n11264), .ZN(n11265) );
  OAI211_X1 U13851 ( .C1(n14010), .C2(n11267), .A(n11266), .B(n11265), .ZN(
        P1_U3230) );
  INV_X1 U13852 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11270) );
  OAI222_X1 U13853 ( .A1(n13839), .A2(n11270), .B1(n13837), .B2(n11269), .C1(
        n11268), .C2(P2_U3088), .ZN(P2_U3307) );
  INV_X1 U13854 ( .A(n11271), .ZN(n11273) );
  OAI222_X1 U13855 ( .A1(P3_U3151), .A2(n11274), .B1(n11825), .B2(n11273), 
        .C1(n11272), .C2(n13130), .ZN(P3_U3271) );
  NAND2_X1 U13856 ( .A1(n11283), .A2(n11275), .ZN(n11276) );
  NAND2_X1 U13857 ( .A1(n11328), .A2(n11327), .ZN(n11326) );
  OR2_X1 U13858 ( .A1(n11486), .A2(n13364), .ZN(n11278) );
  XNOR2_X1 U13859 ( .A(n11379), .B(n11288), .ZN(n11282) );
  NOR2_X1 U13860 ( .A1(n11531), .A2(n13312), .ZN(n11281) );
  NOR2_X1 U13861 ( .A1(n11279), .A2(n13448), .ZN(n11280) );
  OR2_X1 U13862 ( .A1(n11281), .A2(n11280), .ZN(n11357) );
  AOI21_X1 U13863 ( .B1(n11282), .B2(n15048), .A(n11357), .ZN(n14672) );
  NAND2_X1 U13864 ( .A1(n11283), .A2(n13365), .ZN(n11284) );
  NAND2_X1 U13865 ( .A1(n11325), .A2(n13364), .ZN(n11286) );
  XNOR2_X1 U13866 ( .A(n11383), .B(n11288), .ZN(n14674) );
  NAND2_X1 U13867 ( .A1(n14674), .A2(n13609), .ZN(n11292) );
  OAI22_X1 U13868 ( .A1(n13643), .A2(n11651), .B1(n11360), .B2(n15052), .ZN(
        n11290) );
  OAI211_X1 U13869 ( .C1(n7228), .C2(n6718), .A(n7231), .B(n10749), .ZN(n14671) );
  NOR2_X1 U13870 ( .A1(n14671), .A2(n15062), .ZN(n11289) );
  AOI211_X1 U13871 ( .C1(n15055), .C2(n11384), .A(n11290), .B(n11289), .ZN(
        n11291) );
  OAI211_X1 U13872 ( .C1(n15067), .C2(n14672), .A(n11292), .B(n11291), .ZN(
        P2_U3253) );
  XNOR2_X1 U13873 ( .A(n15292), .B(n12435), .ZN(n11578) );
  XNOR2_X1 U13874 ( .A(n15130), .B(n11578), .ZN(n11302) );
  NAND2_X1 U13875 ( .A1(n11294), .A2(n11293), .ZN(n11298) );
  INV_X1 U13876 ( .A(n11295), .ZN(n11296) );
  NAND2_X1 U13877 ( .A1(n11303), .A2(n11296), .ZN(n11297) );
  NAND2_X1 U13878 ( .A1(n11298), .A2(n11297), .ZN(n11301) );
  INV_X1 U13879 ( .A(n11302), .ZN(n11299) );
  INV_X1 U13880 ( .A(n11580), .ZN(n11300) );
  AOI211_X1 U13881 ( .C1(n11302), .C2(n11301), .A(n15146), .B(n11300), .ZN(
        n11309) );
  OR2_X1 U13882 ( .A1(n11303), .A2(n15313), .ZN(n11305) );
  NAND2_X1 U13883 ( .A1(n12497), .A2(n12948), .ZN(n11304) );
  NAND2_X1 U13884 ( .A1(n11305), .A2(n11304), .ZN(n15285) );
  NAND2_X1 U13885 ( .A1(n15285), .A2(n15149), .ZN(n11307) );
  AOI22_X1 U13886 ( .A1(n15140), .A2(n15292), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11306) );
  OAI211_X1 U13887 ( .C1(n15293), .C2(n15159), .A(n11307), .B(n11306), .ZN(
        n11308) );
  OR2_X1 U13888 ( .A1(n11309), .A2(n11308), .ZN(P3_U3179) );
  XNOR2_X1 U13889 ( .A(n11310), .B(n8567), .ZN(n11321) );
  INV_X1 U13890 ( .A(n11321), .ZN(n15360) );
  NAND2_X1 U13891 ( .A1(n11311), .A2(n15328), .ZN(n15357) );
  OAI22_X1 U13892 ( .A1(n11375), .A2(n15357), .B1(n11312), .B2(n15307), .ZN(
        n11323) );
  NAND2_X1 U13893 ( .A1(n11313), .A2(n11870), .ZN(n11314) );
  NAND2_X1 U13894 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  NAND2_X1 U13895 ( .A1(n11316), .A2(n15322), .ZN(n11320) );
  OAI22_X1 U13896 ( .A1(n11317), .A2(n15313), .B1(n15130), .B2(n15315), .ZN(
        n11318) );
  INV_X1 U13897 ( .A(n11318), .ZN(n11319) );
  OAI211_X1 U13898 ( .C1(n11321), .C2(n15289), .A(n11320), .B(n11319), .ZN(
        n15358) );
  MUX2_X1 U13899 ( .A(n15358), .B(P3_REG2_REG_5__SCAN_IN), .S(n15337), .Z(
        n11322) );
  AOI211_X1 U13900 ( .C1(n15360), .C2(n15333), .A(n11323), .B(n11322), .ZN(
        n11324) );
  INV_X1 U13901 ( .A(n11324), .ZN(P3_U3228) );
  XOR2_X1 U13902 ( .A(n11327), .B(n11325), .Z(n11482) );
  OAI21_X1 U13903 ( .B1(n11328), .B2(n11327), .A(n11326), .ZN(n11330) );
  AOI21_X1 U13904 ( .B1(n11330), .B2(n15048), .A(n11329), .ZN(n11331) );
  OAI21_X1 U13905 ( .B1(n11482), .B2(n6873), .A(n11331), .ZN(n11483) );
  NAND2_X1 U13906 ( .A1(n11483), .A2(n13643), .ZN(n11339) );
  AOI211_X1 U13907 ( .C1(n11489), .C2(n11333), .A(n13191), .B(n6718), .ZN(
        n11484) );
  NOR2_X1 U13908 ( .A1(n13678), .A2(n11486), .ZN(n11337) );
  OAI22_X1 U13909 ( .A1(n13643), .A2(n11335), .B1(n11334), .B2(n15052), .ZN(
        n11336) );
  AOI211_X1 U13910 ( .C1(n11484), .C2(n13673), .A(n11337), .B(n11336), .ZN(
        n11338) );
  OAI211_X1 U13911 ( .C1(n11482), .C2(n11340), .A(n11339), .B(n11338), .ZN(
        P2_U3254) );
  INV_X1 U13912 ( .A(n11341), .ZN(n11344) );
  OAI222_X1 U13913 ( .A1(n13839), .A2(n11343), .B1(n13837), .B2(n11344), .C1(
        P2_U3088), .C2(n11342), .ZN(P2_U3306) );
  OAI222_X1 U13914 ( .A1(n14486), .A2(n11345), .B1(n14494), .B2(n11344), .C1(
        P1_U3086), .C2(n12013), .ZN(P1_U3334) );
  XNOR2_X1 U13915 ( .A(n11384), .B(n13186), .ZN(n11348) );
  NAND2_X1 U13916 ( .A1(n13363), .A2(n13191), .ZN(n11349) );
  INV_X1 U13917 ( .A(n11348), .ZN(n11351) );
  INV_X1 U13918 ( .A(n11349), .ZN(n11350) );
  AND2_X1 U13919 ( .A1(n11351), .A2(n11350), .ZN(n11352) );
  INV_X1 U13920 ( .A(n11352), .ZN(n11354) );
  AOI21_X1 U13921 ( .B1(n11355), .B2(n11354), .A(n11353), .ZN(n11356) );
  AOI21_X1 U13922 ( .B1(n11522), .B2(n6723), .A(n11356), .ZN(n11363) );
  NAND2_X1 U13923 ( .A1(n13334), .A2(n11357), .ZN(n11359) );
  OAI211_X1 U13924 ( .C1(n13336), .C2(n11360), .A(n11359), .B(n11358), .ZN(
        n11361) );
  AOI21_X1 U13925 ( .B1(n11384), .B2(n9967), .A(n11361), .ZN(n11362) );
  OAI21_X1 U13926 ( .B1(n11363), .B2(n13339), .A(n11362), .ZN(P2_U3196) );
  NAND2_X1 U13927 ( .A1(n11364), .A2(n11877), .ZN(n15269) );
  NAND2_X1 U13928 ( .A1(n15269), .A2(n15268), .ZN(n11366) );
  NAND2_X1 U13929 ( .A1(n11366), .A2(n11365), .ZN(n11367) );
  XNOR2_X1 U13930 ( .A(n11367), .B(n11979), .ZN(n15371) );
  OAI21_X1 U13931 ( .B1(n11369), .B2(n11979), .A(n11368), .ZN(n11372) );
  INV_X1 U13932 ( .A(n12496), .ZN(n12398) );
  OAI22_X1 U13933 ( .A1(n11370), .A2(n15313), .B1(n12398), .B2(n15315), .ZN(
        n11371) );
  AOI21_X1 U13934 ( .B1(n11372), .B2(n15322), .A(n11371), .ZN(n11373) );
  OAI21_X1 U13935 ( .B1(n15289), .B2(n15371), .A(n11373), .ZN(n15372) );
  NAND2_X1 U13936 ( .A1(n15372), .A2(n15335), .ZN(n11378) );
  AND2_X1 U13937 ( .A1(n12495), .A2(n15328), .ZN(n15373) );
  INV_X1 U13938 ( .A(n15373), .ZN(n11374) );
  OAI22_X1 U13939 ( .A1(n11375), .A2(n11374), .B1(n7765), .B2(n15307), .ZN(
        n11376) );
  AOI21_X1 U13940 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15337), .A(n11376), .ZN(
        n11377) );
  OAI211_X1 U13941 ( .C1(n15371), .C2(n12840), .A(n11378), .B(n11377), .ZN(
        P3_U3225) );
  NAND2_X1 U13942 ( .A1(n11384), .A2(n11381), .ZN(n11380) );
  XNOR2_X1 U13943 ( .A(n11538), .B(n11386), .ZN(n11382) );
  OAI22_X1 U13944 ( .A1(n11560), .A2(n13312), .B1(n11381), .B2(n13448), .ZN(
        n11516) );
  AOI21_X1 U13945 ( .B1(n11382), .B2(n15048), .A(n11516), .ZN(n14667) );
  OR2_X1 U13946 ( .A1(n11384), .A2(n13363), .ZN(n11385) );
  XOR2_X1 U13947 ( .A(n11386), .B(n11545), .Z(n14670) );
  NAND2_X1 U13948 ( .A1(n14670), .A2(n13609), .ZN(n11394) );
  INV_X1 U13949 ( .A(n11387), .ZN(n11518) );
  OAI22_X1 U13950 ( .A1(n13643), .A2(n11388), .B1(n11518), .B2(n15052), .ZN(
        n11392) );
  INV_X1 U13951 ( .A(n11548), .ZN(n11389) );
  OAI211_X1 U13952 ( .C1(n14668), .C2(n11390), .A(n11389), .B(n10749), .ZN(
        n14666) );
  NOR2_X1 U13953 ( .A1(n14666), .A2(n15062), .ZN(n11391) );
  AOI211_X1 U13954 ( .C1(n15055), .C2(n7230), .A(n11392), .B(n11391), .ZN(
        n11393) );
  OAI211_X1 U13955 ( .C1(n15067), .C2(n14667), .A(n11394), .B(n11393), .ZN(
        P2_U3252) );
  INV_X1 U13956 ( .A(n11432), .ZN(n11397) );
  AOI21_X1 U13957 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13829), .A(n11395), 
        .ZN(n11396) );
  OAI21_X1 U13958 ( .B1(n11397), .B2(n13837), .A(n11396), .ZN(P2_U3304) );
  NAND2_X1 U13959 ( .A1(n12052), .A2(n6688), .ZN(n11402) );
  NAND2_X1 U13960 ( .A1(n12378), .A2(n14036), .ZN(n11401) );
  NAND2_X1 U13961 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  XNOR2_X1 U13962 ( .A(n11403), .B(n12376), .ZN(n11436) );
  NAND2_X1 U13963 ( .A1(n12052), .A2(n12378), .ZN(n11404) );
  OAI21_X1 U13964 ( .B1(n12322), .B2(n11405), .A(n11404), .ZN(n11435) );
  XNOR2_X1 U13965 ( .A(n11436), .B(n11435), .ZN(n11439) );
  XNOR2_X1 U13966 ( .A(n11440), .B(n11439), .ZN(n11413) );
  INV_X1 U13967 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11406) );
  OAI22_X1 U13968 ( .A1(n14002), .A2(n11407), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11406), .ZN(n11410) );
  INV_X1 U13969 ( .A(n14007), .ZN(n13944) );
  INV_X1 U13970 ( .A(n13950), .ZN(n14005) );
  OAI22_X1 U13971 ( .A1(n11408), .A2(n13944), .B1(n14005), .B2(n12059), .ZN(
        n11409) );
  AOI211_X1 U13972 ( .C1(n11411), .C2(n13999), .A(n11410), .B(n11409), .ZN(
        n11412) );
  OAI21_X1 U13973 ( .B1(n11413), .B2(n14014), .A(n11412), .ZN(P1_U3239) );
  INV_X1 U13974 ( .A(n11414), .ZN(n11415) );
  OAI222_X1 U13975 ( .A1(n11416), .A2(P3_U3151), .B1(n13130), .B2(n15715), 
        .C1(n11825), .C2(n11415), .ZN(P3_U3270) );
  OAI21_X1 U13976 ( .B1(n11418), .B2(n12214), .A(n11417), .ZN(n11473) );
  INV_X1 U13977 ( .A(n11473), .ZN(n11430) );
  XNOR2_X1 U13978 ( .A(n11419), .B(n11420), .ZN(n11424) );
  NAND2_X1 U13979 ( .A1(n11473), .A2(n11421), .ZN(n11423) );
  AOI22_X1 U13980 ( .A1(n14239), .A2(n14028), .B1(n14031), .B2(n14238), .ZN(
        n11422) );
  OAI211_X1 U13981 ( .C1(n14352), .C2(n11424), .A(n11423), .B(n11422), .ZN(
        n11471) );
  NAND2_X1 U13982 ( .A1(n11471), .A2(n14319), .ZN(n11429) );
  AOI211_X1 U13983 ( .C1(n12246), .C2(n6717), .A(n14423), .B(n6831), .ZN(
        n11472) );
  NOR2_X1 U13984 ( .A1(n13902), .A2(n14300), .ZN(n11427) );
  OAI22_X1 U13985 ( .A1(n14319), .A2(n11425), .B1(n13895), .B2(n14323), .ZN(
        n11426) );
  AOI211_X1 U13986 ( .C1(n11472), .C2(n14333), .A(n11427), .B(n11426), .ZN(
        n11428) );
  OAI211_X1 U13987 ( .C1(n11430), .C2(n14293), .A(n11429), .B(n11428), .ZN(
        P1_U3281) );
  NAND2_X1 U13988 ( .A1(n11432), .A2(n11431), .ZN(n11433) );
  OAI211_X1 U13989 ( .C1(n11434), .C2(n14490), .A(n11433), .B(n12240), .ZN(
        P1_U3332) );
  INV_X1 U13990 ( .A(n11435), .ZN(n11438) );
  INV_X1 U13991 ( .A(n11436), .ZN(n11437) );
  OAI22_X1 U13992 ( .A1(n14846), .A2(n6878), .B1(n12059), .B2(n6683), .ZN(
        n11441) );
  XNOR2_X1 U13993 ( .A(n11441), .B(n12329), .ZN(n11614) );
  OR2_X1 U13994 ( .A1(n14846), .A2(n6683), .ZN(n11443) );
  NAND2_X1 U13995 ( .A1(n12375), .A2(n14035), .ZN(n11442) );
  NAND2_X1 U13996 ( .A1(n11443), .A2(n11442), .ZN(n11615) );
  XNOR2_X1 U13997 ( .A(n11614), .B(n11615), .ZN(n11617) );
  XNOR2_X1 U13998 ( .A(n11444), .B(n11617), .ZN(n11450) );
  AOI22_X1 U13999 ( .A1(n14007), .A2(n14036), .B1(n12060), .B2(n14012), .ZN(
        n11446) );
  OAI211_X1 U14000 ( .C1(n14005), .C2(n11754), .A(n11446), .B(n11445), .ZN(
        n11447) );
  AOI21_X1 U14001 ( .B1(n11448), .B2(n13999), .A(n11447), .ZN(n11449) );
  OAI21_X1 U14002 ( .B1(n11450), .B2(n14014), .A(n11449), .ZN(P1_U3213) );
  XNOR2_X1 U14003 ( .A(n11451), .B(n11456), .ZN(n11452) );
  AOI222_X1 U14004 ( .A1(n14029), .A2(n14238), .B1(n14027), .B2(n14239), .C1(
        n14688), .C2(n11452), .ZN(n14690) );
  INV_X1 U14005 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11453) );
  OAI22_X1 U14006 ( .A1(n14319), .A2(n11453), .B1(n13962), .B2(n14323), .ZN(
        n11455) );
  OAI211_X1 U14007 ( .C1(n6831), .C2(n7122), .A(n14248), .B(n11463), .ZN(
        n14689) );
  NOR2_X1 U14008 ( .A1(n14689), .A2(n14253), .ZN(n11454) );
  AOI211_X1 U14009 ( .C1(n14325), .C2(n13964), .A(n11455), .B(n11454), .ZN(
        n11459) );
  XNOR2_X1 U14010 ( .A(n11457), .B(n11456), .ZN(n14692) );
  NAND2_X1 U14011 ( .A1(n14692), .A2(n14329), .ZN(n11458) );
  OAI211_X1 U14012 ( .C1(n14690), .C2(n14309), .A(n11459), .B(n11458), .ZN(
        P1_U3280) );
  OAI21_X1 U14013 ( .B1(n6829), .B2(n8084), .A(n11460), .ZN(n14685) );
  OAI22_X1 U14014 ( .A1(n14315), .A2(n14395), .B1(n12256), .B2(n14316), .ZN(
        n14679) );
  INV_X1 U14015 ( .A(n13857), .ZN(n11461) );
  AOI22_X1 U14016 ( .A1(n14319), .A2(n14679), .B1(n11461), .B2(n14297), .ZN(
        n11462) );
  OAI21_X1 U14017 ( .B1(n14047), .B2(n14319), .A(n11462), .ZN(n11467) );
  AOI21_X1 U14018 ( .B1(n14681), .B2(n11463), .A(n14423), .ZN(n11465) );
  INV_X1 U14019 ( .A(n11464), .ZN(n11506) );
  NAND2_X1 U14020 ( .A1(n11465), .A2(n11506), .ZN(n14682) );
  NOR2_X1 U14021 ( .A1(n14682), .A2(n14253), .ZN(n11466) );
  AOI211_X1 U14022 ( .C1(n14325), .C2(n14681), .A(n11467), .B(n11466), .ZN(
        n11470) );
  XNOR2_X1 U14023 ( .A(n11468), .B(n8084), .ZN(n14687) );
  NAND2_X1 U14024 ( .A1(n14687), .A2(n14205), .ZN(n11469) );
  OAI211_X1 U14025 ( .C1(n14685), .C2(n14313), .A(n11470), .B(n11469), .ZN(
        P1_U3279) );
  AOI211_X1 U14026 ( .C1(n14842), .C2(n11473), .A(n11472), .B(n11471), .ZN(
        n11478) );
  INV_X1 U14027 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11474) );
  OAI22_X1 U14028 ( .A1(n13902), .A2(n14469), .B1(n14857), .B2(n11474), .ZN(
        n11475) );
  INV_X1 U14029 ( .A(n11475), .ZN(n11476) );
  OAI21_X1 U14030 ( .B1(n11478), .B2(n9673), .A(n11476), .ZN(P1_U3495) );
  AOI22_X1 U14031 ( .A1(n12246), .A2(n14345), .B1(n14861), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11477) );
  OAI21_X1 U14032 ( .B1(n11478), .B2(n14861), .A(n11477), .ZN(P1_U3540) );
  INV_X1 U14033 ( .A(n11479), .ZN(n11480) );
  OAI222_X1 U14034 ( .A1(n11481), .A2(P3_U3151), .B1(n13130), .B2(n15673), 
        .C1(n11825), .C2(n11480), .ZN(P3_U3269) );
  INV_X1 U14035 ( .A(n11482), .ZN(n11485) );
  AOI211_X1 U14036 ( .C1(n9095), .C2(n11485), .A(n11484), .B(n11483), .ZN(
        n11491) );
  OAI22_X1 U14037 ( .A1(n11486), .A2(n13809), .B1(n15119), .B2(n9274), .ZN(
        n11487) );
  INV_X1 U14038 ( .A(n11487), .ZN(n11488) );
  OAI21_X1 U14039 ( .B1(n11491), .B2(n15117), .A(n11488), .ZN(P2_U3463) );
  AOI22_X1 U14040 ( .A1(n11489), .A2(n13766), .B1(n15127), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11490) );
  OAI21_X1 U14041 ( .B1(n11491), .B2(n15127), .A(n11490), .ZN(P2_U3510) );
  NAND2_X1 U14042 ( .A1(n15269), .A2(n11492), .ZN(n11494) );
  NAND2_X1 U14043 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  XNOR2_X1 U14044 ( .A(n11495), .B(n8635), .ZN(n15376) );
  OAI211_X1 U14045 ( .C1(n11496), .C2(n8635), .A(n11602), .B(n15322), .ZN(
        n11499) );
  AOI22_X1 U14046 ( .A1(n11497), .A2(n12946), .B1(n12948), .B2(n12401), .ZN(
        n11498) );
  OAI211_X1 U14047 ( .C1(n15289), .C2(n15376), .A(n11499), .B(n11498), .ZN(
        n15377) );
  NAND2_X1 U14048 ( .A1(n15377), .A2(n15335), .ZN(n11503) );
  AND2_X1 U14049 ( .A1(n11885), .A2(n15328), .ZN(n15378) );
  OAI22_X1 U14050 ( .A1(n15335), .A2(n11500), .B1(n11591), .B2(n15307), .ZN(
        n11501) );
  AOI21_X1 U14051 ( .B1(n15295), .B2(n15378), .A(n11501), .ZN(n11502) );
  OAI211_X1 U14052 ( .C1(n15376), .C2(n12840), .A(n11503), .B(n11502), .ZN(
        P3_U3224) );
  XNOR2_X1 U14053 ( .A(n11504), .B(n12218), .ZN(n14428) );
  XNOR2_X1 U14054 ( .A(n11505), .B(n12218), .ZN(n14426) );
  NAND2_X1 U14055 ( .A1(n14421), .A2(n11506), .ZN(n11507) );
  NAND2_X1 U14056 ( .A1(n14330), .A2(n11507), .ZN(n14424) );
  OAI22_X1 U14057 ( .A1(n14304), .A2(n14395), .B1(n13959), .B2(n14316), .ZN(
        n14420) );
  INV_X1 U14058 ( .A(n14009), .ZN(n11508) );
  AOI22_X1 U14059 ( .A1(n14319), .A2(n14420), .B1(n11508), .B2(n14297), .ZN(
        n11509) );
  OAI21_X1 U14060 ( .B1(n11510), .B2(n14319), .A(n11509), .ZN(n11511) );
  AOI21_X1 U14061 ( .B1(n14421), .B2(n14325), .A(n11511), .ZN(n11512) );
  OAI21_X1 U14062 ( .B1(n14424), .B2(n11513), .A(n11512), .ZN(n11514) );
  AOI21_X1 U14063 ( .B1(n14426), .B2(n14205), .A(n11514), .ZN(n11515) );
  OAI21_X1 U14064 ( .B1(n14428), .B2(n14313), .A(n11515), .ZN(P1_U3278) );
  AOI22_X1 U14065 ( .A1(n13334), .A2(n11516), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11517) );
  OAI21_X1 U14066 ( .B1(n11518), .B2(n13336), .A(n11517), .ZN(n11524) );
  XNOR2_X1 U14067 ( .A(n14668), .B(n13186), .ZN(n11520) );
  NOR2_X1 U14068 ( .A1(n11531), .A2(n10749), .ZN(n11519) );
  NAND2_X1 U14069 ( .A1(n11520), .A2(n11519), .ZN(n11526) );
  OAI21_X1 U14070 ( .B1(n11520), .B2(n11519), .A(n11526), .ZN(n11521) );
  AOI211_X1 U14071 ( .C1(n11522), .C2(n11521), .A(n13339), .B(n11528), .ZN(
        n11523) );
  AOI211_X1 U14072 ( .C1(n7230), .C2(n9967), .A(n11524), .B(n11523), .ZN(
        n11525) );
  INV_X1 U14073 ( .A(n11525), .ZN(P2_U3206) );
  INV_X1 U14074 ( .A(n11526), .ZN(n11527) );
  XNOR2_X1 U14075 ( .A(n11553), .B(n13226), .ZN(n13131) );
  NAND2_X1 U14076 ( .A1(n13361), .A2(n13651), .ZN(n13132) );
  XNOR2_X1 U14077 ( .A(n13131), .B(n13132), .ZN(n11529) );
  OAI21_X1 U14078 ( .B1(n11530), .B2(n11529), .A(n13135), .ZN(n11535) );
  NAND2_X1 U14079 ( .A1(n11553), .A2(n9967), .ZN(n11533) );
  OAI22_X1 U14080 ( .A1(n13137), .A2(n13312), .B1(n11531), .B2(n13448), .ZN(
        n11542) );
  AOI22_X1 U14081 ( .A1(n13334), .A2(n11542), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11532) );
  OAI211_X1 U14082 ( .C1(n13336), .C2(n11551), .A(n11533), .B(n11532), .ZN(
        n11534) );
  AOI21_X1 U14083 ( .B1(n11535), .B2(n13343), .A(n11534), .ZN(n11536) );
  INV_X1 U14084 ( .A(n11536), .ZN(P2_U3187) );
  NOR2_X1 U14085 ( .A1(n14668), .A2(n13362), .ZN(n11537) );
  NAND2_X1 U14086 ( .A1(n14668), .A2(n13362), .ZN(n11539) );
  XNOR2_X1 U14087 ( .A(n11563), .B(n11558), .ZN(n11543) );
  AOI21_X1 U14088 ( .B1(n11543), .B2(n15048), .A(n11542), .ZN(n11641) );
  NAND2_X1 U14089 ( .A1(n11545), .A2(n14668), .ZN(n11544) );
  NAND2_X1 U14090 ( .A1(n11544), .A2(n13362), .ZN(n11547) );
  XNOR2_X1 U14091 ( .A(n11559), .B(n11558), .ZN(n11642) );
  INV_X1 U14092 ( .A(n11642), .ZN(n11556) );
  NOR2_X1 U14093 ( .A1(n11648), .A2(n11548), .ZN(n11549) );
  OR3_X1 U14094 ( .A1(n11568), .A2(n11549), .A3(n13651), .ZN(n11640) );
  NAND2_X1 U14095 ( .A1(n15067), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11550) );
  OAI21_X1 U14096 ( .B1(n15052), .B2(n11551), .A(n11550), .ZN(n11552) );
  AOI21_X1 U14097 ( .B1(n11553), .B2(n15055), .A(n11552), .ZN(n11554) );
  OAI21_X1 U14098 ( .B1(n11640), .B2(n15062), .A(n11554), .ZN(n11555) );
  AOI21_X1 U14099 ( .B1(n11556), .B2(n13609), .A(n11555), .ZN(n11557) );
  OAI21_X1 U14100 ( .B1(n15067), .B2(n11641), .A(n11557), .ZN(P2_U3251) );
  OR2_X1 U14101 ( .A1(n11648), .A2(n11560), .ZN(n11561) );
  XNOR2_X1 U14102 ( .A(n11689), .B(n11688), .ZN(n11716) );
  INV_X1 U14103 ( .A(n11716), .ZN(n11577) );
  AND2_X1 U14104 ( .A1(n11648), .A2(n13361), .ZN(n11562) );
  OR2_X2 U14105 ( .A1(n11563), .A2(n11562), .ZN(n11565) );
  OR2_X1 U14106 ( .A1(n11648), .A2(n13361), .ZN(n11564) );
  INV_X1 U14107 ( .A(n11688), .ZN(n11566) );
  OAI211_X1 U14108 ( .C1(n6823), .C2(n11688), .A(n15048), .B(n11701), .ZN(
        n11567) );
  AOI22_X1 U14109 ( .A1(n13359), .A2(n13409), .B1(n13331), .B2(n13361), .ZN(
        n13347) );
  NAND2_X1 U14110 ( .A1(n11567), .A2(n13347), .ZN(n11714) );
  INV_X1 U14111 ( .A(n11568), .ZN(n11570) );
  INV_X1 U14112 ( .A(n11694), .ZN(n11569) );
  AOI211_X1 U14113 ( .C1(n11571), .C2(n11570), .A(n13191), .B(n11569), .ZN(
        n11715) );
  NAND2_X1 U14114 ( .A1(n11715), .A2(n13673), .ZN(n11574) );
  INV_X1 U14115 ( .A(n11572), .ZN(n13351) );
  AOI22_X1 U14116 ( .A1(n15067), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13351), 
        .B2(n13674), .ZN(n11573) );
  OAI211_X1 U14117 ( .C1(n13355), .C2(n13678), .A(n11574), .B(n11573), .ZN(
        n11575) );
  AOI21_X1 U14118 ( .B1(n13643), .B2(n11714), .A(n11575), .ZN(n11576) );
  OAI21_X1 U14119 ( .B1(n11577), .B2(n15063), .A(n11576), .ZN(P2_U3250) );
  XNOR2_X1 U14120 ( .A(n11885), .B(n12484), .ZN(n12396) );
  XNOR2_X1 U14121 ( .A(n12396), .B(n12496), .ZN(n11590) );
  OR2_X1 U14122 ( .A1(n15130), .A2(n11578), .ZN(n11579) );
  XNOR2_X1 U14123 ( .A(n15272), .B(n12484), .ZN(n15136) );
  INV_X1 U14124 ( .A(n15136), .ZN(n11581) );
  NAND2_X1 U14125 ( .A1(n11581), .A2(n12497), .ZN(n11582) );
  XNOR2_X1 U14126 ( .A(n12495), .B(n12484), .ZN(n11583) );
  XNOR2_X1 U14127 ( .A(n15131), .B(n11583), .ZN(n12493) );
  NAND2_X1 U14128 ( .A1(n12494), .A2(n12493), .ZN(n12492) );
  INV_X1 U14129 ( .A(n11583), .ZN(n11584) );
  OR2_X1 U14130 ( .A1(n15131), .A2(n11584), .ZN(n11585) );
  NAND2_X1 U14131 ( .A1(n12492), .A2(n11585), .ZN(n11589) );
  INV_X1 U14132 ( .A(n11589), .ZN(n11587) );
  INV_X1 U14133 ( .A(n11590), .ZN(n11586) );
  INV_X1 U14134 ( .A(n12400), .ZN(n11588) );
  AOI21_X1 U14135 ( .B1(n11590), .B2(n11589), .A(n11588), .ZN(n11596) );
  NOR2_X1 U14136 ( .A1(n15159), .A2(n11591), .ZN(n11594) );
  AOI22_X1 U14137 ( .A1(n12615), .A2(n12401), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11592) );
  OAI21_X1 U14138 ( .B1(n15131), .B2(n12617), .A(n11592), .ZN(n11593) );
  AOI211_X1 U14139 ( .C1(n15140), .C2(n11885), .A(n11594), .B(n11593), .ZN(
        n11595) );
  OAI21_X1 U14140 ( .B1(n11596), .B2(n15146), .A(n11595), .ZN(P3_U3171) );
  XNOR2_X1 U14141 ( .A(n11598), .B(n11597), .ZN(n11713) );
  INV_X1 U14142 ( .A(n11599), .ZN(n11600) );
  NOR2_X1 U14143 ( .A1(n11982), .A2(n11600), .ZN(n11601) );
  AOI21_X1 U14144 ( .B1(n11602), .B2(n11601), .A(n15311), .ZN(n11605) );
  OR2_X1 U14145 ( .A1(n12583), .A2(n15315), .ZN(n11604) );
  NAND2_X1 U14146 ( .A1(n12496), .A2(n12946), .ZN(n11603) );
  NAND2_X1 U14147 ( .A1(n11604), .A2(n11603), .ZN(n15150) );
  AOI21_X1 U14148 ( .B1(n11606), .B2(n11605), .A(n15150), .ZN(n11708) );
  INV_X1 U14149 ( .A(n11708), .ZN(n11612) );
  INV_X1 U14150 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11607) );
  OAI22_X1 U14151 ( .A1(n13114), .A2(n15153), .B1(n15382), .B2(n11607), .ZN(
        n11608) );
  AOI21_X1 U14152 ( .B1(n11612), .B2(n15382), .A(n11608), .ZN(n11609) );
  OAI21_X1 U14153 ( .B1(n11713), .B2(n13105), .A(n11609), .ZN(P3_U3420) );
  NOR2_X1 U14154 ( .A1(n15394), .A2(n11610), .ZN(n13021) );
  INV_X1 U14155 ( .A(n13021), .ZN(n13019) );
  OAI22_X1 U14156 ( .A1(n13024), .A2(n15153), .B1(n15396), .B2(n11076), .ZN(
        n11611) );
  AOI21_X1 U14157 ( .B1(n11612), .B2(n15396), .A(n11611), .ZN(n11613) );
  OAI21_X1 U14158 ( .B1(n11713), .B2(n13019), .A(n11613), .ZN(P3_U3469) );
  INV_X1 U14159 ( .A(n11614), .ZN(n11616) );
  NAND2_X1 U14160 ( .A1(n12063), .A2(n6688), .ZN(n11620) );
  NAND2_X1 U14161 ( .A1(n12378), .A2(n14034), .ZN(n11619) );
  NAND2_X1 U14162 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  XNOR2_X1 U14163 ( .A(n11621), .B(n12376), .ZN(n11625) );
  NAND2_X1 U14164 ( .A1(n12063), .A2(n12378), .ZN(n11623) );
  NAND2_X1 U14165 ( .A1(n12375), .A2(n14034), .ZN(n11622) );
  NAND2_X1 U14166 ( .A1(n11623), .A2(n11622), .ZN(n11624) );
  NOR2_X1 U14167 ( .A1(n11625), .A2(n11624), .ZN(n11745) );
  AOI21_X1 U14168 ( .B1(n11625), .B2(n11624), .A(n11745), .ZN(n11626) );
  OAI21_X1 U14169 ( .B1(n6841), .B2(n11626), .A(n11746), .ZN(n11627) );
  NAND2_X1 U14170 ( .A1(n11627), .A2(n13991), .ZN(n11633) );
  AOI21_X1 U14171 ( .B1(n13950), .B2(n14033), .A(n11628), .ZN(n11629) );
  OAI21_X1 U14172 ( .B1(n13944), .B2(n12059), .A(n11629), .ZN(n11630) );
  AOI21_X1 U14173 ( .B1(n11631), .B2(n13999), .A(n11630), .ZN(n11632) );
  OAI211_X1 U14174 ( .C1(n11634), .C2(n14002), .A(n11633), .B(n11632), .ZN(
        P1_U3221) );
  INV_X1 U14175 ( .A(n11635), .ZN(n11639) );
  OAI222_X1 U14176 ( .A1(n13839), .A2(n11637), .B1(n13837), .B2(n11639), .C1(
        n11636), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U14177 ( .A(n8376), .ZN(n11638) );
  OAI222_X1 U14178 ( .A1(n14486), .A2(n7602), .B1(n14494), .B2(n11639), .C1(
        n11638), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U14179 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11671) );
  OAI211_X1 U14180 ( .C1(n11642), .C2(n13759), .A(n11641), .B(n11640), .ZN(
        n11643) );
  INV_X1 U14181 ( .A(n11643), .ZN(n11645) );
  MUX2_X1 U14182 ( .A(n11671), .B(n11645), .S(n15129), .Z(n11644) );
  OAI21_X1 U14183 ( .B1(n11648), .B2(n13758), .A(n11644), .ZN(P2_U3513) );
  INV_X1 U14184 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11646) );
  MUX2_X1 U14185 ( .A(n11646), .B(n11645), .S(n15119), .Z(n11647) );
  OAI21_X1 U14186 ( .B1(n11648), .B2(n13809), .A(n11647), .ZN(P2_U3472) );
  NAND2_X1 U14187 ( .A1(n11650), .A2(n11649), .ZN(n11653) );
  NAND2_X1 U14188 ( .A1(n11665), .A2(n11651), .ZN(n11652) );
  NAND2_X1 U14189 ( .A1(n11653), .A2(n11652), .ZN(n14976) );
  XNOR2_X1 U14190 ( .A(n11669), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n14975) );
  NAND2_X1 U14191 ( .A1(n11669), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U14192 ( .A1(n14978), .A2(n11654), .ZN(n11655) );
  NOR2_X1 U14193 ( .A1(n11655), .A2(n11673), .ZN(n11656) );
  NOR2_X1 U14194 ( .A1(n11657), .A2(n11656), .ZN(n14986) );
  AND2_X1 U14195 ( .A1(n14986), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14988) );
  NOR2_X1 U14196 ( .A1(n11657), .A2(n14988), .ZN(n11658) );
  NOR2_X1 U14197 ( .A1(n11658), .A2(n11674), .ZN(n11659) );
  INV_X1 U14198 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n15000) );
  XNOR2_X1 U14199 ( .A(n11674), .B(n11658), .ZN(n15001) );
  NOR2_X1 U14200 ( .A1(n15000), .A2(n15001), .ZN(n14999) );
  NOR2_X1 U14201 ( .A1(n11659), .A2(n14999), .ZN(n15020) );
  XNOR2_X1 U14202 ( .A(n15023), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n15019) );
  OR2_X1 U14203 ( .A1(n15020), .A2(n15019), .ZN(n15016) );
  NAND2_X1 U14204 ( .A1(n15023), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14205 ( .A1(n15016), .A2(n11660), .ZN(n15031) );
  OR2_X1 U14206 ( .A1(n11678), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11661) );
  NAND2_X1 U14207 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n11678), .ZN(n11662) );
  AND2_X1 U14208 ( .A1(n11661), .A2(n11662), .ZN(n15030) );
  NAND2_X1 U14209 ( .A1(n15031), .A2(n15030), .ZN(n15029) );
  NAND2_X1 U14210 ( .A1(n15029), .A2(n11662), .ZN(n13389) );
  XOR2_X1 U14211 ( .A(n13388), .B(n13389), .Z(n11663) );
  NAND2_X1 U14212 ( .A1(n11663), .A2(n9389), .ZN(n13391) );
  OAI21_X1 U14213 ( .B1(n9389), .B2(n11663), .A(n13391), .ZN(n11686) );
  NAND2_X1 U14214 ( .A1(n14864), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U14215 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13323)
         );
  OAI211_X1 U14216 ( .C1(n11679), .C2(n15035), .A(n11664), .B(n13323), .ZN(
        n11685) );
  INV_X1 U14217 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U14218 ( .A1(n11665), .A2(n14675), .ZN(n11666) );
  NAND2_X1 U14219 ( .A1(n11667), .A2(n11666), .ZN(n14972) );
  MUX2_X1 U14220 ( .A(n11668), .B(P2_REG1_REG_13__SCAN_IN), .S(n11669), .Z(
        n14971) );
  NAND2_X1 U14221 ( .A1(n11669), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11670) );
  NAND2_X1 U14222 ( .A1(n14974), .A2(n11670), .ZN(n14991) );
  XNOR2_X1 U14223 ( .A(n11673), .B(n11671), .ZN(n14990) );
  NAND2_X1 U14224 ( .A1(n14991), .A2(n14990), .ZN(n14989) );
  INV_X1 U14225 ( .A(n14989), .ZN(n11672) );
  AOI21_X1 U14226 ( .B1(n11673), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11672), 
        .ZN(n11675) );
  NOR2_X1 U14227 ( .A1(n11675), .A2(n11674), .ZN(n11676) );
  INV_X1 U14228 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15003) );
  XNOR2_X1 U14229 ( .A(n11675), .B(n11674), .ZN(n15004) );
  NOR2_X1 U14230 ( .A1(n15003), .A2(n15004), .ZN(n15002) );
  NOR2_X1 U14231 ( .A1(n11676), .A2(n15002), .ZN(n15015) );
  XNOR2_X1 U14232 ( .A(n15023), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15014) );
  NAND2_X1 U14233 ( .A1(n15023), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11677) );
  NAND2_X1 U14234 ( .A1(n15011), .A2(n11677), .ZN(n15034) );
  XNOR2_X1 U14235 ( .A(n11678), .B(n13756), .ZN(n15033) );
  AOI21_X1 U14236 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n11678), .A(n15037), 
        .ZN(n11680) );
  NOR2_X1 U14237 ( .A1(n11680), .A2(n11679), .ZN(n13393) );
  AOI21_X1 U14238 ( .B1(n11680), .B2(n11679), .A(n13393), .ZN(n11681) );
  INV_X1 U14239 ( .A(n11681), .ZN(n11682) );
  AND2_X1 U14240 ( .A1(n11681), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13394) );
  AOI211_X1 U14241 ( .C1(n11683), .C2(n11682), .A(n15013), .B(n13394), .ZN(
        n11684) );
  AOI211_X1 U14242 ( .C1(n15028), .C2(n11686), .A(n11685), .B(n11684), .ZN(
        n11687) );
  INV_X1 U14243 ( .A(n11687), .ZN(P2_U3232) );
  NAND2_X1 U14244 ( .A1(n13355), .A2(n13137), .ZN(n11690) );
  NAND2_X1 U14245 ( .A1(n11692), .A2(n11698), .ZN(n11693) );
  NAND2_X1 U14246 ( .A1(n13454), .A2(n11693), .ZN(n13760) );
  AOI21_X1 U14247 ( .B1(n11694), .B2(n13813), .A(n13191), .ZN(n11695) );
  AND2_X1 U14248 ( .A1(n11695), .A2(n13671), .ZN(n13761) );
  AOI22_X1 U14249 ( .A1(n15067), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13254), 
        .B2(n13674), .ZN(n11696) );
  OAI21_X1 U14250 ( .B1(n13452), .B2(n13678), .A(n11696), .ZN(n11697) );
  AOI21_X1 U14251 ( .B1(n13761), .B2(n13673), .A(n11697), .ZN(n11706) );
  NAND2_X1 U14252 ( .A1(n13355), .A2(n13360), .ZN(n11699) );
  NAND3_X1 U14253 ( .A1(n11701), .A2(n11700), .A3(n11699), .ZN(n11702) );
  NAND3_X1 U14254 ( .A1(n13666), .A2(n15048), .A3(n11702), .ZN(n11704) );
  OAI22_X1 U14255 ( .A1(n13455), .A2(n13312), .B1(n13137), .B2(n13448), .ZN(
        n13253) );
  INV_X1 U14256 ( .A(n13253), .ZN(n11703) );
  NAND2_X1 U14257 ( .A1(n11704), .A2(n11703), .ZN(n13762) );
  NAND2_X1 U14258 ( .A1(n13762), .A2(n13643), .ZN(n11705) );
  OAI211_X1 U14259 ( .C1(n13760), .C2(n15063), .A(n11706), .B(n11705), .ZN(
        P2_U3249) );
  AND2_X1 U14260 ( .A1(n15289), .A2(n15281), .ZN(n14649) );
  NOR2_X1 U14261 ( .A1(n15337), .A2(n14649), .ZN(n12893) );
  INV_X1 U14262 ( .A(n12893), .ZN(n12957) );
  OAI22_X1 U14263 ( .A1(n15335), .A2(n11707), .B1(n15160), .B2(n15307), .ZN(
        n11710) );
  NOR2_X1 U14264 ( .A1(n11708), .A2(n15337), .ZN(n11709) );
  AOI211_X1 U14265 ( .C1(n12953), .C2(n11711), .A(n11710), .B(n11709), .ZN(
        n11712) );
  OAI21_X1 U14266 ( .B1(n11713), .B2(n12957), .A(n11712), .ZN(P3_U3223) );
  AOI211_X1 U14267 ( .C1(n11716), .C2(n15099), .A(n11715), .B(n11714), .ZN(
        n11718) );
  MUX2_X1 U14268 ( .A(n15003), .B(n11718), .S(n15129), .Z(n11717) );
  OAI21_X1 U14269 ( .B1(n13355), .B2(n13758), .A(n11717), .ZN(P2_U3514) );
  INV_X1 U14270 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11719) );
  MUX2_X1 U14271 ( .A(n11719), .B(n11718), .S(n15119), .Z(n11720) );
  OAI21_X1 U14272 ( .B1(n13355), .B2(n13809), .A(n11720), .ZN(P2_U3475) );
  XNOR2_X1 U14273 ( .A(n11722), .B(n11721), .ZN(n14662) );
  INV_X1 U14274 ( .A(n14662), .ZN(n11731) );
  OAI211_X1 U14275 ( .C1(n11724), .C2(n11985), .A(n6676), .B(n15322), .ZN(
        n11726) );
  OR2_X1 U14276 ( .A1(n12583), .A2(n15313), .ZN(n11725) );
  OAI211_X1 U14277 ( .C1(n12562), .C2(n15315), .A(n11726), .B(n11725), .ZN(
        n14660) );
  NAND2_X1 U14278 ( .A1(n14660), .A2(n15335), .ZN(n11730) );
  NOR2_X1 U14279 ( .A1(n11727), .A2(n15339), .ZN(n14661) );
  INV_X1 U14280 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12664) );
  OAI22_X1 U14281 ( .A1(n15335), .A2(n12664), .B1(n12515), .B2(n15307), .ZN(
        n11728) );
  AOI21_X1 U14282 ( .B1(n15295), .B2(n14661), .A(n11728), .ZN(n11729) );
  OAI211_X1 U14283 ( .C1(n11731), .C2(n12957), .A(n11730), .B(n11729), .ZN(
        P3_U3221) );
  INV_X1 U14284 ( .A(n11984), .ZN(n11733) );
  OAI21_X1 U14285 ( .B1(n6834), .B2(n11733), .A(n11732), .ZN(n14646) );
  OAI21_X1 U14286 ( .B1(n11735), .B2(n11984), .A(n11734), .ZN(n11738) );
  OR2_X1 U14287 ( .A1(n14639), .A2(n15315), .ZN(n11737) );
  NAND2_X1 U14288 ( .A1(n12401), .A2(n12946), .ZN(n11736) );
  NAND2_X1 U14289 ( .A1(n11737), .A2(n11736), .ZN(n12586) );
  AOI21_X1 U14290 ( .B1(n11738), .B2(n15322), .A(n12586), .ZN(n14647) );
  INV_X1 U14291 ( .A(n14647), .ZN(n11739) );
  AOI21_X1 U14292 ( .B1(n15368), .B2(n14646), .A(n11739), .ZN(n11741) );
  MUX2_X1 U14293 ( .A(n8654), .B(n11741), .S(n15396), .Z(n11740) );
  OAI21_X1 U14294 ( .B1(n13024), .B2(n14651), .A(n11740), .ZN(P3_U3470) );
  INV_X1 U14295 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n11742) );
  MUX2_X1 U14296 ( .A(n11742), .B(n11741), .S(n15382), .Z(n11743) );
  OAI21_X1 U14297 ( .B1(n13114), .B2(n14651), .A(n11743), .ZN(P3_U3423) );
  OAI22_X1 U14298 ( .A1(n12068), .A2(n6878), .B1(n12069), .B2(n6683), .ZN(
        n11744) );
  XOR2_X1 U14299 ( .A(n12376), .B(n11744), .Z(n11750) );
  OR2_X1 U14300 ( .A1(n12068), .A2(n6683), .ZN(n11748) );
  NAND2_X1 U14301 ( .A1(n12375), .A2(n14033), .ZN(n11747) );
  NAND2_X1 U14302 ( .A1(n11748), .A2(n11747), .ZN(n11759) );
  OAI21_X1 U14303 ( .B1(n11750), .B2(n11749), .A(n11768), .ZN(n11751) );
  NAND2_X1 U14304 ( .A1(n11751), .A2(n13991), .ZN(n11758) );
  AOI21_X1 U14305 ( .B1(n13950), .B2(n14032), .A(n11752), .ZN(n11753) );
  OAI21_X1 U14306 ( .B1(n13944), .B2(n11754), .A(n11753), .ZN(n11755) );
  AOI21_X1 U14307 ( .B1(n11756), .B2(n13999), .A(n11755), .ZN(n11757) );
  OAI211_X1 U14308 ( .C1(n12068), .C2(n14002), .A(n11758), .B(n11757), .ZN(
        P1_U3231) );
  INV_X1 U14309 ( .A(n11759), .ZN(n11760) );
  NAND2_X1 U14310 ( .A1(n11761), .A2(n11760), .ZN(n11767) );
  AND2_X1 U14311 ( .A1(n11768), .A2(n11767), .ZN(n11770) );
  NAND2_X1 U14312 ( .A1(n12073), .A2(n6688), .ZN(n11763) );
  NAND2_X1 U14313 ( .A1(n12378), .A2(n14032), .ZN(n11762) );
  NAND2_X1 U14314 ( .A1(n11763), .A2(n11762), .ZN(n11764) );
  XNOR2_X1 U14315 ( .A(n11764), .B(n12376), .ZN(n11777) );
  NOR2_X1 U14316 ( .A1(n12322), .A2(n11765), .ZN(n11766) );
  AOI21_X1 U14317 ( .B1(n12073), .B2(n12378), .A(n11766), .ZN(n11778) );
  XNOR2_X1 U14318 ( .A(n11777), .B(n11778), .ZN(n11769) );
  OAI211_X1 U14319 ( .C1(n11770), .C2(n11769), .A(n13991), .B(n11790), .ZN(
        n11776) );
  NOR2_X1 U14320 ( .A1(n14010), .A2(n11771), .ZN(n11774) );
  NAND2_X1 U14321 ( .A1(n13950), .A2(n14031), .ZN(n11772) );
  OAI21_X1 U14322 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n8030), .A(n11772), .ZN(
        n11773) );
  AOI211_X1 U14323 ( .C1(n14007), .C2(n14033), .A(n11774), .B(n11773), .ZN(
        n11775) );
  OAI211_X1 U14324 ( .C1(n7126), .C2(n14002), .A(n11776), .B(n11775), .ZN(
        P1_U3217) );
  INV_X1 U14325 ( .A(n11777), .ZN(n11779) );
  NOR2_X1 U14326 ( .A1(n11779), .A2(n11778), .ZN(n11787) );
  INV_X1 U14327 ( .A(n11787), .ZN(n11786) );
  NAND2_X1 U14328 ( .A1(n12080), .A2(n6688), .ZN(n11781) );
  NAND2_X1 U14329 ( .A1(n12378), .A2(n14031), .ZN(n11780) );
  NAND2_X1 U14330 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  XNOR2_X1 U14331 ( .A(n11782), .B(n12329), .ZN(n12247) );
  NOR2_X1 U14332 ( .A1(n12322), .A2(n11783), .ZN(n11784) );
  AOI21_X1 U14333 ( .B1(n12080), .B2(n12378), .A(n11784), .ZN(n12248) );
  XNOR2_X1 U14334 ( .A(n12247), .B(n12248), .ZN(n11788) );
  INV_X1 U14335 ( .A(n11788), .ZN(n11785) );
  AOI21_X1 U14336 ( .B1(n11790), .B2(n11786), .A(n11785), .ZN(n11791) );
  NOR2_X1 U14337 ( .A1(n11788), .A2(n11787), .ZN(n11789) );
  OAI21_X1 U14338 ( .B1(n11791), .B2(n13892), .A(n13991), .ZN(n11796) );
  NOR2_X1 U14339 ( .A1(n14010), .A2(n11792), .ZN(n11794) );
  NAND2_X1 U14340 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14743)
         );
  OAI21_X1 U14341 ( .B1(n14005), .B2(n12244), .A(n14743), .ZN(n11793) );
  AOI211_X1 U14342 ( .C1(n14007), .C2(n14032), .A(n11794), .B(n11793), .ZN(
        n11795) );
  OAI211_X1 U14343 ( .C1(n14694), .C2(n14002), .A(n11796), .B(n11795), .ZN(
        P1_U3236) );
  AND2_X1 U14344 ( .A1(n11799), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U14345 ( .A1(n11799), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U14346 ( .A1(n11799), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U14347 ( .A1(n11799), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U14348 ( .A1(n11799), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U14349 ( .A1(n11799), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U14350 ( .A1(n11799), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U14351 ( .A1(n11799), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U14352 ( .A1(n11799), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U14353 ( .A1(n11799), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U14354 ( .A1(n11799), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U14355 ( .A1(n11799), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U14356 ( .A1(n11799), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U14357 ( .A1(n11799), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U14358 ( .A1(n11799), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U14359 ( .A1(n11799), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U14360 ( .A1(n11799), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U14361 ( .A1(n11799), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U14362 ( .A1(n11799), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U14363 ( .A1(n11799), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U14364 ( .A1(n11799), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U14365 ( .A1(n11799), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U14366 ( .A1(n11799), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U14367 ( .A1(n11799), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U14368 ( .A1(n11799), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U14369 ( .A1(n11799), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U14370 ( .A1(n11799), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U14371 ( .A1(n11799), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U14372 ( .A1(n11799), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U14373 ( .A1(n11799), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  INV_X1 U14374 ( .A(n11800), .ZN(n11801) );
  OAI222_X1 U14375 ( .A1(n12735), .A2(P3_U3151), .B1(n11825), .B2(n11801), 
        .C1(n15494), .C2(n13130), .ZN(P3_U3268) );
  INV_X1 U14376 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n11802) );
  NOR2_X1 U14377 ( .A1(n7930), .A2(n11802), .ZN(n11803) );
  INV_X1 U14378 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n11816) );
  INV_X1 U14379 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14478) );
  OR2_X1 U14380 ( .A1(n7930), .A2(n14478), .ZN(n11806) );
  INV_X1 U14381 ( .A(n14431), .ZN(n14082) );
  NAND2_X1 U14382 ( .A1(n14082), .A2(n11808), .ZN(n14081) );
  XNOR2_X1 U14383 ( .A(n14081), .B(n12194), .ZN(n11809) );
  NAND2_X1 U14384 ( .A1(n11809), .A2(n14248), .ZN(n14078) );
  INV_X1 U14385 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U14386 ( .A1(n7923), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11813) );
  NAND2_X1 U14387 ( .A1(n6687), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11812) );
  OAI211_X1 U14388 ( .C1(n6899), .C2(n11819), .A(n11813), .B(n11812), .ZN(
        n14016) );
  NAND2_X1 U14389 ( .A1(n11815), .A2(n14016), .ZN(n14338) );
  AND2_X1 U14390 ( .A1(n14078), .A2(n14338), .ZN(n11818) );
  MUX2_X1 U14391 ( .A(n11816), .B(n11818), .S(n14857), .Z(n11817) );
  OAI21_X1 U14392 ( .B1(n12194), .B2(n14469), .A(n11817), .ZN(P1_U3527) );
  MUX2_X1 U14393 ( .A(n11819), .B(n11818), .S(n14863), .Z(n11820) );
  OAI21_X1 U14394 ( .B1(n12194), .B2(n14419), .A(n11820), .ZN(P1_U3559) );
  INV_X1 U14395 ( .A(n11821), .ZN(n13836) );
  OAI222_X1 U14396 ( .A1(n14486), .A2(n11822), .B1(n14494), .B2(n13836), .C1(
        n8375), .C2(P1_U3086), .ZN(P1_U3330) );
  INV_X1 U14397 ( .A(n11823), .ZN(n11824) );
  OAI222_X1 U14398 ( .A1(P3_U3151), .A2(n8926), .B1(n13130), .B2(n15660), .C1(
        n11825), .C2(n11824), .ZN(P3_U3267) );
  INV_X1 U14399 ( .A(n11826), .ZN(n11828) );
  OAI222_X1 U14400 ( .A1(n13839), .A2(n11829), .B1(n13837), .B2(n11828), .C1(
        n11827), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U14401 ( .A(n11830), .ZN(n11831) );
  INV_X1 U14402 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13824) );
  INV_X1 U14403 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11833) );
  XNOR2_X1 U14404 ( .A(n11833), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11836) );
  XNOR2_X1 U14405 ( .A(n11837), .B(n11836), .ZN(n12394) );
  NAND2_X1 U14406 ( .A1(n12394), .A2(n11840), .ZN(n11835) );
  INV_X1 U14407 ( .A(SI_30_), .ZN(n15517) );
  OR2_X1 U14408 ( .A1(n8517), .A2(n15517), .ZN(n11834) );
  NOR2_X1 U14409 ( .A1(n13028), .A2(n11845), .ZN(n11996) );
  OAI22_X1 U14410 ( .A1(n11837), .A2(n11836), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n14478), .ZN(n11839) );
  XNOR2_X1 U14411 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11838) );
  XNOR2_X1 U14412 ( .A(n11839), .B(n11838), .ZN(n13124) );
  NAND2_X1 U14413 ( .A1(n13124), .A2(n11840), .ZN(n11842) );
  INV_X1 U14414 ( .A(SI_31_), .ZN(n13119) );
  OR2_X1 U14415 ( .A1(n8517), .A2(n13119), .ZN(n11841) );
  OR2_X1 U14416 ( .A1(n11849), .A2(n11844), .ZN(n11847) );
  NAND2_X1 U14417 ( .A1(n13028), .A2(n11845), .ZN(n11846) );
  NAND2_X1 U14418 ( .A1(n11847), .A2(n11846), .ZN(n11997) );
  INV_X1 U14419 ( .A(n13028), .ZN(n12757) );
  OAI21_X1 U14420 ( .B1(n12757), .B2(n12752), .A(n11969), .ZN(n11848) );
  INV_X1 U14421 ( .A(n11862), .ZN(n11852) );
  AOI21_X1 U14422 ( .B1(n11853), .B2(n6682), .A(n11852), .ZN(n11864) );
  OAI21_X1 U14423 ( .B1(n11856), .B2(n11855), .A(n11967), .ZN(n11859) );
  OAI21_X1 U14424 ( .B1(n11860), .B2(n11959), .A(n15301), .ZN(n11857) );
  AOI21_X1 U14425 ( .B1(n11861), .B2(n11865), .A(n11959), .ZN(n11863) );
  NAND3_X1 U14426 ( .A1(n11871), .A2(n11870), .A3(n11866), .ZN(n11868) );
  NAND3_X1 U14427 ( .A1(n11871), .A2(n11870), .A3(n11869), .ZN(n11873) );
  NAND3_X1 U14428 ( .A1(n11873), .A2(n11877), .A3(n11872), .ZN(n11875) );
  AND2_X1 U14429 ( .A1(n11875), .A2(n11874), .ZN(n11876) );
  NAND2_X1 U14430 ( .A1(n15139), .A2(n11959), .ZN(n11879) );
  NAND2_X1 U14431 ( .A1(n15276), .A2(n11967), .ZN(n11878) );
  MUX2_X1 U14432 ( .A(n11879), .B(n11878), .S(n12497), .Z(n11880) );
  MUX2_X1 U14433 ( .A(n11883), .B(n11882), .S(n11967), .Z(n11884) );
  NAND2_X1 U14434 ( .A1(n12496), .A2(n11967), .ZN(n11887) );
  NAND2_X1 U14435 ( .A1(n12398), .A2(n11959), .ZN(n11886) );
  MUX2_X1 U14436 ( .A(n11887), .B(n11886), .S(n11885), .Z(n11888) );
  AOI21_X1 U14437 ( .B1(n11889), .B2(n11888), .A(n11982), .ZN(n11893) );
  NOR2_X1 U14438 ( .A1(n12401), .A2(n15153), .ZN(n11891) );
  MUX2_X1 U14439 ( .A(n11891), .B(n7634), .S(n11967), .Z(n11892) );
  NOR3_X1 U14440 ( .A1(n11893), .A2(n11892), .A3(n11984), .ZN(n11903) );
  NAND2_X1 U14441 ( .A1(n11900), .A2(n11894), .ZN(n11897) );
  NAND2_X1 U14442 ( .A1(n11899), .A2(n11895), .ZN(n11896) );
  MUX2_X1 U14443 ( .A(n11897), .B(n11896), .S(n11967), .Z(n11902) );
  INV_X1 U14444 ( .A(n11905), .ZN(n11898) );
  NOR2_X1 U14445 ( .A1(n11904), .A2(n11898), .ZN(n14637) );
  MUX2_X1 U14446 ( .A(n11900), .B(n11899), .S(n11959), .Z(n11901) );
  OAI211_X1 U14447 ( .C1(n11903), .C2(n11902), .A(n14637), .B(n11901), .ZN(
        n11907) );
  INV_X1 U14448 ( .A(n12942), .ZN(n12944) );
  MUX2_X1 U14449 ( .A(n11905), .B(n7613), .S(n11967), .Z(n11906) );
  NAND3_X1 U14450 ( .A1(n11907), .A2(n12944), .A3(n11906), .ZN(n11911) );
  INV_X1 U14451 ( .A(n11911), .ZN(n11909) );
  OAI21_X1 U14452 ( .B1(n11909), .B2(n8993), .A(n12934), .ZN(n11917) );
  NAND3_X1 U14453 ( .A1(n11911), .A2(n11959), .A3(n11910), .ZN(n11915) );
  INV_X1 U14454 ( .A(n11920), .ZN(n11914) );
  INV_X1 U14455 ( .A(n11912), .ZN(n11913) );
  AOI211_X1 U14456 ( .C1(n11915), .C2(n12934), .A(n11914), .B(n11913), .ZN(
        n11916) );
  AOI21_X1 U14457 ( .B1(n11919), .B2(n11918), .A(n11959), .ZN(n11922) );
  MUX2_X1 U14458 ( .A(n11920), .B(n11919), .S(n11959), .Z(n11921) );
  INV_X1 U14459 ( .A(n11923), .ZN(n11926) );
  AND2_X1 U14460 ( .A1(n11924), .A2(n11959), .ZN(n11925) );
  NAND2_X1 U14461 ( .A1(n11934), .A2(n11925), .ZN(n11928) );
  AND3_X1 U14462 ( .A1(n11933), .A2(n11967), .A3(n11929), .ZN(n11932) );
  INV_X1 U14463 ( .A(n11927), .ZN(n11930) );
  AOI21_X1 U14464 ( .B1(n11930), .B2(n11929), .A(n11928), .ZN(n11931) );
  INV_X1 U14465 ( .A(n12877), .ZN(n11990) );
  MUX2_X1 U14466 ( .A(n11934), .B(n11933), .S(n11959), .Z(n11935) );
  NAND3_X1 U14467 ( .A1(n11936), .A2(n11990), .A3(n11935), .ZN(n11940) );
  MUX2_X1 U14468 ( .A(n11938), .B(n11937), .S(n11959), .Z(n11939) );
  AND2_X1 U14469 ( .A1(n11940), .A2(n11939), .ZN(n11944) );
  MUX2_X1 U14470 ( .A(n11942), .B(n11941), .S(n11967), .Z(n11943) );
  OAI21_X1 U14471 ( .B1(n11944), .B2(n12857), .A(n11943), .ZN(n11948) );
  NAND2_X1 U14472 ( .A1(n11945), .A2(n11946), .ZN(n12845) );
  NOR2_X1 U14473 ( .A1(n12846), .A2(n11967), .ZN(n11949) );
  AOI21_X1 U14474 ( .B1(n11951), .B2(n11950), .A(n11959), .ZN(n11953) );
  MUX2_X1 U14475 ( .A(n11959), .B(n11953), .S(n11952), .Z(n11954) );
  INV_X1 U14476 ( .A(n11954), .ZN(n11955) );
  INV_X1 U14477 ( .A(n12811), .ZN(n13051) );
  NAND2_X1 U14478 ( .A1(n13051), .A2(n12821), .ZN(n11956) );
  MUX2_X1 U14479 ( .A(n11957), .B(n11956), .S(n11959), .Z(n11958) );
  MUX2_X1 U14480 ( .A(n11961), .B(n11960), .S(n11959), .Z(n11962) );
  AOI211_X1 U14481 ( .C1(n11970), .C2(n11969), .A(n7629), .B(n11996), .ZN(
        n11971) );
  OAI21_X1 U14482 ( .B1(n11971), .B2(n11997), .A(n6741), .ZN(n11972) );
  INV_X1 U14483 ( .A(n12857), .ZN(n12853) );
  INV_X1 U14484 ( .A(n12889), .ZN(n11989) );
  INV_X1 U14485 ( .A(n12921), .ZN(n12923) );
  NAND4_X1 U14486 ( .A1(n15283), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11978) );
  NOR4_X1 U14487 ( .A1(n11979), .A2(n8567), .A3(n11978), .A4(n15324), .ZN(
        n11981) );
  NAND4_X1 U14488 ( .A1(n11981), .A2(n15308), .A3(n15268), .A4(n11980), .ZN(
        n11983) );
  NOR4_X1 U14489 ( .A1(n11985), .A2(n11984), .A3(n11983), .A4(n11982), .ZN(
        n11986) );
  NAND4_X1 U14490 ( .A1(n12934), .A2(n12944), .A3(n14637), .A4(n11986), .ZN(
        n11987) );
  NOR4_X1 U14491 ( .A1(n12898), .A2(n12911), .A3(n12923), .A4(n11987), .ZN(
        n11988) );
  NAND4_X1 U14492 ( .A1(n12853), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11991) );
  NOR4_X1 U14493 ( .A1(n12820), .A2(n11992), .A3(n12845), .A4(n11991), .ZN(
        n11993) );
  NAND4_X1 U14494 ( .A1(n12776), .A2(n12794), .A3(n11993), .A4(n12802), .ZN(
        n11994) );
  NOR4_X1 U14495 ( .A1(n11996), .A2(n11995), .A3(n12762), .A4(n11994), .ZN(
        n11999) );
  INV_X1 U14496 ( .A(n11997), .ZN(n11998) );
  NAND3_X1 U14497 ( .A1(n11999), .A2(n11998), .A3(n6741), .ZN(n12000) );
  XNOR2_X1 U14498 ( .A(n12000), .B(n12742), .ZN(n12001) );
  NAND2_X1 U14499 ( .A1(n12001), .A2(n6833), .ZN(n12002) );
  NOR3_X1 U14500 ( .A1(n15313), .A2(n8926), .A3(n12003), .ZN(n12006) );
  OAI21_X1 U14501 ( .B1(n12007), .B2(n12004), .A(P3_B_REG_SCAN_IN), .ZN(n12005) );
  OAI21_X1 U14502 ( .B1(n14016), .B2(n12009), .A(n14017), .ZN(n12010) );
  INV_X1 U14503 ( .A(n12010), .ZN(n12015) );
  NAND2_X1 U14504 ( .A1(n12189), .A2(n14287), .ZN(n12011) );
  NAND2_X1 U14505 ( .A1(n12012), .A2(n12011), .ZN(n12181) );
  MUX2_X1 U14506 ( .A(n12014), .B(n12013), .S(n12181), .Z(n12040) );
  MUX2_X1 U14507 ( .A(n14431), .B(n12015), .S(n12067), .Z(n12186) );
  AOI22_X1 U14508 ( .A1(n12018), .A2(n12017), .B1(n14043), .B2(n12016), .ZN(
        n12020) );
  AND2_X1 U14509 ( .A1(n12023), .A2(n12031), .ZN(n12024) );
  MUX2_X1 U14510 ( .A(n12031), .B(n12030), .S(n12026), .Z(n12032) );
  NAND2_X1 U14511 ( .A1(n12026), .A2(n12033), .ZN(n12036) );
  NAND2_X1 U14512 ( .A1(n12040), .A2(n12034), .ZN(n12035) );
  MUX2_X1 U14513 ( .A(n12036), .B(n12035), .S(n6871), .Z(n12037) );
  MUX2_X1 U14514 ( .A(n12039), .B(n12038), .S(n12040), .Z(n12043) );
  MUX2_X1 U14515 ( .A(n12041), .B(n14038), .S(n12040), .Z(n12042) );
  OAI21_X1 U14516 ( .B1(n12044), .B2(n12043), .A(n12042), .ZN(n12046) );
  NAND2_X1 U14517 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  NAND2_X1 U14518 ( .A1(n12046), .A2(n12045), .ZN(n12049) );
  MUX2_X1 U14519 ( .A(n12047), .B(n14037), .S(n12040), .Z(n12050) );
  MUX2_X1 U14520 ( .A(n14037), .B(n12047), .S(n12040), .Z(n12048) );
  INV_X1 U14521 ( .A(n12050), .ZN(n12051) );
  MUX2_X1 U14522 ( .A(n12052), .B(n14036), .S(n12067), .Z(n12056) );
  MUX2_X1 U14523 ( .A(n14036), .B(n12052), .S(n12067), .Z(n12053) );
  NAND2_X1 U14524 ( .A1(n12054), .A2(n12053), .ZN(n12058) );
  MUX2_X1 U14525 ( .A(n12059), .B(n14846), .S(n12195), .Z(n12062) );
  BUF_X1 U14526 ( .A(n12026), .Z(n12067) );
  MUX2_X1 U14527 ( .A(n14035), .B(n12060), .S(n12067), .Z(n12061) );
  MUX2_X1 U14528 ( .A(n14034), .B(n12063), .S(n12195), .Z(n12065) );
  NAND2_X1 U14529 ( .A1(n12063), .A2(n14034), .ZN(n12064) );
  NAND2_X1 U14530 ( .A1(n12065), .A2(n12064), .ZN(n12066) );
  MUX2_X1 U14531 ( .A(n12069), .B(n12068), .S(n12067), .Z(n12072) );
  MUX2_X1 U14532 ( .A(n14033), .B(n12070), .S(n12195), .Z(n12071) );
  MUX2_X1 U14533 ( .A(n14032), .B(n12073), .S(n12195), .Z(n12076) );
  MUX2_X1 U14534 ( .A(n14032), .B(n12073), .S(n12067), .Z(n12074) );
  NAND2_X1 U14535 ( .A1(n12075), .A2(n12074), .ZN(n12079) );
  NAND2_X1 U14536 ( .A1(n12077), .A2(n7189), .ZN(n12078) );
  MUX2_X1 U14537 ( .A(n14031), .B(n12080), .S(n12177), .Z(n12082) );
  MUX2_X1 U14538 ( .A(n14031), .B(n12080), .S(n12195), .Z(n12081) );
  INV_X1 U14539 ( .A(n12082), .ZN(n12083) );
  MUX2_X1 U14540 ( .A(n14029), .B(n12246), .S(n12195), .Z(n12087) );
  MUX2_X1 U14541 ( .A(n14029), .B(n12246), .S(n12177), .Z(n12084) );
  NAND2_X1 U14542 ( .A1(n12085), .A2(n12084), .ZN(n12091) );
  INV_X1 U14543 ( .A(n12086), .ZN(n12089) );
  INV_X1 U14544 ( .A(n12087), .ZN(n12088) );
  NAND2_X1 U14545 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  MUX2_X1 U14546 ( .A(n14028), .B(n13964), .S(n12177), .Z(n12093) );
  MUX2_X1 U14547 ( .A(n14028), .B(n13964), .S(n12195), .Z(n12092) );
  AND2_X1 U14548 ( .A1(n12101), .A2(n12095), .ZN(n12098) );
  AND2_X1 U14549 ( .A1(n12100), .A2(n12096), .ZN(n12097) );
  MUX2_X1 U14550 ( .A(n12098), .B(n12097), .S(n12177), .Z(n12099) );
  MUX2_X1 U14551 ( .A(n12101), .B(n12100), .S(n12195), .Z(n12102) );
  NAND2_X1 U14552 ( .A1(n12120), .A2(n14024), .ZN(n12103) );
  NAND2_X1 U14553 ( .A1(n12177), .A2(n14304), .ZN(n12105) );
  AOI21_X1 U14554 ( .B1(n12103), .B2(n12105), .A(n14301), .ZN(n12109) );
  INV_X1 U14555 ( .A(n14024), .ZN(n14318) );
  NAND2_X1 U14556 ( .A1(n12120), .A2(n14318), .ZN(n12104) );
  OR2_X1 U14557 ( .A1(n14413), .A2(n12067), .ZN(n12110) );
  AOI21_X1 U14558 ( .B1(n12104), .B2(n12110), .A(n14409), .ZN(n12108) );
  NAND2_X1 U14559 ( .A1(n12195), .A2(n14024), .ZN(n12111) );
  OR2_X1 U14560 ( .A1(n14413), .A2(n12111), .ZN(n12107) );
  INV_X1 U14561 ( .A(n12105), .ZN(n12119) );
  NAND2_X1 U14562 ( .A1(n12119), .A2(n14318), .ZN(n12106) );
  NAND2_X1 U14563 ( .A1(n12107), .A2(n12106), .ZN(n12114) );
  INV_X1 U14564 ( .A(n12110), .ZN(n12113) );
  INV_X1 U14565 ( .A(n12111), .ZN(n12112) );
  AOI21_X1 U14566 ( .B1(n12120), .B2(n12113), .A(n12112), .ZN(n12117) );
  INV_X1 U14567 ( .A(n12120), .ZN(n12116) );
  INV_X1 U14568 ( .A(n12114), .ZN(n12115) );
  OAI22_X1 U14569 ( .A1(n12117), .A2(n14409), .B1(n12116), .B2(n12115), .ZN(
        n12118) );
  INV_X1 U14570 ( .A(n12118), .ZN(n12125) );
  NAND2_X1 U14571 ( .A1(n12120), .A2(n12119), .ZN(n12122) );
  NAND2_X1 U14572 ( .A1(n12177), .A2(n14318), .ZN(n12121) );
  AOI21_X1 U14573 ( .B1(n12122), .B2(n12121), .A(n14301), .ZN(n12123) );
  INV_X1 U14574 ( .A(n12123), .ZN(n12124) );
  MUX2_X1 U14575 ( .A(n14305), .B(n14464), .S(n12195), .Z(n12126) );
  OAI21_X1 U14576 ( .B1(n12129), .B2(n12127), .A(n12126), .ZN(n12131) );
  AOI21_X1 U14577 ( .B1(n12129), .B2(n12128), .A(n14262), .ZN(n12130) );
  MUX2_X1 U14578 ( .A(n12133), .B(n12132), .S(n12067), .Z(n12134) );
  MUX2_X1 U14579 ( .A(n14396), .B(n14459), .S(n12067), .Z(n12136) );
  MUX2_X1 U14580 ( .A(n14269), .B(n14251), .S(n12195), .Z(n12135) );
  MUX2_X1 U14581 ( .A(n14240), .B(n14386), .S(n12195), .Z(n12140) );
  MUX2_X1 U14582 ( .A(n14240), .B(n14386), .S(n12177), .Z(n12137) );
  NAND2_X1 U14583 ( .A1(n12138), .A2(n12137), .ZN(n12144) );
  INV_X1 U14584 ( .A(n12139), .ZN(n12142) );
  INV_X1 U14585 ( .A(n12140), .ZN(n12141) );
  NAND2_X1 U14586 ( .A1(n12142), .A2(n12141), .ZN(n12143) );
  MUX2_X1 U14587 ( .A(n14224), .B(n14211), .S(n12067), .Z(n12146) );
  MUX2_X1 U14588 ( .A(n14224), .B(n14211), .S(n12195), .Z(n12145) );
  INV_X1 U14589 ( .A(n12146), .ZN(n12147) );
  MUX2_X1 U14590 ( .A(n14179), .B(n14372), .S(n12177), .Z(n12151) );
  MUX2_X1 U14591 ( .A(n14179), .B(n14372), .S(n12195), .Z(n12148) );
  INV_X1 U14592 ( .A(n12150), .ZN(n12153) );
  INV_X1 U14593 ( .A(n12151), .ZN(n12152) );
  MUX2_X1 U14594 ( .A(n14021), .B(n14185), .S(n12067), .Z(n12155) );
  MUX2_X1 U14595 ( .A(n14021), .B(n14185), .S(n12195), .Z(n12154) );
  MUX2_X1 U14596 ( .A(n14020), .B(n14167), .S(n12195), .Z(n12159) );
  NAND2_X1 U14597 ( .A1(n12156), .A2(n12159), .ZN(n12158) );
  MUX2_X1 U14598 ( .A(n14020), .B(n14167), .S(n12177), .Z(n12157) );
  NAND2_X1 U14599 ( .A1(n12158), .A2(n12157), .ZN(n12163) );
  INV_X1 U14600 ( .A(n12159), .ZN(n12160) );
  NAND2_X1 U14601 ( .A1(n12161), .A2(n12160), .ZN(n12162) );
  MUX2_X1 U14602 ( .A(n14019), .B(n13987), .S(n12067), .Z(n12165) );
  MUX2_X1 U14603 ( .A(n14019), .B(n13987), .S(n12195), .Z(n12164) );
  MUX2_X1 U14604 ( .A(n14104), .B(n14133), .S(n12195), .Z(n12169) );
  NAND2_X1 U14605 ( .A1(n12168), .A2(n12169), .ZN(n12167) );
  MUX2_X1 U14606 ( .A(n14104), .B(n14133), .S(n12177), .Z(n12166) );
  NAND2_X1 U14607 ( .A1(n12167), .A2(n12166), .ZN(n12173) );
  INV_X1 U14608 ( .A(n12168), .ZN(n12171) );
  INV_X1 U14609 ( .A(n12169), .ZN(n12170) );
  NAND2_X1 U14610 ( .A1(n12171), .A2(n12170), .ZN(n12172) );
  MUX2_X1 U14611 ( .A(n14018), .B(n14435), .S(n12067), .Z(n12175) );
  MUX2_X1 U14612 ( .A(n14018), .B(n14435), .S(n12195), .Z(n12174) );
  INV_X1 U14613 ( .A(n12175), .ZN(n12176) );
  MUX2_X1 U14614 ( .A(n14105), .B(n12178), .S(n12040), .Z(n12179) );
  MUX2_X1 U14615 ( .A(n14105), .B(n12178), .S(n12177), .Z(n12180) );
  INV_X1 U14616 ( .A(n12181), .ZN(n12182) );
  NAND2_X1 U14617 ( .A1(n12195), .A2(n14016), .ZN(n12196) );
  OAI21_X1 U14618 ( .B1(n12183), .B2(n12182), .A(n12196), .ZN(n12184) );
  AOI22_X1 U14619 ( .A1(n14431), .A2(n12067), .B1(n14017), .B2(n12184), .ZN(
        n12185) );
  XNOR2_X1 U14620 ( .A(n12194), .B(n14016), .ZN(n12199) );
  NAND2_X1 U14621 ( .A1(n12189), .A2(n12188), .ZN(n12190) );
  NAND2_X1 U14622 ( .A1(n12191), .A2(n12190), .ZN(n12193) );
  NAND2_X1 U14623 ( .A1(n12193), .A2(n12192), .ZN(n12227) );
  NAND2_X1 U14624 ( .A1(n12227), .A2(n12225), .ZN(n12228) );
  INV_X1 U14625 ( .A(n12228), .ZN(n12198) );
  MUX2_X1 U14626 ( .A(n12195), .B(n14016), .S(n12194), .Z(n12197) );
  INV_X1 U14627 ( .A(n12199), .ZN(n12229) );
  NAND4_X1 U14628 ( .A1(n7183), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12206) );
  NOR3_X1 U14629 ( .A1(n12206), .A2(n12205), .A3(n12204), .ZN(n12209) );
  NAND4_X1 U14630 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(
        n12211) );
  NOR4_X1 U14631 ( .A1(n12214), .A2(n12213), .A3(n7398), .A4(n12211), .ZN(
        n12217) );
  NAND4_X1 U14632 ( .A1(n14294), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12219) );
  NOR4_X1 U14633 ( .A1(n12219), .A2(n12218), .A3(n14327), .A4(n8084), .ZN(
        n12220) );
  NAND4_X1 U14634 ( .A1(n14247), .A2(n8324), .A3(n12220), .A4(n14278), .ZN(
        n12221) );
  NOR4_X1 U14635 ( .A1(n14192), .A2(n14209), .A3(n14225), .A4(n12221), .ZN(
        n12222) );
  INV_X1 U14636 ( .A(n12227), .ZN(n12231) );
  NOR2_X1 U14637 ( .A1(n12229), .A2(n12228), .ZN(n12230) );
  MUX2_X1 U14638 ( .A(n12231), .B(n12230), .S(n6745), .Z(n12232) );
  INV_X1 U14639 ( .A(n12232), .ZN(n12233) );
  NAND4_X1 U14640 ( .A1(n12237), .A2(n14238), .A3(n14727), .A4(n12236), .ZN(
        n12238) );
  OAI211_X1 U14641 ( .C1(n14496), .C2(n12240), .A(n12238), .B(P1_B_REG_SCAN_IN), .ZN(n12239) );
  NAND2_X1 U14642 ( .A1(n12246), .A2(n6688), .ZN(n12242) );
  NAND2_X1 U14643 ( .A1(n12378), .A2(n14029), .ZN(n12241) );
  NAND2_X1 U14644 ( .A1(n12242), .A2(n12241), .ZN(n12243) );
  XNOR2_X1 U14645 ( .A(n12243), .B(n12329), .ZN(n12251) );
  NOR2_X1 U14646 ( .A1(n12322), .A2(n12244), .ZN(n12245) );
  AOI21_X1 U14647 ( .B1(n12246), .B2(n12378), .A(n12245), .ZN(n12252) );
  XNOR2_X1 U14648 ( .A(n12251), .B(n12252), .ZN(n13890) );
  INV_X1 U14649 ( .A(n12247), .ZN(n12250) );
  INV_X1 U14650 ( .A(n12248), .ZN(n12249) );
  NOR2_X1 U14651 ( .A1(n12250), .A2(n12249), .ZN(n13891) );
  INV_X1 U14652 ( .A(n12251), .ZN(n12254) );
  INV_X1 U14653 ( .A(n12252), .ZN(n12253) );
  NAND2_X1 U14654 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  NOR2_X1 U14655 ( .A1(n12322), .A2(n12256), .ZN(n12257) );
  AOI21_X1 U14656 ( .B1(n13964), .B2(n12378), .A(n12257), .ZN(n12259) );
  AOI22_X1 U14657 ( .A1(n13964), .A2(n6688), .B1(n12378), .B2(n14028), .ZN(
        n12258) );
  XNOR2_X1 U14658 ( .A(n12258), .B(n12376), .ZN(n12260) );
  XOR2_X1 U14659 ( .A(n12259), .B(n12260), .Z(n13957) );
  NAND2_X1 U14660 ( .A1(n13958), .A2(n13957), .ZN(n12262) );
  OR2_X1 U14661 ( .A1(n12260), .A2(n12259), .ZN(n12261) );
  NAND2_X1 U14662 ( .A1(n14681), .A2(n6688), .ZN(n12264) );
  NAND2_X1 U14663 ( .A1(n12378), .A2(n14027), .ZN(n12263) );
  NAND2_X1 U14664 ( .A1(n12264), .A2(n12263), .ZN(n12265) );
  XNOR2_X1 U14665 ( .A(n12265), .B(n12329), .ZN(n12268) );
  NOR2_X1 U14666 ( .A1(n12322), .A2(n13959), .ZN(n12266) );
  AOI21_X1 U14667 ( .B1(n14681), .B2(n12378), .A(n12266), .ZN(n12267) );
  NAND2_X1 U14668 ( .A1(n12268), .A2(n12267), .ZN(n12269) );
  OAI21_X1 U14669 ( .B1(n12268), .B2(n12267), .A(n12269), .ZN(n13853) );
  NAND2_X1 U14670 ( .A1(n14421), .A2(n6688), .ZN(n12271) );
  NAND2_X1 U14671 ( .A1(n12378), .A2(n14026), .ZN(n12270) );
  NAND2_X1 U14672 ( .A1(n12271), .A2(n12270), .ZN(n12272) );
  XNOR2_X1 U14673 ( .A(n12272), .B(n12376), .ZN(n13916) );
  NAND2_X1 U14674 ( .A1(n14421), .A2(n12378), .ZN(n12274) );
  NAND2_X1 U14675 ( .A1(n12375), .A2(n14026), .ZN(n12273) );
  NAND2_X1 U14676 ( .A1(n12274), .A2(n12273), .ZN(n13915) );
  NAND2_X1 U14677 ( .A1(n14413), .A2(n6688), .ZN(n12276) );
  NAND2_X1 U14678 ( .A1(n12378), .A2(n14025), .ZN(n12275) );
  NAND2_X1 U14679 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  XNOR2_X1 U14680 ( .A(n12277), .B(n12329), .ZN(n12280) );
  NOR2_X1 U14681 ( .A1(n12322), .A2(n14304), .ZN(n12278) );
  AOI21_X1 U14682 ( .B1(n14413), .B2(n12378), .A(n12278), .ZN(n12279) );
  NAND2_X1 U14683 ( .A1(n12280), .A2(n12279), .ZN(n13927) );
  OAI21_X1 U14684 ( .B1(n12280), .B2(n12279), .A(n13927), .ZN(n13919) );
  AOI21_X1 U14685 ( .B1(n13916), .B2(n13915), .A(n13919), .ZN(n12281) );
  NAND2_X1 U14686 ( .A1(n12282), .A2(n12281), .ZN(n13918) );
  NAND2_X1 U14687 ( .A1(n13918), .A2(n13927), .ZN(n12291) );
  OAI22_X1 U14688 ( .A1(n14301), .A2(n6878), .B1(n14318), .B2(n6683), .ZN(
        n12283) );
  XNOR2_X1 U14689 ( .A(n12283), .B(n12329), .ZN(n12286) );
  OR2_X1 U14690 ( .A1(n14301), .A2(n6683), .ZN(n12285) );
  NAND2_X1 U14691 ( .A1(n12375), .A2(n14024), .ZN(n12284) );
  NAND2_X1 U14692 ( .A1(n12286), .A2(n12287), .ZN(n12292) );
  INV_X1 U14693 ( .A(n12286), .ZN(n12289) );
  INV_X1 U14694 ( .A(n12287), .ZN(n12288) );
  NAND2_X1 U14695 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  AND2_X1 U14696 ( .A1(n12292), .A2(n12290), .ZN(n13928) );
  OR2_X1 U14697 ( .A1(n14464), .A2(n6683), .ZN(n12294) );
  NAND2_X1 U14698 ( .A1(n12375), .A2(n14023), .ZN(n12293) );
  NAND2_X1 U14699 ( .A1(n12294), .A2(n12293), .ZN(n12300) );
  OAI22_X1 U14700 ( .A1(n14464), .A2(n6878), .B1(n14305), .B2(n6683), .ZN(
        n12295) );
  XNOR2_X1 U14701 ( .A(n12295), .B(n12376), .ZN(n12301) );
  XOR2_X1 U14702 ( .A(n12300), .B(n12301), .Z(n13981) );
  NAND2_X1 U14703 ( .A1(n14265), .A2(n6688), .ZN(n12297) );
  NAND2_X1 U14704 ( .A1(n12378), .A2(n14237), .ZN(n12296) );
  NAND2_X1 U14705 ( .A1(n12297), .A2(n12296), .ZN(n12298) );
  XNOR2_X1 U14706 ( .A(n12298), .B(n12329), .ZN(n12303) );
  NOR2_X1 U14707 ( .A1(n12322), .A2(n14279), .ZN(n12299) );
  AOI21_X1 U14708 ( .B1(n14265), .B2(n12378), .A(n12299), .ZN(n12304) );
  XNOR2_X1 U14709 ( .A(n12303), .B(n12304), .ZN(n13873) );
  NOR2_X1 U14710 ( .A1(n12301), .A2(n12300), .ZN(n13874) );
  NOR2_X1 U14711 ( .A1(n13873), .A2(n13874), .ZN(n12302) );
  INV_X1 U14712 ( .A(n12303), .ZN(n12306) );
  INV_X1 U14713 ( .A(n12304), .ZN(n12305) );
  NAND2_X1 U14714 ( .A1(n12306), .A2(n12305), .ZN(n12307) );
  OAI22_X1 U14715 ( .A1(n6897), .A2(n6683), .B1(n14396), .B2(n12322), .ZN(
        n12309) );
  OAI22_X1 U14716 ( .A1(n6897), .A2(n6878), .B1(n14396), .B2(n6683), .ZN(
        n12308) );
  XNOR2_X1 U14717 ( .A(n12308), .B(n12376), .ZN(n12310) );
  XOR2_X1 U14718 ( .A(n12309), .B(n12310), .Z(n13948) );
  NAND2_X1 U14719 ( .A1(n12310), .A2(n12309), .ZN(n12311) );
  NAND2_X1 U14720 ( .A1(n14386), .A2(n6688), .ZN(n12313) );
  NAND2_X1 U14721 ( .A1(n14240), .A2(n12378), .ZN(n12312) );
  NAND2_X1 U14722 ( .A1(n12313), .A2(n12312), .ZN(n12314) );
  XNOR2_X1 U14723 ( .A(n12314), .B(n12329), .ZN(n12317) );
  AND2_X1 U14724 ( .A1(n14240), .A2(n12375), .ZN(n12315) );
  AOI21_X1 U14725 ( .B1(n14386), .B2(n12378), .A(n12315), .ZN(n12316) );
  NAND2_X1 U14726 ( .A1(n12317), .A2(n12316), .ZN(n13967) );
  OAI21_X1 U14727 ( .B1(n12317), .B2(n12316), .A(n13967), .ZN(n13883) );
  NAND2_X1 U14728 ( .A1(n14211), .A2(n6688), .ZN(n12319) );
  NAND2_X1 U14729 ( .A1(n12378), .A2(n14224), .ZN(n12318) );
  NAND2_X1 U14730 ( .A1(n12319), .A2(n12318), .ZN(n12320) );
  XNOR2_X1 U14731 ( .A(n12320), .B(n12329), .ZN(n12324) );
  NOR2_X1 U14732 ( .A1(n12322), .A2(n12321), .ZN(n12323) );
  AOI21_X1 U14733 ( .B1(n14211), .B2(n12378), .A(n12323), .ZN(n12325) );
  NAND2_X1 U14734 ( .A1(n12324), .A2(n12325), .ZN(n13866) );
  INV_X1 U14735 ( .A(n12324), .ZN(n12327) );
  INV_X1 U14736 ( .A(n12325), .ZN(n12326) );
  NAND2_X1 U14737 ( .A1(n12327), .A2(n12326), .ZN(n12328) );
  OAI22_X1 U14738 ( .A1(n14372), .A2(n6878), .B1(n14179), .B2(n6683), .ZN(
        n12330) );
  XNOR2_X1 U14739 ( .A(n12330), .B(n12329), .ZN(n12334) );
  INV_X1 U14740 ( .A(n14179), .ZN(n14022) );
  NAND2_X1 U14741 ( .A1(n12375), .A2(n14022), .ZN(n12332) );
  NAND2_X1 U14742 ( .A1(n12334), .A2(n12335), .ZN(n12339) );
  INV_X1 U14743 ( .A(n12334), .ZN(n12337) );
  INV_X1 U14744 ( .A(n12335), .ZN(n12336) );
  NAND2_X1 U14745 ( .A1(n12337), .A2(n12336), .ZN(n12338) );
  NAND2_X1 U14746 ( .A1(n14185), .A2(n6688), .ZN(n12341) );
  NAND2_X1 U14747 ( .A1(n12378), .A2(n14021), .ZN(n12340) );
  NAND2_X1 U14748 ( .A1(n12341), .A2(n12340), .ZN(n12342) );
  XNOR2_X1 U14749 ( .A(n12342), .B(n12376), .ZN(n12346) );
  NAND2_X1 U14750 ( .A1(n14185), .A2(n12378), .ZN(n12344) );
  NAND2_X1 U14751 ( .A1(n12375), .A2(n14021), .ZN(n12343) );
  NAND2_X1 U14752 ( .A1(n12344), .A2(n12343), .ZN(n12345) );
  NOR2_X1 U14753 ( .A1(n12346), .A2(n12345), .ZN(n12347) );
  AOI21_X1 U14754 ( .B1(n12346), .B2(n12345), .A(n12347), .ZN(n13940) );
  INV_X1 U14755 ( .A(n12347), .ZN(n12348) );
  NAND2_X1 U14756 ( .A1(n14167), .A2(n6688), .ZN(n12350) );
  NAND2_X1 U14757 ( .A1(n12378), .A2(n14020), .ZN(n12349) );
  NAND2_X1 U14758 ( .A1(n12350), .A2(n12349), .ZN(n12351) );
  XNOR2_X1 U14759 ( .A(n12351), .B(n12376), .ZN(n12355) );
  NAND2_X1 U14760 ( .A1(n14167), .A2(n12378), .ZN(n12353) );
  NAND2_X1 U14761 ( .A1(n12375), .A2(n14020), .ZN(n12352) );
  NAND2_X1 U14762 ( .A1(n12353), .A2(n12352), .ZN(n12354) );
  NOR2_X1 U14763 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  AOI21_X1 U14764 ( .B1(n12355), .B2(n12354), .A(n12356), .ZN(n13905) );
  INV_X1 U14765 ( .A(n12356), .ZN(n12357) );
  NAND2_X1 U14766 ( .A1(n6884), .A2(n6688), .ZN(n12360) );
  NAND2_X1 U14767 ( .A1(n12378), .A2(n14019), .ZN(n12359) );
  NAND2_X1 U14768 ( .A1(n12360), .A2(n12359), .ZN(n12361) );
  XNOR2_X1 U14769 ( .A(n12361), .B(n12376), .ZN(n12365) );
  NAND2_X1 U14770 ( .A1(n6884), .A2(n12378), .ZN(n12363) );
  NAND2_X1 U14771 ( .A1(n12375), .A2(n14019), .ZN(n12362) );
  NAND2_X1 U14772 ( .A1(n12363), .A2(n12362), .ZN(n12364) );
  NOR2_X1 U14773 ( .A1(n12365), .A2(n12364), .ZN(n12366) );
  AOI21_X1 U14774 ( .B1(n12365), .B2(n12364), .A(n12366), .ZN(n13990) );
  NAND2_X1 U14775 ( .A1(n14133), .A2(n6688), .ZN(n12368) );
  NAND2_X1 U14776 ( .A1(n12378), .A2(n14104), .ZN(n12367) );
  NAND2_X1 U14777 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  XNOR2_X1 U14778 ( .A(n12369), .B(n12376), .ZN(n12373) );
  NAND2_X1 U14779 ( .A1(n14133), .A2(n12378), .ZN(n12371) );
  NAND2_X1 U14780 ( .A1(n12375), .A2(n14104), .ZN(n12370) );
  NAND2_X1 U14781 ( .A1(n12371), .A2(n12370), .ZN(n12372) );
  NOR2_X1 U14782 ( .A1(n12373), .A2(n12372), .ZN(n12374) );
  AOI21_X1 U14783 ( .B1(n12373), .B2(n12372), .A(n12374), .ZN(n13843) );
  AOI22_X1 U14784 ( .A1(n14435), .A2(n12378), .B1(n12375), .B2(n14018), .ZN(
        n12377) );
  XNOR2_X1 U14785 ( .A(n12377), .B(n12376), .ZN(n12380) );
  AOI22_X1 U14786 ( .A1(n14435), .A2(n6688), .B1(n12378), .B2(n14018), .ZN(
        n12379) );
  XNOR2_X1 U14787 ( .A(n12380), .B(n12379), .ZN(n12381) );
  XNOR2_X1 U14788 ( .A(n12382), .B(n12381), .ZN(n12387) );
  AOI22_X1 U14789 ( .A1(n14007), .A2(n14104), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12384) );
  NAND2_X1 U14790 ( .A1(n13950), .A2(n14105), .ZN(n12383) );
  OAI211_X1 U14791 ( .C1(n14010), .C2(n14115), .A(n12384), .B(n12383), .ZN(
        n12385) );
  AOI21_X1 U14792 ( .B1(n14435), .B2(n14012), .A(n12385), .ZN(n12386) );
  OAI21_X1 U14793 ( .B1(n12387), .B2(n14014), .A(n12386), .ZN(P1_U3220) );
  INV_X1 U14794 ( .A(n12388), .ZN(n12389) );
  NAND2_X1 U14795 ( .A1(n12389), .A2(n15332), .ZN(n12753) );
  OAI21_X1 U14796 ( .B1(n12390), .B2(n14652), .A(n12753), .ZN(n12393) );
  INV_X1 U14797 ( .A(n12394), .ZN(n12395) );
  OAI222_X1 U14798 ( .A1(P3_U3151), .A2(n8411), .B1(n13130), .B2(n15517), .C1(
        n11825), .C2(n12395), .ZN(P3_U3265) );
  XNOR2_X1 U14799 ( .A(n12787), .B(n12484), .ZN(n12480) );
  XNOR2_X1 U14800 ( .A(n12480), .B(n12766), .ZN(n12482) );
  INV_X1 U14801 ( .A(n12396), .ZN(n12397) );
  NAND2_X1 U14802 ( .A1(n12398), .A2(n12397), .ZN(n12399) );
  XNOR2_X1 U14803 ( .A(n15153), .B(n12435), .ZN(n12402) );
  XNOR2_X1 U14804 ( .A(n12402), .B(n12401), .ZN(n15147) );
  NAND2_X1 U14805 ( .A1(n12402), .A2(n12401), .ZN(n12403) );
  XNOR2_X1 U14806 ( .A(n12587), .B(n12435), .ZN(n12405) );
  NAND2_X1 U14807 ( .A1(n12584), .A2(n12583), .ZN(n12408) );
  INV_X1 U14808 ( .A(n12404), .ZN(n12406) );
  NAND2_X1 U14809 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  NAND2_X1 U14810 ( .A1(n12408), .A2(n12407), .ZN(n12512) );
  XNOR2_X1 U14811 ( .A(n12517), .B(n12435), .ZN(n12409) );
  XNOR2_X1 U14812 ( .A(n12409), .B(n12566), .ZN(n12511) );
  NAND2_X1 U14813 ( .A1(n12512), .A2(n12511), .ZN(n12411) );
  NAND2_X1 U14814 ( .A1(n12409), .A2(n14639), .ZN(n12410) );
  NAND2_X1 U14815 ( .A1(n12411), .A2(n12410), .ZN(n12565) );
  XNOR2_X1 U14816 ( .A(n14641), .B(n12484), .ZN(n12563) );
  AND2_X1 U14817 ( .A1(n12563), .A2(n12562), .ZN(n12412) );
  OR2_X2 U14818 ( .A1(n12565), .A2(n12412), .ZN(n12415) );
  INV_X1 U14819 ( .A(n12563), .ZN(n12413) );
  NAND2_X1 U14820 ( .A1(n12413), .A2(n12947), .ZN(n12414) );
  XNOR2_X1 U14821 ( .A(n13113), .B(n12435), .ZN(n12416) );
  XNOR2_X1 U14822 ( .A(n12416), .B(n14640), .ZN(n12453) );
  INV_X1 U14823 ( .A(n12416), .ZN(n12417) );
  NAND2_X1 U14824 ( .A1(n12417), .A2(n14640), .ZN(n12418) );
  XNOR2_X1 U14825 ( .A(n13102), .B(n12435), .ZN(n12419) );
  XNOR2_X1 U14826 ( .A(n12419), .B(n12949), .ZN(n12612) );
  INV_X1 U14827 ( .A(n12419), .ZN(n12420) );
  NAND2_X1 U14828 ( .A1(n12420), .A2(n12949), .ZN(n12421) );
  XNOR2_X1 U14829 ( .A(n13095), .B(n12484), .ZN(n12529) );
  XNOR2_X1 U14830 ( .A(n13089), .B(n12435), .ZN(n12422) );
  XNOR2_X1 U14831 ( .A(n12422), .B(n12596), .ZN(n12537) );
  INV_X1 U14832 ( .A(n12422), .ZN(n12424) );
  XNOR2_X1 U14833 ( .A(n13083), .B(n12435), .ZN(n12425) );
  XNOR2_X1 U14834 ( .A(n12425), .B(n12912), .ZN(n12593) );
  INV_X1 U14835 ( .A(n12425), .ZN(n12426) );
  NAND2_X1 U14836 ( .A1(n12426), .A2(n12912), .ZN(n12427) );
  XNOR2_X1 U14837 ( .A(n13080), .B(n12435), .ZN(n12428) );
  XNOR2_X1 U14838 ( .A(n12428), .B(n12597), .ZN(n12472) );
  NAND2_X1 U14839 ( .A1(n12428), .A2(n12868), .ZN(n12429) );
  XNOR2_X1 U14840 ( .A(n12876), .B(n12435), .ZN(n12430) );
  XNOR2_X1 U14841 ( .A(n12430), .B(n12505), .ZN(n12556) );
  INV_X1 U14842 ( .A(n12430), .ZN(n12431) );
  XNOR2_X1 U14843 ( .A(n13070), .B(n12435), .ZN(n12432) );
  XNOR2_X1 U14844 ( .A(n12432), .B(n12869), .ZN(n12503) );
  INV_X1 U14845 ( .A(n12432), .ZN(n12433) );
  NAND2_X1 U14846 ( .A1(n12433), .A2(n12869), .ZN(n12434) );
  XNOR2_X1 U14847 ( .A(n13064), .B(n12435), .ZN(n12460) );
  XNOR2_X1 U14848 ( .A(n13054), .B(n12435), .ZN(n12550) );
  XNOR2_X1 U14849 ( .A(n12987), .B(n12435), .ZN(n12464) );
  OAI22_X1 U14850 ( .A1(n12550), .A2(n12833), .B1(n12579), .B2(n12464), .ZN(
        n12437) );
  INV_X1 U14851 ( .A(n12437), .ZN(n12436) );
  OAI21_X1 U14852 ( .B1(n12832), .B2(n12460), .A(n12436), .ZN(n12442) );
  OAI21_X1 U14853 ( .B1(n12465), .B2(n12846), .A(n12522), .ZN(n12440) );
  NOR3_X1 U14854 ( .A1(n12465), .A2(n12846), .A3(n12522), .ZN(n12439) );
  INV_X1 U14855 ( .A(n12460), .ZN(n12461) );
  NOR3_X1 U14856 ( .A1(n12437), .A2(n12461), .A3(n12573), .ZN(n12438) );
  AOI211_X1 U14857 ( .C1(n12550), .C2(n12440), .A(n12439), .B(n12438), .ZN(
        n12441) );
  OAI21_X2 U14858 ( .B1(n12462), .B2(n12442), .A(n12441), .ZN(n12520) );
  XNOR2_X1 U14859 ( .A(n12811), .B(n12484), .ZN(n12443) );
  XNOR2_X1 U14860 ( .A(n12443), .B(n12605), .ZN(n12521) );
  INV_X1 U14861 ( .A(n12443), .ZN(n12444) );
  XNOR2_X1 U14862 ( .A(n13044), .B(n12484), .ZN(n12445) );
  XNOR2_X1 U14863 ( .A(n12445), .B(n12523), .ZN(n12604) );
  OAI22_X1 U14864 ( .A1(n12603), .A2(n12604), .B1(n12445), .B2(n12523), .ZN(
        n12483) );
  XOR2_X1 U14865 ( .A(n12482), .B(n12483), .Z(n12450) );
  AOI22_X1 U14866 ( .A1(n12523), .A2(n12575), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12447) );
  NAND2_X1 U14867 ( .A1(n12788), .A2(n12619), .ZN(n12446) );
  OAI211_X1 U14868 ( .C1(n12782), .C2(n12578), .A(n12447), .B(n12446), .ZN(
        n12448) );
  AOI21_X1 U14869 ( .B1(n12787), .B2(n15140), .A(n12448), .ZN(n12449) );
  OAI21_X1 U14870 ( .B1(n12450), .B2(n15146), .A(n12449), .ZN(P3_U3154) );
  OAI21_X1 U14871 ( .B1(n12453), .B2(n12452), .A(n12451), .ZN(n12454) );
  NAND2_X1 U14872 ( .A1(n12454), .A2(n15134), .ZN(n12459) );
  INV_X1 U14873 ( .A(n12455), .ZN(n12952) );
  NAND2_X1 U14874 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n15249)
         );
  NAND2_X1 U14875 ( .A1(n12615), .A2(n12949), .ZN(n12456) );
  OAI211_X1 U14876 ( .C1(n12562), .C2(n12617), .A(n15249), .B(n12456), .ZN(
        n12457) );
  AOI21_X1 U14877 ( .B1(n12952), .B2(n12619), .A(n12457), .ZN(n12458) );
  OAI211_X1 U14878 ( .C1(n15154), .C2(n13113), .A(n12459), .B(n12458), .ZN(
        P3_U3155) );
  XNOR2_X1 U14879 ( .A(n12549), .B(n12579), .ZN(n12470) );
  INV_X1 U14880 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15756) );
  OAI22_X1 U14881 ( .A1(n12832), .A2(n12617), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15756), .ZN(n12467) );
  NOR2_X1 U14882 ( .A1(n12833), .A2(n12578), .ZN(n12466) );
  AOI211_X1 U14883 ( .C1(n12837), .C2(n12619), .A(n12467), .B(n12466), .ZN(
        n12469) );
  NAND2_X1 U14884 ( .A1(n12987), .A2(n15140), .ZN(n12468) );
  OAI211_X1 U14885 ( .C1(n12470), .C2(n15146), .A(n12469), .B(n12468), .ZN(
        P3_U3156) );
  OAI211_X1 U14886 ( .C1(n12473), .C2(n12472), .A(n12471), .B(n15134), .ZN(
        n12479) );
  OAI22_X1 U14887 ( .A1(n12474), .A2(n15315), .B1(n12543), .B2(n15313), .ZN(
        n12886) );
  NAND2_X1 U14888 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12730)
         );
  INV_X1 U14889 ( .A(n12730), .ZN(n12477) );
  INV_X1 U14890 ( .A(n12475), .ZN(n12891) );
  NOR2_X1 U14891 ( .A1(n15159), .A2(n12891), .ZN(n12476) );
  AOI211_X1 U14892 ( .C1(n15149), .C2(n12886), .A(n12477), .B(n12476), .ZN(
        n12478) );
  OAI211_X1 U14893 ( .C1(n15154), .C2(n13080), .A(n12479), .B(n12478), .ZN(
        P3_U3159) );
  INV_X1 U14894 ( .A(n12480), .ZN(n12481) );
  AOI22_X1 U14895 ( .A1(n12483), .A2(n12482), .B1(n12766), .B2(n12481), .ZN(
        n12486) );
  XNOR2_X1 U14896 ( .A(n12762), .B(n12484), .ZN(n12485) );
  XNOR2_X1 U14897 ( .A(n12486), .B(n12485), .ZN(n12491) );
  NOR2_X1 U14898 ( .A1(n12767), .A2(n12578), .ZN(n12489) );
  AOI22_X1 U14899 ( .A1(n12773), .A2(n12619), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12487) );
  OAI21_X1 U14900 ( .B1(n12766), .B2(n12617), .A(n12487), .ZN(n12488) );
  AOI211_X1 U14901 ( .C1(n13035), .C2(n15140), .A(n12489), .B(n12488), .ZN(
        n12490) );
  OAI21_X1 U14902 ( .B1(n12491), .B2(n15146), .A(n12490), .ZN(P3_U3160) );
  OAI211_X1 U14903 ( .C1(n12494), .C2(n12493), .A(n12492), .B(n15134), .ZN(
        n12501) );
  AOI22_X1 U14904 ( .A1(n15140), .A2(n12495), .B1(P3_REG3_REG_8__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12500) );
  AOI22_X1 U14905 ( .A1(n12575), .A2(n12497), .B1(n12615), .B2(n12496), .ZN(
        n12499) );
  OR2_X1 U14906 ( .A1(n15159), .A2(n7765), .ZN(n12498) );
  NAND4_X1 U14907 ( .A1(n12501), .A2(n12500), .A3(n12499), .A4(n12498), .ZN(
        P3_U3161) );
  INV_X1 U14908 ( .A(n13070), .ZN(n12510) );
  OAI211_X1 U14909 ( .C1(n12504), .C2(n12503), .A(n12502), .B(n15134), .ZN(
        n12509) );
  AOI22_X1 U14910 ( .A1(n12573), .A2(n12948), .B1(n12505), .B2(n12946), .ZN(
        n12861) );
  INV_X1 U14911 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12506) );
  OAI22_X1 U14912 ( .A1(n12861), .A2(n15143), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12506), .ZN(n12507) );
  AOI21_X1 U14913 ( .B1(n12864), .B2(n12619), .A(n12507), .ZN(n12508) );
  OAI211_X1 U14914 ( .C1(n12510), .C2(n15154), .A(n12509), .B(n12508), .ZN(
        P3_U3163) );
  XOR2_X1 U14915 ( .A(n12512), .B(n12511), .Z(n12519) );
  NAND2_X1 U14916 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n15207)
         );
  OAI21_X1 U14917 ( .B1(n12583), .B2(n12617), .A(n15207), .ZN(n12513) );
  AOI21_X1 U14918 ( .B1(n12615), .B2(n12947), .A(n12513), .ZN(n12514) );
  OAI21_X1 U14919 ( .B1(n12515), .B2(n15159), .A(n12514), .ZN(n12516) );
  AOI21_X1 U14920 ( .B1(n15140), .B2(n12517), .A(n12516), .ZN(n12518) );
  OAI21_X1 U14921 ( .B1(n12519), .B2(n15146), .A(n12518), .ZN(P3_U3164) );
  XOR2_X1 U14922 ( .A(n12521), .B(n12520), .Z(n12527) );
  AOI22_X1 U14923 ( .A1(n12523), .A2(n12948), .B1(n12946), .B2(n12522), .ZN(
        n12808) );
  AOI22_X1 U14924 ( .A1(n12810), .A2(n12619), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12524) );
  OAI21_X1 U14925 ( .B1(n12808), .B2(n15143), .A(n12524), .ZN(n12525) );
  AOI21_X1 U14926 ( .B1(n12811), .B2(n15140), .A(n12525), .ZN(n12526) );
  OAI21_X1 U14927 ( .B1(n12527), .B2(n15146), .A(n12526), .ZN(P3_U3165) );
  XNOR2_X1 U14928 ( .A(n12529), .B(n12528), .ZN(n12530) );
  XNOR2_X1 U14929 ( .A(n6912), .B(n12530), .ZN(n12536) );
  OAI22_X1 U14930 ( .A1(n12532), .A2(n15313), .B1(n12596), .B2(n15315), .ZN(
        n12925) );
  NAND2_X1 U14931 ( .A1(n12925), .A2(n15149), .ZN(n12533) );
  NAND2_X1 U14932 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12657)
         );
  OAI211_X1 U14933 ( .C1(n12928), .C2(n15159), .A(n12533), .B(n12657), .ZN(
        n12534) );
  AOI21_X1 U14934 ( .B1(n13095), .B2(n15140), .A(n12534), .ZN(n12535) );
  OAI21_X1 U14935 ( .B1(n12536), .B2(n15146), .A(n12535), .ZN(P3_U3166) );
  INV_X1 U14936 ( .A(n13089), .ZN(n12547) );
  AOI21_X1 U14937 ( .B1(n12538), .B2(n12537), .A(n15146), .ZN(n12540) );
  NAND2_X1 U14938 ( .A1(n12540), .A2(n12539), .ZN(n12546) );
  INV_X1 U14939 ( .A(n12541), .ZN(n12916) );
  NAND2_X1 U14940 ( .A1(n12937), .A2(n12575), .ZN(n12542) );
  NAND2_X1 U14941 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12691)
         );
  OAI211_X1 U14942 ( .C1(n12578), .C2(n12543), .A(n12542), .B(n12691), .ZN(
        n12544) );
  AOI21_X1 U14943 ( .B1(n12916), .B2(n12619), .A(n12544), .ZN(n12545) );
  OAI211_X1 U14944 ( .C1(n12547), .C2(n15154), .A(n12546), .B(n12545), .ZN(
        P3_U3168) );
  AOI22_X1 U14945 ( .A1(n12821), .A2(n12615), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12552) );
  NAND2_X1 U14946 ( .A1(n12824), .A2(n12619), .ZN(n12551) );
  OAI211_X1 U14947 ( .C1(n12579), .C2(n12617), .A(n12552), .B(n12551), .ZN(
        n12553) );
  AOI21_X1 U14948 ( .B1(n13054), .B2(n15140), .A(n12553), .ZN(n12554) );
  INV_X1 U14949 ( .A(n12876), .ZN(n13003) );
  OAI211_X1 U14950 ( .C1(n12557), .C2(n12556), .A(n12555), .B(n15134), .ZN(
        n12561) );
  AOI22_X1 U14951 ( .A1(n12869), .A2(n12615), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12558) );
  OAI21_X1 U14952 ( .B1(n12597), .B2(n12617), .A(n12558), .ZN(n12559) );
  AOI21_X1 U14953 ( .B1(n12872), .B2(n12619), .A(n12559), .ZN(n12560) );
  OAI211_X1 U14954 ( .C1(n13003), .C2(n15154), .A(n12561), .B(n12560), .ZN(
        P3_U3173) );
  XNOR2_X1 U14955 ( .A(n12563), .B(n12562), .ZN(n12564) );
  XNOR2_X1 U14956 ( .A(n12565), .B(n12564), .ZN(n12572) );
  AOI22_X1 U14957 ( .A1(n12566), .A2(n12575), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12568) );
  NAND2_X1 U14958 ( .A1(n12615), .A2(n12936), .ZN(n12567) );
  OAI211_X1 U14959 ( .C1(n14642), .C2(n15159), .A(n12568), .B(n12567), .ZN(
        n12569) );
  AOI21_X1 U14960 ( .B1(n12570), .B2(n15140), .A(n12569), .ZN(n12571) );
  OAI21_X1 U14961 ( .B1(n12572), .B2(n15146), .A(n12571), .ZN(P3_U3174) );
  XNOR2_X1 U14962 ( .A(n12574), .B(n12573), .ZN(n12582) );
  AOI22_X1 U14963 ( .A1(n12869), .A2(n12575), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12577) );
  NAND2_X1 U14964 ( .A1(n12619), .A2(n12849), .ZN(n12576) );
  OAI211_X1 U14965 ( .C1(n12579), .C2(n12578), .A(n12577), .B(n12576), .ZN(
        n12580) );
  AOI21_X1 U14966 ( .B1(n13064), .B2(n15140), .A(n12580), .ZN(n12581) );
  OAI21_X1 U14967 ( .B1(n12582), .B2(n15146), .A(n12581), .ZN(P3_U3175) );
  XNOR2_X1 U14968 ( .A(n12584), .B(n12583), .ZN(n12585) );
  NAND2_X1 U14969 ( .A1(n12585), .A2(n15134), .ZN(n12591) );
  AOI22_X1 U14970 ( .A1(n12586), .A2(n15149), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12590) );
  NAND2_X1 U14971 ( .A1(n15140), .A2(n12587), .ZN(n12589) );
  OR2_X1 U14972 ( .A1(n15159), .A2(n14656), .ZN(n12588) );
  NAND4_X1 U14973 ( .A1(n12591), .A2(n12590), .A3(n12589), .A4(n12588), .ZN(
        P3_U3176) );
  INV_X1 U14974 ( .A(n13083), .ZN(n12602) );
  OAI211_X1 U14975 ( .C1(n12594), .C2(n12593), .A(n12592), .B(n15134), .ZN(
        n12601) );
  INV_X1 U14976 ( .A(n12595), .ZN(n12903) );
  OAI22_X1 U14977 ( .A1(n12597), .A2(n15315), .B1(n12596), .B2(n15313), .ZN(
        n12900) );
  INV_X1 U14978 ( .A(n12900), .ZN(n12598) );
  NAND2_X1 U14979 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12705)
         );
  OAI21_X1 U14980 ( .B1(n12598), .B2(n15143), .A(n12705), .ZN(n12599) );
  AOI21_X1 U14981 ( .B1(n12903), .B2(n12619), .A(n12599), .ZN(n12600) );
  OAI211_X1 U14982 ( .C1(n12602), .C2(n15154), .A(n12601), .B(n12600), .ZN(
        P3_U3178) );
  XOR2_X1 U14983 ( .A(n12604), .B(n12603), .Z(n12610) );
  OAI22_X1 U14984 ( .A1(n12766), .A2(n15315), .B1(n12605), .B2(n15313), .ZN(
        n12796) );
  INV_X1 U14985 ( .A(n12799), .ZN(n12606) );
  OAI22_X1 U14986 ( .A1(n12606), .A2(n15159), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15555), .ZN(n12607) );
  AOI21_X1 U14987 ( .B1(n12796), .B2(n15149), .A(n12607), .ZN(n12609) );
  NAND2_X1 U14988 ( .A1(n13044), .A2(n15140), .ZN(n12608) );
  OAI211_X1 U14989 ( .C1(n12610), .C2(n15146), .A(n12609), .B(n12608), .ZN(
        P3_U3180) );
  INV_X1 U14990 ( .A(n13102), .ZN(n12622) );
  OAI211_X1 U14991 ( .C1(n12613), .C2(n12612), .A(n12611), .B(n15134), .ZN(
        n12621) );
  INV_X1 U14992 ( .A(n12614), .ZN(n12939) );
  NOR2_X1 U14993 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8388), .ZN(n14617) );
  AOI21_X1 U14994 ( .B1(n12937), .B2(n12615), .A(n14617), .ZN(n12616) );
  OAI21_X1 U14995 ( .B1(n14640), .B2(n12617), .A(n12616), .ZN(n12618) );
  AOI21_X1 U14996 ( .B1(n12939), .B2(n12619), .A(n12618), .ZN(n12620) );
  OAI211_X1 U14997 ( .C1(n12622), .C2(n15154), .A(n12621), .B(n12620), .ZN(
        P3_U3181) );
  MUX2_X1 U14998 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12623), .S(P3_U3897), .Z(
        P3_U3494) );
  XNOR2_X1 U14999 ( .A(n12673), .B(n13013), .ZN(n12637) );
  AND2_X1 U15000 ( .A1(n15248), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12652) );
  INV_X1 U15001 ( .A(n15194), .ZN(n12660) );
  NAND2_X1 U15002 ( .A1(n12625), .A2(n12624), .ZN(n12627) );
  INV_X1 U15003 ( .A(n12627), .ZN(n12626) );
  NOR2_X1 U15004 ( .A1(n12660), .A2(n12626), .ZN(n12628) );
  XNOR2_X1 U15005 ( .A(n12627), .B(n15194), .ZN(n15198) );
  NOR2_X1 U15006 ( .A1(n12628), .A2(n15197), .ZN(n15217) );
  XNOR2_X1 U15007 ( .A(n15214), .B(n12646), .ZN(n15218) );
  NAND2_X1 U15008 ( .A1(n12663), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12629) );
  INV_X1 U15009 ( .A(n12631), .ZN(n12630) );
  INV_X1 U15010 ( .A(n12652), .ZN(n12632) );
  OAI21_X1 U15011 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n15248), .A(n12632), 
        .ZN(n15260) );
  NOR2_X1 U15012 ( .A1(n14626), .A2(n12633), .ZN(n12634) );
  INV_X1 U15013 ( .A(n12683), .ZN(n12635) );
  AOI21_X1 U15014 ( .B1(n12637), .B2(n12636), .A(n12635), .ZN(n12681) );
  MUX2_X1 U15015 ( .A(n12927), .B(n13013), .S(n6684), .Z(n12639) );
  INV_X1 U15016 ( .A(n12639), .ZN(n12638) );
  NOR2_X1 U15017 ( .A1(n12638), .A2(n12692), .ZN(n12688) );
  NOR2_X1 U15018 ( .A1(n12639), .A2(n12673), .ZN(n12685) );
  NOR2_X1 U15019 ( .A1(n12688), .A2(n12685), .ZN(n12655) );
  MUX2_X1 U15020 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12735), .Z(n12649) );
  OAI22_X1 U15021 ( .A1(n12643), .A2(n12642), .B1(n12641), .B2(n12640), .ZN(
        n15191) );
  MUX2_X1 U15022 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12735), .Z(n12644) );
  XNOR2_X1 U15023 ( .A(n12644), .B(n12660), .ZN(n15190) );
  INV_X1 U15024 ( .A(n12644), .ZN(n12645) );
  MUX2_X1 U15025 ( .A(n12664), .B(n12646), .S(n12735), .Z(n12647) );
  NOR2_X1 U15026 ( .A1(n12647), .A2(n15214), .ZN(n15226) );
  AOI21_X1 U15027 ( .B1(n15214), .B2(n12647), .A(n15226), .ZN(n15209) );
  NAND2_X1 U15028 ( .A1(n15210), .A2(n15209), .ZN(n15225) );
  INV_X1 U15029 ( .A(n15226), .ZN(n12648) );
  XNOR2_X1 U15030 ( .A(n12649), .B(n12668), .ZN(n15229) );
  NAND3_X1 U15031 ( .A1(n15225), .A2(n12648), .A3(n15229), .ZN(n15228) );
  OAI21_X1 U15032 ( .B1(n12649), .B2(n15234), .A(n15228), .ZN(n15254) );
  AND2_X1 U15033 ( .A1(n15248), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12670) );
  INV_X1 U15034 ( .A(n12670), .ZN(n12650) );
  OAI21_X1 U15035 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n15248), .A(n12650), 
        .ZN(n15246) );
  MUX2_X1 U15036 ( .A(n15260), .B(n15246), .S(n12651), .Z(n15255) );
  MUX2_X1 U15037 ( .A(n12670), .B(n12652), .S(n12735), .Z(n12653) );
  NOR2_X1 U15038 ( .A1(n15252), .A2(n12653), .ZN(n12654) );
  XNOR2_X1 U15039 ( .A(n12654), .B(n14626), .ZN(n14621) );
  MUX2_X1 U15040 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12735), .Z(n14622) );
  NOR2_X1 U15041 ( .A1(n14621), .A2(n14622), .ZN(n14620) );
  AOI21_X1 U15042 ( .B1(n12654), .B2(n14626), .A(n14620), .ZN(n12686) );
  XOR2_X1 U15043 ( .A(n12655), .B(n12686), .Z(n12679) );
  NAND2_X1 U15044 ( .A1(n15232), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n12656) );
  OAI211_X1 U15045 ( .C1(n15235), .C2(n12692), .A(n12657), .B(n12656), .ZN(
        n12678) );
  NOR2_X1 U15046 ( .A1(n12660), .A2(n12661), .ZN(n12662) );
  NAND2_X1 U15047 ( .A1(n12663), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12666) );
  NAND2_X1 U15048 ( .A1(n15214), .A2(n12664), .ZN(n12665) );
  NAND2_X1 U15049 ( .A1(n12666), .A2(n12665), .ZN(n15205) );
  NOR2_X1 U15050 ( .A1(n12668), .A2(n12667), .ZN(n12669) );
  NOR2_X1 U15051 ( .A1(n14626), .A2(n12671), .ZN(n12672) );
  XNOR2_X1 U15052 ( .A(n12673), .B(n12927), .ZN(n12674) );
  OR2_X2 U15053 ( .A1(n12675), .A2(n12674), .ZN(n12694) );
  NAND2_X1 U15054 ( .A1(n12675), .A2(n12674), .ZN(n12676) );
  AOI21_X1 U15055 ( .B1(n12694), .B2(n12676), .A(n15266), .ZN(n12677) );
  AOI211_X1 U15056 ( .C1(n15237), .C2(n12679), .A(n12678), .B(n12677), .ZN(
        n12680) );
  OAI21_X1 U15057 ( .B1(n12681), .B2(n15241), .A(n12680), .ZN(P3_U3198) );
  NAND2_X1 U15058 ( .A1(n12692), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12682) );
  AOI21_X1 U15059 ( .B1(n13010), .B2(n12684), .A(n12716), .ZN(n12700) );
  MUX2_X1 U15060 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12735), .Z(n12708) );
  XNOR2_X1 U15061 ( .A(n12708), .B(n12718), .ZN(n12687) );
  NOR2_X1 U15062 ( .A1(n12707), .A2(n15253), .ZN(n12699) );
  OAI21_X1 U15063 ( .B1(n12689), .B2(n12688), .A(n12687), .ZN(n12698) );
  NAND2_X1 U15064 ( .A1(n15232), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12690) );
  OAI211_X1 U15065 ( .C1(n15235), .C2(n12718), .A(n12691), .B(n12690), .ZN(
        n12697) );
  NAND2_X1 U15066 ( .A1(n12692), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12693) );
  AOI21_X1 U15067 ( .B1(n12695), .B2(n12915), .A(n12701), .ZN(n12696) );
  NAND2_X1 U15068 ( .A1(n12719), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12726) );
  OAI21_X1 U15069 ( .B1(n12719), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12726), 
        .ZN(n12703) );
  AOI21_X1 U15070 ( .B1(n12704), .B2(n12703), .A(n12728), .ZN(n12725) );
  INV_X1 U15071 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12706) );
  OAI21_X1 U15072 ( .B1(n15251), .B2(n12706), .A(n12705), .ZN(n12714) );
  AOI21_X1 U15073 ( .B1(n12708), .B2(n12718), .A(n12707), .ZN(n12709) );
  NAND2_X1 U15074 ( .A1(n12709), .A2(n12715), .ZN(n12732) );
  OAI21_X1 U15075 ( .B1(n12709), .B2(n12715), .A(n12732), .ZN(n12711) );
  MUX2_X1 U15076 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12735), .Z(n12710) );
  NOR2_X1 U15077 ( .A1(n12711), .A2(n12710), .ZN(n12734) );
  AOI21_X1 U15078 ( .B1(n12711), .B2(n12710), .A(n12734), .ZN(n12712) );
  NOR2_X1 U15079 ( .A1(n12712), .A2(n15253), .ZN(n12713) );
  AOI211_X1 U15080 ( .C1(n15259), .C2(n12715), .A(n12714), .B(n12713), .ZN(
        n12724) );
  NAND2_X1 U15081 ( .A1(n12719), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12743) );
  OAI21_X1 U15082 ( .B1(n12719), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12743), 
        .ZN(n12720) );
  OAI21_X1 U15083 ( .B1(n12745), .B2(n12722), .A(n15262), .ZN(n12723) );
  OAI211_X1 U15084 ( .C1(n12725), .C2(n15266), .A(n12724), .B(n12723), .ZN(
        P3_U3200) );
  INV_X1 U15085 ( .A(n12726), .ZN(n12727) );
  NOR2_X1 U15086 ( .A1(n12728), .A2(n12727), .ZN(n12729) );
  XNOR2_X1 U15087 ( .A(n12742), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12736) );
  XNOR2_X1 U15088 ( .A(n12729), .B(n12736), .ZN(n12749) );
  OAI21_X1 U15089 ( .B1(n15251), .B2(n12731), .A(n12730), .ZN(n12741) );
  INV_X1 U15090 ( .A(n12732), .ZN(n12733) );
  NOR2_X1 U15091 ( .A1(n12734), .A2(n12733), .ZN(n12738) );
  XNOR2_X1 U15092 ( .A(n12742), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12746) );
  MUX2_X1 U15093 ( .A(n12736), .B(n12746), .S(n6684), .Z(n12737) );
  XNOR2_X1 U15094 ( .A(n12738), .B(n12737), .ZN(n12739) );
  NOR2_X1 U15095 ( .A1(n12739), .A2(n15253), .ZN(n12740) );
  INV_X1 U15096 ( .A(n12743), .ZN(n12744) );
  OAI211_X1 U15097 ( .C1(n12749), .C2(n15266), .A(n12748), .B(n12747), .ZN(
        P3_U3201) );
  INV_X1 U15098 ( .A(n12750), .ZN(n12751) );
  NAND2_X1 U15099 ( .A1(n12752), .A2(n12751), .ZN(n13025) );
  AOI21_X1 U15100 ( .B1(n13025), .B2(n12753), .A(n15337), .ZN(n12755) );
  AOI21_X1 U15101 ( .B1(n15337), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12755), 
        .ZN(n12754) );
  OAI21_X1 U15102 ( .B1(n13027), .B2(n14652), .A(n12754), .ZN(P3_U3202) );
  AOI21_X1 U15103 ( .B1(n15337), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12755), 
        .ZN(n12756) );
  OAI21_X1 U15104 ( .B1(n12757), .B2(n14652), .A(n12756), .ZN(P3_U3203) );
  INV_X1 U15105 ( .A(n12779), .ZN(n12759) );
  NAND2_X1 U15106 ( .A1(n12759), .A2(n12758), .ZN(n12760) );
  INV_X1 U15107 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12772) );
  NAND2_X1 U15108 ( .A1(n12780), .A2(n12761), .ZN(n12763) );
  NAND2_X1 U15109 ( .A1(n12763), .A2(n6990), .ZN(n12765) );
  NAND3_X1 U15110 ( .A1(n12765), .A2(n15322), .A3(n12764), .ZN(n12770) );
  OAI22_X1 U15111 ( .A1(n12767), .A2(n15315), .B1(n12766), .B2(n15313), .ZN(
        n12768) );
  INV_X1 U15112 ( .A(n12768), .ZN(n12769) );
  NAND2_X1 U15113 ( .A1(n12770), .A2(n12769), .ZN(n13033) );
  INV_X1 U15114 ( .A(n13033), .ZN(n12771) );
  MUX2_X1 U15115 ( .A(n12772), .B(n12771), .S(n15335), .Z(n12775) );
  AOI22_X1 U15116 ( .A1(n13035), .A2(n12953), .B1(n15332), .B2(n12773), .ZN(
        n12774) );
  OAI211_X1 U15117 ( .C1(n13037), .C2(n12957), .A(n12775), .B(n12774), .ZN(
        P3_U3205) );
  NOR2_X1 U15118 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  INV_X1 U15119 ( .A(n12973), .ZN(n12786) );
  OAI21_X1 U15120 ( .B1(n7755), .B2(n8895), .A(n12780), .ZN(n12784) );
  OAI22_X1 U15121 ( .A1(n12782), .A2(n15315), .B1(n12781), .B2(n15313), .ZN(
        n12783) );
  AOI21_X1 U15122 ( .B1(n12784), .B2(n15322), .A(n12783), .ZN(n12785) );
  INV_X1 U15123 ( .A(n12972), .ZN(n12792) );
  INV_X1 U15124 ( .A(n12787), .ZN(n13041) );
  AOI22_X1 U15125 ( .A1(n12788), .A2(n15332), .B1(n15337), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12789) );
  OAI21_X1 U15126 ( .B1(n13041), .B2(n14652), .A(n12789), .ZN(n12790) );
  AOI21_X1 U15127 ( .B1(n12973), .B2(n15333), .A(n12790), .ZN(n12791) );
  OAI21_X1 U15128 ( .B1(n12792), .B2(n15337), .A(n12791), .ZN(P3_U3206) );
  INV_X1 U15129 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12798) );
  XNOR2_X1 U15130 ( .A(n12795), .B(n12794), .ZN(n12797) );
  MUX2_X1 U15131 ( .A(n12798), .B(n13042), .S(n15335), .Z(n12801) );
  AOI22_X1 U15132 ( .A1(n13044), .A2(n12953), .B1(n15332), .B2(n12799), .ZN(
        n12800) );
  OAI211_X1 U15133 ( .C1(n13047), .C2(n12957), .A(n12801), .B(n12800), .ZN(
        P3_U3207) );
  INV_X1 U15134 ( .A(n12802), .ZN(n12806) );
  INV_X1 U15135 ( .A(n12804), .ZN(n12807) );
  OAI211_X1 U15136 ( .C1(n12807), .C2(n12806), .A(n12805), .B(n15322), .ZN(
        n12809) );
  OAI211_X1 U15137 ( .C1(n15289), .C2(n12979), .A(n12809), .B(n12808), .ZN(
        n12980) );
  AOI22_X1 U15138 ( .A1(n12810), .A2(n15332), .B1(n15337), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U15139 ( .A1(n12811), .A2(n12953), .ZN(n12812) );
  OAI211_X1 U15140 ( .C1(n12979), .C2(n12840), .A(n12813), .B(n12812), .ZN(
        n12814) );
  AOI21_X1 U15141 ( .B1(n12980), .B2(n15335), .A(n12814), .ZN(n12815) );
  INV_X1 U15142 ( .A(n12815), .ZN(P3_U3208) );
  INV_X1 U15143 ( .A(n12816), .ZN(n12817) );
  AOI21_X1 U15144 ( .B1(n12818), .B2(n12820), .A(n12817), .ZN(n13057) );
  INV_X1 U15145 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12823) );
  XOR2_X1 U15146 ( .A(n12820), .B(n12819), .Z(n12822) );
  AOI222_X1 U15147 ( .A1(n15322), .A2(n12822), .B1(n12846), .B2(n12946), .C1(
        n12821), .C2(n12948), .ZN(n13052) );
  MUX2_X1 U15148 ( .A(n12823), .B(n13052), .S(n15335), .Z(n12826) );
  AOI22_X1 U15149 ( .A1(n13054), .A2(n12953), .B1(n15332), .B2(n12824), .ZN(
        n12825) );
  OAI211_X1 U15150 ( .C1(n13057), .C2(n12957), .A(n12826), .B(n12825), .ZN(
        P3_U3209) );
  OR2_X1 U15151 ( .A1(n12827), .A2(n12830), .ZN(n12828) );
  NAND2_X1 U15152 ( .A1(n12829), .A2(n12828), .ZN(n12988) );
  XNOR2_X1 U15153 ( .A(n12831), .B(n12830), .ZN(n12835) );
  OAI22_X1 U15154 ( .A1(n12833), .A2(n15315), .B1(n12832), .B2(n15313), .ZN(
        n12834) );
  AOI21_X1 U15155 ( .B1(n12835), .B2(n15322), .A(n12834), .ZN(n12836) );
  OAI21_X1 U15156 ( .B1(n15289), .B2(n12988), .A(n12836), .ZN(n12989) );
  AOI22_X1 U15157 ( .A1(n12837), .A2(n15332), .B1(P3_REG2_REG_23__SCAN_IN), 
        .B2(n15337), .ZN(n12839) );
  NAND2_X1 U15158 ( .A1(n12987), .A2(n12953), .ZN(n12838) );
  OAI211_X1 U15159 ( .C1(n12988), .C2(n12840), .A(n12839), .B(n12838), .ZN(
        n12841) );
  AOI21_X1 U15160 ( .B1(n12989), .B2(n15335), .A(n12841), .ZN(n12842) );
  INV_X1 U15161 ( .A(n12842), .ZN(P3_U3210) );
  XNOR2_X1 U15162 ( .A(n12843), .B(n12845), .ZN(n13065) );
  INV_X1 U15163 ( .A(n13065), .ZN(n12852) );
  INV_X1 U15164 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12848) );
  XNOR2_X1 U15165 ( .A(n12844), .B(n12845), .ZN(n12847) );
  AOI222_X1 U15166 ( .A1(n15322), .A2(n12847), .B1(n12846), .B2(n12948), .C1(
        n12869), .C2(n12946), .ZN(n13062) );
  MUX2_X1 U15167 ( .A(n12848), .B(n13062), .S(n15335), .Z(n12851) );
  AOI22_X1 U15168 ( .A1(n13064), .A2(n12953), .B1(n15332), .B2(n12849), .ZN(
        n12850) );
  OAI211_X1 U15169 ( .C1(n12852), .C2(n12957), .A(n12851), .B(n12850), .ZN(
        P3_U3211) );
  XNOR2_X1 U15170 ( .A(n12854), .B(n12853), .ZN(n13073) );
  INV_X1 U15171 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12863) );
  INV_X1 U15172 ( .A(n12855), .ZN(n12860) );
  AOI21_X1 U15173 ( .B1(n12856), .B2(n12858), .A(n12857), .ZN(n12859) );
  OAI21_X1 U15174 ( .B1(n12860), .B2(n12859), .A(n15322), .ZN(n12862) );
  MUX2_X1 U15175 ( .A(n12863), .B(n13068), .S(n15335), .Z(n12866) );
  AOI22_X1 U15176 ( .A1(n13070), .A2(n12953), .B1(n15332), .B2(n12864), .ZN(
        n12865) );
  OAI211_X1 U15177 ( .C1(n13073), .C2(n12957), .A(n12866), .B(n12865), .ZN(
        P3_U3212) );
  OAI211_X1 U15178 ( .C1(n12877), .C2(n12867), .A(n12856), .B(n15322), .ZN(
        n12871) );
  AOI22_X1 U15179 ( .A1(n12869), .A2(n12948), .B1(n12946), .B2(n12868), .ZN(
        n12870) );
  INV_X1 U15180 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12874) );
  INV_X1 U15181 ( .A(n12872), .ZN(n12873) );
  OAI22_X1 U15182 ( .A1(n15335), .A2(n12874), .B1(n12873), .B2(n15307), .ZN(
        n12875) );
  AOI21_X1 U15183 ( .B1(n12876), .B2(n12953), .A(n12875), .ZN(n12880) );
  NAND2_X1 U15184 ( .A1(n12878), .A2(n12877), .ZN(n12999) );
  NAND3_X1 U15185 ( .A1(n13000), .A2(n12999), .A3(n12893), .ZN(n12879) );
  OAI211_X1 U15186 ( .C1(n13002), .C2(n15337), .A(n12880), .B(n12879), .ZN(
        P3_U3213) );
  INV_X1 U15187 ( .A(n12881), .ZN(n12885) );
  AOI21_X1 U15188 ( .B1(n12882), .B2(n12883), .A(n12889), .ZN(n12884) );
  NOR3_X1 U15189 ( .A1(n12885), .A2(n12884), .A3(n15311), .ZN(n12887) );
  NOR2_X1 U15190 ( .A1(n12887), .A2(n12886), .ZN(n13075) );
  MUX2_X1 U15191 ( .A(n12888), .B(n13075), .S(n15335), .Z(n12895) );
  XNOR2_X1 U15192 ( .A(n12890), .B(n12889), .ZN(n13077) );
  OAI22_X1 U15193 ( .A1(n13080), .A2(n14652), .B1(n12891), .B2(n15307), .ZN(
        n12892) );
  AOI21_X1 U15194 ( .B1(n13077), .B2(n12893), .A(n12892), .ZN(n12894) );
  NAND2_X1 U15195 ( .A1(n12895), .A2(n12894), .ZN(P3_U3214) );
  XOR2_X1 U15196 ( .A(n12896), .B(n12898), .Z(n13084) );
  INV_X1 U15197 ( .A(n13084), .ZN(n12906) );
  AND2_X1 U15198 ( .A1(n12909), .A2(n12897), .ZN(n12899) );
  OAI21_X1 U15199 ( .B1(n12899), .B2(n12898), .A(n12882), .ZN(n12901) );
  AOI21_X1 U15200 ( .B1(n12901), .B2(n15322), .A(n12900), .ZN(n13081) );
  MUX2_X1 U15201 ( .A(n12902), .B(n13081), .S(n15335), .Z(n12905) );
  AOI22_X1 U15202 ( .A1(n13083), .A2(n12953), .B1(n15332), .B2(n12903), .ZN(
        n12904) );
  OAI211_X1 U15203 ( .C1(n12906), .C2(n12957), .A(n12905), .B(n12904), .ZN(
        P3_U3215) );
  XNOR2_X1 U15204 ( .A(n12908), .B(n12907), .ZN(n13090) );
  INV_X1 U15205 ( .A(n13090), .ZN(n12919) );
  OAI211_X1 U15206 ( .C1(n12911), .C2(n12910), .A(n12909), .B(n15322), .ZN(
        n12914) );
  AOI22_X1 U15207 ( .A1(n12946), .A2(n12937), .B1(n12912), .B2(n12948), .ZN(
        n12913) );
  MUX2_X1 U15208 ( .A(n13088), .B(n12915), .S(n15337), .Z(n12918) );
  AOI22_X1 U15209 ( .A1(n13089), .A2(n12953), .B1(n12916), .B2(n15332), .ZN(
        n12917) );
  OAI211_X1 U15210 ( .C1(n12919), .C2(n12957), .A(n12918), .B(n12917), .ZN(
        P3_U3216) );
  OAI21_X1 U15211 ( .B1(n12922), .B2(n12921), .A(n12920), .ZN(n13096) );
  INV_X1 U15212 ( .A(n13096), .ZN(n12932) );
  XNOR2_X1 U15213 ( .A(n12924), .B(n12923), .ZN(n12926) );
  AOI21_X1 U15214 ( .B1(n12926), .B2(n15322), .A(n12925), .ZN(n13093) );
  MUX2_X1 U15215 ( .A(n12927), .B(n13093), .S(n15335), .Z(n12931) );
  INV_X1 U15216 ( .A(n12928), .ZN(n12929) );
  AOI22_X1 U15217 ( .A1(n13095), .A2(n12953), .B1(n15332), .B2(n12929), .ZN(
        n12930) );
  OAI211_X1 U15218 ( .C1(n12932), .C2(n12957), .A(n12931), .B(n12930), .ZN(
        P3_U3217) );
  XOR2_X1 U15219 ( .A(n12934), .B(n12933), .Z(n13106) );
  XNOR2_X1 U15220 ( .A(n12935), .B(n12934), .ZN(n12938) );
  AOI222_X1 U15221 ( .A1(n15322), .A2(n12938), .B1(n12937), .B2(n12948), .C1(
        n12936), .C2(n12946), .ZN(n13099) );
  MUX2_X1 U15222 ( .A(n14616), .B(n13099), .S(n15335), .Z(n12941) );
  AOI22_X1 U15223 ( .A1(n13102), .A2(n12953), .B1(n15332), .B2(n12939), .ZN(
        n12940) );
  OAI211_X1 U15224 ( .C1(n13106), .C2(n12957), .A(n12941), .B(n12940), .ZN(
        P3_U3218) );
  XNOR2_X1 U15225 ( .A(n12943), .B(n12942), .ZN(n13110) );
  INV_X1 U15226 ( .A(n13110), .ZN(n12958) );
  INV_X1 U15227 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12951) );
  XNOR2_X1 U15228 ( .A(n12945), .B(n12944), .ZN(n12950) );
  AOI222_X1 U15229 ( .A1(n15322), .A2(n12950), .B1(n12949), .B2(n12948), .C1(
        n12947), .C2(n12946), .ZN(n13107) );
  MUX2_X1 U15230 ( .A(n12951), .B(n13107), .S(n15335), .Z(n12956) );
  INV_X1 U15231 ( .A(n13113), .ZN(n12954) );
  AOI22_X1 U15232 ( .A1(n12954), .A2(n12953), .B1(n15332), .B2(n12952), .ZN(
        n12955) );
  OAI211_X1 U15233 ( .C1(n12958), .C2(n12957), .A(n12956), .B(n12955), .ZN(
        P3_U3219) );
  NOR2_X1 U15234 ( .A1(n13025), .A2(n15394), .ZN(n12960) );
  AOI21_X1 U15235 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15394), .A(n12960), 
        .ZN(n12959) );
  OAI21_X1 U15236 ( .B1(n13027), .B2(n13024), .A(n12959), .ZN(P3_U3490) );
  NAND2_X1 U15237 ( .A1(n13028), .A2(n13016), .ZN(n12962) );
  INV_X1 U15238 ( .A(n12960), .ZN(n12961) );
  OAI211_X1 U15239 ( .C1(n15396), .C2(n8923), .A(n12962), .B(n12961), .ZN(
        P3_U3489) );
  AOI22_X1 U15240 ( .A1(n12966), .A2(n13021), .B1(n13016), .B2(n12965), .ZN(
        n12967) );
  NAND2_X1 U15241 ( .A1(n12968), .A2(n12967), .ZN(P3_U3488) );
  MUX2_X1 U15242 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13033), .S(n15396), .Z(
        n12969) );
  AOI21_X1 U15243 ( .B1(n13016), .B2(n13035), .A(n12969), .ZN(n12970) );
  OAI21_X1 U15244 ( .B1(n13019), .B2(n13037), .A(n12970), .ZN(P3_U3487) );
  AOI21_X1 U15245 ( .B1(n15380), .B2(n12973), .A(n12972), .ZN(n13038) );
  MUX2_X1 U15246 ( .A(n12974), .B(n13038), .S(n15396), .Z(n12975) );
  OAI21_X1 U15247 ( .B1(n13041), .B2(n13024), .A(n12975), .ZN(P3_U3486) );
  MUX2_X1 U15248 ( .A(n12976), .B(n13042), .S(n15396), .Z(n12978) );
  NAND2_X1 U15249 ( .A1(n13044), .A2(n13016), .ZN(n12977) );
  OAI211_X1 U15250 ( .C1(n13019), .C2(n13047), .A(n12978), .B(n12977), .ZN(
        P3_U3485) );
  INV_X1 U15251 ( .A(n12979), .ZN(n12981) );
  AOI21_X1 U15252 ( .B1(n15380), .B2(n12981), .A(n12980), .ZN(n13048) );
  MUX2_X1 U15253 ( .A(n12982), .B(n13048), .S(n15396), .Z(n12983) );
  OAI21_X1 U15254 ( .B1(n13051), .B2(n13024), .A(n12983), .ZN(P3_U3484) );
  MUX2_X1 U15255 ( .A(n12984), .B(n13052), .S(n15396), .Z(n12986) );
  NAND2_X1 U15256 ( .A1(n13054), .A2(n13016), .ZN(n12985) );
  OAI211_X1 U15257 ( .C1(n13057), .C2(n13019), .A(n12986), .B(n12985), .ZN(
        P3_U3483) );
  INV_X1 U15258 ( .A(n12987), .ZN(n13061) );
  INV_X1 U15259 ( .A(n12988), .ZN(n12990) );
  AOI21_X1 U15260 ( .B1(n15380), .B2(n12990), .A(n12989), .ZN(n13058) );
  MUX2_X1 U15261 ( .A(n12991), .B(n13058), .S(n15396), .Z(n12992) );
  OAI21_X1 U15262 ( .B1(n13061), .B2(n13024), .A(n12992), .ZN(P3_U3482) );
  INV_X1 U15263 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12993) );
  MUX2_X1 U15264 ( .A(n12993), .B(n13062), .S(n15396), .Z(n12995) );
  AOI22_X1 U15265 ( .A1(n13065), .A2(n13021), .B1(n13016), .B2(n13064), .ZN(
        n12994) );
  NAND2_X1 U15266 ( .A1(n12995), .A2(n12994), .ZN(P3_U3481) );
  INV_X1 U15267 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12996) );
  MUX2_X1 U15268 ( .A(n12996), .B(n13068), .S(n15396), .Z(n12998) );
  NAND2_X1 U15269 ( .A1(n13070), .A2(n13016), .ZN(n12997) );
  OAI211_X1 U15270 ( .C1(n13073), .C2(n13019), .A(n12998), .B(n12997), .ZN(
        P3_U3480) );
  NAND3_X1 U15271 ( .A1(n13000), .A2(n15368), .A3(n12999), .ZN(n13001) );
  OAI211_X1 U15272 ( .C1(n13003), .C2(n15339), .A(n13002), .B(n13001), .ZN(
        n13074) );
  MUX2_X1 U15273 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13074), .S(n15396), .Z(
        P3_U3479) );
  MUX2_X1 U15274 ( .A(n13004), .B(n13075), .S(n15396), .Z(n13006) );
  NAND2_X1 U15275 ( .A1(n13077), .A2(n13021), .ZN(n13005) );
  OAI211_X1 U15276 ( .C1(n13024), .C2(n13080), .A(n13006), .B(n13005), .ZN(
        P3_U3478) );
  MUX2_X1 U15277 ( .A(n13007), .B(n13081), .S(n15396), .Z(n13009) );
  AOI22_X1 U15278 ( .A1(n13084), .A2(n13021), .B1(n13016), .B2(n13083), .ZN(
        n13008) );
  NAND2_X1 U15279 ( .A1(n13009), .A2(n13008), .ZN(P3_U3477) );
  MUX2_X1 U15280 ( .A(n13088), .B(n13010), .S(n15394), .Z(n13012) );
  AOI22_X1 U15281 ( .A1(n13090), .A2(n13021), .B1(n13016), .B2(n13089), .ZN(
        n13011) );
  NAND2_X1 U15282 ( .A1(n13012), .A2(n13011), .ZN(P3_U3476) );
  MUX2_X1 U15283 ( .A(n13013), .B(n13093), .S(n15396), .Z(n13015) );
  AOI22_X1 U15284 ( .A1(n13096), .A2(n13021), .B1(n13016), .B2(n13095), .ZN(
        n13014) );
  NAND2_X1 U15285 ( .A1(n13015), .A2(n13014), .ZN(P3_U3475) );
  MUX2_X1 U15286 ( .A(n14628), .B(n13099), .S(n15396), .Z(n13018) );
  NAND2_X1 U15287 ( .A1(n13102), .A2(n13016), .ZN(n13017) );
  OAI211_X1 U15288 ( .C1(n13019), .C2(n13106), .A(n13018), .B(n13017), .ZN(
        P3_U3474) );
  MUX2_X1 U15289 ( .A(n13020), .B(n13107), .S(n15396), .Z(n13023) );
  NAND2_X1 U15290 ( .A1(n13110), .A2(n13021), .ZN(n13022) );
  OAI211_X1 U15291 ( .C1(n13024), .C2(n13113), .A(n13023), .B(n13022), .ZN(
        P3_U3473) );
  NOR2_X1 U15292 ( .A1(n13025), .A2(n9009), .ZN(n13029) );
  AOI21_X1 U15293 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n9009), .A(n13029), .ZN(
        n13026) );
  OAI21_X1 U15294 ( .B1(n13027), .B2(n13114), .A(n13026), .ZN(P3_U3458) );
  INV_X1 U15295 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13032) );
  NAND2_X1 U15296 ( .A1(n13028), .A2(n13101), .ZN(n13031) );
  INV_X1 U15297 ( .A(n13029), .ZN(n13030) );
  OAI211_X1 U15298 ( .C1(n15382), .C2(n13032), .A(n13031), .B(n13030), .ZN(
        P3_U3457) );
  MUX2_X1 U15299 ( .A(n13033), .B(P3_REG0_REG_28__SCAN_IN), .S(n9009), .Z(
        n13034) );
  AOI21_X1 U15300 ( .B1(n13101), .B2(n13035), .A(n13034), .ZN(n13036) );
  OAI21_X1 U15301 ( .B1(n13105), .B2(n13037), .A(n13036), .ZN(P3_U3455) );
  INV_X1 U15302 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13039) );
  MUX2_X1 U15303 ( .A(n13039), .B(n13038), .S(n15382), .Z(n13040) );
  OAI21_X1 U15304 ( .B1(n13041), .B2(n13114), .A(n13040), .ZN(P3_U3454) );
  INV_X1 U15305 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13043) );
  MUX2_X1 U15306 ( .A(n13043), .B(n13042), .S(n15382), .Z(n13046) );
  NAND2_X1 U15307 ( .A1(n13044), .A2(n13101), .ZN(n13045) );
  OAI211_X1 U15308 ( .C1(n13047), .C2(n13105), .A(n13046), .B(n13045), .ZN(
        P3_U3453) );
  INV_X1 U15309 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13049) );
  MUX2_X1 U15310 ( .A(n13049), .B(n13048), .S(n15382), .Z(n13050) );
  OAI21_X1 U15311 ( .B1(n13051), .B2(n13114), .A(n13050), .ZN(P3_U3452) );
  INV_X1 U15312 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13053) );
  MUX2_X1 U15313 ( .A(n13053), .B(n13052), .S(n15382), .Z(n13056) );
  NAND2_X1 U15314 ( .A1(n13054), .A2(n13101), .ZN(n13055) );
  OAI211_X1 U15315 ( .C1(n13057), .C2(n13105), .A(n13056), .B(n13055), .ZN(
        P3_U3451) );
  INV_X1 U15316 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13059) );
  MUX2_X1 U15317 ( .A(n13059), .B(n13058), .S(n15382), .Z(n13060) );
  OAI21_X1 U15318 ( .B1(n13061), .B2(n13114), .A(n13060), .ZN(P3_U3450) );
  MUX2_X1 U15319 ( .A(n13063), .B(n13062), .S(n15382), .Z(n13067) );
  AOI22_X1 U15320 ( .A1(n13065), .A2(n13109), .B1(n13101), .B2(n13064), .ZN(
        n13066) );
  NAND2_X1 U15321 ( .A1(n13067), .A2(n13066), .ZN(P3_U3449) );
  INV_X1 U15322 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13069) );
  MUX2_X1 U15323 ( .A(n13069), .B(n13068), .S(n15382), .Z(n13072) );
  NAND2_X1 U15324 ( .A1(n13070), .A2(n13101), .ZN(n13071) );
  OAI211_X1 U15325 ( .C1(n13073), .C2(n13105), .A(n13072), .B(n13071), .ZN(
        P3_U3448) );
  MUX2_X1 U15326 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13074), .S(n15382), .Z(
        P3_U3447) );
  MUX2_X1 U15327 ( .A(n13076), .B(n13075), .S(n15382), .Z(n13079) );
  NAND2_X1 U15328 ( .A1(n13077), .A2(n13109), .ZN(n13078) );
  OAI211_X1 U15329 ( .C1(n13114), .C2(n13080), .A(n13079), .B(n13078), .ZN(
        P3_U3446) );
  INV_X1 U15330 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13082) );
  MUX2_X1 U15331 ( .A(n13082), .B(n13081), .S(n15382), .Z(n13086) );
  AOI22_X1 U15332 ( .A1(n13084), .A2(n13109), .B1(n13101), .B2(n13083), .ZN(
        n13085) );
  NAND2_X1 U15333 ( .A1(n13086), .A2(n13085), .ZN(P3_U3444) );
  INV_X1 U15334 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13087) );
  MUX2_X1 U15335 ( .A(n13088), .B(n13087), .S(n9009), .Z(n13092) );
  AOI22_X1 U15336 ( .A1(n13090), .A2(n13109), .B1(n13101), .B2(n13089), .ZN(
        n13091) );
  NAND2_X1 U15337 ( .A1(n13092), .A2(n13091), .ZN(P3_U3441) );
  INV_X1 U15338 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13094) );
  MUX2_X1 U15339 ( .A(n13094), .B(n13093), .S(n15382), .Z(n13098) );
  AOI22_X1 U15340 ( .A1(n13096), .A2(n13109), .B1(n13101), .B2(n13095), .ZN(
        n13097) );
  NAND2_X1 U15341 ( .A1(n13098), .A2(n13097), .ZN(P3_U3438) );
  INV_X1 U15342 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13100) );
  MUX2_X1 U15343 ( .A(n13100), .B(n13099), .S(n15382), .Z(n13104) );
  NAND2_X1 U15344 ( .A1(n13102), .A2(n13101), .ZN(n13103) );
  OAI211_X1 U15345 ( .C1(n13106), .C2(n13105), .A(n13104), .B(n13103), .ZN(
        P3_U3435) );
  MUX2_X1 U15346 ( .A(n13108), .B(n13107), .S(n15382), .Z(n13112) );
  NAND2_X1 U15347 ( .A1(n13110), .A2(n13109), .ZN(n13111) );
  OAI211_X1 U15348 ( .C1(n13114), .C2(n13113), .A(n13112), .B(n13111), .ZN(
        P3_U3432) );
  MUX2_X1 U15349 ( .A(P3_D_REG_0__SCAN_IN), .B(n13116), .S(n13115), .Z(
        P3_U3376) );
  NAND3_X1 U15350 ( .A1(n13117), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13120) );
  OAI22_X1 U15351 ( .A1(n13121), .A2(n13120), .B1(n13119), .B2(n13130), .ZN(
        n13122) );
  AOI21_X1 U15352 ( .B1(n13124), .B2(n13123), .A(n13122), .ZN(n13125) );
  INV_X1 U15353 ( .A(n13125), .ZN(P3_U3264) );
  INV_X1 U15354 ( .A(n13126), .ZN(n13128) );
  OAI222_X1 U15355 ( .A1(n13130), .A2(n13129), .B1(n11825), .B2(n13128), .C1(
        P3_U3151), .C2(n13127), .ZN(P3_U3266) );
  INV_X1 U15356 ( .A(n13131), .ZN(n13133) );
  NAND2_X1 U15357 ( .A1(n13133), .A2(n13132), .ZN(n13134) );
  XNOR2_X1 U15358 ( .A(n13355), .B(n13226), .ZN(n13139) );
  INV_X1 U15359 ( .A(n13139), .ZN(n13136) );
  XNOR2_X1 U15360 ( .A(n13138), .B(n13136), .ZN(n13345) );
  NOR2_X1 U15361 ( .A1(n13137), .A2(n10749), .ZN(n13344) );
  NAND2_X1 U15362 ( .A1(n13345), .A2(n13344), .ZN(n13341) );
  XNOR2_X1 U15363 ( .A(n13452), .B(n13226), .ZN(n13141) );
  NAND2_X1 U15364 ( .A1(n13359), .A2(n13191), .ZN(n13142) );
  XNOR2_X1 U15365 ( .A(n13141), .B(n13142), .ZN(n13252) );
  INV_X1 U15366 ( .A(n13141), .ZN(n13144) );
  INV_X1 U15367 ( .A(n13142), .ZN(n13143) );
  NOR2_X1 U15368 ( .A1(n13144), .A2(n13143), .ZN(n13272) );
  XNOR2_X1 U15369 ( .A(n13810), .B(n13226), .ZN(n13147) );
  NOR2_X1 U15370 ( .A1(n13455), .A2(n10749), .ZN(n13145) );
  XNOR2_X1 U15371 ( .A(n13147), .B(n13145), .ZN(n13271) );
  INV_X1 U15372 ( .A(n13145), .ZN(n13146) );
  INV_X1 U15373 ( .A(n13319), .ZN(n13151) );
  XNOR2_X1 U15374 ( .A(n13656), .B(n13186), .ZN(n13149) );
  NOR2_X1 U15375 ( .A1(n13457), .A2(n10749), .ZN(n13148) );
  NAND2_X1 U15376 ( .A1(n13149), .A2(n13148), .ZN(n13152) );
  OAI21_X1 U15377 ( .B1(n13149), .B2(n13148), .A(n13152), .ZN(n13318) );
  INV_X1 U15378 ( .A(n13318), .ZN(n13150) );
  XNOR2_X1 U15379 ( .A(n13804), .B(n13226), .ZN(n13156) );
  NAND2_X1 U15380 ( .A1(n13428), .A2(n13191), .ZN(n13155) );
  XNOR2_X1 U15381 ( .A(n13156), .B(n13155), .ZN(n13217) );
  NAND2_X1 U15382 ( .A1(n13156), .A2(n13155), .ZN(n13300) );
  XNOR2_X1 U15383 ( .A(n13617), .B(n13226), .ZN(n13160) );
  NOR2_X1 U15384 ( .A1(n13462), .A2(n10749), .ZN(n13158) );
  XNOR2_X1 U15385 ( .A(n13160), .B(n13158), .ZN(n13301) );
  INV_X1 U15386 ( .A(n13171), .ZN(n13302) );
  XNOR2_X1 U15387 ( .A(n13730), .B(n13186), .ZN(n13166) );
  XNOR2_X1 U15388 ( .A(n13799), .B(n13226), .ZN(n13173) );
  INV_X1 U15389 ( .A(n13173), .ZN(n13157) );
  INV_X1 U15390 ( .A(n13465), .ZN(n13432) );
  NAND2_X1 U15391 ( .A1(n13432), .A2(n13191), .ZN(n13161) );
  INV_X1 U15392 ( .A(n13161), .ZN(n13172) );
  NAND2_X1 U15393 ( .A1(n13157), .A2(n13172), .ZN(n13174) );
  INV_X1 U15394 ( .A(n13158), .ZN(n13159) );
  AND2_X1 U15395 ( .A1(n13160), .A2(n13159), .ZN(n13162) );
  AOI211_X1 U15396 ( .C1(n13173), .C2(n13161), .A(n13166), .B(n13162), .ZN(
        n13168) );
  INV_X1 U15397 ( .A(n13166), .ZN(n13175) );
  INV_X1 U15398 ( .A(n13162), .ZN(n13170) );
  OR3_X1 U15399 ( .A1(n13175), .A2(n13172), .A3(n13170), .ZN(n13165) );
  NAND2_X1 U15400 ( .A1(n13170), .A2(n13172), .ZN(n13163) );
  NAND3_X1 U15401 ( .A1(n13163), .A2(n13173), .A3(n13166), .ZN(n13164) );
  OAI211_X1 U15402 ( .C1(n13174), .C2(n13166), .A(n13165), .B(n13164), .ZN(
        n13167) );
  AOI21_X1 U15403 ( .B1(n13171), .B2(n13168), .A(n13167), .ZN(n13169) );
  NOR2_X1 U15404 ( .A1(n13435), .A2(n10749), .ZN(n13309) );
  NAND2_X1 U15405 ( .A1(n13310), .A2(n13309), .ZN(n13308) );
  XNOR2_X1 U15406 ( .A(n13173), .B(n13172), .ZN(n13235) );
  NAND2_X1 U15407 ( .A1(n13236), .A2(n13235), .ZN(n13234) );
  NAND2_X1 U15408 ( .A1(n13234), .A2(n13174), .ZN(n13176) );
  NAND2_X1 U15409 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  XNOR2_X1 U15410 ( .A(n13794), .B(n13226), .ZN(n13178) );
  NOR2_X1 U15411 ( .A1(n13469), .A2(n10749), .ZN(n13209) );
  INV_X1 U15412 ( .A(n13178), .ZN(n13179) );
  NAND2_X1 U15413 ( .A1(n13180), .A2(n13179), .ZN(n13181) );
  XNOR2_X1 U15414 ( .A(n13718), .B(n13186), .ZN(n13183) );
  NAND2_X1 U15415 ( .A1(n13473), .A2(n13191), .ZN(n13182) );
  NOR2_X1 U15416 ( .A1(n13183), .A2(n13182), .ZN(n13184) );
  AOI21_X1 U15417 ( .B1(n13183), .B2(n13182), .A(n13184), .ZN(n13282) );
  INV_X1 U15418 ( .A(n13184), .ZN(n13185) );
  XNOR2_X1 U15419 ( .A(n13788), .B(n13186), .ZN(n13188) );
  NAND2_X1 U15420 ( .A1(n13475), .A2(n13191), .ZN(n13187) );
  NOR2_X1 U15421 ( .A1(n13188), .A2(n13187), .ZN(n13189) );
  AOI21_X1 U15422 ( .B1(n13188), .B2(n13187), .A(n13189), .ZN(n13243) );
  INV_X1 U15423 ( .A(n13189), .ZN(n13190) );
  NAND2_X1 U15424 ( .A1(n13476), .A2(n13191), .ZN(n13193) );
  XNOR2_X1 U15425 ( .A(n13707), .B(n13226), .ZN(n13192) );
  XOR2_X1 U15426 ( .A(n13193), .B(n13192), .Z(n13330) );
  INV_X1 U15427 ( .A(n13192), .ZN(n13194) );
  NAND2_X1 U15428 ( .A1(n13194), .A2(n13193), .ZN(n13195) );
  XNOR2_X1 U15429 ( .A(n13522), .B(n13226), .ZN(n13197) );
  AND2_X1 U15430 ( .A1(n13358), .A2(n13191), .ZN(n13196) );
  NAND2_X1 U15431 ( .A1(n13197), .A2(n13196), .ZN(n13224) );
  OAI21_X1 U15432 ( .B1(n13197), .B2(n13196), .A(n13224), .ZN(n13199) );
  AOI21_X1 U15433 ( .B1(n13198), .B2(n13199), .A(n13339), .ZN(n13207) );
  INV_X1 U15434 ( .A(n13199), .ZN(n13200) );
  NAND2_X1 U15435 ( .A1(n13522), .A2(n9967), .ZN(n13205) );
  NAND2_X1 U15436 ( .A1(n13482), .A2(n13409), .ZN(n13203) );
  NAND2_X1 U15437 ( .A1(n13476), .A2(n13331), .ZN(n13202) );
  NAND2_X1 U15438 ( .A1(n13203), .A2(n13202), .ZN(n13512) );
  AOI22_X1 U15439 ( .A1(n13334), .A2(n13512), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13204) );
  OAI211_X1 U15440 ( .C1(n13336), .C2(n13520), .A(n13205), .B(n13204), .ZN(
        n13206) );
  OAI211_X1 U15441 ( .C1(n13210), .C2(n13209), .A(n13208), .B(n13343), .ZN(
        n13215) );
  INV_X1 U15442 ( .A(n13211), .ZN(n13573) );
  AOI22_X1 U15443 ( .A1(n13467), .A2(n13331), .B1(n13409), .B2(n13473), .ZN(
        n13722) );
  INV_X1 U15444 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13212) );
  OAI22_X1 U15445 ( .A1(n13348), .A2(n13722), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13212), .ZN(n13213) );
  AOI21_X1 U15446 ( .B1(n13573), .B2(n13350), .A(n13213), .ZN(n13214) );
  OAI211_X1 U15447 ( .C1(n13794), .C2(n13354), .A(n13215), .B(n13214), .ZN(
        P2_U3188) );
  AOI21_X1 U15448 ( .B1(n13217), .B2(n13216), .A(n6813), .ZN(n13223) );
  OR2_X1 U15449 ( .A1(n13462), .A2(n13312), .ZN(n13219) );
  NAND2_X1 U15450 ( .A1(n13424), .A2(n13331), .ZN(n13218) );
  NAND2_X1 U15451 ( .A1(n13219), .A2(n13218), .ZN(n13632) );
  NAND2_X1 U15452 ( .A1(n13334), .A2(n13632), .ZN(n13220) );
  NAND2_X1 U15453 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13403)
         );
  OAI211_X1 U15454 ( .C1(n13336), .C2(n13638), .A(n13220), .B(n13403), .ZN(
        n13221) );
  AOI21_X1 U15455 ( .B1(n13637), .B2(n9967), .A(n13221), .ZN(n13222) );
  OAI21_X1 U15456 ( .B1(n13223), .B2(n13339), .A(n13222), .ZN(P2_U3191) );
  NAND2_X1 U15457 ( .A1(n13482), .A2(n13191), .ZN(n13227) );
  XNOR2_X1 U15458 ( .A(n13227), .B(n13226), .ZN(n13228) );
  XNOR2_X1 U15459 ( .A(n13503), .B(n13228), .ZN(n13229) );
  INV_X1 U15460 ( .A(n13358), .ZN(n13480) );
  OAI22_X1 U15461 ( .A1(n13480), .A2(n13448), .B1(n13230), .B2(n13312), .ZN(
        n13497) );
  AOI22_X1 U15462 ( .A1(n13334), .A2(n13497), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13231) );
  OAI21_X1 U15463 ( .B1(n13504), .B2(n13336), .A(n13231), .ZN(n13232) );
  AOI21_X1 U15464 ( .B1(n13503), .B2(n9967), .A(n13232), .ZN(n13233) );
  OAI211_X1 U15465 ( .C1(n13236), .C2(n13235), .A(n13234), .B(n13343), .ZN(
        n13241) );
  OAI22_X1 U15466 ( .A1(n13435), .A2(n13312), .B1(n13462), .B2(n13448), .ZN(
        n13600) );
  AOI22_X1 U15467 ( .A1(n13600), .A2(n13334), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13240) );
  NAND2_X1 U15468 ( .A1(n13237), .A2(n9967), .ZN(n13239) );
  NAND2_X1 U15469 ( .A1(n13350), .A2(n13605), .ZN(n13238) );
  NAND4_X1 U15470 ( .A1(n13241), .A2(n13240), .A3(n13239), .A4(n13238), .ZN(
        P2_U3195) );
  OAI211_X1 U15471 ( .C1(n13244), .C2(n13243), .A(n13242), .B(n13343), .ZN(
        n13250) );
  NAND2_X1 U15472 ( .A1(n13473), .A2(n13331), .ZN(n13246) );
  NAND2_X1 U15473 ( .A1(n13476), .A2(n13409), .ZN(n13245) );
  NAND2_X1 U15474 ( .A1(n13246), .A2(n13245), .ZN(n13542) );
  AOI22_X1 U15475 ( .A1(n13334), .A2(n13542), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13247) );
  OAI21_X1 U15476 ( .B1(n13550), .B2(n13336), .A(n13247), .ZN(n13248) );
  AOI21_X1 U15477 ( .B1(n13788), .B2(n9967), .A(n13248), .ZN(n13249) );
  NAND2_X1 U15478 ( .A1(n13250), .A2(n13249), .ZN(P2_U3197) );
  AOI21_X1 U15479 ( .B1(n13252), .B2(n13251), .A(n13273), .ZN(n13260) );
  NAND2_X1 U15480 ( .A1(n13334), .A2(n13253), .ZN(n13256) );
  NAND2_X1 U15481 ( .A1(n13350), .A2(n13254), .ZN(n13255) );
  OAI211_X1 U15482 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n13257), .A(n13256), .B(
        n13255), .ZN(n13258) );
  AOI21_X1 U15483 ( .B1(n13813), .B2(n9967), .A(n13258), .ZN(n13259) );
  OAI21_X1 U15484 ( .B1(n13260), .B2(n13339), .A(n13259), .ZN(P2_U3198) );
  OAI21_X1 U15485 ( .B1(n13263), .B2(n13262), .A(n13261), .ZN(n13264) );
  NAND2_X1 U15486 ( .A1(n13264), .A2(n13343), .ZN(n13270) );
  NAND2_X1 U15487 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14915) );
  INV_X1 U15488 ( .A(n13265), .ZN(n13266) );
  AOI22_X1 U15489 ( .A1(n9967), .A2(n15078), .B1(n13350), .B2(n13266), .ZN(
        n13269) );
  NAND2_X1 U15490 ( .A1(n13334), .A2(n13267), .ZN(n13268) );
  NAND4_X1 U15491 ( .A1(n13270), .A2(n14915), .A3(n13269), .A4(n13268), .ZN(
        P2_U3199) );
  NOR3_X1 U15492 ( .A1(n13273), .A2(n13272), .A3(n13271), .ZN(n13274) );
  OAI21_X1 U15493 ( .B1(n6820), .B2(n13274), .A(n13343), .ZN(n13280) );
  INV_X1 U15494 ( .A(n13275), .ZN(n13675) );
  NOR2_X1 U15495 ( .A1(n13451), .A2(n13448), .ZN(n13276) );
  AOI21_X1 U15496 ( .B1(n13424), .B2(n13409), .A(n13276), .ZN(n13669) );
  OAI22_X1 U15497 ( .A1(n13348), .A2(n13669), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13277), .ZN(n13278) );
  AOI21_X1 U15498 ( .B1(n13675), .B2(n13350), .A(n13278), .ZN(n13279) );
  OAI211_X1 U15499 ( .C1(n13810), .C2(n13354), .A(n13280), .B(n13279), .ZN(
        P2_U3200) );
  OAI211_X1 U15500 ( .C1(n13283), .C2(n13282), .A(n13281), .B(n13343), .ZN(
        n13288) );
  INV_X1 U15501 ( .A(n13284), .ZN(n13563) );
  AOI22_X1 U15502 ( .A1(n13470), .A2(n13331), .B1(n13409), .B2(n13475), .ZN(
        n13556) );
  OAI22_X1 U15503 ( .A1(n13348), .A2(n13556), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13285), .ZN(n13286) );
  AOI21_X1 U15504 ( .B1(n13563), .B2(n13350), .A(n13286), .ZN(n13287) );
  OAI211_X1 U15505 ( .C1(n7235), .C2(n13354), .A(n13288), .B(n13287), .ZN(
        P2_U3201) );
  OAI21_X1 U15506 ( .B1(n13291), .B2(n13290), .A(n13289), .ZN(n13292) );
  NAND2_X1 U15507 ( .A1(n13292), .A2(n13343), .ZN(n13299) );
  NAND2_X1 U15508 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14902) );
  INV_X1 U15509 ( .A(n13293), .ZN(n13294) );
  AOI22_X1 U15510 ( .A1(n9967), .A2(n13295), .B1(n13350), .B2(n13294), .ZN(
        n13298) );
  NAND2_X1 U15511 ( .A1(n13334), .A2(n13296), .ZN(n13297) );
  NAND4_X1 U15512 ( .A1(n13299), .A2(n14902), .A3(n13298), .A4(n13297), .ZN(
        P2_U3202) );
  NOR3_X1 U15513 ( .A1(n6813), .A2(n7440), .A3(n13301), .ZN(n13303) );
  OAI21_X1 U15514 ( .B1(n13303), .B2(n13302), .A(n13343), .ZN(n13307) );
  AOI22_X1 U15515 ( .A1(n13432), .A2(n13409), .B1(n13331), .B2(n13428), .ZN(
        n13621) );
  OAI22_X1 U15516 ( .A1(n13348), .A2(n13621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13304), .ZN(n13305) );
  AOI21_X1 U15517 ( .B1(n13615), .B2(n13350), .A(n13305), .ZN(n13306) );
  OAI211_X1 U15518 ( .C1(n13617), .C2(n13354), .A(n13307), .B(n13306), .ZN(
        P2_U3205) );
  OAI211_X1 U15519 ( .C1(n13310), .C2(n13309), .A(n13308), .B(n13343), .ZN(
        n13317) );
  INV_X1 U15520 ( .A(n13311), .ZN(n13592) );
  OAI22_X1 U15521 ( .A1(n13465), .A2(n13448), .B1(n13469), .B2(n13312), .ZN(
        n13585) );
  INV_X1 U15522 ( .A(n13585), .ZN(n13314) );
  OAI22_X1 U15523 ( .A1(n13348), .A2(n13314), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13313), .ZN(n13315) );
  AOI21_X1 U15524 ( .B1(n13592), .B2(n13350), .A(n13315), .ZN(n13316) );
  OAI211_X1 U15525 ( .C1(n13595), .C2(n13354), .A(n13317), .B(n13316), .ZN(
        P2_U3207) );
  AOI21_X1 U15526 ( .B1(n13319), .B2(n13318), .A(n13339), .ZN(n13321) );
  NAND2_X1 U15527 ( .A1(n13321), .A2(n13320), .ZN(n13326) );
  NOR2_X1 U15528 ( .A1(n13455), .A2(n13448), .ZN(n13322) );
  AOI21_X1 U15529 ( .B1(n13428), .B2(n13409), .A(n13322), .ZN(n13648) );
  OAI21_X1 U15530 ( .B1(n13348), .B2(n13648), .A(n13323), .ZN(n13324) );
  AOI21_X1 U15531 ( .B1(n13654), .B2(n13350), .A(n13324), .ZN(n13325) );
  OAI211_X1 U15532 ( .C1(n13656), .C2(n13354), .A(n13326), .B(n13325), .ZN(
        P2_U3210) );
  INV_X1 U15533 ( .A(n13327), .ZN(n13328) );
  AOI21_X1 U15534 ( .B1(n13330), .B2(n13329), .A(n13328), .ZN(n13340) );
  NAND2_X1 U15535 ( .A1(n13475), .A2(n13331), .ZN(n13333) );
  NAND2_X1 U15536 ( .A1(n13358), .A2(n13409), .ZN(n13332) );
  NAND2_X1 U15537 ( .A1(n13333), .A2(n13332), .ZN(n13527) );
  AOI22_X1 U15538 ( .A1(n13334), .A2(n13527), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13335) );
  OAI21_X1 U15539 ( .B1(n13531), .B2(n13336), .A(n13335), .ZN(n13337) );
  AOI21_X1 U15540 ( .B1(n13707), .B2(n9967), .A(n13337), .ZN(n13338) );
  OAI21_X1 U15541 ( .B1(n13340), .B2(n13339), .A(n13338), .ZN(P2_U3212) );
  OAI211_X1 U15542 ( .C1(n13345), .C2(n13344), .A(n13342), .B(n13343), .ZN(
        n13353) );
  OAI22_X1 U15543 ( .A1(n13348), .A2(n13347), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13346), .ZN(n13349) );
  AOI21_X1 U15544 ( .B1(n13351), .B2(n13350), .A(n13349), .ZN(n13352) );
  OAI211_X1 U15545 ( .C1(n13355), .C2(n13354), .A(n13353), .B(n13352), .ZN(
        P2_U3213) );
  MUX2_X1 U15546 ( .A(n13410), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13373), .Z(
        P2_U3562) );
  MUX2_X1 U15547 ( .A(n13356), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13373), .Z(
        P2_U3561) );
  MUX2_X1 U15548 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13357), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15549 ( .A(n13482), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13373), .Z(
        P2_U3559) );
  MUX2_X1 U15550 ( .A(n13358), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13373), .Z(
        P2_U3558) );
  MUX2_X1 U15551 ( .A(n13476), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13373), .Z(
        P2_U3557) );
  MUX2_X1 U15552 ( .A(n13475), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13373), .Z(
        P2_U3556) );
  MUX2_X1 U15553 ( .A(n13473), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13373), .Z(
        P2_U3555) );
  MUX2_X1 U15554 ( .A(n13470), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13373), .Z(
        P2_U3554) );
  MUX2_X1 U15555 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13467), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15556 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13432), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15557 ( .A(n13428), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13373), .Z(
        P2_U3550) );
  MUX2_X1 U15558 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13424), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15559 ( .A(n13421), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13373), .Z(
        P2_U3548) );
  MUX2_X1 U15560 ( .A(n13359), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13373), .Z(
        P2_U3547) );
  MUX2_X1 U15561 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13360), .S(P2_U3947), .Z(
        P2_U3546) );
  MUX2_X1 U15562 ( .A(n13361), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13373), .Z(
        P2_U3545) );
  MUX2_X1 U15563 ( .A(n13362), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13373), .Z(
        P2_U3544) );
  MUX2_X1 U15564 ( .A(n13363), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13373), .Z(
        P2_U3543) );
  MUX2_X1 U15565 ( .A(n13364), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13373), .Z(
        P2_U3542) );
  MUX2_X1 U15566 ( .A(n13365), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13373), .Z(
        P2_U3541) );
  MUX2_X1 U15567 ( .A(n13366), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13373), .Z(
        P2_U3540) );
  MUX2_X1 U15568 ( .A(n13367), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13373), .Z(
        P2_U3539) );
  MUX2_X1 U15569 ( .A(n13368), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13373), .Z(
        P2_U3538) );
  MUX2_X1 U15570 ( .A(n7290), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13373), .Z(
        P2_U3537) );
  MUX2_X1 U15571 ( .A(n13369), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13373), .Z(
        P2_U3536) );
  MUX2_X1 U15572 ( .A(n13370), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13373), .Z(
        P2_U3535) );
  MUX2_X1 U15573 ( .A(n13371), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13373), .Z(
        P2_U3534) );
  MUX2_X1 U15574 ( .A(n13372), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13373), .Z(
        P2_U3533) );
  MUX2_X1 U15575 ( .A(n13374), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13373), .Z(
        P2_U3532) );
  MUX2_X1 U15576 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13375), .S(P2_U3947), .Z(
        P2_U3531) );
  OAI22_X1 U15577 ( .A1(n15035), .A2(n13377), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13376), .ZN(n13378) );
  AOI21_X1 U15578 ( .B1(n14864), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n13378), .ZN(
        n13387) );
  OAI211_X1 U15579 ( .C1(n13381), .C2(n13380), .A(n15028), .B(n13379), .ZN(
        n13386) );
  OAI211_X1 U15580 ( .C1(n13384), .C2(n13383), .A(n15032), .B(n13382), .ZN(
        n13385) );
  NAND3_X1 U15581 ( .A1(n13387), .A2(n13386), .A3(n13385), .ZN(P2_U3215) );
  OR2_X1 U15582 ( .A1(n13389), .A2(n13388), .ZN(n13390) );
  NAND2_X1 U15583 ( .A1(n13391), .A2(n13390), .ZN(n13392) );
  XNOR2_X1 U15584 ( .A(n13392), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13399) );
  INV_X1 U15585 ( .A(n13399), .ZN(n13397) );
  NOR2_X1 U15586 ( .A1(n13394), .A2(n13393), .ZN(n13395) );
  XNOR2_X1 U15587 ( .A(n13395), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U15588 ( .B1(n13398), .B2(n15013), .A(n15035), .ZN(n13396) );
  AOI21_X1 U15589 ( .B1(n13397), .B2(n15028), .A(n13396), .ZN(n13402) );
  AOI22_X1 U15590 ( .A1(n13399), .A2(n15028), .B1(n15032), .B2(n13398), .ZN(
        n13401) );
  MUX2_X1 U15591 ( .A(n13402), .B(n13401), .S(n13400), .Z(n13404) );
  OAI211_X1 U15592 ( .C1(n13405), .C2(n15044), .A(n13404), .B(n13403), .ZN(
        P2_U3233) );
  AND2_X1 U15593 ( .A1(n13652), .A2(n13804), .ZN(n13635) );
  NAND2_X1 U15594 ( .A1(n13614), .A2(n13799), .ZN(n13604) );
  OR2_X2 U15595 ( .A1(n13522), .A2(n13529), .ZN(n13517) );
  XNOR2_X1 U15596 ( .A(n13406), .B(n6699), .ZN(n13407) );
  NOR2_X1 U15597 ( .A1(n13407), .A2(n13191), .ZN(n13683) );
  NAND2_X1 U15598 ( .A1(n13683), .A2(n13673), .ZN(n13413) );
  NAND2_X1 U15599 ( .A1(n13830), .A2(P2_B_REG_SCAN_IN), .ZN(n13408) );
  NAND2_X1 U15600 ( .A1(n13409), .A2(n13408), .ZN(n13450) );
  INV_X1 U15601 ( .A(n13450), .ZN(n13411) );
  AND2_X1 U15602 ( .A1(n13411), .A2(n13410), .ZN(n13682) );
  INV_X1 U15603 ( .A(n13682), .ZN(n13686) );
  NOR2_X1 U15604 ( .A1(n15067), .A2(n13686), .ZN(n13416) );
  AOI21_X1 U15605 ( .B1(n15067), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13416), 
        .ZN(n13412) );
  OAI211_X1 U15606 ( .C1(n13771), .C2(n13678), .A(n13413), .B(n13412), .ZN(
        P2_U3234) );
  OAI211_X1 U15607 ( .C1(n13414), .C2(n13775), .A(n10749), .B(n6699), .ZN(
        n13687) );
  NOR2_X1 U15608 ( .A1(n13643), .A2(n13415), .ZN(n13417) );
  AOI211_X1 U15609 ( .C1(n13418), .C2(n15055), .A(n13417), .B(n13416), .ZN(
        n13419) );
  OAI21_X1 U15610 ( .B1(n13687), .B2(n15062), .A(n13419), .ZN(P2_U3235) );
  NAND2_X1 U15611 ( .A1(n13666), .A2(n13664), .ZN(n13420) );
  NAND2_X1 U15612 ( .A1(n13420), .A2(n13662), .ZN(n13668) );
  NAND2_X1 U15613 ( .A1(n13810), .A2(n13421), .ZN(n13422) );
  NAND2_X1 U15614 ( .A1(n13668), .A2(n13422), .ZN(n13647) );
  OR2_X1 U15615 ( .A1(n13656), .A2(n13424), .ZN(n13423) );
  NAND2_X1 U15616 ( .A1(n13647), .A2(n13423), .ZN(n13426) );
  NAND2_X1 U15617 ( .A1(n13656), .A2(n13424), .ZN(n13425) );
  NAND2_X1 U15618 ( .A1(n13426), .A2(n13425), .ZN(n13629) );
  OR2_X1 U15619 ( .A1(n13804), .A2(n13428), .ZN(n13427) );
  NAND2_X1 U15620 ( .A1(n13804), .A2(n13428), .ZN(n13627) );
  OR2_X1 U15621 ( .A1(n13799), .A2(n13432), .ZN(n13431) );
  NAND2_X1 U15622 ( .A1(n13799), .A2(n13432), .ZN(n13433) );
  NAND2_X1 U15623 ( .A1(n13730), .A2(n13435), .ZN(n13436) );
  NAND2_X1 U15624 ( .A1(n13794), .A2(n13470), .ZN(n13437) );
  NAND2_X1 U15625 ( .A1(n13718), .A2(n13438), .ZN(n13439) );
  INV_X1 U15626 ( .A(n13545), .ZN(n13540) );
  NAND2_X1 U15627 ( .A1(n13526), .A2(n13441), .ZN(n13443) );
  NAND2_X1 U15628 ( .A1(n13496), .A2(n13500), .ZN(n13495) );
  NAND2_X1 U15629 ( .A1(n13495), .A2(n13444), .ZN(n13445) );
  OR2_X1 U15630 ( .A1(n13452), .A2(n13451), .ZN(n13453) );
  INV_X1 U15631 ( .A(n13662), .ZN(n13665) );
  OR2_X1 U15632 ( .A1(n13810), .A2(n13455), .ZN(n13456) );
  INV_X1 U15633 ( .A(n13646), .ZN(n13658) );
  NAND2_X1 U15634 ( .A1(n13626), .A2(n13458), .ZN(n13460) );
  AND2_X1 U15635 ( .A1(n13617), .A2(n13462), .ZN(n13461) );
  OR2_X1 U15636 ( .A1(n13617), .A2(n13462), .ZN(n13463) );
  INV_X1 U15637 ( .A(n13602), .ZN(n13464) );
  NAND2_X1 U15638 ( .A1(n13730), .A2(n13467), .ZN(n13468) );
  NOR2_X1 U15639 ( .A1(n13794), .A2(n13469), .ZN(n13472) );
  NAND2_X1 U15640 ( .A1(n13718), .A2(n13473), .ZN(n13474) );
  NOR2_X1 U15641 ( .A1(n13707), .A2(n13476), .ZN(n13478) );
  NAND2_X1 U15642 ( .A1(n13707), .A2(n13476), .ZN(n13477) );
  NAND2_X1 U15643 ( .A1(n13484), .A2(n13483), .ZN(n13486) );
  NAND2_X1 U15644 ( .A1(n15067), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n13488) );
  OAI21_X1 U15645 ( .B1(n15052), .B2(n13489), .A(n13488), .ZN(n13490) );
  AOI21_X1 U15646 ( .B1(n13491), .B2(n15055), .A(n13490), .ZN(n13492) );
  OAI21_X1 U15647 ( .B1(n13691), .B2(n15062), .A(n13492), .ZN(n13493) );
  AOI21_X1 U15648 ( .B1(n13690), .B2(n13609), .A(n13493), .ZN(n13494) );
  OAI21_X1 U15649 ( .B1(n6752), .B2(n15067), .A(n13494), .ZN(P2_U3236) );
  OAI211_X1 U15650 ( .C1(n13496), .C2(n13500), .A(n13495), .B(n15048), .ZN(
        n13499) );
  INV_X1 U15651 ( .A(n13497), .ZN(n13498) );
  NAND2_X1 U15652 ( .A1(n13499), .A2(n13498), .ZN(n13695) );
  INV_X1 U15653 ( .A(n13695), .ZN(n13510) );
  XNOR2_X1 U15654 ( .A(n13501), .B(n13500), .ZN(n13697) );
  NAND2_X1 U15655 ( .A1(n13697), .A2(n13609), .ZN(n13509) );
  AOI211_X1 U15656 ( .C1(n13503), .C2(n13517), .A(n13191), .B(n13502), .ZN(
        n13696) );
  INV_X1 U15657 ( .A(n13504), .ZN(n13505) );
  AOI22_X1 U15658 ( .A1(n15067), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n13505), 
        .B2(n13674), .ZN(n13506) );
  OAI21_X1 U15659 ( .B1(n13780), .B2(n13678), .A(n13506), .ZN(n13507) );
  AOI21_X1 U15660 ( .B1(n13696), .B2(n13673), .A(n13507), .ZN(n13508) );
  OAI211_X1 U15661 ( .C1(n13510), .C2(n15067), .A(n13509), .B(n13508), .ZN(
        P2_U3237) );
  XNOR2_X1 U15662 ( .A(n13511), .B(n13514), .ZN(n13513) );
  AOI21_X1 U15663 ( .B1(n13513), .B2(n15048), .A(n13512), .ZN(n13702) );
  INV_X1 U15664 ( .A(n13514), .ZN(n13515) );
  XNOR2_X1 U15665 ( .A(n13516), .B(n13515), .ZN(n13700) );
  AOI21_X1 U15666 ( .B1(n13522), .B2(n13529), .A(n13191), .ZN(n13518) );
  NAND2_X1 U15667 ( .A1(n13518), .A2(n13517), .ZN(n13701) );
  NAND2_X1 U15668 ( .A1(n15067), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n13519) );
  OAI21_X1 U15669 ( .B1(n15052), .B2(n13520), .A(n13519), .ZN(n13521) );
  AOI21_X1 U15670 ( .B1(n13522), .B2(n15055), .A(n13521), .ZN(n13523) );
  OAI21_X1 U15671 ( .B1(n13701), .B2(n15062), .A(n13523), .ZN(n13524) );
  AOI21_X1 U15672 ( .B1(n13700), .B2(n13609), .A(n13524), .ZN(n13525) );
  OAI21_X1 U15673 ( .B1(n13702), .B2(n15067), .A(n13525), .ZN(P2_U3238) );
  XOR2_X1 U15674 ( .A(n13535), .B(n13526), .Z(n13528) );
  AOI21_X1 U15675 ( .B1(n13528), .B2(n15048), .A(n13527), .ZN(n13709) );
  INV_X1 U15676 ( .A(n13529), .ZN(n13530) );
  AOI211_X1 U15677 ( .C1(n13707), .C2(n13547), .A(n13191), .B(n13530), .ZN(
        n13706) );
  INV_X1 U15678 ( .A(n13531), .ZN(n13532) );
  AOI22_X1 U15679 ( .A1(n15067), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13532), 
        .B2(n13674), .ZN(n13533) );
  OAI21_X1 U15680 ( .B1(n7233), .B2(n13678), .A(n13533), .ZN(n13537) );
  XOR2_X1 U15681 ( .A(n13535), .B(n13534), .Z(n13710) );
  NOR2_X1 U15682 ( .A1(n13710), .A2(n15063), .ZN(n13536) );
  AOI211_X1 U15683 ( .C1(n13706), .C2(n13673), .A(n13537), .B(n13536), .ZN(
        n13538) );
  OAI21_X1 U15684 ( .B1(n15067), .B2(n13709), .A(n13538), .ZN(P2_U3239) );
  OAI21_X1 U15685 ( .B1(n13541), .B2(n13540), .A(n13539), .ZN(n13543) );
  AOI21_X1 U15686 ( .B1(n13543), .B2(n15048), .A(n13542), .ZN(n13713) );
  OAI21_X1 U15687 ( .B1(n13546), .B2(n7330), .A(n13544), .ZN(n13711) );
  AOI21_X1 U15688 ( .B1(n13788), .B2(n13561), .A(n13191), .ZN(n13548) );
  NAND2_X1 U15689 ( .A1(n13548), .A2(n13547), .ZN(n13712) );
  NAND2_X1 U15690 ( .A1(n15067), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13549) );
  OAI21_X1 U15691 ( .B1(n15052), .B2(n13550), .A(n13549), .ZN(n13551) );
  AOI21_X1 U15692 ( .B1(n13788), .B2(n15055), .A(n13551), .ZN(n13552) );
  OAI21_X1 U15693 ( .B1(n13712), .B2(n15062), .A(n13552), .ZN(n13553) );
  AOI21_X1 U15694 ( .B1(n13711), .B2(n13609), .A(n13553), .ZN(n13554) );
  OAI21_X1 U15695 ( .B1(n15067), .B2(n13713), .A(n13554), .ZN(P2_U3240) );
  XNOR2_X1 U15696 ( .A(n13555), .B(n6681), .ZN(n13558) );
  INV_X1 U15697 ( .A(n13556), .ZN(n13557) );
  AOI21_X1 U15698 ( .B1(n13558), .B2(n15048), .A(n13557), .ZN(n13720) );
  OAI21_X1 U15699 ( .B1(n6696), .B2(n6681), .A(n13559), .ZN(n13721) );
  INV_X1 U15700 ( .A(n13721), .ZN(n13567) );
  AOI21_X1 U15701 ( .B1(n13718), .B2(n13574), .A(n13191), .ZN(n13562) );
  AND2_X1 U15702 ( .A1(n13562), .A2(n13561), .ZN(n13717) );
  NAND2_X1 U15703 ( .A1(n13717), .A2(n13673), .ZN(n13565) );
  AOI22_X1 U15704 ( .A1(n15067), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13563), 
        .B2(n13674), .ZN(n13564) );
  OAI211_X1 U15705 ( .C1(n7235), .C2(n13678), .A(n13565), .B(n13564), .ZN(
        n13566) );
  AOI21_X1 U15706 ( .B1(n13567), .B2(n13609), .A(n13566), .ZN(n13568) );
  OAI21_X1 U15707 ( .B1(n15067), .B2(n13720), .A(n13568), .ZN(P2_U3241) );
  INV_X1 U15708 ( .A(n13722), .ZN(n13572) );
  INV_X1 U15709 ( .A(n13569), .ZN(n13570) );
  AOI211_X1 U15710 ( .C1(n13579), .C2(n13571), .A(n13622), .B(n13570), .ZN(
        n13724) );
  AOI211_X1 U15711 ( .C1(n13674), .C2(n13573), .A(n13572), .B(n13724), .ZN(
        n13583) );
  INV_X1 U15712 ( .A(n13590), .ZN(n13575) );
  OAI211_X1 U15713 ( .C1(n13575), .C2(n13794), .A(n10749), .B(n13574), .ZN(
        n13723) );
  INV_X1 U15714 ( .A(n13723), .ZN(n13578) );
  OAI22_X1 U15715 ( .A1(n13794), .A2(n13678), .B1(n13643), .B2(n13576), .ZN(
        n13577) );
  AOI21_X1 U15716 ( .B1(n13578), .B2(n13673), .A(n13577), .ZN(n13582) );
  XOR2_X1 U15717 ( .A(n13580), .B(n13579), .Z(n13726) );
  NAND2_X1 U15718 ( .A1(n13726), .A2(n13609), .ZN(n13581) );
  OAI211_X1 U15719 ( .C1(n13583), .C2(n15067), .A(n13582), .B(n13581), .ZN(
        P2_U3242) );
  XNOR2_X1 U15720 ( .A(n13584), .B(n13588), .ZN(n13586) );
  AOI21_X1 U15721 ( .B1(n13586), .B2(n15048), .A(n13585), .ZN(n13732) );
  OAI21_X1 U15722 ( .B1(n13589), .B2(n13588), .A(n13587), .ZN(n13733) );
  INV_X1 U15723 ( .A(n13733), .ZN(n13597) );
  AOI21_X1 U15724 ( .B1(n13604), .B2(n13730), .A(n13191), .ZN(n13591) );
  AND2_X1 U15725 ( .A1(n13591), .A2(n13590), .ZN(n13729) );
  NAND2_X1 U15726 ( .A1(n13729), .A2(n13673), .ZN(n13594) );
  AOI22_X1 U15727 ( .A1(n15067), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13592), 
        .B2(n13674), .ZN(n13593) );
  OAI211_X1 U15728 ( .C1(n13595), .C2(n13678), .A(n13594), .B(n13593), .ZN(
        n13596) );
  AOI21_X1 U15729 ( .B1(n13597), .B2(n13609), .A(n13596), .ZN(n13598) );
  OAI21_X1 U15730 ( .B1(n15067), .B2(n13732), .A(n13598), .ZN(P2_U3243) );
  XNOR2_X1 U15731 ( .A(n13599), .B(n13602), .ZN(n13601) );
  AOI21_X1 U15732 ( .B1(n13601), .B2(n15048), .A(n13600), .ZN(n13735) );
  XNOR2_X1 U15733 ( .A(n13603), .B(n13602), .ZN(n13736) );
  INV_X1 U15734 ( .A(n13736), .ZN(n13610) );
  OAI211_X1 U15735 ( .C1(n13614), .C2(n13799), .A(n10749), .B(n13604), .ZN(
        n13734) );
  NOR2_X1 U15736 ( .A1(n13734), .A2(n15062), .ZN(n13608) );
  AOI22_X1 U15737 ( .A1(n15067), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13605), 
        .B2(n13674), .ZN(n13606) );
  OAI21_X1 U15738 ( .B1(n13799), .B2(n13678), .A(n13606), .ZN(n13607) );
  AOI211_X1 U15739 ( .C1(n13610), .C2(n13609), .A(n13608), .B(n13607), .ZN(
        n13611) );
  OAI21_X1 U15740 ( .B1(n15067), .B2(n13735), .A(n13611), .ZN(P2_U3244) );
  XOR2_X1 U15741 ( .A(n13620), .B(n13612), .Z(n13743) );
  NOR2_X1 U15742 ( .A1(n13617), .A2(n13635), .ZN(n13613) );
  AOI22_X1 U15743 ( .A1(n15067), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13615), 
        .B2(n13674), .ZN(n13616) );
  OAI21_X1 U15744 ( .B1(n13617), .B2(n13678), .A(n13616), .ZN(n13618) );
  AOI21_X1 U15745 ( .B1(n6815), .B2(n13673), .A(n13618), .ZN(n13625) );
  XOR2_X1 U15746 ( .A(n13620), .B(n13619), .Z(n13623) );
  OAI21_X1 U15747 ( .B1(n13623), .B2(n13622), .A(n13621), .ZN(n13740) );
  NAND2_X1 U15748 ( .A1(n13740), .A2(n13643), .ZN(n13624) );
  OAI211_X1 U15749 ( .C1(n13743), .C2(n15063), .A(n13625), .B(n13624), .ZN(
        P2_U3245) );
  XNOR2_X1 U15750 ( .A(n13626), .B(n13628), .ZN(n13746) );
  INV_X1 U15751 ( .A(n13746), .ZN(n13645) );
  OR2_X1 U15752 ( .A1(n13629), .A2(n7084), .ZN(n13630) );
  OAI211_X1 U15753 ( .C1(n13631), .C2(n7300), .A(n15048), .B(n13630), .ZN(
        n13634) );
  INV_X1 U15754 ( .A(n13632), .ZN(n13633) );
  NAND2_X1 U15755 ( .A1(n13634), .A2(n13633), .ZN(n13744) );
  INV_X1 U15756 ( .A(n13652), .ZN(n13636) );
  AOI211_X1 U15757 ( .C1(n13637), .C2(n13636), .A(n13191), .B(n13635), .ZN(
        n13745) );
  NAND2_X1 U15758 ( .A1(n13745), .A2(n13673), .ZN(n13641) );
  INV_X1 U15759 ( .A(n13638), .ZN(n13639) );
  AOI22_X1 U15760 ( .A1(n15067), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13639), 
        .B2(n13674), .ZN(n13640) );
  OAI211_X1 U15761 ( .C1(n13804), .C2(n13678), .A(n13641), .B(n13640), .ZN(
        n13642) );
  AOI21_X1 U15762 ( .B1(n13744), .B2(n13643), .A(n13642), .ZN(n13644) );
  OAI21_X1 U15763 ( .B1(n13645), .B2(n15063), .A(n13644), .ZN(P2_U3246) );
  XNOR2_X1 U15764 ( .A(n13647), .B(n13646), .ZN(n13650) );
  INV_X1 U15765 ( .A(n13648), .ZN(n13649) );
  AOI21_X1 U15766 ( .B1(n13650), .B2(n15048), .A(n13649), .ZN(n13751) );
  NOR2_X1 U15767 ( .A1(n6814), .A2(n13656), .ZN(n13653) );
  AOI22_X1 U15768 ( .A1(n15067), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13654), 
        .B2(n13674), .ZN(n13655) );
  OAI21_X1 U15769 ( .B1(n13656), .B2(n13678), .A(n13655), .ZN(n13660) );
  AOI21_X1 U15770 ( .B1(n13658), .B2(n13657), .A(n6762), .ZN(n13752) );
  NOR2_X1 U15771 ( .A1(n13752), .A2(n15063), .ZN(n13659) );
  AOI211_X1 U15772 ( .C1(n7756), .C2(n13673), .A(n13660), .B(n13659), .ZN(
        n13661) );
  OAI21_X1 U15773 ( .B1(n15067), .B2(n13751), .A(n13661), .ZN(P2_U3247) );
  XNOR2_X1 U15774 ( .A(n13663), .B(n13662), .ZN(n13755) );
  INV_X1 U15775 ( .A(n13755), .ZN(n13681) );
  NAND3_X1 U15776 ( .A1(n13666), .A2(n13665), .A3(n13664), .ZN(n13667) );
  NAND3_X1 U15777 ( .A1(n13668), .A2(n15048), .A3(n13667), .ZN(n13670) );
  NAND2_X1 U15778 ( .A1(n13670), .A2(n13669), .ZN(n13753) );
  AOI211_X1 U15779 ( .C1(n13672), .C2(n13671), .A(n13191), .B(n6814), .ZN(
        n13754) );
  NAND2_X1 U15780 ( .A1(n13754), .A2(n13673), .ZN(n13677) );
  AOI22_X1 U15781 ( .A1(n15067), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13675), 
        .B2(n13674), .ZN(n13676) );
  OAI211_X1 U15782 ( .C1(n13810), .C2(n13678), .A(n13677), .B(n13676), .ZN(
        n13679) );
  AOI21_X1 U15783 ( .B1(n13643), .B2(n13753), .A(n13679), .ZN(n13680) );
  OAI21_X1 U15784 ( .B1(n13681), .B2(n15063), .A(n13680), .ZN(P2_U3248) );
  NOR2_X1 U15785 ( .A1(n13683), .A2(n13682), .ZN(n13768) );
  MUX2_X1 U15786 ( .A(n13684), .B(n13768), .S(n15129), .Z(n13685) );
  OAI21_X1 U15787 ( .B1(n13771), .B2(n13758), .A(n13685), .ZN(P2_U3530) );
  AND2_X1 U15788 ( .A1(n13687), .A2(n13686), .ZN(n13772) );
  MUX2_X1 U15789 ( .A(n13688), .B(n13772), .S(n15129), .Z(n13689) );
  OAI21_X1 U15790 ( .B1(n13775), .B2(n13758), .A(n13689), .ZN(P2_U3529) );
  NAND2_X1 U15791 ( .A1(n13690), .A2(n15099), .ZN(n13694) );
  OAI21_X1 U15792 ( .B1(n13692), .B2(n15111), .A(n13691), .ZN(n13693) );
  INV_X1 U15793 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n13698) );
  MUX2_X1 U15794 ( .A(n13698), .B(n13777), .S(n15129), .Z(n13699) );
  NAND2_X1 U15795 ( .A1(n13700), .A2(n15099), .ZN(n13703) );
  NAND3_X1 U15796 ( .A1(n13703), .A2(n13702), .A3(n13701), .ZN(n13781) );
  MUX2_X1 U15797 ( .A(n13781), .B(P2_REG1_REG_27__SCAN_IN), .S(n15127), .Z(
        n13704) );
  INV_X1 U15798 ( .A(n13704), .ZN(n13705) );
  OAI21_X1 U15799 ( .B1(n13784), .B2(n13758), .A(n13705), .ZN(P2_U3526) );
  AOI21_X1 U15800 ( .B1(n15079), .B2(n13707), .A(n13706), .ZN(n13708) );
  OAI211_X1 U15801 ( .C1(n13710), .C2(n13759), .A(n13709), .B(n13708), .ZN(
        n13785) );
  MUX2_X1 U15802 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13785), .S(n15129), .Z(
        P2_U3525) );
  NAND2_X1 U15803 ( .A1(n13711), .A2(n15099), .ZN(n13714) );
  NAND3_X1 U15804 ( .A1(n13714), .A2(n13713), .A3(n13712), .ZN(n13786) );
  MUX2_X1 U15805 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13786), .S(n15129), .Z(
        n13715) );
  AOI21_X1 U15806 ( .B1(n13766), .B2(n13788), .A(n13715), .ZN(n13716) );
  INV_X1 U15807 ( .A(n13716), .ZN(P2_U3524) );
  AOI21_X1 U15808 ( .B1(n15079), .B2(n13718), .A(n13717), .ZN(n13719) );
  OAI211_X1 U15809 ( .C1(n13721), .C2(n13759), .A(n13720), .B(n13719), .ZN(
        n13790) );
  MUX2_X1 U15810 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13790), .S(n15129), .Z(
        P2_U3523) );
  INV_X1 U15811 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13727) );
  NAND2_X1 U15812 ( .A1(n13723), .A2(n13722), .ZN(n13725) );
  AOI211_X1 U15813 ( .C1(n13726), .C2(n15099), .A(n13725), .B(n13724), .ZN(
        n13791) );
  MUX2_X1 U15814 ( .A(n13727), .B(n13791), .S(n15129), .Z(n13728) );
  OAI21_X1 U15815 ( .B1(n13794), .B2(n13758), .A(n13728), .ZN(P2_U3522) );
  AOI21_X1 U15816 ( .B1(n15079), .B2(n13730), .A(n13729), .ZN(n13731) );
  OAI211_X1 U15817 ( .C1(n13733), .C2(n13759), .A(n13732), .B(n13731), .ZN(
        n13795) );
  MUX2_X1 U15818 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13795), .S(n15129), .Z(
        P2_U3521) );
  OAI211_X1 U15819 ( .C1(n13736), .C2(n13759), .A(n13735), .B(n13734), .ZN(
        n13737) );
  INV_X1 U15820 ( .A(n13737), .ZN(n13796) );
  MUX2_X1 U15821 ( .A(n13738), .B(n13796), .S(n15129), .Z(n13739) );
  OAI21_X1 U15822 ( .B1(n13799), .B2(n13758), .A(n13739), .ZN(P2_U3520) );
  AOI211_X1 U15823 ( .C1(n15079), .C2(n13741), .A(n6815), .B(n13740), .ZN(
        n13742) );
  OAI21_X1 U15824 ( .B1(n13743), .B2(n13759), .A(n13742), .ZN(n13800) );
  MUX2_X1 U15825 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13800), .S(n15129), .Z(
        P2_U3519) );
  AOI211_X1 U15826 ( .C1(n13746), .C2(n15099), .A(n13745), .B(n13744), .ZN(
        n13801) );
  MUX2_X1 U15827 ( .A(n13747), .B(n13801), .S(n15129), .Z(n13748) );
  OAI21_X1 U15828 ( .B1(n13804), .B2(n13758), .A(n13748), .ZN(P2_U3518) );
  AOI21_X1 U15829 ( .B1(n15079), .B2(n13749), .A(n7756), .ZN(n13750) );
  OAI211_X1 U15830 ( .C1(n13752), .C2(n13759), .A(n13751), .B(n13750), .ZN(
        n13805) );
  MUX2_X1 U15831 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13805), .S(n15129), .Z(
        P2_U3517) );
  AOI211_X1 U15832 ( .C1(n13755), .C2(n15099), .A(n13754), .B(n13753), .ZN(
        n13806) );
  MUX2_X1 U15833 ( .A(n13756), .B(n13806), .S(n15129), .Z(n13757) );
  OAI21_X1 U15834 ( .B1(n13810), .B2(n13758), .A(n13757), .ZN(P2_U3516) );
  OR2_X1 U15835 ( .A1(n13760), .A2(n13759), .ZN(n13764) );
  NOR2_X1 U15836 ( .A1(n13762), .A2(n13761), .ZN(n13763) );
  NAND2_X1 U15837 ( .A1(n13764), .A2(n13763), .ZN(n13811) );
  MUX2_X1 U15838 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13811), .S(n15129), .Z(
        n13765) );
  AOI21_X1 U15839 ( .B1(n13766), .B2(n13813), .A(n13765), .ZN(n13767) );
  INV_X1 U15840 ( .A(n13767), .ZN(P2_U3515) );
  INV_X1 U15841 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13769) );
  MUX2_X1 U15842 ( .A(n13769), .B(n13768), .S(n15119), .Z(n13770) );
  OAI21_X1 U15843 ( .B1(n13771), .B2(n13809), .A(n13770), .ZN(P2_U3498) );
  MUX2_X1 U15844 ( .A(n13773), .B(n13772), .S(n15119), .Z(n13774) );
  OAI21_X1 U15845 ( .B1(n13775), .B2(n13809), .A(n13774), .ZN(P2_U3497) );
  MUX2_X1 U15846 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13776), .S(n15119), .Z(
        P2_U3496) );
  INV_X1 U15847 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n13778) );
  MUX2_X1 U15848 ( .A(n13778), .B(n13777), .S(n15119), .Z(n13779) );
  MUX2_X1 U15849 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13781), .S(n15119), .Z(
        n13782) );
  INV_X1 U15850 ( .A(n13782), .ZN(n13783) );
  OAI21_X1 U15851 ( .B1(n13784), .B2(n13809), .A(n13783), .ZN(P2_U3494) );
  MUX2_X1 U15852 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13785), .S(n15119), .Z(
        P2_U3493) );
  INV_X1 U15853 ( .A(n13809), .ZN(n13814) );
  MUX2_X1 U15854 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13786), .S(n15119), .Z(
        n13787) );
  AOI21_X1 U15855 ( .B1(n13814), .B2(n13788), .A(n13787), .ZN(n13789) );
  INV_X1 U15856 ( .A(n13789), .ZN(P2_U3492) );
  MUX2_X1 U15857 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13790), .S(n15119), .Z(
        P2_U3491) );
  MUX2_X1 U15858 ( .A(n13792), .B(n13791), .S(n15119), .Z(n13793) );
  OAI21_X1 U15859 ( .B1(n13794), .B2(n13809), .A(n13793), .ZN(P2_U3490) );
  MUX2_X1 U15860 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13795), .S(n15119), .Z(
        P2_U3489) );
  INV_X1 U15861 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13797) );
  MUX2_X1 U15862 ( .A(n13797), .B(n13796), .S(n15119), .Z(n13798) );
  OAI21_X1 U15863 ( .B1(n13799), .B2(n13809), .A(n13798), .ZN(P2_U3488) );
  MUX2_X1 U15864 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13800), .S(n15119), .Z(
        P2_U3487) );
  INV_X1 U15865 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13802) );
  MUX2_X1 U15866 ( .A(n13802), .B(n13801), .S(n15119), .Z(n13803) );
  OAI21_X1 U15867 ( .B1(n13804), .B2(n13809), .A(n13803), .ZN(P2_U3486) );
  MUX2_X1 U15868 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13805), .S(n15119), .Z(
        P2_U3484) );
  INV_X1 U15869 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13807) );
  MUX2_X1 U15870 ( .A(n13807), .B(n13806), .S(n15119), .Z(n13808) );
  OAI21_X1 U15871 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(P2_U3481) );
  MUX2_X1 U15872 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13811), .S(n15119), .Z(
        n13812) );
  AOI21_X1 U15873 ( .B1(n13814), .B2(n13813), .A(n13812), .ZN(n13815) );
  INV_X1 U15874 ( .A(n13815), .ZN(P2_U3478) );
  INV_X1 U15875 ( .A(n13816), .ZN(n14476) );
  NOR4_X1 U15876 ( .A1(n13818), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9143), .A4(
        P2_U3088), .ZN(n13819) );
  AOI21_X1 U15877 ( .B1(n13829), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13819), 
        .ZN(n13820) );
  OAI21_X1 U15878 ( .B1(n14476), .B2(n13837), .A(n13820), .ZN(P2_U3296) );
  AOI22_X1 U15879 ( .A1(n13821), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n13829), .ZN(n13822) );
  OAI21_X1 U15880 ( .B1(n14479), .B2(n13837), .A(n13822), .ZN(P2_U3297) );
  INV_X1 U15881 ( .A(n13823), .ZN(n14482) );
  OAI222_X1 U15882 ( .A1(n13839), .A2(n13824), .B1(n13837), .B2(n14482), .C1(
        n7378), .C2(P2_U3088), .ZN(P2_U3298) );
  INV_X1 U15883 ( .A(n13825), .ZN(n14484) );
  NAND2_X1 U15884 ( .A1(n13829), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13826) );
  OAI211_X1 U15885 ( .C1(n14484), .C2(n13837), .A(n13827), .B(n13826), .ZN(
        P2_U3299) );
  INV_X1 U15886 ( .A(n13828), .ZN(n14489) );
  AOI22_X1 U15887 ( .A1(n13830), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n13829), .ZN(n13831) );
  OAI21_X1 U15888 ( .B1(n14489), .B2(n13837), .A(n13831), .ZN(P2_U3300) );
  INV_X1 U15889 ( .A(n13832), .ZN(n14493) );
  OAI222_X1 U15890 ( .A1(n13834), .A2(P2_U3088), .B1(n13837), .B2(n14493), 
        .C1(n13833), .C2(n13839), .ZN(P2_U3301) );
  OAI222_X1 U15891 ( .A1(n13839), .A2(n13838), .B1(n13837), .B2(n13836), .C1(
        n13835), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15892 ( .A(n13840), .ZN(n13841) );
  MUX2_X1 U15893 ( .A(n13841), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15894 ( .A(n13844), .ZN(n14134) );
  NAND2_X1 U15895 ( .A1(n14239), .A2(n14018), .ZN(n13846) );
  NAND2_X1 U15896 ( .A1(n14019), .A2(n14238), .ZN(n13845) );
  AND2_X1 U15897 ( .A1(n13846), .A2(n13845), .ZN(n14131) );
  OAI22_X1 U15898 ( .A1(n13996), .A2(n14131), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13847), .ZN(n13848) );
  AOI21_X1 U15899 ( .B1(n13999), .B2(n14134), .A(n13848), .ZN(n13849) );
  INV_X1 U15900 ( .A(n13850), .ZN(n13851) );
  AOI21_X1 U15901 ( .B1(n13853), .B2(n13852), .A(n13851), .ZN(n13860) );
  NAND2_X1 U15902 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14768)
         );
  INV_X1 U15903 ( .A(n14768), .ZN(n13854) );
  AOI21_X1 U15904 ( .B1(n13950), .B2(n14026), .A(n13854), .ZN(n13856) );
  NAND2_X1 U15905 ( .A1(n14007), .A2(n14028), .ZN(n13855) );
  OAI211_X1 U15906 ( .C1(n14010), .C2(n13857), .A(n13856), .B(n13855), .ZN(
        n13858) );
  AOI21_X1 U15907 ( .B1(n14681), .B2(n14012), .A(n13858), .ZN(n13859) );
  OAI21_X1 U15908 ( .B1(n13860), .B2(n14014), .A(n13859), .ZN(P1_U3215) );
  NAND2_X1 U15909 ( .A1(n14239), .A2(n14021), .ZN(n13862) );
  NAND2_X1 U15910 ( .A1(n14224), .A2(n14238), .ZN(n13861) );
  NAND2_X1 U15911 ( .A1(n13862), .A2(n13861), .ZN(n14198) );
  AOI22_X1 U15912 ( .A1(n13863), .A2(n14198), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13864) );
  OAI21_X1 U15913 ( .B1(n14010), .B2(n14199), .A(n13864), .ZN(n13870) );
  NAND3_X1 U15914 ( .A1(n6940), .A2(n13866), .A3(n7731), .ZN(n13867) );
  AOI21_X1 U15915 ( .B1(n13868), .B2(n13867), .A(n14014), .ZN(n13869) );
  AOI211_X1 U15916 ( .C1(n14202), .C2(n14012), .A(n13870), .B(n13869), .ZN(
        n13871) );
  INV_X1 U15917 ( .A(n13871), .ZN(P1_U3216) );
  INV_X1 U15918 ( .A(n14265), .ZN(n14397) );
  INV_X1 U15919 ( .A(n13872), .ZN(n13875) );
  OAI21_X1 U15920 ( .B1(n13875), .B2(n13874), .A(n13873), .ZN(n13877) );
  NAND3_X1 U15921 ( .A1(n13877), .A2(n13991), .A3(n13876), .ZN(n13881) );
  NOR2_X1 U15922 ( .A1(n14010), .A2(n14266), .ZN(n13879) );
  NAND2_X1 U15923 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14074)
         );
  OAI21_X1 U15924 ( .B1(n14005), .B2(n14396), .A(n14074), .ZN(n13878) );
  AOI211_X1 U15925 ( .C1(n14007), .C2(n14023), .A(n13879), .B(n13878), .ZN(
        n13880) );
  OAI211_X1 U15926 ( .C1(n14397), .C2(n14002), .A(n13881), .B(n13880), .ZN(
        P1_U3219) );
  INV_X1 U15927 ( .A(n13882), .ZN(n13970) );
  AOI21_X1 U15928 ( .B1(n13884), .B2(n13883), .A(n13970), .ZN(n13889) );
  AOI22_X1 U15929 ( .A1(n13950), .A2(n14224), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13886) );
  NAND2_X1 U15930 ( .A1(n13999), .A2(n14229), .ZN(n13885) );
  OAI211_X1 U15931 ( .C1(n13944), .C2(n14396), .A(n13886), .B(n13885), .ZN(
        n13887) );
  AOI21_X1 U15932 ( .B1(n14386), .B2(n14012), .A(n13887), .ZN(n13888) );
  OAI21_X1 U15933 ( .B1(n13889), .B2(n14014), .A(n13888), .ZN(P1_U3223) );
  OAI21_X1 U15934 ( .B1(n13892), .B2(n13891), .A(n13890), .ZN(n13894) );
  NAND3_X1 U15935 ( .A1(n13894), .A2(n13991), .A3(n13893), .ZN(n13901) );
  NOR2_X1 U15936 ( .A1(n14010), .A2(n13895), .ZN(n13899) );
  NAND2_X1 U15937 ( .A1(n13950), .A2(n14028), .ZN(n13897) );
  NAND2_X1 U15938 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  AOI211_X1 U15939 ( .C1(n14007), .C2(n14031), .A(n13899), .B(n13898), .ZN(
        n13900) );
  OAI211_X1 U15940 ( .C1(n13902), .C2(n14002), .A(n13901), .B(n13900), .ZN(
        P1_U3224) );
  OAI21_X1 U15941 ( .B1(n13905), .B2(n13904), .A(n13903), .ZN(n13906) );
  NAND2_X1 U15942 ( .A1(n13906), .A2(n13991), .ZN(n13913) );
  INV_X1 U15943 ( .A(n14162), .ZN(n13911) );
  NAND2_X1 U15944 ( .A1(n14239), .A2(n14019), .ZN(n13908) );
  NAND2_X1 U15945 ( .A1(n14021), .A2(n14238), .ZN(n13907) );
  AND2_X1 U15946 ( .A1(n13908), .A2(n13907), .ZN(n14358) );
  OAI22_X1 U15947 ( .A1(n13996), .A2(n14358), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13909), .ZN(n13910) );
  AOI21_X1 U15948 ( .B1(n13999), .B2(n13911), .A(n13910), .ZN(n13912) );
  OAI211_X1 U15949 ( .C1(n7131), .C2(n14002), .A(n13913), .B(n13912), .ZN(
        P1_U3225) );
  XOR2_X1 U15950 ( .A(n13916), .B(n13914), .Z(n14004) );
  INV_X1 U15951 ( .A(n13915), .ZN(n14003) );
  INV_X1 U15952 ( .A(n13916), .ZN(n13917) );
  OAI22_X1 U15953 ( .A1(n14004), .A2(n14003), .B1(n13917), .B2(n13914), .ZN(
        n13920) );
  INV_X1 U15954 ( .A(n13918), .ZN(n13930) );
  AOI21_X1 U15955 ( .B1(n13920), .B2(n13919), .A(n13930), .ZN(n13926) );
  NAND2_X1 U15956 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14797)
         );
  INV_X1 U15957 ( .A(n14797), .ZN(n13921) );
  AOI21_X1 U15958 ( .B1(n13950), .B2(n14024), .A(n13921), .ZN(n13923) );
  NAND2_X1 U15959 ( .A1(n14007), .A2(n14026), .ZN(n13922) );
  OAI211_X1 U15960 ( .C1(n14010), .C2(n14322), .A(n13923), .B(n13922), .ZN(
        n13924) );
  AOI21_X1 U15961 ( .B1(n14413), .B2(n14012), .A(n13924), .ZN(n13925) );
  OAI21_X1 U15962 ( .B1(n13926), .B2(n14014), .A(n13925), .ZN(P1_U3226) );
  INV_X1 U15963 ( .A(n13927), .ZN(n13929) );
  NOR3_X1 U15964 ( .A1(n13930), .A2(n13929), .A3(n13928), .ZN(n13933) );
  INV_X1 U15965 ( .A(n13931), .ZN(n13932) );
  OAI21_X1 U15966 ( .B1(n13933), .B2(n13932), .A(n13991), .ZN(n13937) );
  NAND2_X1 U15967 ( .A1(n14007), .A2(n14025), .ZN(n13934) );
  NAND2_X1 U15968 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14812)
         );
  OAI211_X1 U15969 ( .C1(n14305), .C2(n14005), .A(n13934), .B(n14812), .ZN(
        n13935) );
  AOI21_X1 U15970 ( .B1(n14298), .B2(n13999), .A(n13935), .ZN(n13936) );
  OAI211_X1 U15971 ( .C1(n14301), .C2(n14002), .A(n13937), .B(n13936), .ZN(
        P1_U3228) );
  INV_X1 U15972 ( .A(n14185), .ZN(n14449) );
  OAI21_X1 U15973 ( .B1(n13940), .B2(n13939), .A(n13938), .ZN(n13941) );
  NAND2_X1 U15974 ( .A1(n13941), .A2(n13991), .ZN(n13947) );
  INV_X1 U15975 ( .A(n13942), .ZN(n14186) );
  AOI22_X1 U15976 ( .A1(n13950), .A2(n14020), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13943) );
  OAI21_X1 U15977 ( .B1(n14179), .B2(n13944), .A(n13943), .ZN(n13945) );
  AOI21_X1 U15978 ( .B1(n14186), .B2(n13999), .A(n13945), .ZN(n13946) );
  OAI211_X1 U15979 ( .C1(n14449), .C2(n14002), .A(n13947), .B(n13946), .ZN(
        P1_U3229) );
  XNOR2_X1 U15980 ( .A(n13949), .B(n13948), .ZN(n13956) );
  AOI22_X1 U15981 ( .A1(n13950), .A2(n14240), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13952) );
  NAND2_X1 U15982 ( .A1(n14007), .A2(n14237), .ZN(n13951) );
  OAI211_X1 U15983 ( .C1(n14010), .C2(n13953), .A(n13952), .B(n13951), .ZN(
        n13954) );
  AOI21_X1 U15984 ( .B1(n14251), .B2(n14012), .A(n13954), .ZN(n13955) );
  OAI21_X1 U15985 ( .B1(n13956), .B2(n14014), .A(n13955), .ZN(P1_U3233) );
  XNOR2_X1 U15986 ( .A(n13958), .B(n13957), .ZN(n13966) );
  NAND2_X1 U15987 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14755)
         );
  OAI21_X1 U15988 ( .B1(n14005), .B2(n13959), .A(n14755), .ZN(n13960) );
  AOI21_X1 U15989 ( .B1(n14007), .B2(n14029), .A(n13960), .ZN(n13961) );
  OAI21_X1 U15990 ( .B1(n14010), .B2(n13962), .A(n13961), .ZN(n13963) );
  AOI21_X1 U15991 ( .B1(n13964), .B2(n14012), .A(n13963), .ZN(n13965) );
  OAI21_X1 U15992 ( .B1(n13966), .B2(n14014), .A(n13965), .ZN(P1_U3234) );
  INV_X1 U15993 ( .A(n13967), .ZN(n13969) );
  NOR3_X1 U15994 ( .A1(n13970), .A2(n13969), .A3(n13968), .ZN(n13973) );
  INV_X1 U15995 ( .A(n6940), .ZN(n13972) );
  OAI21_X1 U15996 ( .B1(n13973), .B2(n13972), .A(n13991), .ZN(n13979) );
  INV_X1 U15997 ( .A(n14214), .ZN(n13977) );
  NOR2_X1 U15998 ( .A1(n14395), .A2(n14179), .ZN(n13974) );
  AOI21_X1 U15999 ( .B1(n14240), .B2(n14238), .A(n13974), .ZN(n14379) );
  INV_X1 U16000 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13975) );
  OAI22_X1 U16001 ( .A1(n13996), .A2(n14379), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13975), .ZN(n13976) );
  AOI21_X1 U16002 ( .B1(n13999), .B2(n13977), .A(n13976), .ZN(n13978) );
  OAI211_X1 U16003 ( .C1(n14002), .C2(n14454), .A(n13979), .B(n13978), .ZN(
        P1_U3235) );
  OAI21_X1 U16004 ( .B1(n13981), .B2(n13980), .A(n13872), .ZN(n13982) );
  NAND2_X1 U16005 ( .A1(n13982), .A2(n13991), .ZN(n13986) );
  NOR2_X1 U16006 ( .A1(n14010), .A2(n14286), .ZN(n13984) );
  NAND2_X1 U16007 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14830)
         );
  OAI21_X1 U16008 ( .B1(n14005), .B2(n14279), .A(n14830), .ZN(n13983) );
  AOI211_X1 U16009 ( .C1(n14007), .C2(n14024), .A(n13984), .B(n13983), .ZN(
        n13985) );
  OAI211_X1 U16010 ( .C1(n14464), .C2(n14002), .A(n13986), .B(n13985), .ZN(
        P1_U3238) );
  INV_X1 U16011 ( .A(n6884), .ZN(n14444) );
  OAI21_X1 U16012 ( .B1(n13990), .B2(n13989), .A(n13988), .ZN(n13992) );
  NAND2_X1 U16013 ( .A1(n13992), .A2(n13991), .ZN(n14001) );
  INV_X1 U16014 ( .A(n14148), .ZN(n13998) );
  NAND2_X1 U16015 ( .A1(n14239), .A2(n14104), .ZN(n13994) );
  NAND2_X1 U16016 ( .A1(n14020), .A2(n14238), .ZN(n13993) );
  AND2_X1 U16017 ( .A1(n13994), .A2(n13993), .ZN(n14351) );
  OAI22_X1 U16018 ( .A1(n13996), .A2(n14351), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13995), .ZN(n13997) );
  AOI21_X1 U16019 ( .B1(n13999), .B2(n13998), .A(n13997), .ZN(n14000) );
  OAI211_X1 U16020 ( .C1(n14444), .C2(n14002), .A(n14001), .B(n14000), .ZN(
        P1_U3240) );
  XNOR2_X1 U16021 ( .A(n14004), .B(n14003), .ZN(n14015) );
  NAND2_X1 U16022 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14782)
         );
  OAI21_X1 U16023 ( .B1(n14005), .B2(n14304), .A(n14782), .ZN(n14006) );
  AOI21_X1 U16024 ( .B1(n14007), .B2(n14027), .A(n14006), .ZN(n14008) );
  OAI21_X1 U16025 ( .B1(n14010), .B2(n14009), .A(n14008), .ZN(n14011) );
  AOI21_X1 U16026 ( .B1(n14421), .B2(n14012), .A(n14011), .ZN(n14013) );
  OAI21_X1 U16027 ( .B1(n14015), .B2(n14014), .A(n14013), .ZN(P1_U3241) );
  MUX2_X1 U16028 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14016), .S(n14042), .Z(
        P1_U3591) );
  MUX2_X1 U16029 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14017), .S(n14042), .Z(
        P1_U3590) );
  MUX2_X1 U16030 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14105), .S(n14042), .Z(
        P1_U3589) );
  MUX2_X1 U16031 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14018), .S(n14042), .Z(
        P1_U3588) );
  MUX2_X1 U16032 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14104), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16033 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14019), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16034 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14020), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16035 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14021), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16036 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14022), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16037 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14224), .S(n14042), .Z(
        P1_U3582) );
  MUX2_X1 U16038 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14240), .S(n14042), .Z(
        P1_U3581) );
  MUX2_X1 U16039 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14269), .S(n14042), .Z(
        P1_U3580) );
  MUX2_X1 U16040 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14237), .S(n14042), .Z(
        P1_U3579) );
  MUX2_X1 U16041 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14023), .S(n14042), .Z(
        P1_U3578) );
  MUX2_X1 U16042 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14024), .S(n14042), .Z(
        P1_U3577) );
  MUX2_X1 U16043 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14025), .S(n14042), .Z(
        P1_U3576) );
  MUX2_X1 U16044 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14026), .S(n14042), .Z(
        P1_U3575) );
  MUX2_X1 U16045 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14027), .S(n14042), .Z(
        P1_U3574) );
  MUX2_X1 U16046 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14028), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16047 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14029), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16048 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14031), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16049 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14032), .S(n14042), .Z(
        P1_U3570) );
  MUX2_X1 U16050 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14033), .S(n14042), .Z(
        P1_U3569) );
  MUX2_X1 U16051 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14034), .S(n14042), .Z(
        P1_U3568) );
  MUX2_X1 U16052 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14035), .S(n14042), .Z(
        P1_U3567) );
  MUX2_X1 U16053 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14036), .S(n14042), .Z(
        P1_U3566) );
  MUX2_X1 U16054 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14037), .S(n14042), .Z(
        P1_U3565) );
  MUX2_X1 U16055 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14038), .S(n14042), .Z(
        P1_U3564) );
  MUX2_X1 U16056 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n6871), .S(n14042), .Z(
        P1_U3563) );
  MUX2_X1 U16057 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14040), .S(n14042), .Z(
        P1_U3562) );
  MUX2_X1 U16058 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14041), .S(n14042), .Z(
        P1_U3561) );
  MUX2_X1 U16059 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14043), .S(n14042), .Z(
        P1_U3560) );
  NAND2_X1 U16060 ( .A1(n14795), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14044) );
  OAI21_X1 U16061 ( .B1(n14795), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14044), 
        .ZN(n14791) );
  OAI21_X1 U16062 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n14058), .A(n14045), 
        .ZN(n14751) );
  NAND2_X1 U16063 ( .A1(n14754), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n14046) );
  OAI21_X1 U16064 ( .B1(n14754), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14046), 
        .ZN(n14750) );
  NOR2_X1 U16065 ( .A1(n14751), .A2(n14750), .ZN(n14749) );
  MUX2_X1 U16066 ( .A(n14047), .B(P1_REG2_REG_14__SCAN_IN), .S(n14060), .Z(
        n14763) );
  NAND2_X1 U16067 ( .A1(n14048), .A2(n14780), .ZN(n14050) );
  XNOR2_X1 U16068 ( .A(n14780), .B(n14049), .ZN(n14776) );
  NOR2_X1 U16069 ( .A1(n14791), .A2(n14792), .ZN(n14790) );
  OR2_X1 U16070 ( .A1(n14063), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14052) );
  NAND2_X1 U16071 ( .A1(n14063), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14051) );
  NAND2_X1 U16072 ( .A1(n14052), .A2(n14051), .ZN(n14805) );
  NOR2_X1 U16073 ( .A1(n14806), .A2(n14805), .ZN(n14804) );
  NOR2_X1 U16074 ( .A1(n14053), .A2(n14827), .ZN(n14054) );
  XNOR2_X1 U16075 ( .A(n14827), .B(n14053), .ZN(n14822) );
  NOR2_X1 U16076 ( .A1(n14054), .A2(n14820), .ZN(n14055) );
  XNOR2_X1 U16077 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14055), .ZN(n14070) );
  XNOR2_X1 U16078 ( .A(n14795), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14787) );
  MUX2_X1 U16079 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14056), .S(n14060), .Z(
        n14759) );
  INV_X1 U16080 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14059) );
  MUX2_X1 U16081 ( .A(n14059), .B(P1_REG1_REG_13__SCAN_IN), .S(n14754), .Z(
        n14748) );
  NOR2_X1 U16082 ( .A1(n14747), .A2(n14748), .ZN(n14746) );
  NAND2_X1 U16083 ( .A1(n14759), .A2(n14760), .ZN(n14758) );
  NAND2_X1 U16084 ( .A1(n14780), .A2(n14061), .ZN(n14062) );
  NAND2_X1 U16085 ( .A1(n14773), .A2(n14772), .ZN(n14771) );
  NAND2_X1 U16086 ( .A1(n14062), .A2(n14771), .ZN(n14788) );
  NOR2_X1 U16087 ( .A1(n14787), .A2(n14788), .ZN(n14786) );
  XNOR2_X1 U16088 ( .A(n14063), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14801) );
  NOR2_X1 U16089 ( .A1(n14802), .A2(n14801), .ZN(n14800) );
  NOR2_X1 U16090 ( .A1(n14064), .A2(n14827), .ZN(n14065) );
  XNOR2_X1 U16091 ( .A(n14827), .B(n14064), .ZN(n14817) );
  NOR2_X1 U16092 ( .A1(n14065), .A2(n14815), .ZN(n14066) );
  XNOR2_X1 U16093 ( .A(n14066), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14069) );
  INV_X1 U16094 ( .A(n14069), .ZN(n14067) );
  NAND2_X1 U16095 ( .A1(n14067), .A2(n14819), .ZN(n14068) );
  AOI22_X1 U16096 ( .A1(n14070), .A2(n14824), .B1(n14819), .B2(n14069), .ZN(
        n14072) );
  NOR2_X1 U16097 ( .A1(n14309), .A2(n14338), .ZN(n14084) );
  NOR2_X1 U16098 ( .A1(n12194), .A2(n14300), .ZN(n14076) );
  AOI211_X1 U16099 ( .C1(n14309), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14084), 
        .B(n14076), .ZN(n14077) );
  OAI21_X1 U16100 ( .B1(n14078), .B2(n14253), .A(n14077), .ZN(P1_U3263) );
  AOI21_X1 U16101 ( .B1(n14431), .B2(n14079), .A(n14423), .ZN(n14080) );
  NAND2_X1 U16102 ( .A1(n14081), .A2(n14080), .ZN(n14339) );
  NOR2_X1 U16103 ( .A1(n14082), .A2(n14300), .ZN(n14083) );
  AOI211_X1 U16104 ( .C1(n14309), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14084), 
        .B(n14083), .ZN(n14085) );
  OAI21_X1 U16105 ( .B1(n14253), .B2(n14339), .A(n14085), .ZN(P1_U3264) );
  NAND2_X1 U16106 ( .A1(n14088), .A2(n14333), .ZN(n14096) );
  OAI22_X1 U16107 ( .A1(n14091), .A2(n14090), .B1(n14089), .B2(n14323), .ZN(
        n14094) );
  NOR2_X1 U16108 ( .A1(n14309), .A2(n14092), .ZN(n14093) );
  AOI211_X1 U16109 ( .C1(n14320), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14094), 
        .B(n14093), .ZN(n14095) );
  OAI211_X1 U16110 ( .C1(n14097), .C2(n14300), .A(n14096), .B(n14095), .ZN(
        n14098) );
  AOI21_X1 U16111 ( .B1(n14087), .B2(n14329), .A(n14098), .ZN(n14099) );
  OAI21_X1 U16112 ( .B1(n14100), .B2(n14220), .A(n14099), .ZN(P1_U3356) );
  OAI21_X1 U16113 ( .B1(n14107), .B2(n14102), .A(n14101), .ZN(n14103) );
  AOI22_X1 U16114 ( .A1(n14239), .A2(n14105), .B1(n14104), .B2(n14238), .ZN(
        n14106) );
  AND2_X1 U16115 ( .A1(n14108), .A2(n14107), .ZN(n14109) );
  INV_X1 U16116 ( .A(n14344), .ZN(n14119) );
  AOI21_X1 U16117 ( .B1(n14435), .B2(n14132), .A(n14423), .ZN(n14113) );
  NAND2_X1 U16118 ( .A1(n14113), .A2(n14112), .ZN(n14342) );
  NAND2_X1 U16119 ( .A1(n14320), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14114) );
  OAI21_X1 U16120 ( .B1(n14323), .B2(n14115), .A(n14114), .ZN(n14116) );
  AOI21_X1 U16121 ( .B1(n14435), .B2(n14325), .A(n14116), .ZN(n14117) );
  OAI21_X1 U16122 ( .B1(n14342), .B2(n14253), .A(n14117), .ZN(n14118) );
  AOI21_X1 U16123 ( .B1(n14119), .B2(n14329), .A(n14118), .ZN(n14120) );
  OAI21_X1 U16124 ( .B1(n14343), .B2(n14309), .A(n14120), .ZN(P1_U3265) );
  INV_X1 U16125 ( .A(n14122), .ZN(n14123) );
  INV_X1 U16126 ( .A(n14125), .ZN(n14129) );
  OAI21_X1 U16127 ( .B1(n14129), .B2(n14128), .A(n14688), .ZN(n14130) );
  AOI211_X1 U16128 ( .C1(n14133), .C2(n14146), .A(n14423), .B(n14111), .ZN(
        n14347) );
  AOI22_X1 U16129 ( .A1(n14320), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14134), 
        .B2(n14297), .ZN(n14135) );
  OAI21_X1 U16130 ( .B1(n14440), .B2(n14300), .A(n14135), .ZN(n14136) );
  AOI21_X1 U16131 ( .B1(n14347), .B2(n14333), .A(n14136), .ZN(n14137) );
  OAI211_X1 U16132 ( .C1(n14346), .C2(n14293), .A(n14138), .B(n14137), .ZN(
        P1_U3266) );
  INV_X1 U16133 ( .A(n14139), .ZN(n14143) );
  INV_X1 U16134 ( .A(n14140), .ZN(n14141) );
  AOI21_X1 U16135 ( .B1(n14143), .B2(n14142), .A(n14141), .ZN(n14353) );
  XNOR2_X1 U16136 ( .A(n14145), .B(n14144), .ZN(n14355) );
  NAND2_X1 U16137 ( .A1(n14355), .A2(n14329), .ZN(n14154) );
  INV_X1 U16138 ( .A(n14160), .ZN(n14147) );
  OAI211_X1 U16139 ( .C1(n14444), .C2(n14147), .A(n14248), .B(n14146), .ZN(
        n14350) );
  INV_X1 U16140 ( .A(n14350), .ZN(n14152) );
  OAI22_X1 U16141 ( .A1(n14320), .A2(n14351), .B1(n14148), .B2(n14323), .ZN(
        n14149) );
  AOI21_X1 U16142 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n14309), .A(n14149), 
        .ZN(n14150) );
  OAI21_X1 U16143 ( .B1(n14444), .B2(n14300), .A(n14150), .ZN(n14151) );
  AOI21_X1 U16144 ( .B1(n14152), .B2(n14333), .A(n14151), .ZN(n14153) );
  OAI211_X1 U16145 ( .C1(n14353), .C2(n14220), .A(n14154), .B(n14153), .ZN(
        P1_U3267) );
  OAI21_X1 U16146 ( .B1(n14156), .B2(n14157), .A(n14155), .ZN(n14361) );
  INV_X1 U16147 ( .A(n14361), .ZN(n14172) );
  INV_X1 U16148 ( .A(n14157), .ZN(n14159) );
  OAI21_X1 U16149 ( .B1(n14159), .B2(n6781), .A(n14158), .ZN(n14363) );
  INV_X1 U16150 ( .A(n14363), .ZN(n14170) );
  AOI21_X1 U16151 ( .B1(n14167), .B2(n14184), .A(n14423), .ZN(n14161) );
  NAND2_X1 U16152 ( .A1(n14161), .A2(n14160), .ZN(n14359) );
  OAI21_X1 U16153 ( .B1(n14323), .B2(n14162), .A(n14358), .ZN(n14163) );
  INV_X1 U16154 ( .A(n14163), .ZN(n14165) );
  NAND2_X1 U16155 ( .A1(n14320), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14164) );
  OAI21_X1 U16156 ( .B1(n14320), .B2(n14165), .A(n14164), .ZN(n14166) );
  AOI21_X1 U16157 ( .B1(n14167), .B2(n14325), .A(n14166), .ZN(n14168) );
  OAI21_X1 U16158 ( .B1(n14359), .B2(n14253), .A(n14168), .ZN(n14169) );
  AOI21_X1 U16159 ( .B1(n14170), .B2(n14329), .A(n14169), .ZN(n14171) );
  OAI21_X1 U16160 ( .B1(n14172), .B2(n14220), .A(n14171), .ZN(P1_U3268) );
  INV_X1 U16161 ( .A(n14173), .ZN(n14174) );
  AOI21_X1 U16162 ( .B1(n14177), .B2(n14175), .A(n14174), .ZN(n14364) );
  OAI21_X1 U16163 ( .B1(n14178), .B2(n14177), .A(n14176), .ZN(n14182) );
  OAI22_X1 U16164 ( .A1(n14180), .A2(n14395), .B1(n14179), .B2(n14316), .ZN(
        n14181) );
  AOI21_X1 U16165 ( .B1(n14182), .B2(n14688), .A(n14181), .ZN(n14183) );
  OAI21_X1 U16166 ( .B1(n14364), .B2(n14283), .A(n14183), .ZN(n14365) );
  NAND2_X1 U16167 ( .A1(n14365), .A2(n14319), .ZN(n14190) );
  AOI211_X1 U16168 ( .C1(n14185), .C2(n14196), .A(n14423), .B(n7132), .ZN(
        n14366) );
  AOI22_X1 U16169 ( .A1(n14320), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14186), 
        .B2(n14297), .ZN(n14187) );
  OAI21_X1 U16170 ( .B1(n14449), .B2(n14300), .A(n14187), .ZN(n14188) );
  AOI21_X1 U16171 ( .B1(n14366), .B2(n14333), .A(n14188), .ZN(n14189) );
  OAI211_X1 U16172 ( .C1(n14364), .C2(n14293), .A(n14190), .B(n14189), .ZN(
        P1_U3269) );
  OAI21_X1 U16173 ( .B1(n6722), .B2(n14192), .A(n14191), .ZN(n14376) );
  OAI21_X1 U16174 ( .B1(n14195), .B2(n14194), .A(n14193), .ZN(n14374) );
  OAI211_X1 U16175 ( .C1(n14213), .C2(n14372), .A(n14196), .B(n14248), .ZN(
        n14371) );
  NOR2_X1 U16176 ( .A1(n14319), .A2(n14197), .ZN(n14201) );
  INV_X1 U16177 ( .A(n14198), .ZN(n14370) );
  OAI22_X1 U16178 ( .A1(n14320), .A2(n14370), .B1(n14199), .B2(n14323), .ZN(
        n14200) );
  AOI211_X1 U16179 ( .C1(n14202), .C2(n14325), .A(n14201), .B(n14200), .ZN(
        n14203) );
  OAI21_X1 U16180 ( .B1(n14371), .B2(n14253), .A(n14203), .ZN(n14204) );
  AOI21_X1 U16181 ( .B1(n14374), .B2(n14205), .A(n14204), .ZN(n14206) );
  OAI21_X1 U16182 ( .B1(n14376), .B2(n14313), .A(n14206), .ZN(P1_U3270) );
  XNOR2_X1 U16183 ( .A(n14207), .B(n14209), .ZN(n14382) );
  INV_X1 U16184 ( .A(n14382), .ZN(n14221) );
  OAI21_X1 U16185 ( .B1(n14210), .B2(n14209), .A(n14208), .ZN(n14377) );
  AND2_X1 U16186 ( .A1(n14227), .A2(n14211), .ZN(n14212) );
  OR3_X1 U16187 ( .A1(n14213), .A2(n14212), .A3(n14423), .ZN(n14378) );
  OAI22_X1 U16188 ( .A1(n14320), .A2(n14379), .B1(n14214), .B2(n14323), .ZN(
        n14216) );
  NOR2_X1 U16189 ( .A1(n14454), .A2(n14300), .ZN(n14215) );
  AOI211_X1 U16190 ( .C1(n14320), .C2(P1_REG2_REG_22__SCAN_IN), .A(n14216), 
        .B(n14215), .ZN(n14217) );
  OAI21_X1 U16191 ( .B1(n14253), .B2(n14378), .A(n14217), .ZN(n14218) );
  AOI21_X1 U16192 ( .B1(n14377), .B2(n14329), .A(n14218), .ZN(n14219) );
  OAI21_X1 U16193 ( .B1(n14221), .B2(n14220), .A(n14219), .ZN(P1_U3271) );
  XNOR2_X1 U16194 ( .A(n14222), .B(n14225), .ZN(n14223) );
  AOI222_X1 U16195 ( .A1(n14269), .A2(n14238), .B1(n14224), .B2(n14239), .C1(
        n14688), .C2(n14223), .ZN(n14388) );
  XNOR2_X1 U16196 ( .A(n14226), .B(n14225), .ZN(n14389) );
  INV_X1 U16197 ( .A(n14389), .ZN(n14234) );
  INV_X1 U16198 ( .A(n14386), .ZN(n14232) );
  AOI21_X1 U16199 ( .B1(n14250), .B2(n14386), .A(n14423), .ZN(n14228) );
  AND2_X1 U16200 ( .A1(n14228), .A2(n14227), .ZN(n14385) );
  NAND2_X1 U16201 ( .A1(n14385), .A2(n14333), .ZN(n14231) );
  AOI22_X1 U16202 ( .A1(n14320), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14229), 
        .B2(n14297), .ZN(n14230) );
  OAI211_X1 U16203 ( .C1(n14232), .C2(n14300), .A(n14231), .B(n14230), .ZN(
        n14233) );
  AOI21_X1 U16204 ( .B1(n14234), .B2(n14329), .A(n14233), .ZN(n14235) );
  OAI21_X1 U16205 ( .B1(n14388), .B2(n14309), .A(n14235), .ZN(P1_U3272) );
  OAI211_X1 U16206 ( .C1(n6799), .C2(n14247), .A(n14236), .B(n14688), .ZN(
        n14242) );
  AOI22_X1 U16207 ( .A1(n14240), .A2(n14239), .B1(n14238), .B2(n14237), .ZN(
        n14241) );
  NAND2_X1 U16208 ( .A1(n14242), .A2(n14241), .ZN(n14390) );
  AOI21_X1 U16209 ( .B1(n14243), .B2(n14297), .A(n14390), .ZN(n14257) );
  INV_X1 U16210 ( .A(n14244), .ZN(n14245) );
  AOI21_X1 U16211 ( .B1(n14247), .B2(n14246), .A(n14245), .ZN(n14392) );
  OR2_X1 U16212 ( .A1(n6897), .A2(n14264), .ZN(n14249) );
  AND3_X1 U16213 ( .A1(n14250), .A2(n14249), .A3(n14248), .ZN(n14391) );
  INV_X1 U16214 ( .A(n14391), .ZN(n14254) );
  AOI22_X1 U16215 ( .A1(n14251), .A2(n14325), .B1(n14320), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14252) );
  OAI21_X1 U16216 ( .B1(n14254), .B2(n14253), .A(n14252), .ZN(n14255) );
  AOI21_X1 U16217 ( .B1(n14392), .B2(n14329), .A(n14255), .ZN(n14256) );
  OAI21_X1 U16218 ( .B1(n14309), .B2(n14257), .A(n14256), .ZN(P1_U3273) );
  XNOR2_X1 U16219 ( .A(n14258), .B(n8324), .ZN(n14402) );
  INV_X1 U16220 ( .A(n14259), .ZN(n14260) );
  AOI21_X1 U16221 ( .B1(n14262), .B2(n14261), .A(n14260), .ZN(n14263) );
  OAI22_X1 U16222 ( .A1(n14263), .A2(n14352), .B1(n14305), .B2(n14316), .ZN(
        n14400) );
  AOI211_X1 U16223 ( .C1(n14265), .C2(n14284), .A(n14423), .B(n14264), .ZN(
        n14399) );
  NAND2_X1 U16224 ( .A1(n14399), .A2(n14333), .ZN(n14272) );
  INV_X1 U16225 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14267) );
  OAI22_X1 U16226 ( .A1(n14319), .A2(n14267), .B1(n14266), .B2(n14323), .ZN(
        n14268) );
  AOI21_X1 U16227 ( .B1(n14270), .B2(n14269), .A(n14268), .ZN(n14271) );
  OAI211_X1 U16228 ( .C1(n14397), .C2(n14300), .A(n14272), .B(n14271), .ZN(
        n14273) );
  AOI21_X1 U16229 ( .B1(n14400), .B2(n14319), .A(n14273), .ZN(n14274) );
  OAI21_X1 U16230 ( .B1(n14402), .B2(n14313), .A(n14274), .ZN(P1_U3274) );
  INV_X1 U16231 ( .A(n14278), .ZN(n14275) );
  XNOR2_X1 U16232 ( .A(n14276), .B(n14275), .ZN(n14403) );
  XOR2_X1 U16233 ( .A(n14277), .B(n14278), .Z(n14281) );
  OAI22_X1 U16234 ( .A1(n14279), .A2(n14395), .B1(n14318), .B2(n14316), .ZN(
        n14280) );
  AOI21_X1 U16235 ( .B1(n14281), .B2(n14688), .A(n14280), .ZN(n14282) );
  OAI21_X1 U16236 ( .B1(n14403), .B2(n14283), .A(n14282), .ZN(n14404) );
  INV_X1 U16237 ( .A(n14284), .ZN(n14285) );
  AOI211_X1 U16238 ( .C1(n14290), .C2(n7130), .A(n14423), .B(n14285), .ZN(
        n14405) );
  INV_X1 U16239 ( .A(n14405), .ZN(n14288) );
  OAI22_X1 U16240 ( .A1(n14288), .A2(n14287), .B1(n14323), .B2(n14286), .ZN(
        n14289) );
  OAI21_X1 U16241 ( .B1(n14404), .B2(n14289), .A(n14319), .ZN(n14292) );
  AOI22_X1 U16242 ( .A1(n14290), .A2(n14325), .B1(P1_REG2_REG_18__SCAN_IN), 
        .B2(n14309), .ZN(n14291) );
  OAI211_X1 U16243 ( .C1(n14403), .C2(n14293), .A(n14292), .B(n14291), .ZN(
        P1_U3275) );
  XNOR2_X1 U16244 ( .A(n14295), .B(n14294), .ZN(n14412) );
  AOI211_X1 U16245 ( .C1(n14409), .C2(n14332), .A(n14423), .B(n14296), .ZN(
        n14408) );
  AOI22_X1 U16246 ( .A1(n14320), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14298), 
        .B2(n14297), .ZN(n14299) );
  OAI21_X1 U16247 ( .B1(n14301), .B2(n14300), .A(n14299), .ZN(n14311) );
  AOI21_X1 U16248 ( .B1(n14303), .B2(n14302), .A(n14352), .ZN(n14308) );
  OAI22_X1 U16249 ( .A1(n14305), .A2(n14395), .B1(n14304), .B2(n14316), .ZN(
        n14306) );
  AOI21_X1 U16250 ( .B1(n14308), .B2(n14307), .A(n14306), .ZN(n14411) );
  NOR2_X1 U16251 ( .A1(n14411), .A2(n14309), .ZN(n14310) );
  AOI211_X1 U16252 ( .C1(n14408), .C2(n14333), .A(n14311), .B(n14310), .ZN(
        n14312) );
  OAI21_X1 U16253 ( .B1(n14313), .B2(n14412), .A(n14312), .ZN(P1_U3276) );
  XOR2_X1 U16254 ( .A(n14314), .B(n14327), .Z(n14317) );
  OAI222_X1 U16255 ( .A1(n14395), .A2(n14318), .B1(n14317), .B2(n14352), .C1(
        n14316), .C2(n14315), .ZN(n14414) );
  NAND2_X1 U16256 ( .A1(n14414), .A2(n14319), .ZN(n14337) );
  NAND2_X1 U16257 ( .A1(n14320), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14321) );
  OAI21_X1 U16258 ( .B1(n14323), .B2(n14322), .A(n14321), .ZN(n14324) );
  AOI21_X1 U16259 ( .B1(n14413), .B2(n14325), .A(n14324), .ZN(n14336) );
  OAI21_X1 U16260 ( .B1(n14328), .B2(n14327), .A(n14326), .ZN(n14416) );
  NAND2_X1 U16261 ( .A1(n14416), .A2(n14329), .ZN(n14335) );
  AOI21_X1 U16262 ( .B1(n14330), .B2(n14413), .A(n14423), .ZN(n14331) );
  AND2_X1 U16263 ( .A1(n14332), .A2(n14331), .ZN(n14415) );
  NAND2_X1 U16264 ( .A1(n14415), .A2(n14333), .ZN(n14334) );
  NAND4_X1 U16265 ( .A1(n14337), .A2(n14336), .A3(n14335), .A4(n14334), .ZN(
        P1_U3277) );
  NAND2_X1 U16266 ( .A1(n14339), .A2(n14338), .ZN(n14429) );
  MUX2_X1 U16267 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14429), .S(n14863), .Z(
        n14340) );
  AOI21_X1 U16268 ( .B1(n14345), .B2(n14431), .A(n14340), .ZN(n14341) );
  INV_X1 U16269 ( .A(n14341), .ZN(P1_U3558) );
  INV_X1 U16270 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14349) );
  INV_X1 U16271 ( .A(n14346), .ZN(n14348) );
  INV_X1 U16272 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n14356) );
  OAI211_X1 U16273 ( .C1(n14353), .C2(n14352), .A(n14351), .B(n14350), .ZN(
        n14354) );
  AOI21_X1 U16274 ( .B1(n14855), .B2(n14355), .A(n14354), .ZN(n14441) );
  MUX2_X1 U16275 ( .A(n14356), .B(n14441), .S(n14863), .Z(n14357) );
  OAI21_X1 U16276 ( .B1(n14444), .B2(n14419), .A(n14357), .ZN(P1_U3554) );
  OAI211_X1 U16277 ( .C1(n7131), .C2(n14852), .A(n14359), .B(n14358), .ZN(
        n14360) );
  AOI21_X1 U16278 ( .B1(n14361), .B2(n14688), .A(n14360), .ZN(n14362) );
  OAI21_X1 U16279 ( .B1(n14363), .B2(n14684), .A(n14362), .ZN(n14445) );
  MUX2_X1 U16280 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14445), .S(n14863), .Z(
        P1_U3553) );
  INV_X1 U16281 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14368) );
  INV_X1 U16282 ( .A(n14364), .ZN(n14367) );
  AOI211_X1 U16283 ( .C1(n14842), .C2(n14367), .A(n14366), .B(n14365), .ZN(
        n14446) );
  MUX2_X1 U16284 ( .A(n14368), .B(n14446), .S(n14863), .Z(n14369) );
  OAI21_X1 U16285 ( .B1(n14449), .B2(n14419), .A(n14369), .ZN(P1_U3552) );
  OAI211_X1 U16286 ( .C1(n14372), .C2(n14852), .A(n14371), .B(n14370), .ZN(
        n14373) );
  AOI21_X1 U16287 ( .B1(n14374), .B2(n14688), .A(n14373), .ZN(n14375) );
  OAI21_X1 U16288 ( .B1(n14376), .B2(n14684), .A(n14375), .ZN(n14450) );
  MUX2_X1 U16289 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14450), .S(n14863), .Z(
        P1_U3551) );
  INV_X1 U16290 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n14383) );
  INV_X1 U16291 ( .A(n14377), .ZN(n14380) );
  OAI211_X1 U16292 ( .C1(n14380), .C2(n14684), .A(n14379), .B(n14378), .ZN(
        n14381) );
  AOI21_X1 U16293 ( .B1(n14688), .B2(n14382), .A(n14381), .ZN(n14451) );
  MUX2_X1 U16294 ( .A(n14383), .B(n14451), .S(n14863), .Z(n14384) );
  OAI21_X1 U16295 ( .B1(n14419), .B2(n14454), .A(n14384), .ZN(P1_U3550) );
  AOI21_X1 U16296 ( .B1(n14386), .B2(n14680), .A(n14385), .ZN(n14387) );
  OAI211_X1 U16297 ( .C1(n14684), .C2(n14389), .A(n14388), .B(n14387), .ZN(
        n14455) );
  MUX2_X1 U16298 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14455), .S(n14863), .Z(
        P1_U3549) );
  AOI211_X1 U16299 ( .C1(n14392), .C2(n14855), .A(n14391), .B(n14390), .ZN(
        n14456) );
  MUX2_X1 U16300 ( .A(n14393), .B(n14456), .S(n14863), .Z(n14394) );
  OAI21_X1 U16301 ( .B1(n6897), .B2(n14419), .A(n14394), .ZN(P1_U3548) );
  OAI22_X1 U16302 ( .A1(n14397), .A2(n14852), .B1(n14396), .B2(n14395), .ZN(
        n14398) );
  NOR3_X1 U16303 ( .A1(n14400), .A2(n14399), .A3(n14398), .ZN(n14401) );
  OAI21_X1 U16304 ( .B1(n14684), .B2(n14402), .A(n14401), .ZN(n14460) );
  MUX2_X1 U16305 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14460), .S(n14863), .Z(
        P1_U3547) );
  INV_X1 U16306 ( .A(n14403), .ZN(n14406) );
  AOI211_X1 U16307 ( .C1(n14842), .C2(n14406), .A(n14405), .B(n14404), .ZN(
        n14461) );
  MUX2_X1 U16308 ( .A(n14816), .B(n14461), .S(n14863), .Z(n14407) );
  OAI21_X1 U16309 ( .B1(n14464), .B2(n14419), .A(n14407), .ZN(P1_U3546) );
  AOI21_X1 U16310 ( .B1(n14409), .B2(n14680), .A(n14408), .ZN(n14410) );
  OAI211_X1 U16311 ( .C1(n14412), .C2(n14684), .A(n14411), .B(n14410), .ZN(
        n14465) );
  MUX2_X1 U16312 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14465), .S(n14863), .Z(
        P1_U3545) );
  INV_X1 U16313 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14417) );
  AOI211_X1 U16314 ( .C1(n14855), .C2(n14416), .A(n14415), .B(n14414), .ZN(
        n14466) );
  MUX2_X1 U16315 ( .A(n14417), .B(n14466), .S(n14863), .Z(n14418) );
  OAI21_X1 U16316 ( .B1(n7129), .B2(n14419), .A(n14418), .ZN(P1_U3544) );
  AOI21_X1 U16317 ( .B1(n14421), .B2(n14680), .A(n14420), .ZN(n14422) );
  OAI21_X1 U16318 ( .B1(n14424), .B2(n14423), .A(n14422), .ZN(n14425) );
  AOI21_X1 U16319 ( .B1(n14426), .B2(n14688), .A(n14425), .ZN(n14427) );
  OAI21_X1 U16320 ( .B1(n14428), .B2(n14684), .A(n14427), .ZN(n14470) );
  MUX2_X1 U16321 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14470), .S(n14863), .Z(
        P1_U3543) );
  MUX2_X1 U16322 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14429), .S(n14857), .Z(
        n14430) );
  AOI21_X1 U16323 ( .B1(n14436), .B2(n14431), .A(n14430), .ZN(n14432) );
  INV_X1 U16324 ( .A(n14432), .ZN(P1_U3526) );
  AOI21_X1 U16325 ( .B1(n14436), .B2(n14435), .A(n14434), .ZN(n14437) );
  INV_X1 U16326 ( .A(n14437), .ZN(P1_U3524) );
  INV_X1 U16327 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14439) );
  INV_X1 U16328 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n14442) );
  MUX2_X1 U16329 ( .A(n14442), .B(n14441), .S(n14857), .Z(n14443) );
  OAI21_X1 U16330 ( .B1(n14444), .B2(n14469), .A(n14443), .ZN(P1_U3522) );
  MUX2_X1 U16331 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14445), .S(n14857), .Z(
        P1_U3521) );
  INV_X1 U16332 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14447) );
  MUX2_X1 U16333 ( .A(n14447), .B(n14446), .S(n14857), .Z(n14448) );
  OAI21_X1 U16334 ( .B1(n14449), .B2(n14469), .A(n14448), .ZN(P1_U3520) );
  MUX2_X1 U16335 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14450), .S(n14857), .Z(
        P1_U3519) );
  INV_X1 U16336 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n14452) );
  MUX2_X1 U16337 ( .A(n14452), .B(n14451), .S(n14857), .Z(n14453) );
  OAI21_X1 U16338 ( .B1(n14469), .B2(n14454), .A(n14453), .ZN(P1_U3518) );
  MUX2_X1 U16339 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14455), .S(n14857), .Z(
        P1_U3517) );
  INV_X1 U16340 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14457) );
  MUX2_X1 U16341 ( .A(n14457), .B(n14456), .S(n14857), .Z(n14458) );
  OAI21_X1 U16342 ( .B1(n6897), .B2(n14469), .A(n14458), .ZN(P1_U3516) );
  MUX2_X1 U16343 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14460), .S(n14857), .Z(
        P1_U3515) );
  INV_X1 U16344 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14462) );
  MUX2_X1 U16345 ( .A(n14462), .B(n14461), .S(n14857), .Z(n14463) );
  OAI21_X1 U16346 ( .B1(n14464), .B2(n14469), .A(n14463), .ZN(P1_U3513) );
  MUX2_X1 U16347 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14465), .S(n14857), .Z(
        P1_U3510) );
  INV_X1 U16348 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14467) );
  MUX2_X1 U16349 ( .A(n14467), .B(n14466), .S(n14857), .Z(n14468) );
  OAI21_X1 U16350 ( .B1(n7129), .B2(n14469), .A(n14468), .ZN(P1_U3507) );
  MUX2_X1 U16351 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14470), .S(n14857), .Z(
        P1_U3504) );
  INV_X1 U16352 ( .A(n14471), .ZN(n14472) );
  NOR4_X1 U16353 ( .A1(n14472), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n8290), .ZN(n14473) );
  AOI21_X1 U16354 ( .B1(n14474), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14473), 
        .ZN(n14475) );
  OAI21_X1 U16355 ( .B1(n14476), .B2(n14494), .A(n14475), .ZN(P1_U3324) );
  OAI222_X1 U16356 ( .A1(n14494), .A2(n14479), .B1(n14477), .B2(P1_U3086), 
        .C1(n14478), .C2(n14486), .ZN(P1_U3325) );
  OAI222_X1 U16357 ( .A1(n14494), .A2(n14482), .B1(n14481), .B2(P1_U3086), 
        .C1(n14480), .C2(n14490), .ZN(P1_U3326) );
  OAI222_X1 U16358 ( .A1(n14486), .A2(n14485), .B1(n14494), .B2(n14484), .C1(
        P1_U3086), .C2(n14483), .ZN(P1_U3327) );
  OAI222_X1 U16359 ( .A1(n14494), .A2(n14489), .B1(n14488), .B2(P1_U3086), 
        .C1(n14487), .C2(n14490), .ZN(P1_U3328) );
  OAI222_X1 U16360 ( .A1(n14494), .A2(n14493), .B1(P1_U3086), .B2(n14492), 
        .C1(n14491), .C2(n14490), .ZN(P1_U3329) );
  MUX2_X1 U16361 ( .A(n14496), .B(n14495), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16362 ( .A(n14497), .ZN(n14498) );
  MUX2_X1 U16363 ( .A(n14498), .B(n6889), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U16364 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15045) );
  INV_X1 U16365 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15027) );
  INV_X1 U16366 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14784) );
  OR2_X1 U16367 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14784), .ZN(n14527) );
  INV_X1 U16368 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14770) );
  XNOR2_X1 U16369 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14529) );
  INV_X1 U16370 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14757) );
  INV_X1 U16371 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15208) );
  XNOR2_X1 U16372 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n14572) );
  INV_X1 U16373 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14521) );
  XNOR2_X1 U16374 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P3_ADDR_REG_11__SCAN_IN), 
        .ZN(n14569) );
  INV_X1 U16375 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14516) );
  INV_X1 U16376 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15187) );
  XNOR2_X1 U16377 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), 
        .ZN(n14563) );
  INV_X1 U16378 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15687) );
  XNOR2_X1 U16379 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n14557) );
  INV_X1 U16380 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15500) );
  XOR2_X1 U16381 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n15500), .Z(n14550) );
  XNOR2_X1 U16382 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14534) );
  NAND2_X1 U16383 ( .A1(n14536), .A2(n14535), .ZN(n14499) );
  NAND2_X1 U16384 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14502), .ZN(n14503) );
  NAND2_X1 U16385 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14504), .ZN(n14506) );
  NAND2_X1 U16386 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14507), .ZN(n14509) );
  INV_X1 U16387 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14544) );
  NAND2_X1 U16388 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14511), .ZN(n14513) );
  XNOR2_X1 U16389 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14511), .ZN(n14554) );
  NAND2_X1 U16390 ( .A1(n14557), .A2(n14558), .ZN(n14514) );
  NAND2_X1 U16391 ( .A1(n14563), .A2(n14562), .ZN(n14515) );
  NAND2_X1 U16392 ( .A1(n14516), .A2(n14517), .ZN(n14519) );
  XNOR2_X1 U16393 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14517), .ZN(n14566) );
  NAND2_X1 U16394 ( .A1(n14566), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n14518) );
  NAND2_X1 U16395 ( .A1(n14569), .A2(n14568), .ZN(n14520) );
  NAND2_X1 U16396 ( .A1(n14572), .A2(n14571), .ZN(n14522) );
  INV_X1 U16397 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14523) );
  NAND2_X1 U16398 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14523), .ZN(n14524) );
  AOI22_X1 U16399 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14757), .B1(n14530), 
        .B2(n14524), .ZN(n14528) );
  NAND2_X1 U16400 ( .A1(n14529), .A2(n14528), .ZN(n14525) );
  OAI21_X1 U16401 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14770), .A(n14525), 
        .ZN(n14526) );
  INV_X1 U16402 ( .A(n14526), .ZN(n14577) );
  AOI22_X1 U16403 ( .A1(n14784), .A2(P3_ADDR_REG_15__SCAN_IN), .B1(n14527), 
        .B2(n14577), .ZN(n14581) );
  XNOR2_X1 U16404 ( .A(n14581), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n14582) );
  XOR2_X1 U16405 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n14582), .Z(n14723) );
  INV_X1 U16406 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15010) );
  INV_X1 U16407 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14998) );
  XOR2_X1 U16408 ( .A(n14529), .B(n14528), .Z(n14715) );
  INV_X1 U16409 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14985) );
  XNOR2_X1 U16410 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n14531) );
  XNOR2_X1 U16411 ( .A(n14531), .B(n14530), .ZN(n14711) );
  INV_X1 U16412 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14707) );
  INV_X1 U16413 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14970) );
  NAND2_X1 U16414 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14541), .ZN(n14542) );
  INV_X1 U16415 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15796) );
  INV_X1 U16416 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14597) );
  XNOR2_X1 U16417 ( .A(n14534), .B(n14533), .ZN(n14595) );
  NAND2_X1 U16418 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14537), .ZN(n14538) );
  AOI21_X1 U16419 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15514), .A(n14536), .ZN(
        n15790) );
  INV_X1 U16420 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15789) );
  NOR2_X1 U16421 ( .A1(n15790), .A2(n15789), .ZN(n15799) );
  XNOR2_X1 U16422 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14539), .ZN(n15794) );
  NAND2_X1 U16423 ( .A1(n15795), .A2(n15794), .ZN(n14540) );
  NOR2_X1 U16424 ( .A1(n15795), .A2(n15794), .ZN(n15793) );
  INV_X1 U16425 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14904) );
  XNOR2_X1 U16426 ( .A(n14541), .B(n14904), .ZN(n15786) );
  NOR2_X1 U16427 ( .A1(n14546), .A2(n14545), .ZN(n14548) );
  XNOR2_X1 U16428 ( .A(n14545), .B(n14546), .ZN(n15788) );
  NOR2_X1 U16429 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15788), .ZN(n14547) );
  NAND2_X1 U16430 ( .A1(n14549), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14552) );
  XNOR2_X1 U16431 ( .A(n14551), .B(n14550), .ZN(n14599) );
  NOR2_X1 U16432 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14553), .ZN(n14556) );
  XNOR2_X1 U16433 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14554), .ZN(n15791) );
  NOR2_X1 U16434 ( .A1(n15792), .A2(n15791), .ZN(n14555) );
  XNOR2_X1 U16435 ( .A(n14558), .B(n14557), .ZN(n14560) );
  NAND2_X1 U16436 ( .A1(n14559), .A2(n14560), .ZN(n14561) );
  XNOR2_X1 U16437 ( .A(n14563), .B(n14562), .ZN(n14603) );
  NOR2_X1 U16438 ( .A1(n14604), .A2(n14603), .ZN(n14565) );
  INV_X1 U16439 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14564) );
  NAND2_X1 U16440 ( .A1(n14604), .A2(n14603), .ZN(n14602) );
  OAI21_X2 U16441 ( .B1(n14565), .B2(n14564), .A(n14602), .ZN(n14607) );
  XNOR2_X1 U16442 ( .A(n14566), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14608) );
  NAND2_X1 U16443 ( .A1(n14607), .A2(n14608), .ZN(n14567) );
  NOR2_X1 U16444 ( .A1(n14607), .A2(n14608), .ZN(n14606) );
  XNOR2_X1 U16445 ( .A(n14569), .B(n14568), .ZN(n14705) );
  NAND2_X1 U16446 ( .A1(n14706), .A2(n14705), .ZN(n14570) );
  XNOR2_X1 U16447 ( .A(n14572), .B(n14571), .ZN(n14574) );
  NAND2_X1 U16448 ( .A1(n14711), .A2(n14712), .ZN(n14575) );
  AOI21_X2 U16449 ( .B1(n14985), .B2(n14575), .A(n14710), .ZN(n14716) );
  NAND2_X1 U16450 ( .A1(n14715), .A2(n14716), .ZN(n14576) );
  XNOR2_X1 U16451 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n14578) );
  XNOR2_X1 U16452 ( .A(n14578), .B(n14577), .ZN(n14719) );
  NAND2_X1 U16453 ( .A1(n14720), .A2(n14719), .ZN(n14579) );
  AOI21_X2 U16454 ( .B1(n15010), .B2(n14579), .A(n14718), .ZN(n14724) );
  NAND2_X1 U16455 ( .A1(n14723), .A2(n14724), .ZN(n14580) );
  AND2_X1 U16456 ( .A1(n14581), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14584) );
  NOR2_X1 U16457 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14582), .ZN(n14583) );
  NOR2_X1 U16458 ( .A1(n14584), .A2(n14583), .ZN(n14586) );
  XNOR2_X1 U16459 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14586), .ZN(n14587) );
  XNOR2_X1 U16460 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14587), .ZN(n14611) );
  NAND2_X1 U16461 ( .A1(n14612), .A2(n14611), .ZN(n14585) );
  NOR2_X1 U16462 ( .A1(n14612), .A2(n14611), .ZN(n14610) );
  XNOR2_X1 U16463 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n14590) );
  INV_X1 U16464 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14814) );
  NAND2_X1 U16465 ( .A1(n14586), .A2(n14814), .ZN(n14589) );
  NAND2_X1 U16466 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14587), .ZN(n14588) );
  NAND2_X1 U16467 ( .A1(n14589), .A2(n14588), .ZN(n15398) );
  XOR2_X1 U16468 ( .A(n14590), .B(n15398), .Z(n14591) );
  AOI21_X1 U16469 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14593) );
  OAI21_X1 U16470 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14593), 
        .ZN(U28) );
  INV_X1 U16471 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15682) );
  OAI221_X1 U16472 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7035), .C2(n7771), .A(n15682), .ZN(U29) );
  AOI21_X1 U16473 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n14598) );
  XNOR2_X1 U16474 ( .A(n14598), .B(n14597), .ZN(SUB_1596_U61) );
  XOR2_X1 U16475 ( .A(n14600), .B(n14599), .Z(SUB_1596_U57) );
  INV_X1 U16476 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14955) );
  XNOR2_X1 U16477 ( .A(n14601), .B(n14955), .ZN(SUB_1596_U55) );
  OAI21_X1 U16478 ( .B1(n14604), .B2(n14603), .A(n14602), .ZN(n14605) );
  XNOR2_X1 U16479 ( .A(n14605), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  AOI21_X1 U16480 ( .B1(n14608), .B2(n14607), .A(n14606), .ZN(n14609) );
  XNOR2_X1 U16481 ( .A(n14609), .B(n14970), .ZN(SUB_1596_U70) );
  AOI21_X1 U16482 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14613) );
  XNOR2_X1 U16483 ( .A(n14613), .B(n15045), .ZN(SUB_1596_U63) );
  AOI21_X1 U16484 ( .B1(n14616), .B2(n14615), .A(n14614), .ZN(n14633) );
  INV_X1 U16485 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14619) );
  INV_X1 U16486 ( .A(n14617), .ZN(n14618) );
  OAI21_X1 U16487 ( .B1(n15251), .B2(n14619), .A(n14618), .ZN(n14625) );
  AOI21_X1 U16488 ( .B1(n14622), .B2(n14621), .A(n14620), .ZN(n14623) );
  NOR2_X1 U16489 ( .A1(n14623), .A2(n15253), .ZN(n14624) );
  AOI211_X1 U16490 ( .C1(n15259), .C2(n14626), .A(n14625), .B(n14624), .ZN(
        n14632) );
  AOI21_X1 U16491 ( .B1(n14629), .B2(n14628), .A(n14627), .ZN(n14630) );
  OR2_X1 U16492 ( .A1(n15241), .A2(n14630), .ZN(n14631) );
  OAI211_X1 U16493 ( .C1(n14633), .C2(n15266), .A(n14632), .B(n14631), .ZN(
        P3_U3197) );
  XNOR2_X1 U16494 ( .A(n14634), .B(n14637), .ZN(n14659) );
  INV_X1 U16495 ( .A(n14649), .ZN(n15317) );
  NAND2_X1 U16496 ( .A1(n6676), .A2(n14635), .ZN(n14636) );
  XOR2_X1 U16497 ( .A(n14637), .B(n14636), .Z(n14638) );
  OAI222_X1 U16498 ( .A1(n15315), .A2(n14640), .B1(n15313), .B2(n14639), .C1(
        n14638), .C2(n15311), .ZN(n14657) );
  AOI21_X1 U16499 ( .B1(n14659), .B2(n15317), .A(n14657), .ZN(n14645) );
  NOR2_X1 U16500 ( .A1(n14641), .A2(n15339), .ZN(n14658) );
  INV_X1 U16501 ( .A(n14642), .ZN(n14643) );
  AOI22_X1 U16502 ( .A1(n14658), .A2(n15295), .B1(n15332), .B2(n14643), .ZN(
        n14644) );
  OAI221_X1 U16503 ( .B1(n15337), .B2(n14645), .C1(n15335), .C2(n8694), .A(
        n14644), .ZN(P3_U3220) );
  INV_X1 U16504 ( .A(n14646), .ZN(n14648) );
  OAI21_X1 U16505 ( .B1(n14649), .B2(n14648), .A(n14647), .ZN(n14654) );
  OAI22_X1 U16506 ( .A1(n14652), .A2(n14651), .B1(n15335), .B2(n14650), .ZN(
        n14653) );
  AOI21_X1 U16507 ( .B1(n14654), .B2(n15335), .A(n14653), .ZN(n14655) );
  OAI21_X1 U16508 ( .B1(n14656), .B2(n15307), .A(n14655), .ZN(P3_U3222) );
  AOI211_X1 U16509 ( .C1(n14659), .C2(n15368), .A(n14658), .B(n14657), .ZN(
        n14664) );
  AOI22_X1 U16510 ( .A1(n15396), .A2(n14664), .B1(n8695), .B2(n15394), .ZN(
        P3_U3472) );
  AOI211_X1 U16511 ( .C1(n14662), .C2(n15368), .A(n14661), .B(n14660), .ZN(
        n14665) );
  AOI22_X1 U16512 ( .A1(n15396), .A2(n14665), .B1(n12646), .B2(n15394), .ZN(
        P3_U3471) );
  INV_X1 U16513 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14663) );
  AOI22_X1 U16514 ( .A1(n15382), .A2(n14664), .B1(n14663), .B2(n9009), .ZN(
        P3_U3429) );
  AOI22_X1 U16515 ( .A1(n15382), .A2(n14665), .B1(n8671), .B2(n9009), .ZN(
        P3_U3426) );
  OAI211_X1 U16516 ( .C1(n14668), .C2(n15111), .A(n14667), .B(n14666), .ZN(
        n14669) );
  AOI21_X1 U16517 ( .B1(n14670), .B2(n15099), .A(n14669), .ZN(n14676) );
  AOI22_X1 U16518 ( .A1(n15129), .A2(n14676), .B1(n11668), .B2(n15127), .ZN(
        P2_U3512) );
  OAI211_X1 U16519 ( .C1(n7228), .C2(n15111), .A(n14672), .B(n14671), .ZN(
        n14673) );
  AOI21_X1 U16520 ( .B1(n15099), .B2(n14674), .A(n14673), .ZN(n14678) );
  AOI22_X1 U16521 ( .A1(n15129), .A2(n14678), .B1(n14675), .B2(n15127), .ZN(
        P2_U3511) );
  AOI22_X1 U16522 ( .A1(n15119), .A2(n14676), .B1(n9312), .B2(n15117), .ZN(
        P2_U3469) );
  INV_X1 U16523 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14677) );
  AOI22_X1 U16524 ( .A1(n15119), .A2(n14678), .B1(n14677), .B2(n15117), .ZN(
        P2_U3466) );
  AOI21_X1 U16525 ( .B1(n14681), .B2(n14680), .A(n14679), .ZN(n14683) );
  OAI211_X1 U16526 ( .C1(n14685), .C2(n14684), .A(n14683), .B(n14682), .ZN(
        n14686) );
  AOI21_X1 U16527 ( .B1(n14688), .B2(n14687), .A(n14686), .ZN(n14699) );
  AOI22_X1 U16528 ( .A1(n14863), .A2(n14699), .B1(n14056), .B2(n14861), .ZN(
        P1_U3542) );
  OAI211_X1 U16529 ( .C1(n7122), .C2(n14852), .A(n14690), .B(n14689), .ZN(
        n14691) );
  AOI21_X1 U16530 ( .B1(n14692), .B2(n14855), .A(n14691), .ZN(n14701) );
  AOI22_X1 U16531 ( .A1(n14863), .A2(n14701), .B1(n14059), .B2(n14861), .ZN(
        P1_U3541) );
  OAI21_X1 U16532 ( .B1(n14694), .B2(n14852), .A(n14693), .ZN(n14696) );
  AOI211_X1 U16533 ( .C1(n14855), .C2(n14697), .A(n14696), .B(n14695), .ZN(
        n14703) );
  AOI22_X1 U16534 ( .A1(n14863), .A2(n14703), .B1(n11175), .B2(n14861), .ZN(
        P1_U3539) );
  INV_X1 U16535 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U16536 ( .A1(n14857), .A2(n14699), .B1(n14698), .B2(n9673), .ZN(
        P1_U3501) );
  INV_X1 U16537 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14700) );
  AOI22_X1 U16538 ( .A1(n14857), .A2(n14701), .B1(n14700), .B2(n9673), .ZN(
        P1_U3498) );
  INV_X1 U16539 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14702) );
  AOI22_X1 U16540 ( .A1(n14857), .A2(n14703), .B1(n14702), .B2(n9673), .ZN(
        P1_U3492) );
  AOI21_X1 U16541 ( .B1(n14706), .B2(n14705), .A(n14704), .ZN(n14708) );
  XNOR2_X1 U16542 ( .A(n14708), .B(n14707), .ZN(SUB_1596_U69) );
  XNOR2_X1 U16543 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14709), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16544 ( .B1(n14712), .B2(n14711), .A(n14710), .ZN(n14713) );
  XNOR2_X1 U16545 ( .A(n14713), .B(n14985), .ZN(SUB_1596_U67) );
  AOI21_X1 U16546 ( .B1(n14716), .B2(n14715), .A(n14714), .ZN(n14717) );
  XNOR2_X1 U16547 ( .A(n14717), .B(n14998), .ZN(SUB_1596_U66) );
  AOI21_X1 U16548 ( .B1(n14720), .B2(n14719), .A(n14718), .ZN(n14721) );
  XNOR2_X1 U16549 ( .A(n14721), .B(n15010), .ZN(SUB_1596_U65) );
  AOI21_X1 U16550 ( .B1(n14724), .B2(n14723), .A(n14722), .ZN(n14725) );
  XNOR2_X1 U16551 ( .A(n14725), .B(n15027), .ZN(SUB_1596_U64) );
  OAI21_X1 U16552 ( .B1(n14727), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14726), .ZN(
        n14728) );
  XNOR2_X1 U16553 ( .A(n14728), .B(n7684), .ZN(n14732) );
  AOI22_X1 U16554 ( .A1(n14729), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14730) );
  OAI21_X1 U16555 ( .B1(n14732), .B2(n14731), .A(n14730), .ZN(P1_U3243) );
  INV_X1 U16556 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14745) );
  OAI21_X1 U16557 ( .B1(n14735), .B2(n14734), .A(n14733), .ZN(n14742) );
  NOR2_X1 U16558 ( .A1(n14828), .A2(n14736), .ZN(n14741) );
  AOI211_X1 U16559 ( .C1(n14739), .C2(n14738), .A(n14789), .B(n14737), .ZN(
        n14740) );
  AOI211_X1 U16560 ( .C1(n14819), .C2(n14742), .A(n14741), .B(n14740), .ZN(
        n14744) );
  OAI211_X1 U16561 ( .C1(n14745), .C2(n14832), .A(n14744), .B(n14743), .ZN(
        P1_U3254) );
  AOI211_X1 U16562 ( .C1(n14748), .C2(n14747), .A(n14785), .B(n14746), .ZN(
        n14753) );
  AOI211_X1 U16563 ( .C1(n14751), .C2(n14750), .A(n14789), .B(n14749), .ZN(
        n14752) );
  AOI211_X1 U16564 ( .C1(n14796), .C2(n14754), .A(n14753), .B(n14752), .ZN(
        n14756) );
  OAI211_X1 U16565 ( .C1(n14757), .C2(n14832), .A(n14756), .B(n14755), .ZN(
        P1_U3256) );
  OAI21_X1 U16566 ( .B1(n14760), .B2(n14759), .A(n14758), .ZN(n14767) );
  NOR2_X1 U16567 ( .A1(n14828), .A2(n14761), .ZN(n14766) );
  AOI211_X1 U16568 ( .C1(n14764), .C2(n14763), .A(n14762), .B(n14789), .ZN(
        n14765) );
  AOI211_X1 U16569 ( .C1(n14819), .C2(n14767), .A(n14766), .B(n14765), .ZN(
        n14769) );
  OAI211_X1 U16570 ( .C1(n14770), .C2(n14832), .A(n14769), .B(n14768), .ZN(
        P1_U3257) );
  OAI21_X1 U16571 ( .B1(n14773), .B2(n14772), .A(n14771), .ZN(n14774) );
  NAND2_X1 U16572 ( .A1(n14819), .A2(n14774), .ZN(n14779) );
  OAI21_X1 U16573 ( .B1(n14776), .B2(n11510), .A(n14775), .ZN(n14777) );
  NAND2_X1 U16574 ( .A1(n14824), .A2(n14777), .ZN(n14778) );
  OAI211_X1 U16575 ( .C1(n14828), .C2(n14780), .A(n14779), .B(n14778), .ZN(
        n14781) );
  INV_X1 U16576 ( .A(n14781), .ZN(n14783) );
  OAI211_X1 U16577 ( .C1(n14784), .C2(n14832), .A(n14783), .B(n14782), .ZN(
        P1_U3258) );
  INV_X1 U16578 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14799) );
  AOI211_X1 U16579 ( .C1(n14788), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n14794) );
  AOI211_X1 U16580 ( .C1(n14792), .C2(n14791), .A(n14790), .B(n14789), .ZN(
        n14793) );
  AOI211_X1 U16581 ( .C1(n14796), .C2(n14795), .A(n14794), .B(n14793), .ZN(
        n14798) );
  OAI211_X1 U16582 ( .C1(n14799), .C2(n14832), .A(n14798), .B(n14797), .ZN(
        P1_U3259) );
  AOI21_X1 U16583 ( .B1(n14802), .B2(n14801), .A(n14800), .ZN(n14803) );
  NAND2_X1 U16584 ( .A1(n14819), .A2(n14803), .ZN(n14809) );
  AOI21_X1 U16585 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n14807) );
  NAND2_X1 U16586 ( .A1(n14824), .A2(n14807), .ZN(n14808) );
  OAI211_X1 U16587 ( .C1(n14828), .C2(n14810), .A(n14809), .B(n14808), .ZN(
        n14811) );
  INV_X1 U16588 ( .A(n14811), .ZN(n14813) );
  OAI211_X1 U16589 ( .C1(n14814), .C2(n14832), .A(n14813), .B(n14812), .ZN(
        P1_U3260) );
  INV_X1 U16590 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15399) );
  AOI21_X1 U16591 ( .B1(n14817), .B2(n14816), .A(n14815), .ZN(n14818) );
  NAND2_X1 U16592 ( .A1(n14819), .A2(n14818), .ZN(n14826) );
  AOI21_X1 U16593 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(n14823) );
  NAND2_X1 U16594 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  OAI211_X1 U16595 ( .C1(n14828), .C2(n14827), .A(n14826), .B(n14825), .ZN(
        n14829) );
  INV_X1 U16596 ( .A(n14829), .ZN(n14831) );
  OAI211_X1 U16597 ( .C1(n15399), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        P1_U3261) );
  AND2_X1 U16598 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14833), .ZN(P1_U3294) );
  AND2_X1 U16599 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14833), .ZN(P1_U3295) );
  AND2_X1 U16600 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14833), .ZN(P1_U3296) );
  AND2_X1 U16601 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14833), .ZN(P1_U3297) );
  AND2_X1 U16602 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14833), .ZN(P1_U3298) );
  AND2_X1 U16603 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14833), .ZN(P1_U3299) );
  AND2_X1 U16604 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14833), .ZN(P1_U3300) );
  AND2_X1 U16605 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14833), .ZN(P1_U3301) );
  AND2_X1 U16606 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14833), .ZN(P1_U3302) );
  AND2_X1 U16607 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14833), .ZN(P1_U3303) );
  AND2_X1 U16608 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14833), .ZN(P1_U3304) );
  AND2_X1 U16609 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14833), .ZN(P1_U3305) );
  AND2_X1 U16610 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14833), .ZN(P1_U3306) );
  AND2_X1 U16611 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14833), .ZN(P1_U3307) );
  AND2_X1 U16612 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14833), .ZN(P1_U3308) );
  AND2_X1 U16613 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14833), .ZN(P1_U3309) );
  AND2_X1 U16614 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14833), .ZN(P1_U3310) );
  AND2_X1 U16615 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14833), .ZN(P1_U3311) );
  AND2_X1 U16616 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14833), .ZN(P1_U3312) );
  AND2_X1 U16617 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14833), .ZN(P1_U3313) );
  AND2_X1 U16618 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14833), .ZN(P1_U3314) );
  AND2_X1 U16619 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14833), .ZN(P1_U3315) );
  AND2_X1 U16620 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14833), .ZN(P1_U3316) );
  AND2_X1 U16621 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14833), .ZN(P1_U3317) );
  AND2_X1 U16622 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14833), .ZN(P1_U3318) );
  AND2_X1 U16623 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14833), .ZN(P1_U3319) );
  AND2_X1 U16624 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14833), .ZN(P1_U3320) );
  AND2_X1 U16625 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14833), .ZN(P1_U3321) );
  AND2_X1 U16626 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14833), .ZN(P1_U3322) );
  AND2_X1 U16627 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14833), .ZN(P1_U3323) );
  INV_X1 U16628 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14834) );
  AOI22_X1 U16629 ( .A1(n14857), .A2(n14835), .B1(n14834), .B2(n9673), .ZN(
        P1_U3459) );
  OAI21_X1 U16630 ( .B1(n14837), .B2(n14852), .A(n14836), .ZN(n14839) );
  AOI211_X1 U16631 ( .C1(n14842), .C2(n14840), .A(n14839), .B(n14838), .ZN(
        n14859) );
  INV_X1 U16632 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14841) );
  AOI22_X1 U16633 ( .A1(n14857), .A2(n14859), .B1(n14841), .B2(n9673), .ZN(
        P1_U3474) );
  NAND2_X1 U16634 ( .A1(n14843), .A2(n14842), .ZN(n14845) );
  OAI211_X1 U16635 ( .C1(n14846), .C2(n14852), .A(n14845), .B(n14844), .ZN(
        n14847) );
  NOR2_X1 U16636 ( .A1(n14848), .A2(n14847), .ZN(n14860) );
  INV_X1 U16637 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14849) );
  AOI22_X1 U16638 ( .A1(n14857), .A2(n14860), .B1(n14849), .B2(n9673), .ZN(
        P1_U3480) );
  OAI211_X1 U16639 ( .C1(n7126), .C2(n14852), .A(n14851), .B(n14850), .ZN(
        n14853) );
  AOI21_X1 U16640 ( .B1(n14855), .B2(n14854), .A(n14853), .ZN(n14862) );
  INV_X1 U16641 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14856) );
  AOI22_X1 U16642 ( .A1(n14857), .A2(n14862), .B1(n14856), .B2(n9673), .ZN(
        P1_U3489) );
  INV_X1 U16643 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14858) );
  AOI22_X1 U16644 ( .A1(n14863), .A2(n14859), .B1(n14858), .B2(n14861), .ZN(
        P1_U3533) );
  AOI22_X1 U16645 ( .A1(n14863), .A2(n14860), .B1(n7982), .B2(n14861), .ZN(
        P1_U3535) );
  AOI22_X1 U16646 ( .A1(n14863), .A2(n14862), .B1(n10730), .B2(n14861), .ZN(
        P1_U3538) );
  NOR2_X1 U16647 ( .A1(n14864), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16648 ( .A1(n14864), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14877) );
  OAI211_X1 U16649 ( .C1(n14867), .C2(n14866), .A(n15028), .B(n14865), .ZN(
        n14873) );
  OAI21_X1 U16650 ( .B1(n14870), .B2(n14869), .A(n14868), .ZN(n14871) );
  OR2_X1 U16651 ( .A1(n15013), .A2(n14871), .ZN(n14872) );
  OAI211_X1 U16652 ( .C1(n15035), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14875) );
  INV_X1 U16653 ( .A(n14875), .ZN(n14876) );
  NAND2_X1 U16654 ( .A1(n14877), .A2(n14876), .ZN(P2_U3216) );
  OAI211_X1 U16655 ( .C1(n14880), .C2(n14879), .A(n15028), .B(n14878), .ZN(
        n14886) );
  OAI21_X1 U16656 ( .B1(n14883), .B2(n14882), .A(n14881), .ZN(n14884) );
  OR2_X1 U16657 ( .A1(n15013), .A2(n14884), .ZN(n14885) );
  OAI211_X1 U16658 ( .C1(n15035), .C2(n14887), .A(n14886), .B(n14885), .ZN(
        n14888) );
  INV_X1 U16659 ( .A(n14888), .ZN(n14890) );
  NAND2_X1 U16660 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n14889) );
  OAI211_X1 U16661 ( .C1(n15044), .C2(n15796), .A(n14890), .B(n14889), .ZN(
        P2_U3217) );
  OAI211_X1 U16662 ( .C1(n14893), .C2(n14892), .A(n15028), .B(n14891), .ZN(
        n14899) );
  OAI21_X1 U16663 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14897) );
  OR2_X1 U16664 ( .A1(n15013), .A2(n14897), .ZN(n14898) );
  OAI211_X1 U16665 ( .C1(n15035), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        n14901) );
  INV_X1 U16666 ( .A(n14901), .ZN(n14903) );
  OAI211_X1 U16667 ( .C1(n15044), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        P2_U3218) );
  INV_X1 U16668 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n14917) );
  OAI211_X1 U16669 ( .C1(n14907), .C2(n14906), .A(n15032), .B(n14905), .ZN(
        n14912) );
  OAI211_X1 U16670 ( .C1(n14910), .C2(n14909), .A(n15028), .B(n14908), .ZN(
        n14911) );
  OAI211_X1 U16671 ( .C1(n15035), .C2(n14913), .A(n14912), .B(n14911), .ZN(
        n14914) );
  INV_X1 U16672 ( .A(n14914), .ZN(n14916) );
  OAI211_X1 U16673 ( .C1(n15044), .C2(n14917), .A(n14916), .B(n14915), .ZN(
        P2_U3219) );
  OAI211_X1 U16674 ( .C1(n14920), .C2(n14919), .A(n15032), .B(n14918), .ZN(
        n14925) );
  OAI211_X1 U16675 ( .C1(n14923), .C2(n14922), .A(n15028), .B(n14921), .ZN(
        n14924) );
  OAI211_X1 U16676 ( .C1(n15035), .C2(n14926), .A(n14925), .B(n14924), .ZN(
        n14927) );
  INV_X1 U16677 ( .A(n14927), .ZN(n14929) );
  OAI211_X1 U16678 ( .C1(n15044), .C2(n7239), .A(n14929), .B(n14928), .ZN(
        P2_U3220) );
  INV_X1 U16679 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14942) );
  OAI211_X1 U16680 ( .C1(n14932), .C2(n14931), .A(n14930), .B(n15032), .ZN(
        n14937) );
  OAI211_X1 U16681 ( .C1(n14935), .C2(n14934), .A(n14933), .B(n15028), .ZN(
        n14936) );
  OAI211_X1 U16682 ( .C1(n15035), .C2(n14938), .A(n14937), .B(n14936), .ZN(
        n14939) );
  INV_X1 U16683 ( .A(n14939), .ZN(n14941) );
  NAND2_X1 U16684 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n14940) );
  OAI211_X1 U16685 ( .C1(n14942), .C2(n15044), .A(n14941), .B(n14940), .ZN(
        P2_U3221) );
  OAI211_X1 U16686 ( .C1(n14945), .C2(n14944), .A(n14943), .B(n15028), .ZN(
        n14950) );
  OAI211_X1 U16687 ( .C1(n14948), .C2(n14947), .A(n14946), .B(n15032), .ZN(
        n14949) );
  OAI211_X1 U16688 ( .C1(n15035), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14952) );
  INV_X1 U16689 ( .A(n14952), .ZN(n14954) );
  OAI211_X1 U16690 ( .C1(n14955), .C2(n15044), .A(n14954), .B(n14953), .ZN(
        P2_U3222) );
  NAND2_X1 U16691 ( .A1(n14957), .A2(n14956), .ZN(n14958) );
  NAND3_X1 U16692 ( .A1(n14959), .A2(n15028), .A3(n14958), .ZN(n14965) );
  NAND2_X1 U16693 ( .A1(n14961), .A2(n14960), .ZN(n14962) );
  NAND3_X1 U16694 ( .A1(n14963), .A2(n15032), .A3(n14962), .ZN(n14964) );
  OAI211_X1 U16695 ( .C1(n15035), .C2(n14966), .A(n14965), .B(n14964), .ZN(
        n14967) );
  INV_X1 U16696 ( .A(n14967), .ZN(n14969) );
  OAI211_X1 U16697 ( .C1(n14970), .C2(n15044), .A(n14969), .B(n14968), .ZN(
        P2_U3224) );
  NAND2_X1 U16698 ( .A1(n14972), .A2(n14971), .ZN(n14973) );
  NAND3_X1 U16699 ( .A1(n14974), .A2(n15032), .A3(n14973), .ZN(n14980) );
  NAND2_X1 U16700 ( .A1(n14976), .A2(n14975), .ZN(n14977) );
  NAND3_X1 U16701 ( .A1(n14978), .A2(n15028), .A3(n14977), .ZN(n14979) );
  OAI211_X1 U16702 ( .C1(n15035), .C2(n14981), .A(n14980), .B(n14979), .ZN(
        n14982) );
  INV_X1 U16703 ( .A(n14982), .ZN(n14984) );
  NAND2_X1 U16704 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14983)
         );
  OAI211_X1 U16705 ( .C1(n14985), .C2(n15044), .A(n14984), .B(n14983), .ZN(
        P2_U3227) );
  OAI21_X1 U16706 ( .B1(n14986), .B2(P2_REG2_REG_14__SCAN_IN), .A(n15028), 
        .ZN(n14987) );
  OR2_X1 U16707 ( .A1(n14988), .A2(n14987), .ZN(n14993) );
  OAI211_X1 U16708 ( .C1(n14991), .C2(n14990), .A(n14989), .B(n15032), .ZN(
        n14992) );
  OAI211_X1 U16709 ( .C1(n15035), .C2(n14994), .A(n14993), .B(n14992), .ZN(
        n14995) );
  INV_X1 U16710 ( .A(n14995), .ZN(n14997) );
  NAND2_X1 U16711 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14996)
         );
  OAI211_X1 U16712 ( .C1(n14998), .C2(n15044), .A(n14997), .B(n14996), .ZN(
        P2_U3228) );
  INV_X1 U16713 ( .A(n15035), .ZN(n15024) );
  AOI211_X1 U16714 ( .C1(n15001), .C2(n15000), .A(n14999), .B(n15018), .ZN(
        n15006) );
  AOI211_X1 U16715 ( .C1(n15004), .C2(n15003), .A(n15002), .B(n15013), .ZN(
        n15005) );
  AOI211_X1 U16716 ( .C1(n15024), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        n15009) );
  NAND2_X1 U16717 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15008)
         );
  OAI211_X1 U16718 ( .C1(n15010), .C2(n15044), .A(n15009), .B(n15008), .ZN(
        P2_U3229) );
  INV_X1 U16719 ( .A(n15011), .ZN(n15012) );
  AOI211_X1 U16720 ( .C1(n15015), .C2(n15014), .A(n15013), .B(n15012), .ZN(
        n15022) );
  INV_X1 U16721 ( .A(n15016), .ZN(n15017) );
  AOI211_X1 U16722 ( .C1(n15020), .C2(n15019), .A(n15018), .B(n15017), .ZN(
        n15021) );
  AOI211_X1 U16723 ( .C1(n15024), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15026) );
  NAND2_X1 U16724 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n15025)
         );
  OAI211_X1 U16725 ( .C1(n15027), .C2(n15044), .A(n15026), .B(n15025), .ZN(
        P2_U3230) );
  OAI211_X1 U16726 ( .C1(n15031), .C2(n15030), .A(n15029), .B(n15028), .ZN(
        n15041) );
  OAI21_X1 U16727 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15038) );
  OAI22_X1 U16728 ( .A1(n15038), .A2(n15037), .B1(n15036), .B2(n15035), .ZN(
        n15039) );
  INV_X1 U16729 ( .A(n15039), .ZN(n15040) );
  AND2_X1 U16730 ( .A1(n15041), .A2(n15040), .ZN(n15043) );
  NAND2_X1 U16731 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15042)
         );
  OAI211_X1 U16732 ( .C1(n15045), .C2(n15044), .A(n15043), .B(n15042), .ZN(
        P2_U3231) );
  XNOR2_X1 U16733 ( .A(n15046), .B(n15056), .ZN(n15049) );
  AOI21_X1 U16734 ( .B1(n15049), .B2(n15048), .A(n15047), .ZN(n15090) );
  NAND2_X1 U16735 ( .A1(n15067), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n15050) );
  OAI21_X1 U16736 ( .B1(n15052), .B2(n15051), .A(n15050), .ZN(n15053) );
  AOI21_X1 U16737 ( .B1(n15055), .B2(n15054), .A(n15053), .ZN(n15066) );
  NAND2_X1 U16738 ( .A1(n15057), .A2(n15056), .ZN(n15058) );
  NAND2_X1 U16739 ( .A1(n15059), .A2(n15058), .ZN(n15087) );
  OAI211_X1 U16740 ( .C1(n15061), .C2(n15089), .A(n10749), .B(n15060), .ZN(
        n15088) );
  OAI22_X1 U16741 ( .A1(n15063), .A2(n15087), .B1(n15088), .B2(n15062), .ZN(
        n15064) );
  INV_X1 U16742 ( .A(n15064), .ZN(n15065) );
  OAI211_X1 U16743 ( .C1(n15067), .C2(n15090), .A(n15066), .B(n15065), .ZN(
        P2_U3259) );
  NAND2_X1 U16744 ( .A1(n15072), .A2(n15068), .ZN(n15069) );
  AND2_X1 U16745 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15069), .ZN(P2_U3266) );
  AND2_X1 U16746 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15069), .ZN(P2_U3267) );
  AND2_X1 U16747 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15069), .ZN(P2_U3268) );
  AND2_X1 U16748 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15069), .ZN(P2_U3269) );
  AND2_X1 U16749 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15069), .ZN(P2_U3270) );
  AND2_X1 U16750 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15069), .ZN(P2_U3271) );
  AND2_X1 U16751 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15069), .ZN(P2_U3272) );
  AND2_X1 U16752 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15069), .ZN(P2_U3273) );
  AND2_X1 U16753 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15069), .ZN(P2_U3274) );
  AND2_X1 U16754 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15069), .ZN(P2_U3275) );
  AND2_X1 U16755 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15069), .ZN(P2_U3276) );
  AND2_X1 U16756 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15069), .ZN(P2_U3277) );
  AND2_X1 U16757 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15069), .ZN(P2_U3278) );
  AND2_X1 U16758 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15069), .ZN(P2_U3279) );
  AND2_X1 U16759 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15069), .ZN(P2_U3280) );
  AND2_X1 U16760 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15069), .ZN(P2_U3281) );
  AND2_X1 U16761 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15069), .ZN(P2_U3282) );
  AND2_X1 U16762 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15069), .ZN(P2_U3283) );
  AND2_X1 U16763 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15069), .ZN(P2_U3284) );
  AND2_X1 U16764 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15069), .ZN(P2_U3285) );
  AND2_X1 U16765 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15069), .ZN(P2_U3286) );
  AND2_X1 U16766 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15069), .ZN(P2_U3287) );
  AND2_X1 U16767 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15069), .ZN(P2_U3288) );
  AND2_X1 U16768 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15069), .ZN(P2_U3289) );
  AND2_X1 U16769 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15069), .ZN(P2_U3290) );
  AND2_X1 U16770 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15069), .ZN(P2_U3291) );
  AND2_X1 U16771 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15069), .ZN(P2_U3292) );
  AND2_X1 U16772 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15069), .ZN(P2_U3293) );
  AND2_X1 U16773 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15069), .ZN(P2_U3294) );
  AND2_X1 U16774 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15069), .ZN(P2_U3295) );
  INV_X1 U16775 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U16776 ( .A1(n15072), .A2(n15071), .B1(n15070), .B2(n15074), .ZN(
        P2_U3416) );
  AOI21_X1 U16777 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n15074), .A(n15073), .ZN(
        n15075) );
  INV_X1 U16778 ( .A(n15075), .ZN(P2_U3417) );
  AOI22_X1 U16779 ( .A1(n15119), .A2(n15076), .B1(n9080), .B2(n15117), .ZN(
        P2_U3430) );
  INV_X1 U16780 ( .A(n15082), .ZN(n15085) );
  AOI21_X1 U16781 ( .B1(n15079), .B2(n15078), .A(n15077), .ZN(n15081) );
  OAI211_X1 U16782 ( .C1(n15083), .C2(n15082), .A(n15081), .B(n15080), .ZN(
        n15084) );
  AOI21_X1 U16783 ( .B1(n15106), .B2(n15085), .A(n15084), .ZN(n15121) );
  INV_X1 U16784 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15086) );
  AOI22_X1 U16785 ( .A1(n15119), .A2(n15121), .B1(n15086), .B2(n15117), .ZN(
        P2_U3445) );
  INV_X1 U16786 ( .A(n15087), .ZN(n15093) );
  OAI21_X1 U16787 ( .B1(n15089), .B2(n15111), .A(n15088), .ZN(n15092) );
  INV_X1 U16788 ( .A(n15090), .ZN(n15091) );
  AOI211_X1 U16789 ( .C1(n15093), .C2(n15099), .A(n15092), .B(n15091), .ZN(
        n15123) );
  AOI22_X1 U16790 ( .A1(n15119), .A2(n15123), .B1(n9185), .B2(n15117), .ZN(
        P2_U3448) );
  INV_X1 U16791 ( .A(n15094), .ZN(n15100) );
  OAI21_X1 U16792 ( .B1(n15096), .B2(n15111), .A(n15095), .ZN(n15098) );
  AOI211_X1 U16793 ( .C1(n15100), .C2(n15099), .A(n15098), .B(n15097), .ZN(
        n15125) );
  INV_X1 U16794 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U16795 ( .A1(n15119), .A2(n15125), .B1(n15101), .B2(n15117), .ZN(
        P2_U3451) );
  OAI21_X1 U16796 ( .B1(n15103), .B2(n15111), .A(n15102), .ZN(n15104) );
  AOI21_X1 U16797 ( .B1(n15107), .B2(n9095), .A(n15104), .ZN(n15109) );
  AOI21_X1 U16798 ( .B1(n15107), .B2(n15106), .A(n15105), .ZN(n15108) );
  AND2_X1 U16799 ( .A1(n15109), .A2(n15108), .ZN(n15126) );
  AOI22_X1 U16800 ( .A1(n15119), .A2(n15126), .B1(n9224), .B2(n15117), .ZN(
        P2_U3454) );
  OAI21_X1 U16801 ( .B1(n15112), .B2(n15111), .A(n15110), .ZN(n15113) );
  AOI21_X1 U16802 ( .B1(n15114), .B2(n9095), .A(n15113), .ZN(n15115) );
  AND2_X1 U16803 ( .A1(n15116), .A2(n15115), .ZN(n15128) );
  INV_X1 U16804 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15118) );
  AOI22_X1 U16805 ( .A1(n15119), .A2(n15128), .B1(n15118), .B2(n15117), .ZN(
        P2_U3460) );
  AOI22_X1 U16806 ( .A1(n15129), .A2(n15121), .B1(n15120), .B2(n15127), .ZN(
        P2_U3504) );
  AOI22_X1 U16807 ( .A1(n15129), .A2(n15123), .B1(n15122), .B2(n15127), .ZN(
        P2_U3505) );
  AOI22_X1 U16808 ( .A1(n15129), .A2(n15125), .B1(n15124), .B2(n15127), .ZN(
        P2_U3506) );
  AOI22_X1 U16809 ( .A1(n15129), .A2(n15126), .B1(n9220), .B2(n15127), .ZN(
        P2_U3507) );
  AOI22_X1 U16810 ( .A1(n15129), .A2(n15128), .B1(n10001), .B2(n15127), .ZN(
        P2_U3509) );
  NOR2_X1 U16811 ( .A1(P3_U3897), .A2(n15232), .ZN(P3_U3150) );
  OR2_X1 U16812 ( .A1(n15130), .A2(n15313), .ZN(n15133) );
  OR2_X1 U16813 ( .A1(n15131), .A2(n15315), .ZN(n15132) );
  AND2_X1 U16814 ( .A1(n15133), .A2(n15132), .ZN(n15274) );
  OAI211_X1 U16815 ( .C1(n15137), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        n15142) );
  AOI21_X1 U16816 ( .B1(n15140), .B2(n15139), .A(n15138), .ZN(n15141) );
  OAI211_X1 U16817 ( .C1(n15274), .C2(n15143), .A(n15142), .B(n15141), .ZN(
        n15144) );
  INV_X1 U16818 ( .A(n15144), .ZN(n15145) );
  OAI21_X1 U16819 ( .B1(n15277), .B2(n15159), .A(n15145), .ZN(P3_U3153) );
  AOI21_X1 U16820 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(n15157) );
  NAND2_X1 U16821 ( .A1(n15150), .A2(n15149), .ZN(n15152) );
  OAI211_X1 U16822 ( .C1(n15154), .C2(n15153), .A(n15152), .B(n15151), .ZN(
        n15155) );
  AOI21_X1 U16823 ( .B1(n15157), .B2(n15156), .A(n15155), .ZN(n15158) );
  OAI21_X1 U16824 ( .B1(n15160), .B2(n15159), .A(n15158), .ZN(P3_U3157) );
  NAND3_X1 U16825 ( .A1(n15241), .A2(n15266), .A3(n15253), .ZN(n15164) );
  NAND2_X1 U16826 ( .A1(n15164), .A2(n15163), .ZN(n15167) );
  OAI211_X1 U16827 ( .C1(n15514), .C2(n15251), .A(n15167), .B(n15166), .ZN(
        P3_U3182) );
  AOI21_X1 U16828 ( .B1(n11500), .B2(n15169), .A(n15168), .ZN(n15170) );
  OR2_X1 U16829 ( .A1(n15170), .A2(n15266), .ZN(n15184) );
  AOI21_X1 U16830 ( .B1(n11058), .B2(n15172), .A(n15171), .ZN(n15173) );
  OR2_X1 U16831 ( .A1(n15173), .A2(n15241), .ZN(n15183) );
  INV_X1 U16832 ( .A(n15174), .ZN(n15176) );
  NOR2_X1 U16833 ( .A1(n15176), .A2(n15175), .ZN(n15177) );
  XNOR2_X1 U16834 ( .A(n15178), .B(n15177), .ZN(n15179) );
  NAND2_X1 U16835 ( .A1(n15179), .A2(n15237), .ZN(n15182) );
  NAND2_X1 U16836 ( .A1(n15259), .A2(n15180), .ZN(n15181) );
  AND4_X1 U16837 ( .A1(n15184), .A2(n15183), .A3(n15182), .A4(n15181), .ZN(
        n15186) );
  NAND2_X1 U16838 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15185) );
  OAI211_X1 U16839 ( .C1(n15187), .C2(n15251), .A(n15186), .B(n15185), .ZN(
        P3_U3191) );
  AOI21_X1 U16840 ( .B1(n14650), .B2(n15189), .A(n15188), .ZN(n15202) );
  XNOR2_X1 U16841 ( .A(n15191), .B(n15190), .ZN(n15196) );
  INV_X1 U16842 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15747) );
  NOR2_X1 U16843 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15747), .ZN(n15192) );
  AOI21_X1 U16844 ( .B1(n15232), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n15192), 
        .ZN(n15193) );
  OAI21_X1 U16845 ( .B1(n15235), .B2(n15194), .A(n15193), .ZN(n15195) );
  AOI21_X1 U16846 ( .B1(n15196), .B2(n15237), .A(n15195), .ZN(n15201) );
  AOI21_X1 U16847 ( .B1(n15198), .B2(n8654), .A(n15197), .ZN(n15199) );
  OR2_X1 U16848 ( .A1(n15199), .A2(n15241), .ZN(n15200) );
  OAI211_X1 U16849 ( .C1(n15202), .C2(n15266), .A(n15201), .B(n15200), .ZN(
        P3_U3193) );
  INV_X1 U16850 ( .A(n15203), .ZN(n15204) );
  AOI21_X1 U16851 ( .B1(n15206), .B2(n15205), .A(n15204), .ZN(n15222) );
  OAI21_X1 U16852 ( .B1(n15251), .B2(n15208), .A(n15207), .ZN(n15213) );
  OAI211_X1 U16853 ( .C1(n15210), .C2(n15209), .A(n15225), .B(n15237), .ZN(
        n15211) );
  INV_X1 U16854 ( .A(n15211), .ZN(n15212) );
  AOI211_X1 U16855 ( .C1(n15259), .C2(n15214), .A(n15213), .B(n15212), .ZN(
        n15221) );
  INV_X1 U16856 ( .A(n15215), .ZN(n15216) );
  AOI21_X1 U16857 ( .B1(n15218), .B2(n15217), .A(n15216), .ZN(n15219) );
  OR2_X1 U16858 ( .A1(n15219), .A2(n15241), .ZN(n15220) );
  OAI211_X1 U16859 ( .C1(n15222), .C2(n15266), .A(n15221), .B(n15220), .ZN(
        P3_U3194) );
  AOI21_X1 U16860 ( .B1(n8694), .B2(n15224), .A(n15223), .ZN(n15245) );
  INV_X1 U16861 ( .A(n15225), .ZN(n15227) );
  NOR2_X1 U16862 ( .A1(n15227), .A2(n15226), .ZN(n15230) );
  OAI21_X1 U16863 ( .B1(n15230), .B2(n15229), .A(n15228), .ZN(n15238) );
  NOR2_X1 U16864 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8386), .ZN(n15231) );
  AOI21_X1 U16865 ( .B1(n15232), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15231), 
        .ZN(n15233) );
  OAI21_X1 U16866 ( .B1(n15235), .B2(n15234), .A(n15233), .ZN(n15236) );
  AOI21_X1 U16867 ( .B1(n15238), .B2(n15237), .A(n15236), .ZN(n15244) );
  AOI21_X1 U16868 ( .B1(n15240), .B2(n8695), .A(n15239), .ZN(n15242) );
  OR2_X1 U16869 ( .A1(n15242), .A2(n15241), .ZN(n15243) );
  OAI211_X1 U16870 ( .C1(n15245), .C2(n15266), .A(n15244), .B(n15243), .ZN(
        P3_U3195) );
  AOI21_X1 U16871 ( .B1(n15247), .B2(n15246), .A(n6822), .ZN(n15267) );
  INV_X1 U16872 ( .A(n15248), .ZN(n15258) );
  INV_X1 U16873 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15250) );
  OAI21_X1 U16874 ( .B1(n15251), .B2(n15250), .A(n15249), .ZN(n15257) );
  AOI211_X1 U16875 ( .C1(n15255), .C2(n15254), .A(n15253), .B(n15252), .ZN(
        n15256) );
  AOI211_X1 U16876 ( .C1(n15259), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        n15265) );
  XNOR2_X1 U16877 ( .A(n15261), .B(n15260), .ZN(n15263) );
  NAND2_X1 U16878 ( .A1(n15263), .A2(n15262), .ZN(n15264) );
  OAI211_X1 U16879 ( .C1(n15267), .C2(n15266), .A(n15265), .B(n15264), .ZN(
        P3_U3196) );
  XNOR2_X1 U16880 ( .A(n15269), .B(n15268), .ZN(n15369) );
  OR2_X1 U16881 ( .A1(n15284), .A2(n15283), .ZN(n15286) );
  NAND2_X1 U16882 ( .A1(n15286), .A2(n15270), .ZN(n15273) );
  NAND2_X1 U16883 ( .A1(n15273), .A2(n15272), .ZN(n15271) );
  OAI211_X1 U16884 ( .C1(n15273), .C2(n15272), .A(n15271), .B(n15322), .ZN(
        n15275) );
  NAND2_X1 U16885 ( .A1(n15275), .A2(n15274), .ZN(n15366) );
  AOI21_X1 U16886 ( .B1(n15369), .B2(n15317), .A(n15366), .ZN(n15280) );
  NOR2_X1 U16887 ( .A1(n15276), .A2(n15339), .ZN(n15367) );
  INV_X1 U16888 ( .A(n15277), .ZN(n15278) );
  AOI22_X1 U16889 ( .A1(n15295), .A2(n15367), .B1(n15332), .B2(n15278), .ZN(
        n15279) );
  OAI221_X1 U16890 ( .B1(n15337), .B2(n15280), .C1(n15335), .C2(n9744), .A(
        n15279), .ZN(P3_U3226) );
  INV_X1 U16891 ( .A(n15281), .ZN(n15291) );
  XOR2_X1 U16892 ( .A(n15282), .B(n15283), .Z(n15290) );
  INV_X1 U16893 ( .A(n15290), .ZN(n15364) );
  AOI21_X1 U16894 ( .B1(n15284), .B2(n15283), .A(n15311), .ZN(n15287) );
  AOI21_X1 U16895 ( .B1(n15287), .B2(n15286), .A(n15285), .ZN(n15288) );
  OAI21_X1 U16896 ( .B1(n15290), .B2(n15289), .A(n15288), .ZN(n15362) );
  AOI21_X1 U16897 ( .B1(n15291), .B2(n15364), .A(n15362), .ZN(n15298) );
  AND2_X1 U16898 ( .A1(n15292), .A2(n15328), .ZN(n15363) );
  INV_X1 U16899 ( .A(n15293), .ZN(n15294) );
  AOI22_X1 U16900 ( .A1(n15295), .A2(n15363), .B1(n15332), .B2(n15294), .ZN(
        n15296) );
  OAI221_X1 U16901 ( .B1(n15337), .B2(n15298), .C1(n15335), .C2(n15297), .A(
        n15296), .ZN(P3_U3227) );
  INV_X1 U16902 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15319) );
  INV_X1 U16903 ( .A(n15299), .ZN(n15300) );
  NAND2_X1 U16904 ( .A1(n15300), .A2(n15301), .ZN(n15302) );
  MUX2_X1 U16905 ( .A(n15302), .B(n15301), .S(n15308), .Z(n15304) );
  NAND2_X1 U16906 ( .A1(n15304), .A2(n15303), .ZN(n15346) );
  NOR2_X1 U16907 ( .A1(n6682), .A2(n15339), .ZN(n15345) );
  NAND2_X1 U16908 ( .A1(n15345), .A2(n15327), .ZN(n15306) );
  OAI21_X1 U16909 ( .B1(n8508), .B2(n15307), .A(n15306), .ZN(n15316) );
  XNOR2_X1 U16910 ( .A(n15309), .B(n15308), .ZN(n15310) );
  OAI222_X1 U16911 ( .A1(n15315), .A2(n15314), .B1(n15313), .B2(n15312), .C1(
        n15311), .C2(n15310), .ZN(n15344) );
  AOI211_X1 U16912 ( .C1(n15317), .C2(n15346), .A(n15316), .B(n15344), .ZN(
        n15318) );
  AOI22_X1 U16913 ( .A1(n15337), .A2(n15319), .B1(n15318), .B2(n15335), .ZN(
        P3_U3231) );
  XNOR2_X1 U16914 ( .A(n15324), .B(n15320), .ZN(n15323) );
  AOI21_X1 U16915 ( .B1(n15323), .B2(n15322), .A(n15321), .ZN(n15338) );
  XNOR2_X1 U16916 ( .A(n15325), .B(n15324), .ZN(n15342) );
  NAND2_X1 U16917 ( .A1(n15342), .A2(n15326), .ZN(n15331) );
  NAND3_X1 U16918 ( .A1(n15329), .A2(n15328), .A3(n15327), .ZN(n15330) );
  AND3_X1 U16919 ( .A1(n15338), .A2(n15331), .A3(n15330), .ZN(n15336) );
  AOI22_X1 U16920 ( .A1(n15342), .A2(n15333), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15332), .ZN(n15334) );
  OAI221_X1 U16921 ( .B1(n15337), .B2(n15336), .C1(n15335), .C2(n9711), .A(
        n15334), .ZN(P3_U3232) );
  OAI21_X1 U16922 ( .B1(n15340), .B2(n15339), .A(n15338), .ZN(n15341) );
  AOI21_X1 U16923 ( .B1(n15368), .B2(n15342), .A(n15341), .ZN(n15383) );
  INV_X1 U16924 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15343) );
  AOI22_X1 U16925 ( .A1(n15382), .A2(n15383), .B1(n15343), .B2(n9009), .ZN(
        P3_U3393) );
  AOI211_X1 U16926 ( .C1(n15368), .C2(n15346), .A(n15345), .B(n15344), .ZN(
        n15384) );
  AOI22_X1 U16927 ( .A1(n15382), .A2(n15384), .B1(n8509), .B2(n9009), .ZN(
        P3_U3396) );
  INV_X1 U16928 ( .A(n15347), .ZN(n15348) );
  AOI211_X1 U16929 ( .C1(n15380), .C2(n15350), .A(n15349), .B(n15348), .ZN(
        n15385) );
  INV_X1 U16930 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15351) );
  AOI22_X1 U16931 ( .A1(n15382), .A2(n15385), .B1(n15351), .B2(n9009), .ZN(
        P3_U3399) );
  AOI21_X1 U16932 ( .B1(n15353), .B2(n15380), .A(n15352), .ZN(n15354) );
  AND2_X1 U16933 ( .A1(n15355), .A2(n15354), .ZN(n15387) );
  INV_X1 U16934 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15356) );
  AOI22_X1 U16935 ( .A1(n15382), .A2(n15387), .B1(n15356), .B2(n9009), .ZN(
        P3_U3402) );
  INV_X1 U16936 ( .A(n15357), .ZN(n15359) );
  AOI211_X1 U16937 ( .C1(n15360), .C2(n15380), .A(n15359), .B(n15358), .ZN(
        n15388) );
  INV_X1 U16938 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15361) );
  AOI22_X1 U16939 ( .A1(n15382), .A2(n15388), .B1(n15361), .B2(n9009), .ZN(
        P3_U3405) );
  AOI211_X1 U16940 ( .C1(n15364), .C2(n15380), .A(n15363), .B(n15362), .ZN(
        n15390) );
  INV_X1 U16941 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U16942 ( .A1(n15382), .A2(n15390), .B1(n15365), .B2(n9009), .ZN(
        P3_U3408) );
  AOI211_X1 U16943 ( .C1(n15369), .C2(n15368), .A(n15367), .B(n15366), .ZN(
        n15391) );
  INV_X1 U16944 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15370) );
  AOI22_X1 U16945 ( .A1(n15382), .A2(n15391), .B1(n15370), .B2(n9009), .ZN(
        P3_U3411) );
  INV_X1 U16946 ( .A(n15371), .ZN(n15374) );
  AOI211_X1 U16947 ( .C1(n15374), .C2(n15380), .A(n15373), .B(n15372), .ZN(
        n15393) );
  INV_X1 U16948 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15375) );
  AOI22_X1 U16949 ( .A1(n15382), .A2(n15393), .B1(n15375), .B2(n9009), .ZN(
        P3_U3414) );
  INV_X1 U16950 ( .A(n15376), .ZN(n15379) );
  AOI211_X1 U16951 ( .C1(n15380), .C2(n15379), .A(n15378), .B(n15377), .ZN(
        n15395) );
  INV_X1 U16952 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15381) );
  AOI22_X1 U16953 ( .A1(n15382), .A2(n15395), .B1(n15381), .B2(n9009), .ZN(
        P3_U3417) );
  AOI22_X1 U16954 ( .A1(n15396), .A2(n15383), .B1(n9710), .B2(n15394), .ZN(
        P3_U3460) );
  AOI22_X1 U16955 ( .A1(n15396), .A2(n15384), .B1(n9717), .B2(n15394), .ZN(
        P3_U3461) );
  AOI22_X1 U16956 ( .A1(n15396), .A2(n15385), .B1(n9723), .B2(n15394), .ZN(
        P3_U3462) );
  AOI22_X1 U16957 ( .A1(n15396), .A2(n15387), .B1(n15386), .B2(n15394), .ZN(
        P3_U3463) );
  AOI22_X1 U16958 ( .A1(n15396), .A2(n15388), .B1(n9733), .B2(n15394), .ZN(
        P3_U3464) );
  AOI22_X1 U16959 ( .A1(n15396), .A2(n15390), .B1(n15389), .B2(n15394), .ZN(
        P3_U3465) );
  AOI22_X1 U16960 ( .A1(n15396), .A2(n15391), .B1(n9743), .B2(n15394), .ZN(
        P3_U3466) );
  AOI22_X1 U16961 ( .A1(n15396), .A2(n15393), .B1(n15392), .B2(n15394), .ZN(
        P3_U3467) );
  AOI22_X1 U16962 ( .A1(n15396), .A2(n15395), .B1(n11058), .B2(n15394), .ZN(
        P3_U3468) );
  OR2_X1 U16963 ( .A1(n15399), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n15397) );
  AOI22_X1 U16964 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n15399), .B1(n15398), 
        .B2(n15397), .ZN(n15785) );
  XNOR2_X1 U16965 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15400) );
  XNOR2_X1 U16966 ( .A(n15400), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n15782) );
  OAI22_X1 U16967 ( .A1(SI_25_), .A2(keyinput_g7), .B1(SI_2_), .B2(
        keyinput_g30), .ZN(n15401) );
  AOI221_X1 U16968 ( .B1(SI_25_), .B2(keyinput_g7), .C1(keyinput_g30), .C2(
        SI_2_), .A(n15401), .ZN(n15408) );
  OAI22_X1 U16969 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(
        P3_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .ZN(n15402) );
  AOI221_X1 U16970 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        keyinput_g78), .C2(P3_DATAO_REG_18__SCAN_IN), .A(n15402), .ZN(n15407)
         );
  OAI22_X1 U16971 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(keyinput_g52), .B1(
        P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .ZN(n15403) );
  AOI221_X1 U16972 ( .B1(P3_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g85), .C2(P3_DATAO_REG_11__SCAN_IN), .A(n15403), .ZN(n15406)
         );
  OAI22_X1 U16973 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P3_DATAO_REG_3__SCAN_IN), .B2(keyinput_g93), .ZN(n15404) );
  AOI221_X1 U16974 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g93), .C2(P3_DATAO_REG_3__SCAN_IN), .A(n15404), .ZN(n15405)
         );
  NAND4_X1 U16975 ( .A1(n15408), .A2(n15407), .A3(n15406), .A4(n15405), .ZN(
        n15438) );
  OAI22_X1 U16976 ( .A1(SI_31_), .A2(keyinput_g1), .B1(keyinput_g75), .B2(
        P3_DATAO_REG_21__SCAN_IN), .ZN(n15409) );
  AOI221_X1 U16977 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P3_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n15409), .ZN(n15416)
         );
  OAI22_X1 U16978 ( .A1(SI_11_), .A2(keyinput_g21), .B1(keyinput_g79), .B2(
        P3_DATAO_REG_17__SCAN_IN), .ZN(n15410) );
  AOI221_X1 U16979 ( .B1(SI_11_), .B2(keyinput_g21), .C1(
        P3_DATAO_REG_17__SCAN_IN), .C2(keyinput_g79), .A(n15410), .ZN(n15415)
         );
  OAI22_X1 U16980 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(keyinput_g105), .B1(
        P3_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .ZN(n15411) );
  AOI221_X1 U16981 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(keyinput_g105), .C1(
        keyinput_g82), .C2(P3_DATAO_REG_14__SCAN_IN), .A(n15411), .ZN(n15414)
         );
  OAI22_X1 U16982 ( .A1(P3_DATAO_REG_31__SCAN_IN), .A2(keyinput_g65), .B1(
        P3_DATAO_REG_6__SCAN_IN), .B2(keyinput_g90), .ZN(n15412) );
  AOI221_X1 U16983 ( .B1(P3_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .C1(
        keyinput_g90), .C2(P3_DATAO_REG_6__SCAN_IN), .A(n15412), .ZN(n15413)
         );
  NAND4_X1 U16984 ( .A1(n15416), .A2(n15415), .A3(n15414), .A4(n15413), .ZN(
        n15437) );
  OAI22_X1 U16985 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .ZN(n15417) );
  AOI221_X1 U16986 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        keyinput_g44), .C2(P3_REG3_REG_1__SCAN_IN), .A(n15417), .ZN(n15424) );
  OAI22_X1 U16987 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(keyinput_g100), .B1(
        P3_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .ZN(n15418) );
  AOI221_X1 U16988 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_g100), .C1(
        keyinput_g83), .C2(P3_DATAO_REG_13__SCAN_IN), .A(n15418), .ZN(n15423)
         );
  OAI22_X1 U16989 ( .A1(SI_6_), .A2(keyinput_g26), .B1(keyinput_g99), .B2(
        P3_ADDR_REG_2__SCAN_IN), .ZN(n15419) );
  AOI221_X1 U16990 ( .B1(SI_6_), .B2(keyinput_g26), .C1(P3_ADDR_REG_2__SCAN_IN), .C2(keyinput_g99), .A(n15419), .ZN(n15422) );
  OAI22_X1 U16991 ( .A1(SI_24_), .A2(keyinput_g8), .B1(keyinput_g94), .B2(
        P3_DATAO_REG_2__SCAN_IN), .ZN(n15420) );
  AOI221_X1 U16992 ( .B1(SI_24_), .B2(keyinput_g8), .C1(
        P3_DATAO_REG_2__SCAN_IN), .C2(keyinput_g94), .A(n15420), .ZN(n15421)
         );
  NAND4_X1 U16993 ( .A1(n15424), .A2(n15423), .A3(n15422), .A4(n15421), .ZN(
        n15436) );
  OAI22_X1 U16994 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        keyinput_g56), .B2(P3_REG3_REG_13__SCAN_IN), .ZN(n15425) );
  AOI221_X1 U16995 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n15425), .ZN(n15434)
         );
  OAI22_X1 U16996 ( .A1(SI_29_), .A2(keyinput_g3), .B1(keyinput_g110), .B2(
        P1_IR_REG_3__SCAN_IN), .ZN(n15426) );
  AOI221_X1 U16997 ( .B1(SI_29_), .B2(keyinput_g3), .C1(P1_IR_REG_3__SCAN_IN), 
        .C2(keyinput_g110), .A(n15426), .ZN(n15433) );
  OAI22_X1 U16998 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(SI_8_), .B2(keyinput_g24), .ZN(n15427) );
  AOI221_X1 U16999 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        keyinput_g24), .C2(SI_8_), .A(n15427), .ZN(n15432) );
  XNOR2_X1 U17000 ( .A(n15428), .B(keyinput_g109), .ZN(n15430) );
  XNOR2_X1 U17001 ( .A(SI_20_), .B(keyinput_g12), .ZN(n15429) );
  NOR2_X1 U17002 ( .A1(n15430), .A2(n15429), .ZN(n15431) );
  NAND4_X1 U17003 ( .A1(n15434), .A2(n15433), .A3(n15432), .A4(n15431), .ZN(
        n15435) );
  NOR4_X1 U17004 ( .A1(n15438), .A2(n15437), .A3(n15436), .A4(n15435), .ZN(
        n15780) );
  OAI22_X1 U17005 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_g124), .ZN(n15439) );
  AOI221_X1 U17006 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        keyinput_g124), .C2(P1_IR_REG_17__SCAN_IN), .A(n15439), .ZN(n15446) );
  OAI22_X1 U17007 ( .A1(SI_18_), .A2(keyinput_g14), .B1(P1_IR_REG_12__SCAN_IN), 
        .B2(keyinput_g119), .ZN(n15440) );
  AOI221_X1 U17008 ( .B1(SI_18_), .B2(keyinput_g14), .C1(keyinput_g119), .C2(
        P1_IR_REG_12__SCAN_IN), .A(n15440), .ZN(n15445) );
  OAI22_X1 U17009 ( .A1(SI_19_), .A2(keyinput_g13), .B1(keyinput_g87), .B2(
        P3_DATAO_REG_9__SCAN_IN), .ZN(n15441) );
  AOI221_X1 U17010 ( .B1(SI_19_), .B2(keyinput_g13), .C1(
        P3_DATAO_REG_9__SCAN_IN), .C2(keyinput_g87), .A(n15441), .ZN(n15444)
         );
  OAI22_X1 U17011 ( .A1(P3_DATAO_REG_1__SCAN_IN), .A2(keyinput_g95), .B1(
        keyinput_g86), .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n15442) );
  AOI221_X1 U17012 ( .B1(P3_DATAO_REG_1__SCAN_IN), .B2(keyinput_g95), .C1(
        P3_DATAO_REG_10__SCAN_IN), .C2(keyinput_g86), .A(n15442), .ZN(n15443)
         );
  NAND4_X1 U17013 ( .A1(n15446), .A2(n15445), .A3(n15444), .A4(n15443), .ZN(
        n15583) );
  OAI22_X1 U17014 ( .A1(P3_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        keyinput_g33), .B2(P3_RD_REG_SCAN_IN), .ZN(n15447) );
  AOI221_X1 U17015 ( .B1(P3_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        P3_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n15447), .ZN(n15473) );
  OAI22_X1 U17016 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        keyinput_g17), .B2(SI_15_), .ZN(n15448) );
  AOI221_X1 U17017 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        SI_15_), .C2(keyinput_g17), .A(n15448), .ZN(n15451) );
  OAI22_X1 U17018 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_g113), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_g112), .ZN(n15449) );
  AOI221_X1 U17019 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_g113), .C1(
        keyinput_g112), .C2(P1_IR_REG_5__SCAN_IN), .A(n15449), .ZN(n15450) );
  OAI211_X1 U17020 ( .C1(n15453), .C2(keyinput_g16), .A(n15451), .B(n15450), 
        .ZN(n15452) );
  AOI21_X1 U17021 ( .B1(n15453), .B2(keyinput_g16), .A(n15452), .ZN(n15472) );
  AOI22_X1 U17022 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_g104), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n15454) );
  OAI221_X1 U17023 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_g104), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n15454), .ZN(n15461)
         );
  AOI22_X1 U17024 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(n6889), .B2(keyinput_g107), .ZN(n15455) );
  OAI221_X1 U17025 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        n6889), .C2(keyinput_g107), .A(n15455), .ZN(n15460) );
  AOI22_X1 U17026 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g120), .B1(
        P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n15456) );
  OAI221_X1 U17027 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g120), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n15456), .ZN(n15459) );
  AOI22_X1 U17028 ( .A1(P3_DATAO_REG_7__SCAN_IN), .A2(keyinput_g89), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .ZN(n15457) );
  OAI221_X1 U17029 ( .B1(P3_DATAO_REG_7__SCAN_IN), .B2(keyinput_g89), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_g35), .A(n15457), .ZN(n15458) );
  NOR4_X1 U17030 ( .A1(n15461), .A2(n15460), .A3(n15459), .A4(n15458), .ZN(
        n15471) );
  AOI22_X1 U17031 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_g111), .B1(SI_21_), 
        .B2(keyinput_g11), .ZN(n15462) );
  OAI221_X1 U17032 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_g111), .C1(SI_21_), .C2(keyinput_g11), .A(n15462), .ZN(n15469) );
  AOI22_X1 U17033 ( .A1(P3_DATAO_REG_12__SCAN_IN), .A2(keyinput_g84), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_g114), .ZN(n15463) );
  OAI221_X1 U17034 ( .B1(P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_g114), .A(n15463), .ZN(n15468) );
  AOI22_X1 U17035 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(keyinput_g106), .B1(SI_4_), .B2(keyinput_g28), .ZN(n15464) );
  OAI221_X1 U17036 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(keyinput_g106), .C1(
        SI_4_), .C2(keyinput_g28), .A(n15464), .ZN(n15467) );
  AOI22_X1 U17037 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(keyinput_g66), .B1(
        SI_7_), .B2(keyinput_g25), .ZN(n15465) );
  OAI221_X1 U17038 ( .B1(P3_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .C1(
        SI_7_), .C2(keyinput_g25), .A(n15465), .ZN(n15466) );
  NOR4_X1 U17039 ( .A1(n15469), .A2(n15468), .A3(n15467), .A4(n15466), .ZN(
        n15470) );
  NAND4_X1 U17040 ( .A1(n15473), .A2(n15472), .A3(n15471), .A4(n15470), .ZN(
        n15582) );
  AOI22_X1 U17041 ( .A1(n15475), .A2(keyinput_g98), .B1(keyinput_g92), .B2(
        n15744), .ZN(n15474) );
  OAI221_X1 U17042 ( .B1(n15475), .B2(keyinput_g98), .C1(n15744), .C2(
        keyinput_g92), .A(n15474), .ZN(n15487) );
  AOI22_X1 U17043 ( .A1(n15478), .A2(keyinput_g9), .B1(keyinput_g69), .B2(
        n15477), .ZN(n15476) );
  OAI221_X1 U17044 ( .B1(n15478), .B2(keyinput_g9), .C1(n15477), .C2(
        keyinput_g69), .A(n15476), .ZN(n15486) );
  AOI22_X1 U17045 ( .A1(n15481), .A2(keyinput_g46), .B1(keyinput_g20), .B2(
        n15480), .ZN(n15479) );
  OAI221_X1 U17046 ( .B1(n15481), .B2(keyinput_g46), .C1(n15480), .C2(
        keyinput_g20), .A(n15479), .ZN(n15485) );
  XOR2_X1 U17047 ( .A(n8101), .B(keyinput_g122), .Z(n15483) );
  XNOR2_X1 U17048 ( .A(SI_5_), .B(keyinput_g27), .ZN(n15482) );
  NAND2_X1 U17049 ( .A1(n15483), .A2(n15482), .ZN(n15484) );
  NOR4_X1 U17050 ( .A1(n15487), .A2(n15486), .A3(n15485), .A4(n15484), .ZN(
        n15525) );
  AOI22_X1 U17051 ( .A1(n15489), .A2(keyinput_g96), .B1(n8550), .B2(
        keyinput_g49), .ZN(n15488) );
  OAI221_X1 U17052 ( .B1(n15489), .B2(keyinput_g96), .C1(n8550), .C2(
        keyinput_g49), .A(n15488), .ZN(n15498) );
  AOI22_X1 U17053 ( .A1(n15491), .A2(keyinput_g67), .B1(n8508), .B2(
        keyinput_g59), .ZN(n15490) );
  OAI221_X1 U17054 ( .B1(n15491), .B2(keyinput_g67), .C1(n8508), .C2(
        keyinput_g59), .A(n15490), .ZN(n15497) );
  AOI22_X1 U17055 ( .A1(n15732), .A2(keyinput_g72), .B1(n15706), .B2(
        keyinput_g80), .ZN(n15492) );
  OAI221_X1 U17056 ( .B1(n15732), .B2(keyinput_g72), .C1(n15706), .C2(
        keyinput_g80), .A(n15492), .ZN(n15496) );
  AOI22_X1 U17057 ( .A1(n8388), .A2(keyinput_g63), .B1(keyinput_g5), .B2(
        n15494), .ZN(n15493) );
  OAI221_X1 U17058 ( .B1(n8388), .B2(keyinput_g63), .C1(n15494), .C2(
        keyinput_g5), .A(n15493), .ZN(n15495) );
  NOR4_X1 U17059 ( .A1(n15498), .A2(n15497), .A3(n15496), .A4(n15495), .ZN(
        n15524) );
  INV_X1 U17060 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15701) );
  AOI22_X1 U17061 ( .A1(n15701), .A2(keyinput_g101), .B1(n15500), .B2(
        keyinput_g103), .ZN(n15499) );
  OAI221_X1 U17062 ( .B1(n15701), .B2(keyinput_g101), .C1(n15500), .C2(
        keyinput_g103), .A(n15499), .ZN(n15510) );
  AOI22_X1 U17063 ( .A1(n15503), .A2(keyinput_g22), .B1(keyinput_g68), .B2(
        n15502), .ZN(n15501) );
  OAI221_X1 U17064 ( .B1(n15503), .B2(keyinput_g22), .C1(n15502), .C2(
        keyinput_g68), .A(n15501), .ZN(n15509) );
  AOI22_X1 U17065 ( .A1(n15660), .A2(keyinput_g4), .B1(n15658), .B2(
        keyinput_g55), .ZN(n15504) );
  OAI221_X1 U17066 ( .B1(n15660), .B2(keyinput_g4), .C1(n15658), .C2(
        keyinput_g55), .A(n15504), .ZN(n15508) );
  XNOR2_X1 U17067 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g127), .ZN(n15506)
         );
  XNOR2_X1 U17068 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_g34), .ZN(n15505) );
  NAND2_X1 U17069 ( .A1(n15506), .A2(n15505), .ZN(n15507) );
  NOR4_X1 U17070 ( .A1(n15510), .A2(n15509), .A3(n15508), .A4(n15507), .ZN(
        n15523) );
  INV_X1 U17071 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15662) );
  AOI22_X1 U17072 ( .A1(n15662), .A2(keyinput_g39), .B1(keyinput_g32), .B2(
        n9808), .ZN(n15511) );
  OAI221_X1 U17073 ( .B1(n15662), .B2(keyinput_g39), .C1(n9808), .C2(
        keyinput_g32), .A(n15511), .ZN(n15521) );
  AOI22_X1 U17074 ( .A1(n15724), .A2(keyinput_g77), .B1(n15673), .B2(
        keyinput_g6), .ZN(n15512) );
  OAI221_X1 U17075 ( .B1(n15724), .B2(keyinput_g77), .C1(n15673), .C2(
        keyinput_g6), .A(n15512), .ZN(n15520) );
  AOI22_X1 U17076 ( .A1(n15514), .A2(keyinput_g97), .B1(n15756), .B2(
        keyinput_g38), .ZN(n15513) );
  OAI221_X1 U17077 ( .B1(n15514), .B2(keyinput_g97), .C1(n15756), .C2(
        keyinput_g38), .A(n15513), .ZN(n15519) );
  INV_X1 U17078 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U17079 ( .A1(n15517), .A2(keyinput_g2), .B1(n15516), .B2(
        keyinput_g60), .ZN(n15515) );
  OAI221_X1 U17080 ( .B1(n15517), .B2(keyinput_g2), .C1(n15516), .C2(
        keyinput_g60), .A(n15515), .ZN(n15518) );
  NOR4_X1 U17081 ( .A1(n15521), .A2(n15520), .A3(n15519), .A4(n15518), .ZN(
        n15522) );
  NAND4_X1 U17082 ( .A1(n15525), .A2(n15524), .A3(n15523), .A4(n15522), .ZN(
        n15581) );
  AOI22_X1 U17083 ( .A1(n15723), .A2(keyinput_g19), .B1(keyinput_g115), .B2(
        n8003), .ZN(n15526) );
  OAI221_X1 U17084 ( .B1(n15723), .B2(keyinput_g19), .C1(n8003), .C2(
        keyinput_g115), .A(n15526), .ZN(n15537) );
  INV_X1 U17085 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15528) );
  AOI22_X1 U17086 ( .A1(n15528), .A2(keyinput_g0), .B1(keyinput_g81), .B2(
        n15731), .ZN(n15527) );
  OAI221_X1 U17087 ( .B1(n15528), .B2(keyinput_g0), .C1(n15731), .C2(
        keyinput_g81), .A(n15527), .ZN(n15536) );
  INV_X1 U17088 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15531) );
  AOI22_X1 U17089 ( .A1(n15531), .A2(keyinput_g37), .B1(keyinput_g91), .B2(
        n15530), .ZN(n15529) );
  OAI221_X1 U17090 ( .B1(n15531), .B2(keyinput_g37), .C1(n15530), .C2(
        keyinput_g91), .A(n15529), .ZN(n15535) );
  INV_X1 U17091 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15746) );
  AOI22_X1 U17092 ( .A1(n15533), .A2(keyinput_g70), .B1(n15746), .B2(
        keyinput_g41), .ZN(n15532) );
  OAI221_X1 U17093 ( .B1(n15533), .B2(keyinput_g70), .C1(n15746), .C2(
        keyinput_g41), .A(n15532), .ZN(n15534) );
  NOR4_X1 U17094 ( .A1(n15537), .A2(n15536), .A3(n15535), .A4(n15534), .ZN(
        n15579) );
  AOI22_X1 U17095 ( .A1(n15539), .A2(keyinput_g117), .B1(n8621), .B2(
        keyinput_g53), .ZN(n15538) );
  OAI221_X1 U17096 ( .B1(n15539), .B2(keyinput_g117), .C1(n8621), .C2(
        keyinput_g53), .A(n15538), .ZN(n15551) );
  AOI22_X1 U17097 ( .A1(n15542), .A2(keyinput_g18), .B1(keyinput_g118), .B2(
        n15541), .ZN(n15540) );
  OAI221_X1 U17098 ( .B1(n15542), .B2(keyinput_g18), .C1(n15541), .C2(
        keyinput_g118), .A(n15540), .ZN(n15550) );
  INV_X1 U17099 ( .A(P3_B_REG_SCAN_IN), .ZN(n15544) );
  AOI22_X1 U17100 ( .A1(n15545), .A2(keyinput_g15), .B1(n15544), .B2(
        keyinput_g64), .ZN(n15543) );
  OAI221_X1 U17101 ( .B1(n15545), .B2(keyinput_g15), .C1(n15544), .C2(
        keyinput_g64), .A(n15543), .ZN(n15549) );
  XOR2_X1 U17102 ( .A(n6979), .B(keyinput_g102), .Z(n15547) );
  XNOR2_X1 U17103 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g125), .ZN(n15546)
         );
  NAND2_X1 U17104 ( .A1(n15547), .A2(n15546), .ZN(n15548) );
  NOR4_X1 U17105 ( .A1(n15551), .A2(n15550), .A3(n15549), .A4(n15548), .ZN(
        n15578) );
  AOI22_X1 U17106 ( .A1(n15553), .A2(keyinput_g116), .B1(n8289), .B2(
        keyinput_g126), .ZN(n15552) );
  OAI221_X1 U17107 ( .B1(n15553), .B2(keyinput_g116), .C1(n8289), .C2(
        keyinput_g126), .A(n15552), .ZN(n15563) );
  AOI22_X1 U17108 ( .A1(n15556), .A2(keyinput_g42), .B1(keyinput_g62), .B2(
        n15555), .ZN(n15554) );
  OAI221_X1 U17109 ( .B1(n15556), .B2(keyinput_g42), .C1(n15555), .C2(
        keyinput_g62), .A(n15554), .ZN(n15562) );
  XNOR2_X1 U17110 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g108), .ZN(n15560)
         );
  XNOR2_X1 U17111 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_g121), .ZN(n15559)
         );
  XNOR2_X1 U17112 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_g123), .ZN(n15558)
         );
  XNOR2_X1 U17113 ( .A(SI_3_), .B(keyinput_g29), .ZN(n15557) );
  NAND4_X1 U17114 ( .A1(n15560), .A2(n15559), .A3(n15558), .A4(n15557), .ZN(
        n15561) );
  NOR3_X1 U17115 ( .A1(n15563), .A2(n15562), .A3(n15561), .ZN(n15577) );
  AOI22_X1 U17116 ( .A1(n15566), .A2(keyinput_g73), .B1(n15565), .B2(
        keyinput_g71), .ZN(n15564) );
  OAI221_X1 U17117 ( .B1(n15566), .B2(keyinput_g73), .C1(n15565), .C2(
        keyinput_g71), .A(n15564), .ZN(n15575) );
  AOI22_X1 U17118 ( .A1(n15749), .A2(keyinput_g43), .B1(keyinput_g74), .B2(
        n15674), .ZN(n15567) );
  OAI221_X1 U17119 ( .B1(n15749), .B2(keyinput_g43), .C1(n15674), .C2(
        keyinput_g74), .A(n15567), .ZN(n15574) );
  INV_X1 U17120 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15569) );
  AOI22_X1 U17121 ( .A1(n15742), .A2(keyinput_g10), .B1(n15569), .B2(
        keyinput_g36), .ZN(n15568) );
  OAI221_X1 U17122 ( .B1(n15742), .B2(keyinput_g10), .C1(n15569), .C2(
        keyinput_g36), .A(n15568), .ZN(n15573) );
  XNOR2_X1 U17123 ( .A(SI_1_), .B(keyinput_g31), .ZN(n15571) );
  XNOR2_X1 U17124 ( .A(SI_9_), .B(keyinput_g23), .ZN(n15570) );
  NAND2_X1 U17125 ( .A1(n15571), .A2(n15570), .ZN(n15572) );
  NOR4_X1 U17126 ( .A1(n15575), .A2(n15574), .A3(n15573), .A4(n15572), .ZN(
        n15576) );
  NAND4_X1 U17127 ( .A1(n15579), .A2(n15578), .A3(n15577), .A4(n15576), .ZN(
        n15580) );
  NOR4_X1 U17128 ( .A1(n15583), .A2(n15582), .A3(n15581), .A4(n15580), .ZN(
        n15779) );
  XOR2_X1 U17129 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_f93), .Z(n15590)
         );
  AOI22_X1 U17130 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(keyinput_f103), .B1(
        P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n15584) );
  OAI221_X1 U17131 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_f103), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n15584), .ZN(n15589) );
  AOI22_X1 U17132 ( .A1(n6889), .A2(keyinput_f107), .B1(P1_IR_REG_4__SCAN_IN), 
        .B2(keyinput_f111), .ZN(n15585) );
  OAI221_X1 U17133 ( .B1(n6889), .B2(keyinput_f107), .C1(P1_IR_REG_4__SCAN_IN), 
        .C2(keyinput_f111), .A(n15585), .ZN(n15588) );
  AOI22_X1 U17134 ( .A1(keyinput_f82), .A2(P3_DATAO_REG_14__SCAN_IN), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_f126), .ZN(n15586) );
  OAI221_X1 U17135 ( .B1(keyinput_f82), .B2(P3_DATAO_REG_14__SCAN_IN), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_f126), .A(n15586), .ZN(n15587) );
  NOR4_X1 U17136 ( .A1(n15590), .A2(n15589), .A3(n15588), .A4(n15587), .ZN(
        n15618) );
  AOI22_X1 U17137 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f113), .B1(SI_12_), 
        .B2(keyinput_f20), .ZN(n15591) );
  OAI221_X1 U17138 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f113), .C1(SI_12_), .C2(keyinput_f20), .A(n15591), .ZN(n15598) );
  AOI22_X1 U17139 ( .A1(SI_9_), .A2(keyinput_f23), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n15592) );
  OAI221_X1 U17140 ( .B1(SI_9_), .B2(keyinput_f23), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n15592), .ZN(n15597) );
  AOI22_X1 U17141 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(keyinput_f102), .B1(
        P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_f99), .ZN(n15593) );
  OAI221_X1 U17142 ( .B1(P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_f102), .C1(
        P3_ADDR_REG_2__SCAN_IN), .C2(keyinput_f99), .A(n15593), .ZN(n15596) );
  AOI22_X1 U17143 ( .A1(keyinput_f91), .A2(P3_DATAO_REG_5__SCAN_IN), .B1(
        SI_11_), .B2(keyinput_f21), .ZN(n15594) );
  OAI221_X1 U17144 ( .B1(keyinput_f91), .B2(P3_DATAO_REG_5__SCAN_IN), .C1(
        SI_11_), .C2(keyinput_f21), .A(n15594), .ZN(n15595) );
  NOR4_X1 U17145 ( .A1(n15598), .A2(n15597), .A3(n15596), .A4(n15595), .ZN(
        n15617) );
  AOI22_X1 U17146 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(keyinput_f69), .B1(
        keyinput_f68), .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n15599) );
  OAI221_X1 U17147 ( .B1(P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .C1(
        keyinput_f68), .C2(P3_DATAO_REG_28__SCAN_IN), .A(n15599), .ZN(n15606)
         );
  AOI22_X1 U17148 ( .A1(keyinput_f71), .A2(P3_DATAO_REG_25__SCAN_IN), .B1(
        keyinput_f88), .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n15600) );
  OAI221_X1 U17149 ( .B1(keyinput_f71), .B2(P3_DATAO_REG_25__SCAN_IN), .C1(
        keyinput_f88), .C2(P3_DATAO_REG_8__SCAN_IN), .A(n15600), .ZN(n15605)
         );
  AOI22_X1 U17150 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_f117), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_f109), .ZN(n15601) );
  OAI221_X1 U17151 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_f117), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput_f109), .A(n15601), .ZN(n15604) );
  AOI22_X1 U17152 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_f114), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n15602) );
  OAI221_X1 U17153 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_f114), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n15602), .ZN(n15603)
         );
  NOR4_X1 U17154 ( .A1(n15606), .A2(n15605), .A3(n15604), .A4(n15603), .ZN(
        n15616) );
  AOI22_X1 U17155 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f120), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n15607) );
  OAI221_X1 U17156 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f120), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n15607), .ZN(n15614)
         );
  AOI22_X1 U17157 ( .A1(SI_21_), .A2(keyinput_f11), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n15608) );
  OAI221_X1 U17158 ( .B1(SI_21_), .B2(keyinput_f11), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n15608), .ZN(n15613)
         );
  AOI22_X1 U17159 ( .A1(SI_16_), .A2(keyinput_f16), .B1(SI_10_), .B2(
        keyinput_f22), .ZN(n15609) );
  OAI221_X1 U17160 ( .B1(SI_16_), .B2(keyinput_f16), .C1(SI_10_), .C2(
        keyinput_f22), .A(n15609), .ZN(n15612) );
  AOI22_X1 U17161 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_14_), .B2(
        keyinput_f18), .ZN(n15610) );
  OAI221_X1 U17162 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_14_), .C2(
        keyinput_f18), .A(n15610), .ZN(n15611) );
  NOR4_X1 U17163 ( .A1(n15614), .A2(n15613), .A3(n15612), .A4(n15611), .ZN(
        n15615) );
  NAND4_X1 U17164 ( .A1(n15618), .A2(n15617), .A3(n15616), .A4(n15615), .ZN(
        n15773) );
  AOI22_X1 U17165 ( .A1(keyinput_f95), .A2(P3_DATAO_REG_1__SCAN_IN), .B1(
        keyinput_f73), .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n15619) );
  OAI221_X1 U17166 ( .B1(keyinput_f95), .B2(P3_DATAO_REG_1__SCAN_IN), .C1(
        keyinput_f73), .C2(P3_DATAO_REG_23__SCAN_IN), .A(n15619), .ZN(n15626)
         );
  AOI22_X1 U17167 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P3_B_REG_SCAN_IN), .B2(
        keyinput_f64), .ZN(n15620) );
  OAI221_X1 U17168 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P3_B_REG_SCAN_IN), 
        .C2(keyinput_f64), .A(n15620), .ZN(n15625) );
  AOI22_X1 U17169 ( .A1(keyinput_f86), .A2(P3_DATAO_REG_10__SCAN_IN), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n15621) );
  OAI221_X1 U17170 ( .B1(keyinput_f86), .B2(P3_DATAO_REG_10__SCAN_IN), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n15621), .ZN(n15624)
         );
  AOI22_X1 U17171 ( .A1(keyinput_f67), .A2(P3_DATAO_REG_29__SCAN_IN), .B1(
        SI_8_), .B2(keyinput_f24), .ZN(n15622) );
  OAI221_X1 U17172 ( .B1(keyinput_f67), .B2(P3_DATAO_REG_29__SCAN_IN), .C1(
        SI_8_), .C2(keyinput_f24), .A(n15622), .ZN(n15623) );
  NOR4_X1 U17173 ( .A1(n15626), .A2(n15625), .A3(n15624), .A4(n15623), .ZN(
        n15654) );
  AOI22_X1 U17174 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f118), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n15627) );
  OAI221_X1 U17175 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f118), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n15627), .ZN(n15634)
         );
  AOI22_X1 U17176 ( .A1(keyinput_f70), .A2(P3_DATAO_REG_26__SCAN_IN), .B1(
        SI_0_), .B2(keyinput_f32), .ZN(n15628) );
  OAI221_X1 U17177 ( .B1(keyinput_f70), .B2(P3_DATAO_REG_26__SCAN_IN), .C1(
        SI_0_), .C2(keyinput_f32), .A(n15628), .ZN(n15633) );
  AOI22_X1 U17178 ( .A1(keyinput_f94), .A2(P3_DATAO_REG_2__SCAN_IN), .B1(
        SI_18_), .B2(keyinput_f14), .ZN(n15629) );
  OAI221_X1 U17179 ( .B1(keyinput_f94), .B2(P3_DATAO_REG_2__SCAN_IN), .C1(
        SI_18_), .C2(keyinput_f14), .A(n15629), .ZN(n15632) );
  AOI22_X1 U17180 ( .A1(keyinput_f79), .A2(P3_DATAO_REG_17__SCAN_IN), .B1(
        SI_15_), .B2(keyinput_f17), .ZN(n15630) );
  OAI221_X1 U17181 ( .B1(keyinput_f79), .B2(P3_DATAO_REG_17__SCAN_IN), .C1(
        SI_15_), .C2(keyinput_f17), .A(n15630), .ZN(n15631) );
  NOR4_X1 U17182 ( .A1(n15634), .A2(n15633), .A3(n15632), .A4(n15631), .ZN(
        n15653) );
  AOI22_X1 U17183 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput_f98), .B1(SI_19_), .B2(keyinput_f13), .ZN(n15635) );
  OAI221_X1 U17184 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput_f98), .C1(
        SI_19_), .C2(keyinput_f13), .A(n15635), .ZN(n15642) );
  AOI22_X1 U17185 ( .A1(keyinput_f87), .A2(P3_DATAO_REG_9__SCAN_IN), .B1(
        SI_23_), .B2(keyinput_f9), .ZN(n15636) );
  OAI221_X1 U17186 ( .B1(keyinput_f87), .B2(P3_DATAO_REG_9__SCAN_IN), .C1(
        SI_23_), .C2(keyinput_f9), .A(n15636), .ZN(n15641) );
  AOI22_X1 U17187 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(keyinput_f106), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n15637) );
  OAI221_X1 U17188 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(keyinput_f106), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n15637), .ZN(n15640)
         );
  AOI22_X1 U17189 ( .A1(keyinput_f76), .A2(P3_DATAO_REG_20__SCAN_IN), .B1(
        keyinput_f65), .B2(P3_DATAO_REG_31__SCAN_IN), .ZN(n15638) );
  OAI221_X1 U17190 ( .B1(keyinput_f76), .B2(P3_DATAO_REG_20__SCAN_IN), .C1(
        keyinput_f65), .C2(P3_DATAO_REG_31__SCAN_IN), .A(n15638), .ZN(n15639)
         );
  NOR4_X1 U17191 ( .A1(n15642), .A2(n15641), .A3(n15640), .A4(n15639), .ZN(
        n15652) );
  AOI22_X1 U17192 ( .A1(SI_17_), .A2(keyinput_f15), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n15643) );
  OAI221_X1 U17193 ( .B1(SI_17_), .B2(keyinput_f15), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n15643), .ZN(n15650)
         );
  AOI22_X1 U17194 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(keyinput_f97), .B1(SI_20_), .B2(keyinput_f12), .ZN(n15644) );
  OAI221_X1 U17195 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(keyinput_f97), .C1(
        SI_20_), .C2(keyinput_f12), .A(n15644), .ZN(n15649) );
  AOI22_X1 U17196 ( .A1(keyinput_f96), .A2(P3_DATAO_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n15645) );
  OAI221_X1 U17197 ( .B1(keyinput_f96), .B2(P3_DATAO_REG_0__SCAN_IN), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n15645), .ZN(n15648)
         );
  AOI22_X1 U17198 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .ZN(n15646) );
  OAI221_X1 U17199 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n15646), .ZN(n15647)
         );
  NOR4_X1 U17200 ( .A1(n15650), .A2(n15649), .A3(n15648), .A4(n15647), .ZN(
        n15651) );
  NAND4_X1 U17201 ( .A1(n15654), .A2(n15653), .A3(n15652), .A4(n15651), .ZN(
        n15772) );
  AOI22_X1 U17202 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_f116), .B1(
        P3_U3151), .B2(keyinput_f34), .ZN(n15655) );
  OAI221_X1 U17203 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_f116), .C1(
        P3_U3151), .C2(keyinput_f34), .A(n15655), .ZN(n15667) );
  INV_X1 U17204 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U17205 ( .A1(n15658), .A2(keyinput_f55), .B1(keyinput_f104), .B2(
        n15657), .ZN(n15656) );
  OAI221_X1 U17206 ( .B1(n15658), .B2(keyinput_f55), .C1(n15657), .C2(
        keyinput_f104), .A(n15656), .ZN(n15666) );
  AOI22_X1 U17207 ( .A1(n11272), .A2(keyinput_f8), .B1(n15660), .B2(
        keyinput_f4), .ZN(n15659) );
  OAI221_X1 U17208 ( .B1(n11272), .B2(keyinput_f8), .C1(n15660), .C2(
        keyinput_f4), .A(n15659), .ZN(n15665) );
  INV_X1 U17209 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n15663) );
  AOI22_X1 U17210 ( .A1(n15663), .A2(keyinput_f119), .B1(n15662), .B2(
        keyinput_f39), .ZN(n15661) );
  OAI221_X1 U17211 ( .B1(n15663), .B2(keyinput_f119), .C1(n15662), .C2(
        keyinput_f39), .A(n15661), .ZN(n15664) );
  NOR4_X1 U17212 ( .A1(n15667), .A2(n15666), .A3(n15665), .A4(n15664), .ZN(
        n15713) );
  INV_X1 U17213 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15669) );
  AOI22_X1 U17214 ( .A1(n15669), .A2(keyinput_f100), .B1(n8101), .B2(
        keyinput_f122), .ZN(n15668) );
  OAI221_X1 U17215 ( .B1(n15669), .B2(keyinput_f100), .C1(n8101), .C2(
        keyinput_f122), .A(n15668), .ZN(n15680) );
  AOI22_X1 U17216 ( .A1(n15671), .A2(keyinput_f83), .B1(n6854), .B2(
        keyinput_f124), .ZN(n15670) );
  OAI221_X1 U17217 ( .B1(n15671), .B2(keyinput_f83), .C1(n6854), .C2(
        keyinput_f124), .A(n15670), .ZN(n15679) );
  AOI22_X1 U17218 ( .A1(n15674), .A2(keyinput_f74), .B1(n15673), .B2(
        keyinput_f6), .ZN(n15672) );
  OAI221_X1 U17219 ( .B1(n15674), .B2(keyinput_f74), .C1(n15673), .C2(
        keyinput_f6), .A(n15672), .ZN(n15678) );
  XNOR2_X1 U17220 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_f112), .ZN(n15676)
         );
  XNOR2_X1 U17221 ( .A(SI_4_), .B(keyinput_f28), .ZN(n15675) );
  NAND2_X1 U17222 ( .A1(n15676), .A2(n15675), .ZN(n15677) );
  NOR4_X1 U17223 ( .A1(n15680), .A2(n15679), .A3(n15678), .A4(n15677), .ZN(
        n15712) );
  AOI22_X1 U17224 ( .A1(n15682), .A2(keyinput_f33), .B1(n10509), .B2(
        keyinput_f44), .ZN(n15681) );
  OAI221_X1 U17225 ( .B1(n15682), .B2(keyinput_f33), .C1(n10509), .C2(
        keyinput_f44), .A(n15681), .ZN(n15694) );
  AOI22_X1 U17226 ( .A1(n15685), .A2(keyinput_f85), .B1(keyinput_f66), .B2(
        n15684), .ZN(n15683) );
  OAI221_X1 U17227 ( .B1(n15685), .B2(keyinput_f85), .C1(n15684), .C2(
        keyinput_f66), .A(n15683), .ZN(n15693) );
  AOI22_X1 U17228 ( .A1(n8388), .A2(keyinput_f63), .B1(keyinput_f105), .B2(
        n15687), .ZN(n15686) );
  OAI221_X1 U17229 ( .B1(n8388), .B2(keyinput_f63), .C1(n15687), .C2(
        keyinput_f105), .A(n15686), .ZN(n15692) );
  AOI22_X1 U17230 ( .A1(n15690), .A2(keyinput_f84), .B1(n15689), .B2(
        keyinput_f30), .ZN(n15688) );
  OAI221_X1 U17231 ( .B1(n15690), .B2(keyinput_f84), .C1(n15689), .C2(
        keyinput_f30), .A(n15688), .ZN(n15691) );
  NOR4_X1 U17232 ( .A1(n15694), .A2(n15693), .A3(n15692), .A4(n15691), .ZN(
        n15711) );
  AOI22_X1 U17233 ( .A1(n15697), .A2(keyinput_f75), .B1(keyinput_f90), .B2(
        n15696), .ZN(n15695) );
  OAI221_X1 U17234 ( .B1(n15697), .B2(keyinput_f75), .C1(n15696), .C2(
        keyinput_f90), .A(n15695), .ZN(n15709) );
  XOR2_X1 U17235 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_f51), .Z(n15700)
         );
  XNOR2_X1 U17236 ( .A(n15698), .B(keyinput_f123), .ZN(n15699) );
  NOR2_X1 U17237 ( .A1(n15700), .A2(n15699), .ZN(n15705) );
  XNOR2_X1 U17238 ( .A(keyinput_f101), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n15704)
         );
  XNOR2_X1 U17239 ( .A(SI_1_), .B(keyinput_f31), .ZN(n15703) );
  XNOR2_X1 U17240 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f108), .ZN(n15702)
         );
  NAND4_X1 U17241 ( .A1(n15705), .A2(n15704), .A3(n15703), .A4(n15702), .ZN(
        n15708) );
  XNOR2_X1 U17242 ( .A(n15706), .B(keyinput_f80), .ZN(n15707) );
  NOR3_X1 U17243 ( .A1(n15709), .A2(n15708), .A3(n15707), .ZN(n15710) );
  NAND4_X1 U17244 ( .A1(n15713), .A2(n15712), .A3(n15711), .A4(n15710), .ZN(
        n15771) );
  AOI22_X1 U17245 ( .A1(n15716), .A2(keyinput_f78), .B1(n15715), .B2(
        keyinput_f7), .ZN(n15714) );
  OAI221_X1 U17246 ( .B1(n15716), .B2(keyinput_f78), .C1(n15715), .C2(
        keyinput_f7), .A(n15714), .ZN(n15720) );
  XNOR2_X1 U17247 ( .A(n15717), .B(keyinput_f89), .ZN(n15719) );
  XOR2_X1 U17248 ( .A(SI_3_), .B(keyinput_f29), .Z(n15718) );
  OR3_X1 U17249 ( .A1(n15720), .A2(n15719), .A3(n15718), .ZN(n15727) );
  AOI22_X1 U17250 ( .A1(n8003), .A2(keyinput_f115), .B1(n13129), .B2(
        keyinput_f3), .ZN(n15721) );
  OAI221_X1 U17251 ( .B1(n8003), .B2(keyinput_f115), .C1(n13129), .C2(
        keyinput_f3), .A(n15721), .ZN(n15726) );
  AOI22_X1 U17252 ( .A1(n15724), .A2(keyinput_f77), .B1(n15723), .B2(
        keyinput_f19), .ZN(n15722) );
  OAI221_X1 U17253 ( .B1(n15724), .B2(keyinput_f77), .C1(n15723), .C2(
        keyinput_f19), .A(n15722), .ZN(n15725) );
  NOR3_X1 U17254 ( .A1(n15727), .A2(n15726), .A3(n15725), .ZN(n15769) );
  INV_X1 U17255 ( .A(keyinput_f0), .ZN(n15729) );
  AOI22_X1 U17256 ( .A1(n15730), .A2(keyinput_f35), .B1(P3_WR_REG_SCAN_IN), 
        .B2(n15729), .ZN(n15728) );
  OAI221_X1 U17257 ( .B1(n15730), .B2(keyinput_f35), .C1(n15729), .C2(
        P3_WR_REG_SCAN_IN), .A(n15728), .ZN(n15740) );
  XNOR2_X1 U17258 ( .A(n15731), .B(keyinput_f81), .ZN(n15739) );
  XNOR2_X1 U17259 ( .A(n15732), .B(keyinput_f72), .ZN(n15738) );
  XNOR2_X1 U17260 ( .A(SI_5_), .B(keyinput_f27), .ZN(n15736) );
  XNOR2_X1 U17261 ( .A(SI_27_), .B(keyinput_f5), .ZN(n15735) );
  XNOR2_X1 U17262 ( .A(SI_6_), .B(keyinput_f26), .ZN(n15734) );
  XNOR2_X1 U17263 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_f121), .ZN(n15733)
         );
  NAND4_X1 U17264 ( .A1(n15736), .A2(n15735), .A3(n15734), .A4(n15733), .ZN(
        n15737) );
  NOR4_X1 U17265 ( .A1(n15740), .A2(n15739), .A3(n15738), .A4(n15737), .ZN(
        n15768) );
  AOI22_X1 U17266 ( .A1(n8508), .A2(keyinput_f59), .B1(n15742), .B2(
        keyinput_f10), .ZN(n15741) );
  OAI221_X1 U17267 ( .B1(n8508), .B2(keyinput_f59), .C1(n15742), .C2(
        keyinput_f10), .A(n15741), .ZN(n15754) );
  AOI22_X1 U17268 ( .A1(n8386), .A2(keyinput_f56), .B1(keyinput_f92), .B2(
        n15744), .ZN(n15743) );
  OAI221_X1 U17269 ( .B1(n8386), .B2(keyinput_f56), .C1(n15744), .C2(
        keyinput_f92), .A(n15743), .ZN(n15753) );
  AOI22_X1 U17270 ( .A1(n15747), .A2(keyinput_f58), .B1(n15746), .B2(
        keyinput_f41), .ZN(n15745) );
  OAI221_X1 U17271 ( .B1(n15747), .B2(keyinput_f58), .C1(n15746), .C2(
        keyinput_f41), .A(n15745), .ZN(n15752) );
  AOI22_X1 U17272 ( .A1(n15750), .A2(keyinput_f52), .B1(n15749), .B2(
        keyinput_f43), .ZN(n15748) );
  OAI221_X1 U17273 ( .B1(n15750), .B2(keyinput_f52), .C1(n15749), .C2(
        keyinput_f43), .A(n15748), .ZN(n15751) );
  NOR4_X1 U17274 ( .A1(n15754), .A2(n15753), .A3(n15752), .A4(n15751), .ZN(
        n15767) );
  AOI22_X1 U17275 ( .A1(n8493), .A2(keyinput_f54), .B1(n15756), .B2(
        keyinput_f38), .ZN(n15755) );
  OAI221_X1 U17276 ( .B1(n8493), .B2(keyinput_f54), .C1(n15756), .C2(
        keyinput_f38), .A(n15755), .ZN(n15765) );
  XNOR2_X1 U17277 ( .A(n15757), .B(keyinput_f110), .ZN(n15764) );
  XNOR2_X1 U17278 ( .A(keyinput_f53), .B(n8621), .ZN(n15763) );
  XNOR2_X1 U17279 ( .A(SI_30_), .B(keyinput_f2), .ZN(n15761) );
  XNOR2_X1 U17280 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_f125), .ZN(n15760)
         );
  XNOR2_X1 U17281 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_f50), .ZN(n15759)
         );
  XNOR2_X1 U17282 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f127), .ZN(n15758)
         );
  NAND4_X1 U17283 ( .A1(n15761), .A2(n15760), .A3(n15759), .A4(n15758), .ZN(
        n15762) );
  NOR4_X1 U17284 ( .A1(n15765), .A2(n15764), .A3(n15763), .A4(n15762), .ZN(
        n15766) );
  NAND4_X1 U17285 ( .A1(n15769), .A2(n15768), .A3(n15767), .A4(n15766), .ZN(
        n15770) );
  OR4_X1 U17286 ( .A1(n15773), .A2(n15772), .A3(n15771), .A4(n15770), .ZN(
        n15775) );
  AOI21_X1 U17287 ( .B1(keyinput_f45), .B2(n15775), .A(keyinput_g45), .ZN(
        n15777) );
  INV_X1 U17288 ( .A(keyinput_f45), .ZN(n15774) );
  AOI21_X1 U17289 ( .B1(n15775), .B2(n15774), .A(n12506), .ZN(n15776) );
  AOI22_X1 U17290 ( .A1(n12506), .A2(n15777), .B1(keyinput_g45), .B2(n15776), 
        .ZN(n15778) );
  AOI21_X1 U17291 ( .B1(n15780), .B2(n15779), .A(n15778), .ZN(n15781) );
  XOR2_X1 U17292 ( .A(n15782), .B(n15781), .Z(n15784) );
  XOR2_X1 U17293 ( .A(n15787), .B(n15786), .Z(SUB_1596_U59) );
  XNOR2_X1 U17294 ( .A(n15788), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17295 ( .B1(n15790), .B2(n15789), .A(n15799), .ZN(SUB_1596_U53) );
  XNOR2_X1 U17296 ( .A(n15792), .B(n15791), .ZN(SUB_1596_U56) );
  AOI21_X1 U17297 ( .B1(n15795), .B2(n15794), .A(n15793), .ZN(n15797) );
  XNOR2_X1 U17298 ( .A(n15797), .B(n15796), .ZN(SUB_1596_U60) );
  XOR2_X1 U17299 ( .A(n15798), .B(n15799), .Z(SUB_1596_U5) );
  XNOR2_X1 U7768 ( .A(n8355), .B(n7387), .ZN(n8375) );
  OR2_X1 U9930 ( .A1(n14110), .A2(n14109), .ZN(n14344) );
  INV_X1 U10258 ( .A(n8267), .ZN(n8195) );
  CLKBUF_X2 U7432 ( .A(n9170), .Z(n9594) );
  CLKBUF_X1 U7433 ( .A(n11247), .Z(n6688) );
  CLKBUF_X1 U7438 ( .A(n13560), .Z(n6681) );
  CLKBUF_X1 U7440 ( .A(n9255), .Z(n9398) );
  CLKBUF_X2 U7451 ( .A(n9063), .Z(n9579) );
  CLKBUF_X1 U7473 ( .A(n13971), .Z(n6940) );
  NAND2_X1 U7504 ( .A1(n7220), .A2(n7219), .ZN(n11073) );
  CLKBUF_X2 U7542 ( .A(n7941), .Z(n11804) );
  CLKBUF_X1 U7913 ( .A(n14459), .Z(n6897) );
endmodule

